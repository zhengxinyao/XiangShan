module ICacheMainPipe(
  input          clock,
  input          reset,
  input          io_metaArray_toIMeta_ready,
  output         io_metaArray_toIMeta_valid,
  output         io_metaArray_toIMeta_bits_isDoubleLine,
  output [5:0]   io_metaArray_toIMeta_bits_vSetIdx_0,
  output [5:0]   io_metaArray_toIMeta_bits_vSetIdx_1,
  input  [1:0]   io_metaArray_fromIMeta_metaData_0_0_coh_state,
  input  [23:0]  io_metaArray_fromIMeta_metaData_0_0_tag,
  input  [1:0]   io_metaArray_fromIMeta_metaData_0_1_coh_state,
  input  [23:0]  io_metaArray_fromIMeta_metaData_0_1_tag,
  input  [1:0]   io_metaArray_fromIMeta_metaData_0_2_coh_state,
  input  [23:0]  io_metaArray_fromIMeta_metaData_0_2_tag,
  input  [1:0]   io_metaArray_fromIMeta_metaData_0_3_coh_state,
  input  [23:0]  io_metaArray_fromIMeta_metaData_0_3_tag,
  input  [1:0]   io_metaArray_fromIMeta_metaData_0_4_coh_state,
  input  [23:0]  io_metaArray_fromIMeta_metaData_0_4_tag,
  input  [1:0]   io_metaArray_fromIMeta_metaData_0_5_coh_state,
  input  [23:0]  io_metaArray_fromIMeta_metaData_0_5_tag,
  input  [1:0]   io_metaArray_fromIMeta_metaData_0_6_coh_state,
  input  [23:0]  io_metaArray_fromIMeta_metaData_0_6_tag,
  input  [1:0]   io_metaArray_fromIMeta_metaData_0_7_coh_state,
  input  [23:0]  io_metaArray_fromIMeta_metaData_0_7_tag,
  input  [1:0]   io_metaArray_fromIMeta_metaData_1_0_coh_state,
  input  [23:0]  io_metaArray_fromIMeta_metaData_1_0_tag,
  input  [1:0]   io_metaArray_fromIMeta_metaData_1_1_coh_state,
  input  [23:0]  io_metaArray_fromIMeta_metaData_1_1_tag,
  input  [1:0]   io_metaArray_fromIMeta_metaData_1_2_coh_state,
  input  [23:0]  io_metaArray_fromIMeta_metaData_1_2_tag,
  input  [1:0]   io_metaArray_fromIMeta_metaData_1_3_coh_state,
  input  [23:0]  io_metaArray_fromIMeta_metaData_1_3_tag,
  input  [1:0]   io_metaArray_fromIMeta_metaData_1_4_coh_state,
  input  [23:0]  io_metaArray_fromIMeta_metaData_1_4_tag,
  input  [1:0]   io_metaArray_fromIMeta_metaData_1_5_coh_state,
  input  [23:0]  io_metaArray_fromIMeta_metaData_1_5_tag,
  input  [1:0]   io_metaArray_fromIMeta_metaData_1_6_coh_state,
  input  [23:0]  io_metaArray_fromIMeta_metaData_1_6_tag,
  input  [1:0]   io_metaArray_fromIMeta_metaData_1_7_coh_state,
  input  [23:0]  io_metaArray_fromIMeta_metaData_1_7_tag,
  input          io_metaArray_fromIMeta_errors_0_0,
  input          io_metaArray_fromIMeta_errors_0_1,
  input          io_metaArray_fromIMeta_errors_0_2,
  input          io_metaArray_fromIMeta_errors_0_3,
  input          io_metaArray_fromIMeta_errors_0_4,
  input          io_metaArray_fromIMeta_errors_0_5,
  input          io_metaArray_fromIMeta_errors_0_6,
  input          io_metaArray_fromIMeta_errors_0_7,
  input          io_metaArray_fromIMeta_errors_1_0,
  input          io_metaArray_fromIMeta_errors_1_1,
  input          io_metaArray_fromIMeta_errors_1_2,
  input          io_metaArray_fromIMeta_errors_1_3,
  input          io_metaArray_fromIMeta_errors_1_4,
  input          io_metaArray_fromIMeta_errors_1_5,
  input          io_metaArray_fromIMeta_errors_1_6,
  input          io_metaArray_fromIMeta_errors_1_7,
  input          io_dataArray_toIData_ready,
  output         io_dataArray_toIData_valid,
  output         io_dataArray_toIData_bits_0_isDoubleLine,
  output [5:0]   io_dataArray_toIData_bits_0_vSetIdx_0,
  output [5:0]   io_dataArray_toIData_bits_0_vSetIdx_1,
  output         io_dataArray_toIData_bits_1_isDoubleLine,
  output [5:0]   io_dataArray_toIData_bits_1_vSetIdx_0,
  output [5:0]   io_dataArray_toIData_bits_1_vSetIdx_1,
  output         io_dataArray_toIData_bits_2_isDoubleLine,
  output [5:0]   io_dataArray_toIData_bits_2_vSetIdx_0,
  output [5:0]   io_dataArray_toIData_bits_2_vSetIdx_1,
  output         io_dataArray_toIData_bits_3_isDoubleLine,
  output [5:0]   io_dataArray_toIData_bits_3_vSetIdx_0,
  output [5:0]   io_dataArray_toIData_bits_3_vSetIdx_1,
  input  [511:0] io_dataArray_fromIData_datas_0_0,
  input  [511:0] io_dataArray_fromIData_datas_0_1,
  input  [511:0] io_dataArray_fromIData_datas_0_2,
  input  [511:0] io_dataArray_fromIData_datas_0_3,
  input  [511:0] io_dataArray_fromIData_datas_0_4,
  input  [511:0] io_dataArray_fromIData_datas_0_5,
  input  [511:0] io_dataArray_fromIData_datas_0_6,
  input  [511:0] io_dataArray_fromIData_datas_0_7,
  input  [511:0] io_dataArray_fromIData_datas_1_0,
  input  [511:0] io_dataArray_fromIData_datas_1_1,
  input  [511:0] io_dataArray_fromIData_datas_1_2,
  input  [511:0] io_dataArray_fromIData_datas_1_3,
  input  [511:0] io_dataArray_fromIData_datas_1_4,
  input  [511:0] io_dataArray_fromIData_datas_1_5,
  input  [511:0] io_dataArray_fromIData_datas_1_6,
  input  [511:0] io_dataArray_fromIData_datas_1_7,
  input  [31:0]  io_dataArray_fromIData_codes_0_0,
  input  [31:0]  io_dataArray_fromIData_codes_0_1,
  input  [31:0]  io_dataArray_fromIData_codes_0_2,
  input  [31:0]  io_dataArray_fromIData_codes_0_3,
  input  [31:0]  io_dataArray_fromIData_codes_0_4,
  input  [31:0]  io_dataArray_fromIData_codes_0_5,
  input  [31:0]  io_dataArray_fromIData_codes_0_6,
  input  [31:0]  io_dataArray_fromIData_codes_0_7,
  input  [31:0]  io_dataArray_fromIData_codes_1_0,
  input  [31:0]  io_dataArray_fromIData_codes_1_1,
  input  [31:0]  io_dataArray_fromIData_codes_1_2,
  input  [31:0]  io_dataArray_fromIData_codes_1_3,
  input  [31:0]  io_dataArray_fromIData_codes_1_4,
  input  [31:0]  io_dataArray_fromIData_codes_1_5,
  input  [31:0]  io_dataArray_fromIData_codes_1_6,
  input  [31:0]  io_dataArray_fromIData_codes_1_7,
  input          io_mshr_0_toMSHR_ready,
  output         io_mshr_0_toMSHR_valid,
  output [35:0]  io_mshr_0_toMSHR_bits_paddr,
  output [38:0]  io_mshr_0_toMSHR_bits_vaddr,
  output [7:0]   io_mshr_0_toMSHR_bits_waymask,
  input          io_mshr_0_fromMSHR_valid,
  input  [511:0] io_mshr_0_fromMSHR_bits_data,
  input          io_mshr_0_fromMSHR_bits_corrupt,
  input          io_mshr_1_toMSHR_ready,
  output         io_mshr_1_toMSHR_valid,
  output [35:0]  io_mshr_1_toMSHR_bits_paddr,
  output [38:0]  io_mshr_1_toMSHR_bits_vaddr,
  output [7:0]   io_mshr_1_toMSHR_bits_waymask,
  input          io_mshr_1_fromMSHR_valid,
  input  [511:0] io_mshr_1_fromMSHR_bits_data,
  input          io_mshr_1_fromMSHR_bits_corrupt,
  output         io_errors_0_source_tag,
  output         io_errors_0_source_data,
  output         io_errors_0_source_l2,
  output [35:0]  io_errors_0_paddr,
  output         io_errors_0_report_to_beu,
  output         io_errors_0_valid,
  output         io_errors_1_source_tag,
  output         io_errors_1_source_data,
  output         io_errors_1_source_l2,
  output [35:0]  io_errors_1_paddr,
  output         io_errors_1_report_to_beu,
  output         io_errors_1_valid,
  output         io_fetch_req_ready,
  input          io_fetch_req_valid,
  input  [38:0]  io_fetch_req_bits_pcMemRead_0_startAddr,
  input  [38:0]  io_fetch_req_bits_pcMemRead_0_nextlineStart,
  input  [38:0]  io_fetch_req_bits_pcMemRead_1_startAddr,
  input  [38:0]  io_fetch_req_bits_pcMemRead_1_nextlineStart,
  input  [38:0]  io_fetch_req_bits_pcMemRead_2_startAddr,
  input  [38:0]  io_fetch_req_bits_pcMemRead_2_nextlineStart,
  input  [38:0]  io_fetch_req_bits_pcMemRead_3_startAddr,
  input  [38:0]  io_fetch_req_bits_pcMemRead_3_nextlineStart,
  input  [38:0]  io_fetch_req_bits_pcMemRead_4_startAddr,
  input  [38:0]  io_fetch_req_bits_pcMemRead_4_nextlineStart,
  input          io_fetch_req_bits_readValid_0,
  input          io_fetch_req_bits_readValid_1,
  input          io_fetch_req_bits_readValid_2,
  input          io_fetch_req_bits_readValid_3,
  input          io_fetch_req_bits_readValid_4,
  output         io_fetch_resp_0_valid,
  output [38:0]  io_fetch_resp_0_bits_vaddr,
  output [511:0] io_fetch_resp_0_bits_registerData,
  output [511:0] io_fetch_resp_0_bits_sramData,
  output         io_fetch_resp_0_bits_select,
  output [35:0]  io_fetch_resp_0_bits_paddr,
  output         io_fetch_resp_0_bits_tlbExcp_pageFault,
  output         io_fetch_resp_0_bits_tlbExcp_accessFault,
  output         io_fetch_resp_0_bits_tlbExcp_mmio,
  output         io_fetch_resp_1_valid,
  output [38:0]  io_fetch_resp_1_bits_vaddr,
  output [511:0] io_fetch_resp_1_bits_registerData,
  output [511:0] io_fetch_resp_1_bits_sramData,
  output         io_fetch_resp_1_bits_select,
  output         io_fetch_resp_1_bits_tlbExcp_pageFault,
  output         io_fetch_resp_1_bits_tlbExcp_accessFault,
  output [35:0]  io_pmp_0_req_bits_addr,
  input          io_pmp_0_resp_instr,
  input          io_pmp_0_resp_mmio,
  output [35:0]  io_pmp_1_req_bits_addr,
  input          io_pmp_1_resp_instr,
  input          io_itlb_0_req_ready,
  output         io_itlb_0_req_valid,
  output [38:0]  io_itlb_0_req_bits_vaddr,
  output         io_itlb_0_req_bits_kill,
  output         io_itlb_0_resp_ready,
  input          io_itlb_0_resp_valid,
  input  [35:0]  io_itlb_0_resp_bits_paddr_0,
  input          io_itlb_0_resp_bits_excp_0_pf_instr,
  input          io_itlb_0_resp_bits_excp_0_af_instr,
  input          io_itlb_1_req_ready,
  output         io_itlb_1_req_valid,
  output [38:0]  io_itlb_1_req_bits_vaddr,
  output         io_itlb_1_req_bits_kill,
  output         io_itlb_1_resp_ready,
  input          io_itlb_1_resp_valid,
  input  [35:0]  io_itlb_1_resp_bits_paddr_0,
  input          io_itlb_1_resp_bits_excp_0_pf_instr,
  input          io_itlb_1_resp_bits_excp_0_af_instr,
  input          io_respStall,
  output         io_perfInfo_only_0_hit,
  output         io_perfInfo_only_0_miss,
  output         io_perfInfo_hit_0_hit_1,
  output         io_perfInfo_hit_0_miss_1,
  output         io_perfInfo_miss_0_hit_1,
  output         io_perfInfo_miss_0_miss_1,
  output         io_perfInfo_hit_0_except_1,
  output         io_perfInfo_miss_0_except_1,
  output         io_perfInfo_except_0,
  output         io_perfInfo_bank_hit_1,
  output         io_perfInfo_hit,
  input          io_csr_parity_enable
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [63:0] _RAND_39;
  reg [63:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [63:0] _RAND_44;
  reg [63:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [511:0] _RAND_102;
  reg [511:0] _RAND_103;
  reg [511:0] _RAND_104;
  reg [511:0] _RAND_105;
  reg [511:0] _RAND_106;
  reg [511:0] _RAND_107;
  reg [511:0] _RAND_108;
  reg [511:0] _RAND_109;
  reg [511:0] _RAND_110;
  reg [511:0] _RAND_111;
  reg [511:0] _RAND_112;
  reg [511:0] _RAND_113;
  reg [511:0] _RAND_114;
  reg [511:0] _RAND_115;
  reg [511:0] _RAND_116;
  reg [511:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [63:0] _RAND_222;
  reg [63:0] _RAND_223;
  reg [63:0] _RAND_224;
  reg [63:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [511:0] _RAND_258;
  reg [511:0] _RAND_259;
  reg [511:0] _RAND_260;
  reg [511:0] _RAND_261;
  reg [511:0] _RAND_262;
  reg [511:0] _RAND_263;
  reg [511:0] _RAND_264;
  reg [511:0] _RAND_265;
  reg [511:0] _RAND_266;
  reg [511:0] _RAND_267;
  reg [511:0] _RAND_268;
  reg [511:0] _RAND_269;
  reg [511:0] _RAND_270;
  reg [511:0] _RAND_271;
  reg [511:0] _RAND_272;
  reg [511:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
  reg [31:0] _RAND_726;
  reg [31:0] _RAND_727;
  reg [31:0] _RAND_728;
  reg [31:0] _RAND_729;
  reg [31:0] _RAND_730;
  reg [31:0] _RAND_731;
  reg [31:0] _RAND_732;
  reg [31:0] _RAND_733;
  reg [31:0] _RAND_734;
  reg [31:0] _RAND_735;
  reg [31:0] _RAND_736;
  reg [31:0] _RAND_737;
  reg [31:0] _RAND_738;
  reg [31:0] _RAND_739;
  reg [31:0] _RAND_740;
  reg [31:0] _RAND_741;
  reg [31:0] _RAND_742;
  reg [31:0] _RAND_743;
  reg [31:0] _RAND_744;
  reg [31:0] _RAND_745;
  reg [31:0] _RAND_746;
  reg [31:0] _RAND_747;
  reg [31:0] _RAND_748;
  reg [31:0] _RAND_749;
  reg [31:0] _RAND_750;
  reg [31:0] _RAND_751;
  reg [31:0] _RAND_752;
  reg [31:0] _RAND_753;
  reg [31:0] _RAND_754;
  reg [31:0] _RAND_755;
  reg [31:0] _RAND_756;
  reg [31:0] _RAND_757;
  reg [31:0] _RAND_758;
  reg [31:0] _RAND_759;
  reg [31:0] _RAND_760;
  reg [31:0] _RAND_761;
  reg [31:0] _RAND_762;
  reg [31:0] _RAND_763;
  reg [31:0] _RAND_764;
  reg [31:0] _RAND_765;
  reg [31:0] _RAND_766;
  reg [31:0] _RAND_767;
  reg [31:0] _RAND_768;
  reg [31:0] _RAND_769;
  reg [31:0] _RAND_770;
  reg [31:0] _RAND_771;
  reg [31:0] _RAND_772;
  reg [31:0] _RAND_773;
  reg [31:0] _RAND_774;
  reg [31:0] _RAND_775;
  reg [31:0] _RAND_776;
  reg [31:0] _RAND_777;
  reg [31:0] _RAND_778;
  reg [31:0] _RAND_779;
  reg [31:0] _RAND_780;
  reg [31:0] _RAND_781;
  reg [31:0] _RAND_782;
  reg [31:0] _RAND_783;
  reg [31:0] _RAND_784;
  reg [31:0] _RAND_785;
  reg [31:0] _RAND_786;
  reg [31:0] _RAND_787;
  reg [31:0] _RAND_788;
  reg [31:0] _RAND_789;
  reg [31:0] _RAND_790;
  reg [31:0] _RAND_791;
  reg [31:0] _RAND_792;
  reg [31:0] _RAND_793;
  reg [31:0] _RAND_794;
  reg [31:0] _RAND_795;
  reg [31:0] _RAND_796;
  reg [31:0] _RAND_797;
  reg [31:0] _RAND_798;
  reg [31:0] _RAND_799;
  reg [31:0] _RAND_800;
  reg [31:0] _RAND_801;
  reg [31:0] _RAND_802;
  reg [31:0] _RAND_803;
  reg [31:0] _RAND_804;
  reg [31:0] _RAND_805;
  reg [31:0] _RAND_806;
  reg [31:0] _RAND_807;
  reg [31:0] _RAND_808;
  reg [31:0] _RAND_809;
  reg [31:0] _RAND_810;
  reg [31:0] _RAND_811;
  reg [31:0] _RAND_812;
  reg [31:0] _RAND_813;
  reg [31:0] _RAND_814;
  reg [31:0] _RAND_815;
  reg [31:0] _RAND_816;
  reg [31:0] _RAND_817;
  reg [31:0] _RAND_818;
  reg [31:0] _RAND_819;
  reg [31:0] _RAND_820;
  reg [31:0] _RAND_821;
  reg [31:0] _RAND_822;
  reg [31:0] _RAND_823;
  reg [31:0] _RAND_824;
  reg [31:0] _RAND_825;
  reg [31:0] _RAND_826;
  reg [31:0] _RAND_827;
  reg [31:0] _RAND_828;
  reg [31:0] _RAND_829;
  reg [31:0] _RAND_830;
  reg [31:0] _RAND_831;
  reg [31:0] _RAND_832;
  reg [31:0] _RAND_833;
  reg [31:0] _RAND_834;
  reg [31:0] _RAND_835;
  reg [31:0] _RAND_836;
  reg [31:0] _RAND_837;
  reg [31:0] _RAND_838;
  reg [31:0] _RAND_839;
  reg [31:0] _RAND_840;
  reg [31:0] _RAND_841;
  reg [63:0] _RAND_842;
  reg [63:0] _RAND_843;
  reg [31:0] _RAND_844;
  reg [31:0] _RAND_845;
  reg [31:0] _RAND_846;
  reg [31:0] _RAND_847;
  reg [31:0] _RAND_848;
  reg [31:0] _RAND_849;
  reg [31:0] _RAND_850;
  reg [31:0] _RAND_851;
  reg [31:0] _RAND_852;
  reg [63:0] _RAND_853;
  reg [63:0] _RAND_854;
  reg [31:0] _RAND_855;
  reg [31:0] _RAND_856;
  reg [31:0] _RAND_857;
  reg [31:0] _RAND_858;
  reg [31:0] _RAND_859;
  reg [31:0] _RAND_860;
  reg [31:0] _RAND_861;
  reg [31:0] _RAND_862;
  reg [31:0] _RAND_863;
  reg [31:0] _RAND_864;
  reg [31:0] _RAND_865;
  reg [31:0] _RAND_866;
  reg [511:0] _RAND_867;
  reg [31:0] _RAND_868;
  reg [31:0] _RAND_869;
  reg [31:0] _RAND_870;
  reg [511:0] _RAND_871;
  reg [31:0] _RAND_872;
  reg [31:0] _RAND_873;
  reg [31:0] _RAND_874;
  reg [31:0] _RAND_875;
  reg [31:0] _RAND_876;
  reg [31:0] _RAND_877;
  reg [31:0] _RAND_878;
  reg [31:0] _RAND_879;
  reg [31:0] _RAND_880;
  reg [31:0] _RAND_881;
  reg [31:0] _RAND_882;
  reg [31:0] _RAND_883;
  reg [31:0] _RAND_884;
  reg [31:0] _RAND_885;
  reg [31:0] _RAND_886;
  reg [511:0] _RAND_887;
  reg [511:0] _RAND_888;
  reg [31:0] _RAND_889;
  reg [63:0] _RAND_890;
  reg [31:0] _RAND_891;
  reg [63:0] _RAND_892;
`endif // RANDOMIZE_REG_INIT
  reg  missSwitchBit; // @[ICacheMainPipe.scala 133:30]
  wire [5:0] ftq_req_to_data_vset_idx_0_0 = io_fetch_req_bits_pcMemRead_0_startAddr[11:6]; // @[L1Cache.scala 81:33]
  wire [5:0] ftq_req_to_data_vset_idx_0_1 = io_fetch_req_bits_pcMemRead_0_nextlineStart[11:6]; // @[L1Cache.scala 81:33]
  wire  ftq_req_to_data_doubleline_0 = io_fetch_req_bits_readValid_0 & io_fetch_req_bits_pcMemRead_0_startAddr[5]; // @[ICacheMainPipe.scala 152:84]
  wire  ftq_req_to_itlb_doubleline = io_fetch_req_bits_readValid_4 & io_fetch_req_bits_pcMemRead_4_startAddr[5]; // @[ICacheMainPipe.scala 152:84]
  wire  _io_dataArray_toIData_valid_T = ~missSwitchBit; // @[ICacheMainPipe.scala 176:66]
  wire  itlb_can_go = io_itlb_0_req_ready & io_itlb_1_req_ready; // @[ICacheMainPipe.scala 211:40]
  wire  icache_can_go = io_dataArray_toIData_ready & io_metaArray_toIMeta_ready; // @[ICacheMainPipe.scala 212:37]
  reg  s2_valid; // @[ICache.scala 98:25]
  reg  s2_port_hit_0; // @[Reg.scala 16:16]
  reg  miss_0_s2_0_latch_bit; // @[ICacheMainPipe.scala 478:22]
  reg  miss_0_s2_0_REG; // @[ICacheMainPipe.scala 504:12]
  reg  miss_0_s2_0_REG_1; // @[ICacheMainPipe.scala 505:12]
  wire  _miss_0_s2_0_T_1 = miss_0_s2_0_REG & miss_0_s2_0_REG_1; // @[ICacheMainPipe.scala 504:22]
  reg  miss_0_s2_0_REG_2; // @[ICacheMainPipe.scala 506:12]
  wire  _miss_0_s2_0_T_3 = _miss_0_s2_0_T_1 & miss_0_s2_0_REG_2; // @[ICacheMainPipe.scala 505:70]
  wire  _miss_0_s2_0_T_4 = ~s2_port_hit_0; // @[ICacheMainPipe.scala 507:5]
  wire  _miss_0_s2_0_T_5 = _miss_0_s2_0_T_3 & _miss_0_s2_0_T_4; // @[ICacheMainPipe.scala 506:66]
  reg [2:0] missStateQueue_0; // @[ICacheMainPipe.scala 449:31]
  wire  _miss_0_s2_0_T_6 = missStateQueue_0 == 3'h4; // @[ICacheMainPipe.scala 501:60]
  wire  miss_0_s2_0 = _miss_0_s2_0_T_5 & _miss_0_s2_0_T_6; // @[ICacheMainPipe.scala 507:28]
  wire  miss_0_s2_0_latch = miss_0_s2_0_latch_bit | miss_0_s2_0; // @[ICacheMainPipe.scala 482:9]
  reg  miss_1_s2_0_latch_bit; // @[ICacheMainPipe.scala 478:22]
  reg  miss_1_s2_0_REG; // @[ICacheMainPipe.scala 504:12]
  reg  miss_1_s2_0_REG_1; // @[ICacheMainPipe.scala 505:12]
  wire  _miss_1_s2_0_T_1 = miss_1_s2_0_REG & miss_1_s2_0_REG_1; // @[ICacheMainPipe.scala 504:22]
  reg  miss_1_s2_0_REG_2; // @[ICacheMainPipe.scala 506:12]
  wire  _miss_1_s2_0_T_3 = _miss_1_s2_0_T_1 & miss_1_s2_0_REG_2; // @[ICacheMainPipe.scala 505:70]
  wire  _miss_1_s2_0_T_5 = _miss_1_s2_0_T_3 & _miss_0_s2_0_T_4; // @[ICacheMainPipe.scala 506:66]
  reg [2:0] missStateQueue_1; // @[ICacheMainPipe.scala 449:31]
  wire  _miss_1_s2_0_T_6 = missStateQueue_1 == 3'h4; // @[ICacheMainPipe.scala 501:60]
  wire  miss_1_s2_0 = _miss_1_s2_0_T_5 & _miss_1_s2_0_T_6; // @[ICacheMainPipe.scala 507:28]
  wire  miss_1_s2_0_latch = miss_1_s2_0_latch_bit | miss_1_s2_0; // @[ICacheMainPipe.scala 482:9]
  wire  sec_meet_0_miss = miss_0_s2_0_latch | miss_1_s2_0_latch; // @[ICacheMainPipe.scala 455:41]
  wire  s2_fixed_hit_vec_0 = s2_port_hit_0 | sec_meet_0_miss; // @[ICacheMainPipe.scala 359:70]
  reg  s2_port_hit_1; // @[Reg.scala 16:16]
  reg  miss_0_s2_1_latch_bit; // @[ICacheMainPipe.scala 478:22]
  reg  miss_0_s2_1_REG; // @[ICacheMainPipe.scala 504:12]
  reg  miss_0_s2_1_REG_1; // @[ICacheMainPipe.scala 505:12]
  wire  _miss_0_s2_1_T_1 = miss_0_s2_1_REG & miss_0_s2_1_REG_1; // @[ICacheMainPipe.scala 504:22]
  reg  miss_0_s2_1_REG_2; // @[ICacheMainPipe.scala 506:12]
  wire  _miss_0_s2_1_T_3 = _miss_0_s2_1_T_1 & miss_0_s2_1_REG_2; // @[ICacheMainPipe.scala 505:70]
  wire  _miss_0_s2_1_T_4 = ~s2_port_hit_1; // @[ICacheMainPipe.scala 507:5]
  wire  _miss_0_s2_1_T_5 = _miss_0_s2_1_T_3 & _miss_0_s2_1_T_4; // @[ICacheMainPipe.scala 506:66]
  wire  miss_0_s2_1 = _miss_0_s2_1_T_5 & _miss_0_s2_0_T_6; // @[ICacheMainPipe.scala 507:28]
  wire  miss_0_s2_1_latch = miss_0_s2_1_latch_bit | miss_0_s2_1; // @[ICacheMainPipe.scala 482:9]
  reg  miss_1_s2_1_latch_bit; // @[ICacheMainPipe.scala 478:22]
  reg  miss_1_s2_1_REG; // @[ICacheMainPipe.scala 504:12]
  reg  miss_1_s2_1_REG_1; // @[ICacheMainPipe.scala 505:12]
  wire  _miss_1_s2_1_T_1 = miss_1_s2_1_REG & miss_1_s2_1_REG_1; // @[ICacheMainPipe.scala 504:22]
  reg  miss_1_s2_1_REG_2; // @[ICacheMainPipe.scala 506:12]
  wire  _miss_1_s2_1_T_3 = _miss_1_s2_1_T_1 & miss_1_s2_1_REG_2; // @[ICacheMainPipe.scala 505:70]
  wire  _miss_1_s2_1_T_5 = _miss_1_s2_1_T_3 & _miss_0_s2_1_T_4; // @[ICacheMainPipe.scala 506:66]
  wire  miss_1_s2_1 = _miss_1_s2_1_T_5 & _miss_1_s2_0_T_6; // @[ICacheMainPipe.scala 507:28]
  wire  miss_1_s2_1_latch = miss_1_s2_1_latch_bit | miss_1_s2_1; // @[ICacheMainPipe.scala 482:9]
  wire  sec_meet_1_miss = miss_0_s2_1_latch | miss_1_s2_1_latch; // @[ICacheMainPipe.scala 456:41]
  wire  s2_fixed_hit_vec_1 = s2_port_hit_1 | sec_meet_1_miss; // @[ICacheMainPipe.scala 359:70]
  reg  s2_double_line; // @[Reg.scala 16:16]
  wire  _s2_fixed_hit_T_4 = ~s2_double_line; // @[ICacheMainPipe.scala 360:136]
  wire  s2_fixed_hit = s2_valid & s2_fixed_hit_vec_0 & s2_fixed_hit_vec_1 & s2_double_line | s2_valid &
    s2_fixed_hit_vec_0 & ~s2_double_line; // @[ICacheMainPipe.scala 360:97]
  reg [3:0] wait_state; // @[ICacheMainPipe.scala 435:27]
  wire  miss_all_fix = wait_state == 4'h7; // @[ICacheMainPipe.scala 665:40]
  reg  hit_0_except_1_latch_bit; // @[ICacheMainPipe.scala 478:22]
  reg  hit_0_except_1_REG; // @[ICacheMainPipe.scala 473:34]
  reg  s2_except_pf_0; // @[Reg.scala 16:16]
  reg  s2_except_tlb_af_0; // @[Reg.scala 16:16]
  wire  s2_except_0 = s2_except_pf_0 | s2_except_tlb_af_0; // @[ICacheMainPipe.scala 420:67]
  wire  _hit_0_except_1_T_1 = ~s2_except_0; // @[ICacheMainPipe.scala 473:66]
  reg  s2_except_pf_1; // @[Reg.scala 16:16]
  reg  s2_except_tlb_af_1; // @[Reg.scala 16:16]
  wire  s2_except_1 = s2_except_pf_1 | s2_except_tlb_af_1; // @[ICacheMainPipe.scala 420:67]
  wire  hit_0_except_1 = hit_0_except_1_REG & s2_double_line & ~s2_except_0 & s2_except_1 & s2_fixed_hit_vec_0; // @[ICacheMainPipe.scala 473:97]
  wire  hit_0_except_1_latch = hit_0_except_1_latch_bit | hit_0_except_1; // @[ICacheMainPipe.scala 482:9]
  reg  except_0_latch_bit; // @[ICacheMainPipe.scala 478:22]
  reg  except_0_REG; // @[ICacheMainPipe.scala 475:34]
  wire  except_0 = except_0_REG & s2_except_0; // @[ICacheMainPipe.scala 475:44]
  wire  except_0_latch = except_0_latch_bit | except_0; // @[ICacheMainPipe.scala 482:9]
  wire  s2_fetch_finish = s2_valid & s2_fixed_hit | miss_all_fix | hit_0_except_1_latch | except_0_latch; // @[ICacheMainPipe.scala 667:97]
  wire  _s2_ready_T = s2_valid & s2_fetch_finish; // @[ICacheMainPipe.scala 337:30]
  wire  _s2_ready_T_1 = ~io_respStall; // @[ICacheMainPipe.scala 337:52]
  wire  _s2_ready_T_2 = s2_valid & s2_fetch_finish & ~io_respStall; // @[ICacheMainPipe.scala 337:49]
  wire  _s2_miss_available_T = missStateQueue_0 == 3'h0; // @[ICacheMainPipe.scala 452:67]
  wire  _s2_miss_available_T_3 = missStateQueue_1 == 3'h0; // @[ICacheMainPipe.scala 452:67]
  wire  s2_miss_available = (missStateQueue_0 == 3'h0 | _miss_0_s2_0_T_6) & (missStateQueue_1 == 3'h0 | _miss_1_s2_0_T_6
    ); // @[ICacheMainPipe.scala 452:121]
  wire  s2_ready = s2_valid & s2_fetch_finish & ~io_respStall | ~s2_valid & s2_miss_available; // @[ICacheMainPipe.scala 337:67]
  reg  tlb_need_back_valid; // @[Hold.scala 40:24]
  reg  tlb_already_recv_0; // @[ICacheMainPipe.scala 243:33]
  reg  tlb_ready_recv_REG; // @[ICacheMainPipe.scala 244:69]
  reg  s1_valid; // @[ICache.scala 98:25]
  wire  tlb_ready_recv_0 = tlb_ready_recv_REG | s1_valid & ~tlb_already_recv_0; // @[ICacheMainPipe.scala 244:88]
  wire  tlb_back_0 = io_itlb_0_resp_ready & io_itlb_0_resp_valid; // @[Decoupled.scala 50:35]
  wire  tlb_resp_valid_0 = tlb_already_recv_0 | tlb_ready_recv_0 & tlb_back_0; // @[ICacheMainPipe.scala 247:46]
  wire  _tlbRespAllValid_T_1 = ~tlb_need_back_valid | tlb_resp_valid_0; // @[ICacheMainPipe.scala 268:77]
  reg  tlb_need_back_valid_1; // @[Hold.scala 40:24]
  reg  tlb_already_recv_1; // @[ICacheMainPipe.scala 243:33]
  reg  tlb_ready_recv_REG_1; // @[ICacheMainPipe.scala 244:69]
  wire  tlb_ready_recv_1 = tlb_ready_recv_REG_1 | s1_valid & ~tlb_already_recv_1; // @[ICacheMainPipe.scala 244:88]
  wire  tlb_back_1 = io_itlb_1_resp_ready & io_itlb_1_resp_valid; // @[Decoupled.scala 50:35]
  wire  tlb_resp_valid_1 = tlb_already_recv_1 | tlb_ready_recv_1 & tlb_back_1; // @[ICacheMainPipe.scala 247:46]
  wire  _tlbRespAllValid_T_3 = ~tlb_need_back_valid_1 | tlb_resp_valid_1; // @[ICacheMainPipe.scala 268:77]
  wire [1:0] _tlbRespAllValid_T_4 = {_tlbRespAllValid_T_1,_tlbRespAllValid_T_3}; // @[Cat.scala 31:58]
  wire  tlbRespAllValid = &_tlbRespAllValid_T_4; // @[ICacheMainPipe.scala 268:100]
  wire  s1_ready = s2_ready & tlbRespAllValid | ~s1_valid; // @[ICacheMainPipe.scala 269:44]
  wire  pipe_can_go = _io_dataArray_toIData_valid_T & s1_ready; // @[ICacheMainPipe.scala 213:39]
  wire  s0_can_go = itlb_can_go & icache_can_go & pipe_can_go; // @[ICacheMainPipe.scala 214:53]
  wire  s0_fetch_fire = io_fetch_req_valid & s0_can_go; // @[ICacheMainPipe.scala 215:33]
  wire  s1_fire = s1_valid & tlbRespAllValid & s2_ready; // @[ICacheMainPipe.scala 270:43]
  wire  _GEN_0 = s1_fire ? 1'h0 : s1_valid; // @[ICache.scala 101:{43,51} 98:25]
  reg [38:0] s1_req_vaddr_0; // @[Reg.scala 16:16]
  reg [38:0] s1_req_vaddr_1; // @[Reg.scala 16:16]
  reg [5:0] s1_req_vsetIdx_0; // @[Reg.scala 16:16]
  reg [5:0] s1_req_vsetIdx_1; // @[Reg.scala 16:16]
  reg  s1_double_line; // @[Reg.scala 16:16]
  wire  _tlb_need_back_T = io_itlb_0_req_ready & io_itlb_0_req_valid; // @[Decoupled.scala 50:35]
  wire  _tlb_need_back_T_1 = s0_fetch_fire & _tlb_need_back_T; // @[ICacheMainPipe.scala 242:79]
  wire  _GEN_9 = s1_fire ? 1'h0 : tlb_need_back_valid; // @[Hold.scala 41:20 40:24 41:28]
  wire  _tlb_need_back_T_2 = io_itlb_1_req_ready & io_itlb_1_req_valid; // @[Decoupled.scala 50:35]
  wire  _tlb_need_back_T_3 = s0_fetch_fire & _tlb_need_back_T_2; // @[ICacheMainPipe.scala 242:79]
  wire  _GEN_12 = s1_fire ? 1'h0 : tlb_need_back_valid_1; // @[Hold.scala 41:20 40:24 41:28]
  wire  _GEN_15 = tlb_already_recv_0 & s1_fire ? 1'h0 : tlb_already_recv_0; // @[ICacheMainPipe.scala 248:43 249:27 243:33]
  wire  _GEN_17 = tlb_already_recv_1 & s1_fire ? 1'h0 : tlb_already_recv_1; // @[ICacheMainPipe.scala 248:43 249:27 243:33]
  reg [35:0] tlbRespPAddr_r; // @[Reg.scala 16:16]
  wire [35:0] _GEN_19 = tlb_back_0 ? io_itlb_0_resp_bits_paddr_0 : tlbRespPAddr_r; // @[Reg.scala 16:16 17:{18,22}]
  reg [35:0] tlbRespPAddr_r1; // @[Reg.scala 16:16]
  wire [35:0] _GEN_20 = tlb_back_1 ? io_itlb_1_resp_bits_paddr_0 : tlbRespPAddr_r1; // @[Reg.scala 16:16 17:{18,22}]
  reg  tlbExcpPF_r; // @[Reg.scala 16:16]
  wire  _GEN_21 = tlb_back_0 ? io_itlb_0_resp_bits_excp_0_pf_instr : tlbExcpPF_r; // @[Reg.scala 16:16 17:{18,22}]
  wire  tlbExcpPF_0 = _GEN_21 & tlb_need_back_valid; // @[ICacheMainPipe.scala 264:137]
  reg  tlbExcpPF_r1; // @[Reg.scala 16:16]
  wire  _GEN_22 = tlb_back_1 ? io_itlb_1_resp_bits_excp_0_pf_instr : tlbExcpPF_r1; // @[Reg.scala 16:16 17:{18,22}]
  wire  tlbExcpPF_1 = _GEN_22 & tlb_need_back_valid_1; // @[ICacheMainPipe.scala 264:137]
  reg  tlbExcpAF_r; // @[Reg.scala 16:16]
  wire  _GEN_23 = tlb_back_0 ? io_itlb_0_resp_bits_excp_0_af_instr : tlbExcpAF_r; // @[Reg.scala 16:16 17:{18,22}]
  wire  tlbExcpAF_0 = _GEN_23 & tlb_need_back_valid; // @[ICacheMainPipe.scala 265:137]
  reg  tlbExcpAF_r1; // @[Reg.scala 16:16]
  wire  _GEN_24 = tlb_back_1 ? io_itlb_1_resp_bits_excp_0_af_instr : tlbExcpAF_r1; // @[Reg.scala 16:16 17:{18,22}]
  wire  tlbExcpAF_1 = _GEN_24 & tlb_need_back_valid_1; // @[ICacheMainPipe.scala 265:137]
  wire [23:0] s1_req_ptags_0 = _GEN_19[35:12]; // @[L1Cache.scala 79:41]
  wire [23:0] s1_req_ptags_1 = _GEN_20[35:12]; // @[L1Cache.scala 79:41]
  reg  s1_meta_ptags_REG; // @[ICacheMainPipe.scala 276:90]
  reg [23:0] s1_meta_ptags_r0_0; // @[Reg.scala 16:16]
  reg [23:0] s1_meta_ptags_r0_1; // @[Reg.scala 16:16]
  reg [23:0] s1_meta_ptags_r0_2; // @[Reg.scala 16:16]
  reg [23:0] s1_meta_ptags_r0_3; // @[Reg.scala 16:16]
  reg [23:0] s1_meta_ptags_r0_4; // @[Reg.scala 16:16]
  reg [23:0] s1_meta_ptags_r0_5; // @[Reg.scala 16:16]
  reg [23:0] s1_meta_ptags_r0_6; // @[Reg.scala 16:16]
  reg [23:0] s1_meta_ptags_r0_7; // @[Reg.scala 16:16]
  reg [23:0] s1_meta_ptags_r1_0; // @[Reg.scala 16:16]
  reg [23:0] s1_meta_ptags_r1_1; // @[Reg.scala 16:16]
  reg [23:0] s1_meta_ptags_r1_2; // @[Reg.scala 16:16]
  reg [23:0] s1_meta_ptags_r1_3; // @[Reg.scala 16:16]
  reg [23:0] s1_meta_ptags_r1_4; // @[Reg.scala 16:16]
  reg [23:0] s1_meta_ptags_r1_5; // @[Reg.scala 16:16]
  reg [23:0] s1_meta_ptags_r1_6; // @[Reg.scala 16:16]
  reg [23:0] s1_meta_ptags_r1_7; // @[Reg.scala 16:16]
  wire [23:0] _GEN_25 = s1_meta_ptags_REG ? io_metaArray_fromIMeta_metaData_0_0_tag : s1_meta_ptags_r0_0; // @[Reg.scala 16:16 17:{18,22}]
  wire [23:0] _GEN_26 = s1_meta_ptags_REG ? io_metaArray_fromIMeta_metaData_0_1_tag : s1_meta_ptags_r0_1; // @[Reg.scala 16:16 17:{18,22}]
  wire [23:0] _GEN_27 = s1_meta_ptags_REG ? io_metaArray_fromIMeta_metaData_0_2_tag : s1_meta_ptags_r0_2; // @[Reg.scala 16:16 17:{18,22}]
  wire [23:0] _GEN_28 = s1_meta_ptags_REG ? io_metaArray_fromIMeta_metaData_0_3_tag : s1_meta_ptags_r0_3; // @[Reg.scala 16:16 17:{18,22}]
  wire [23:0] _GEN_29 = s1_meta_ptags_REG ? io_metaArray_fromIMeta_metaData_0_4_tag : s1_meta_ptags_r0_4; // @[Reg.scala 16:16 17:{18,22}]
  wire [23:0] _GEN_30 = s1_meta_ptags_REG ? io_metaArray_fromIMeta_metaData_0_5_tag : s1_meta_ptags_r0_5; // @[Reg.scala 16:16 17:{18,22}]
  wire [23:0] _GEN_31 = s1_meta_ptags_REG ? io_metaArray_fromIMeta_metaData_0_6_tag : s1_meta_ptags_r0_6; // @[Reg.scala 16:16 17:{18,22}]
  wire [23:0] _GEN_32 = s1_meta_ptags_REG ? io_metaArray_fromIMeta_metaData_0_7_tag : s1_meta_ptags_r0_7; // @[Reg.scala 16:16 17:{18,22}]
  wire [23:0] _GEN_33 = s1_meta_ptags_REG ? io_metaArray_fromIMeta_metaData_1_0_tag : s1_meta_ptags_r1_0; // @[Reg.scala 16:16 17:{18,22}]
  wire [23:0] _GEN_34 = s1_meta_ptags_REG ? io_metaArray_fromIMeta_metaData_1_1_tag : s1_meta_ptags_r1_1; // @[Reg.scala 16:16 17:{18,22}]
  wire [23:0] _GEN_35 = s1_meta_ptags_REG ? io_metaArray_fromIMeta_metaData_1_2_tag : s1_meta_ptags_r1_2; // @[Reg.scala 16:16 17:{18,22}]
  wire [23:0] _GEN_36 = s1_meta_ptags_REG ? io_metaArray_fromIMeta_metaData_1_3_tag : s1_meta_ptags_r1_3; // @[Reg.scala 16:16 17:{18,22}]
  wire [23:0] _GEN_37 = s1_meta_ptags_REG ? io_metaArray_fromIMeta_metaData_1_4_tag : s1_meta_ptags_r1_4; // @[Reg.scala 16:16 17:{18,22}]
  wire [23:0] _GEN_38 = s1_meta_ptags_REG ? io_metaArray_fromIMeta_metaData_1_5_tag : s1_meta_ptags_r1_5; // @[Reg.scala 16:16 17:{18,22}]
  wire [23:0] _GEN_39 = s1_meta_ptags_REG ? io_metaArray_fromIMeta_metaData_1_6_tag : s1_meta_ptags_r1_6; // @[Reg.scala 16:16 17:{18,22}]
  wire [23:0] _GEN_40 = s1_meta_ptags_REG ? io_metaArray_fromIMeta_metaData_1_7_tag : s1_meta_ptags_r1_7; // @[Reg.scala 16:16 17:{18,22}]
  reg  s1_meta_cohs_REG; // @[ICacheMainPipe.scala 277:90]
  reg [1:0] s1_meta_cohs_r0_0_state; // @[Reg.scala 16:16]
  reg [1:0] s1_meta_cohs_r0_1_state; // @[Reg.scala 16:16]
  reg [1:0] s1_meta_cohs_r0_2_state; // @[Reg.scala 16:16]
  reg [1:0] s1_meta_cohs_r0_3_state; // @[Reg.scala 16:16]
  reg [1:0] s1_meta_cohs_r0_4_state; // @[Reg.scala 16:16]
  reg [1:0] s1_meta_cohs_r0_5_state; // @[Reg.scala 16:16]
  reg [1:0] s1_meta_cohs_r0_6_state; // @[Reg.scala 16:16]
  reg [1:0] s1_meta_cohs_r0_7_state; // @[Reg.scala 16:16]
  reg [1:0] s1_meta_cohs_r1_0_state; // @[Reg.scala 16:16]
  reg [1:0] s1_meta_cohs_r1_1_state; // @[Reg.scala 16:16]
  reg [1:0] s1_meta_cohs_r1_2_state; // @[Reg.scala 16:16]
  reg [1:0] s1_meta_cohs_r1_3_state; // @[Reg.scala 16:16]
  reg [1:0] s1_meta_cohs_r1_4_state; // @[Reg.scala 16:16]
  reg [1:0] s1_meta_cohs_r1_5_state; // @[Reg.scala 16:16]
  reg [1:0] s1_meta_cohs_r1_6_state; // @[Reg.scala 16:16]
  reg [1:0] s1_meta_cohs_r1_7_state; // @[Reg.scala 16:16]
  wire [1:0] _GEN_41 = s1_meta_cohs_REG ? io_metaArray_fromIMeta_metaData_0_0_coh_state : s1_meta_cohs_r0_0_state; // @[Reg.scala 16:16 17:{18,22}]
  wire [1:0] _GEN_42 = s1_meta_cohs_REG ? io_metaArray_fromIMeta_metaData_0_1_coh_state : s1_meta_cohs_r0_1_state; // @[Reg.scala 16:16 17:{18,22}]
  wire [1:0] _GEN_43 = s1_meta_cohs_REG ? io_metaArray_fromIMeta_metaData_0_2_coh_state : s1_meta_cohs_r0_2_state; // @[Reg.scala 16:16 17:{18,22}]
  wire [1:0] _GEN_44 = s1_meta_cohs_REG ? io_metaArray_fromIMeta_metaData_0_3_coh_state : s1_meta_cohs_r0_3_state; // @[Reg.scala 16:16 17:{18,22}]
  wire [1:0] _GEN_45 = s1_meta_cohs_REG ? io_metaArray_fromIMeta_metaData_0_4_coh_state : s1_meta_cohs_r0_4_state; // @[Reg.scala 16:16 17:{18,22}]
  wire [1:0] _GEN_46 = s1_meta_cohs_REG ? io_metaArray_fromIMeta_metaData_0_5_coh_state : s1_meta_cohs_r0_5_state; // @[Reg.scala 16:16 17:{18,22}]
  wire [1:0] _GEN_47 = s1_meta_cohs_REG ? io_metaArray_fromIMeta_metaData_0_6_coh_state : s1_meta_cohs_r0_6_state; // @[Reg.scala 16:16 17:{18,22}]
  wire [1:0] _GEN_48 = s1_meta_cohs_REG ? io_metaArray_fromIMeta_metaData_0_7_coh_state : s1_meta_cohs_r0_7_state; // @[Reg.scala 16:16 17:{18,22}]
  wire [1:0] _GEN_49 = s1_meta_cohs_REG ? io_metaArray_fromIMeta_metaData_1_0_coh_state : s1_meta_cohs_r1_0_state; // @[Reg.scala 16:16 17:{18,22}]
  wire [1:0] _GEN_50 = s1_meta_cohs_REG ? io_metaArray_fromIMeta_metaData_1_1_coh_state : s1_meta_cohs_r1_1_state; // @[Reg.scala 16:16 17:{18,22}]
  wire [1:0] _GEN_51 = s1_meta_cohs_REG ? io_metaArray_fromIMeta_metaData_1_2_coh_state : s1_meta_cohs_r1_2_state; // @[Reg.scala 16:16 17:{18,22}]
  wire [1:0] _GEN_52 = s1_meta_cohs_REG ? io_metaArray_fromIMeta_metaData_1_3_coh_state : s1_meta_cohs_r1_3_state; // @[Reg.scala 16:16 17:{18,22}]
  wire [1:0] _GEN_53 = s1_meta_cohs_REG ? io_metaArray_fromIMeta_metaData_1_4_coh_state : s1_meta_cohs_r1_4_state; // @[Reg.scala 16:16 17:{18,22}]
  wire [1:0] _GEN_54 = s1_meta_cohs_REG ? io_metaArray_fromIMeta_metaData_1_5_coh_state : s1_meta_cohs_r1_5_state; // @[Reg.scala 16:16 17:{18,22}]
  wire [1:0] _GEN_55 = s1_meta_cohs_REG ? io_metaArray_fromIMeta_metaData_1_6_coh_state : s1_meta_cohs_r1_6_state; // @[Reg.scala 16:16 17:{18,22}]
  wire [1:0] _GEN_56 = s1_meta_cohs_REG ? io_metaArray_fromIMeta_metaData_1_7_coh_state : s1_meta_cohs_r1_7_state; // @[Reg.scala 16:16 17:{18,22}]
  reg  s1_meta_errors_REG; // @[ICacheMainPipe.scala 278:92]
  reg  s1_meta_errors_r0_0; // @[Reg.scala 16:16]
  reg  s1_meta_errors_r0_1; // @[Reg.scala 16:16]
  reg  s1_meta_errors_r0_2; // @[Reg.scala 16:16]
  reg  s1_meta_errors_r0_3; // @[Reg.scala 16:16]
  reg  s1_meta_errors_r0_4; // @[Reg.scala 16:16]
  reg  s1_meta_errors_r0_5; // @[Reg.scala 16:16]
  reg  s1_meta_errors_r0_6; // @[Reg.scala 16:16]
  reg  s1_meta_errors_r0_7; // @[Reg.scala 16:16]
  reg  s1_meta_errors_r1_0; // @[Reg.scala 16:16]
  reg  s1_meta_errors_r1_1; // @[Reg.scala 16:16]
  reg  s1_meta_errors_r1_2; // @[Reg.scala 16:16]
  reg  s1_meta_errors_r1_3; // @[Reg.scala 16:16]
  reg  s1_meta_errors_r1_4; // @[Reg.scala 16:16]
  reg  s1_meta_errors_r1_5; // @[Reg.scala 16:16]
  reg  s1_meta_errors_r1_6; // @[Reg.scala 16:16]
  reg  s1_meta_errors_r1_7; // @[Reg.scala 16:16]
  reg  s1_data_cacheline_REG; // @[ICacheMainPipe.scala 280:91]
  reg [511:0] s1_data_cacheline_r0_0; // @[Reg.scala 16:16]
  reg [511:0] s1_data_cacheline_r0_1; // @[Reg.scala 16:16]
  reg [511:0] s1_data_cacheline_r0_2; // @[Reg.scala 16:16]
  reg [511:0] s1_data_cacheline_r0_3; // @[Reg.scala 16:16]
  reg [511:0] s1_data_cacheline_r0_4; // @[Reg.scala 16:16]
  reg [511:0] s1_data_cacheline_r0_5; // @[Reg.scala 16:16]
  reg [511:0] s1_data_cacheline_r0_6; // @[Reg.scala 16:16]
  reg [511:0] s1_data_cacheline_r0_7; // @[Reg.scala 16:16]
  reg [511:0] s1_data_cacheline_r1_0; // @[Reg.scala 16:16]
  reg [511:0] s1_data_cacheline_r1_1; // @[Reg.scala 16:16]
  reg [511:0] s1_data_cacheline_r1_2; // @[Reg.scala 16:16]
  reg [511:0] s1_data_cacheline_r1_3; // @[Reg.scala 16:16]
  reg [511:0] s1_data_cacheline_r1_4; // @[Reg.scala 16:16]
  reg [511:0] s1_data_cacheline_r1_5; // @[Reg.scala 16:16]
  reg [511:0] s1_data_cacheline_r1_6; // @[Reg.scala 16:16]
  reg [511:0] s1_data_cacheline_r1_7; // @[Reg.scala 16:16]
  reg  s1_data_errorBits_REG; // @[ICacheMainPipe.scala 281:91]
  reg [31:0] s1_data_errorBits_r0_0; // @[Reg.scala 16:16]
  reg [31:0] s1_data_errorBits_r0_1; // @[Reg.scala 16:16]
  reg [31:0] s1_data_errorBits_r0_2; // @[Reg.scala 16:16]
  reg [31:0] s1_data_errorBits_r0_3; // @[Reg.scala 16:16]
  reg [31:0] s1_data_errorBits_r0_4; // @[Reg.scala 16:16]
  reg [31:0] s1_data_errorBits_r0_5; // @[Reg.scala 16:16]
  reg [31:0] s1_data_errorBits_r0_6; // @[Reg.scala 16:16]
  reg [31:0] s1_data_errorBits_r0_7; // @[Reg.scala 16:16]
  reg [31:0] s1_data_errorBits_r1_0; // @[Reg.scala 16:16]
  reg [31:0] s1_data_errorBits_r1_1; // @[Reg.scala 16:16]
  reg [31:0] s1_data_errorBits_r1_2; // @[Reg.scala 16:16]
  reg [31:0] s1_data_errorBits_r1_3; // @[Reg.scala 16:16]
  reg [31:0] s1_data_errorBits_r1_4; // @[Reg.scala 16:16]
  reg [31:0] s1_data_errorBits_r1_5; // @[Reg.scala 16:16]
  reg [31:0] s1_data_errorBits_r1_6; // @[Reg.scala 16:16]
  reg [31:0] s1_data_errorBits_r1_7; // @[Reg.scala 16:16]
  wire  s1_tag_eq_vec_0_0 = _GEN_25 == s1_req_ptags_0; // @[ICacheMainPipe.scala 283:124]
  wire  s1_tag_eq_vec_0_1 = _GEN_26 == s1_req_ptags_0; // @[ICacheMainPipe.scala 283:124]
  wire  s1_tag_eq_vec_0_2 = _GEN_27 == s1_req_ptags_0; // @[ICacheMainPipe.scala 283:124]
  wire  s1_tag_eq_vec_0_3 = _GEN_28 == s1_req_ptags_0; // @[ICacheMainPipe.scala 283:124]
  wire  s1_tag_eq_vec_0_4 = _GEN_29 == s1_req_ptags_0; // @[ICacheMainPipe.scala 283:124]
  wire  s1_tag_eq_vec_0_5 = _GEN_30 == s1_req_ptags_0; // @[ICacheMainPipe.scala 283:124]
  wire  s1_tag_eq_vec_0_6 = _GEN_31 == s1_req_ptags_0; // @[ICacheMainPipe.scala 283:124]
  wire  s1_tag_eq_vec_0_7 = _GEN_32 == s1_req_ptags_0; // @[ICacheMainPipe.scala 283:124]
  wire  s1_tag_eq_vec_1_0 = _GEN_33 == s1_req_ptags_1; // @[ICacheMainPipe.scala 283:124]
  wire  s1_tag_eq_vec_1_1 = _GEN_34 == s1_req_ptags_1; // @[ICacheMainPipe.scala 283:124]
  wire  s1_tag_eq_vec_1_2 = _GEN_35 == s1_req_ptags_1; // @[ICacheMainPipe.scala 283:124]
  wire  s1_tag_eq_vec_1_3 = _GEN_36 == s1_req_ptags_1; // @[ICacheMainPipe.scala 283:124]
  wire  s1_tag_eq_vec_1_4 = _GEN_37 == s1_req_ptags_1; // @[ICacheMainPipe.scala 283:124]
  wire  s1_tag_eq_vec_1_5 = _GEN_38 == s1_req_ptags_1; // @[ICacheMainPipe.scala 283:124]
  wire  s1_tag_eq_vec_1_6 = _GEN_39 == s1_req_ptags_1; // @[ICacheMainPipe.scala 283:124]
  wire  s1_tag_eq_vec_1_7 = _GEN_40 == s1_req_ptags_1; // @[ICacheMainPipe.scala 283:124]
  wire  _s1_tag_match_vec_T = _GEN_41 > 2'h0; // @[Metadata.scala 49:45]
  wire  s1_tag_match_vec_0_0 = s1_tag_eq_vec_0_0 & _s1_tag_match_vec_T; // @[ICacheMainPipe.scala 284:146]
  wire  _s1_tag_match_vec_T_2 = _GEN_42 > 2'h0; // @[Metadata.scala 49:45]
  wire  s1_tag_match_vec_0_1 = s1_tag_eq_vec_0_1 & _s1_tag_match_vec_T_2; // @[ICacheMainPipe.scala 284:146]
  wire  _s1_tag_match_vec_T_4 = _GEN_43 > 2'h0; // @[Metadata.scala 49:45]
  wire  s1_tag_match_vec_0_2 = s1_tag_eq_vec_0_2 & _s1_tag_match_vec_T_4; // @[ICacheMainPipe.scala 284:146]
  wire  _s1_tag_match_vec_T_6 = _GEN_44 > 2'h0; // @[Metadata.scala 49:45]
  wire  s1_tag_match_vec_0_3 = s1_tag_eq_vec_0_3 & _s1_tag_match_vec_T_6; // @[ICacheMainPipe.scala 284:146]
  wire  _s1_tag_match_vec_T_8 = _GEN_45 > 2'h0; // @[Metadata.scala 49:45]
  wire  s1_tag_match_vec_0_4 = s1_tag_eq_vec_0_4 & _s1_tag_match_vec_T_8; // @[ICacheMainPipe.scala 284:146]
  wire  _s1_tag_match_vec_T_10 = _GEN_46 > 2'h0; // @[Metadata.scala 49:45]
  wire  s1_tag_match_vec_0_5 = s1_tag_eq_vec_0_5 & _s1_tag_match_vec_T_10; // @[ICacheMainPipe.scala 284:146]
  wire  _s1_tag_match_vec_T_12 = _GEN_47 > 2'h0; // @[Metadata.scala 49:45]
  wire  s1_tag_match_vec_0_6 = s1_tag_eq_vec_0_6 & _s1_tag_match_vec_T_12; // @[ICacheMainPipe.scala 284:146]
  wire  _s1_tag_match_vec_T_14 = _GEN_48 > 2'h0; // @[Metadata.scala 49:45]
  wire  s1_tag_match_vec_0_7 = s1_tag_eq_vec_0_7 & _s1_tag_match_vec_T_14; // @[ICacheMainPipe.scala 284:146]
  wire  _s1_tag_match_vec_T_16 = _GEN_49 > 2'h0; // @[Metadata.scala 49:45]
  wire  s1_tag_match_vec_1_0 = s1_tag_eq_vec_1_0 & _s1_tag_match_vec_T_16; // @[ICacheMainPipe.scala 284:146]
  wire  _s1_tag_match_vec_T_18 = _GEN_50 > 2'h0; // @[Metadata.scala 49:45]
  wire  s1_tag_match_vec_1_1 = s1_tag_eq_vec_1_1 & _s1_tag_match_vec_T_18; // @[ICacheMainPipe.scala 284:146]
  wire  _s1_tag_match_vec_T_20 = _GEN_51 > 2'h0; // @[Metadata.scala 49:45]
  wire  s1_tag_match_vec_1_2 = s1_tag_eq_vec_1_2 & _s1_tag_match_vec_T_20; // @[ICacheMainPipe.scala 284:146]
  wire  _s1_tag_match_vec_T_22 = _GEN_52 > 2'h0; // @[Metadata.scala 49:45]
  wire  s1_tag_match_vec_1_3 = s1_tag_eq_vec_1_3 & _s1_tag_match_vec_T_22; // @[ICacheMainPipe.scala 284:146]
  wire  _s1_tag_match_vec_T_24 = _GEN_53 > 2'h0; // @[Metadata.scala 49:45]
  wire  s1_tag_match_vec_1_4 = s1_tag_eq_vec_1_4 & _s1_tag_match_vec_T_24; // @[ICacheMainPipe.scala 284:146]
  wire  _s1_tag_match_vec_T_26 = _GEN_54 > 2'h0; // @[Metadata.scala 49:45]
  wire  s1_tag_match_vec_1_5 = s1_tag_eq_vec_1_5 & _s1_tag_match_vec_T_26; // @[ICacheMainPipe.scala 284:146]
  wire  _s1_tag_match_vec_T_28 = _GEN_55 > 2'h0; // @[Metadata.scala 49:45]
  wire  s1_tag_match_vec_1_6 = s1_tag_eq_vec_1_6 & _s1_tag_match_vec_T_28; // @[ICacheMainPipe.scala 284:146]
  wire  _s1_tag_match_vec_T_30 = _GEN_56 > 2'h0; // @[Metadata.scala 49:45]
  wire  s1_tag_match_vec_1_7 = s1_tag_eq_vec_1_7 & _s1_tag_match_vec_T_30; // @[ICacheMainPipe.scala 284:146]
  wire  s1_tag_match_0 = s1_tag_match_vec_0_0 | s1_tag_match_vec_0_1 | (s1_tag_match_vec_0_2 | s1_tag_match_vec_0_3) | (
    s1_tag_match_vec_0_4 | s1_tag_match_vec_0_5 | (s1_tag_match_vec_0_6 | s1_tag_match_vec_0_7)); // @[ParallelMux.scala 36:53]
  wire  s1_tag_match_1 = s1_tag_match_vec_1_0 | s1_tag_match_vec_1_1 | (s1_tag_match_vec_1_2 | s1_tag_match_vec_1_3) | (
    s1_tag_match_vec_1_4 | s1_tag_match_vec_1_5 | (s1_tag_match_vec_1_6 | s1_tag_match_vec_1_7)); // @[ParallelMux.scala 36:53]
  wire  s1_port_hit_0 = s1_tag_match_0 & s1_valid & ~tlbExcpPF_0; // @[ICacheMainPipe.scala 287:71]
  wire  s1_port_hit_1 = s1_tag_match_1 & s1_valid & s1_double_line & ~tlbExcpPF_1; // @[ICacheMainPipe.scala 287:134]
  reg [6:0] state_vec__0; // @[Replacement.scala 305:17]
  reg [6:0] state_vec__1; // @[Replacement.scala 305:17]
  reg [6:0] state_vec__2; // @[Replacement.scala 305:17]
  reg [6:0] state_vec__3; // @[Replacement.scala 305:17]
  reg [6:0] state_vec__4; // @[Replacement.scala 305:17]
  reg [6:0] state_vec__5; // @[Replacement.scala 305:17]
  reg [6:0] state_vec__6; // @[Replacement.scala 305:17]
  reg [6:0] state_vec__7; // @[Replacement.scala 305:17]
  reg [6:0] state_vec__8; // @[Replacement.scala 305:17]
  reg [6:0] state_vec__9; // @[Replacement.scala 305:17]
  reg [6:0] state_vec__10; // @[Replacement.scala 305:17]
  reg [6:0] state_vec__11; // @[Replacement.scala 305:17]
  reg [6:0] state_vec__12; // @[Replacement.scala 305:17]
  reg [6:0] state_vec__13; // @[Replacement.scala 305:17]
  reg [6:0] state_vec__14; // @[Replacement.scala 305:17]
  reg [6:0] state_vec__15; // @[Replacement.scala 305:17]
  reg [6:0] state_vec__16; // @[Replacement.scala 305:17]
  reg [6:0] state_vec__17; // @[Replacement.scala 305:17]
  reg [6:0] state_vec__18; // @[Replacement.scala 305:17]
  reg [6:0] state_vec__19; // @[Replacement.scala 305:17]
  reg [6:0] state_vec__20; // @[Replacement.scala 305:17]
  reg [6:0] state_vec__21; // @[Replacement.scala 305:17]
  reg [6:0] state_vec__22; // @[Replacement.scala 305:17]
  reg [6:0] state_vec__23; // @[Replacement.scala 305:17]
  reg [6:0] state_vec__24; // @[Replacement.scala 305:17]
  reg [6:0] state_vec__25; // @[Replacement.scala 305:17]
  reg [6:0] state_vec__26; // @[Replacement.scala 305:17]
  reg [6:0] state_vec__27; // @[Replacement.scala 305:17]
  reg [6:0] state_vec__28; // @[Replacement.scala 305:17]
  reg [6:0] state_vec__29; // @[Replacement.scala 305:17]
  reg [6:0] state_vec__30; // @[Replacement.scala 305:17]
  reg [6:0] state_vec__31; // @[Replacement.scala 305:17]
  reg [6:0] state_vec_1_0; // @[Replacement.scala 305:17]
  reg [6:0] state_vec_1_1; // @[Replacement.scala 305:17]
  reg [6:0] state_vec_1_2; // @[Replacement.scala 305:17]
  reg [6:0] state_vec_1_3; // @[Replacement.scala 305:17]
  reg [6:0] state_vec_1_4; // @[Replacement.scala 305:17]
  reg [6:0] state_vec_1_5; // @[Replacement.scala 305:17]
  reg [6:0] state_vec_1_6; // @[Replacement.scala 305:17]
  reg [6:0] state_vec_1_7; // @[Replacement.scala 305:17]
  reg [6:0] state_vec_1_8; // @[Replacement.scala 305:17]
  reg [6:0] state_vec_1_9; // @[Replacement.scala 305:17]
  reg [6:0] state_vec_1_10; // @[Replacement.scala 305:17]
  reg [6:0] state_vec_1_11; // @[Replacement.scala 305:17]
  reg [6:0] state_vec_1_12; // @[Replacement.scala 305:17]
  reg [6:0] state_vec_1_13; // @[Replacement.scala 305:17]
  reg [6:0] state_vec_1_14; // @[Replacement.scala 305:17]
  reg [6:0] state_vec_1_15; // @[Replacement.scala 305:17]
  reg [6:0] state_vec_1_16; // @[Replacement.scala 305:17]
  reg [6:0] state_vec_1_17; // @[Replacement.scala 305:17]
  reg [6:0] state_vec_1_18; // @[Replacement.scala 305:17]
  reg [6:0] state_vec_1_19; // @[Replacement.scala 305:17]
  reg [6:0] state_vec_1_20; // @[Replacement.scala 305:17]
  reg [6:0] state_vec_1_21; // @[Replacement.scala 305:17]
  reg [6:0] state_vec_1_22; // @[Replacement.scala 305:17]
  reg [6:0] state_vec_1_23; // @[Replacement.scala 305:17]
  reg [6:0] state_vec_1_24; // @[Replacement.scala 305:17]
  reg [6:0] state_vec_1_25; // @[Replacement.scala 305:17]
  reg [6:0] state_vec_1_26; // @[Replacement.scala 305:17]
  reg [6:0] state_vec_1_27; // @[Replacement.scala 305:17]
  reg [6:0] state_vec_1_28; // @[Replacement.scala 305:17]
  reg [6:0] state_vec_1_29; // @[Replacement.scala 305:17]
  reg [6:0] state_vec_1_30; // @[Replacement.scala 305:17]
  reg [6:0] state_vec_1_31; // @[Replacement.scala 305:17]
  wire [6:0] _GEN_106 = 5'h1 == s1_req_vsetIdx_0[4:0] ? state_vec__1 : state_vec__0; // @[Replacement.scala 243:{38,38}]
  wire [6:0] _GEN_107 = 5'h2 == s1_req_vsetIdx_0[4:0] ? state_vec__2 : _GEN_106; // @[Replacement.scala 243:{38,38}]
  wire [6:0] _GEN_108 = 5'h3 == s1_req_vsetIdx_0[4:0] ? state_vec__3 : _GEN_107; // @[Replacement.scala 243:{38,38}]
  wire [6:0] _GEN_109 = 5'h4 == s1_req_vsetIdx_0[4:0] ? state_vec__4 : _GEN_108; // @[Replacement.scala 243:{38,38}]
  wire [6:0] _GEN_110 = 5'h5 == s1_req_vsetIdx_0[4:0] ? state_vec__5 : _GEN_109; // @[Replacement.scala 243:{38,38}]
  wire [6:0] _GEN_111 = 5'h6 == s1_req_vsetIdx_0[4:0] ? state_vec__6 : _GEN_110; // @[Replacement.scala 243:{38,38}]
  wire [6:0] _GEN_112 = 5'h7 == s1_req_vsetIdx_0[4:0] ? state_vec__7 : _GEN_111; // @[Replacement.scala 243:{38,38}]
  wire [6:0] _GEN_113 = 5'h8 == s1_req_vsetIdx_0[4:0] ? state_vec__8 : _GEN_112; // @[Replacement.scala 243:{38,38}]
  wire [6:0] _GEN_114 = 5'h9 == s1_req_vsetIdx_0[4:0] ? state_vec__9 : _GEN_113; // @[Replacement.scala 243:{38,38}]
  wire [6:0] _GEN_115 = 5'ha == s1_req_vsetIdx_0[4:0] ? state_vec__10 : _GEN_114; // @[Replacement.scala 243:{38,38}]
  wire [6:0] _GEN_116 = 5'hb == s1_req_vsetIdx_0[4:0] ? state_vec__11 : _GEN_115; // @[Replacement.scala 243:{38,38}]
  wire [6:0] _GEN_117 = 5'hc == s1_req_vsetIdx_0[4:0] ? state_vec__12 : _GEN_116; // @[Replacement.scala 243:{38,38}]
  wire [6:0] _GEN_118 = 5'hd == s1_req_vsetIdx_0[4:0] ? state_vec__13 : _GEN_117; // @[Replacement.scala 243:{38,38}]
  wire [6:0] _GEN_119 = 5'he == s1_req_vsetIdx_0[4:0] ? state_vec__14 : _GEN_118; // @[Replacement.scala 243:{38,38}]
  wire [6:0] _GEN_120 = 5'hf == s1_req_vsetIdx_0[4:0] ? state_vec__15 : _GEN_119; // @[Replacement.scala 243:{38,38}]
  wire [6:0] _GEN_121 = 5'h10 == s1_req_vsetIdx_0[4:0] ? state_vec__16 : _GEN_120; // @[Replacement.scala 243:{38,38}]
  wire [6:0] _GEN_122 = 5'h11 == s1_req_vsetIdx_0[4:0] ? state_vec__17 : _GEN_121; // @[Replacement.scala 243:{38,38}]
  wire [6:0] _GEN_123 = 5'h12 == s1_req_vsetIdx_0[4:0] ? state_vec__18 : _GEN_122; // @[Replacement.scala 243:{38,38}]
  wire [6:0] _GEN_124 = 5'h13 == s1_req_vsetIdx_0[4:0] ? state_vec__19 : _GEN_123; // @[Replacement.scala 243:{38,38}]
  wire [6:0] _GEN_125 = 5'h14 == s1_req_vsetIdx_0[4:0] ? state_vec__20 : _GEN_124; // @[Replacement.scala 243:{38,38}]
  wire [6:0] _GEN_126 = 5'h15 == s1_req_vsetIdx_0[4:0] ? state_vec__21 : _GEN_125; // @[Replacement.scala 243:{38,38}]
  wire [6:0] _GEN_127 = 5'h16 == s1_req_vsetIdx_0[4:0] ? state_vec__22 : _GEN_126; // @[Replacement.scala 243:{38,38}]
  wire [6:0] _GEN_128 = 5'h17 == s1_req_vsetIdx_0[4:0] ? state_vec__23 : _GEN_127; // @[Replacement.scala 243:{38,38}]
  wire [6:0] _GEN_129 = 5'h18 == s1_req_vsetIdx_0[4:0] ? state_vec__24 : _GEN_128; // @[Replacement.scala 243:{38,38}]
  wire [6:0] _GEN_130 = 5'h19 == s1_req_vsetIdx_0[4:0] ? state_vec__25 : _GEN_129; // @[Replacement.scala 243:{38,38}]
  wire [6:0] _GEN_131 = 5'h1a == s1_req_vsetIdx_0[4:0] ? state_vec__26 : _GEN_130; // @[Replacement.scala 243:{38,38}]
  wire [6:0] _GEN_132 = 5'h1b == s1_req_vsetIdx_0[4:0] ? state_vec__27 : _GEN_131; // @[Replacement.scala 243:{38,38}]
  wire [6:0] _GEN_133 = 5'h1c == s1_req_vsetIdx_0[4:0] ? state_vec__28 : _GEN_132; // @[Replacement.scala 243:{38,38}]
  wire [6:0] _GEN_134 = 5'h1d == s1_req_vsetIdx_0[4:0] ? state_vec__29 : _GEN_133; // @[Replacement.scala 243:{38,38}]
  wire [6:0] _GEN_135 = 5'h1e == s1_req_vsetIdx_0[4:0] ? state_vec__30 : _GEN_134; // @[Replacement.scala 243:{38,38}]
  wire [6:0] _GEN_136 = 5'h1f == s1_req_vsetIdx_0[4:0] ? state_vec__31 : _GEN_135; // @[Replacement.scala 243:{38,38}]
  wire  s1_victim_oh_left_subtree_older = _GEN_136[6]; // @[Replacement.scala 243:38]
  wire [2:0] s1_victim_oh_left_subtree_state = _GEN_136[5:3]; // @[package.scala 154:13]
  wire [2:0] s1_victim_oh_right_subtree_state = _GEN_136[2:0]; // @[Replacement.scala 245:38]
  wire  s1_victim_oh_left_subtree_older_1 = s1_victim_oh_left_subtree_state[2]; // @[Replacement.scala 243:38]
  wire  s1_victim_oh_left_subtree_state_1 = s1_victim_oh_left_subtree_state[1]; // @[package.scala 154:13]
  wire  s1_victim_oh_right_subtree_state_1 = s1_victim_oh_left_subtree_state[0]; // @[Replacement.scala 245:38]
  wire  _s1_victim_oh_T_3 = s1_victim_oh_left_subtree_older_1 ? s1_victim_oh_left_subtree_state_1 :
    s1_victim_oh_right_subtree_state_1; // @[Replacement.scala 250:16]
  wire [1:0] _s1_victim_oh_T_4 = {s1_victim_oh_left_subtree_older_1,_s1_victim_oh_T_3}; // @[Cat.scala 31:58]
  wire  s1_victim_oh_left_subtree_older_2 = s1_victim_oh_right_subtree_state[2]; // @[Replacement.scala 243:38]
  wire  s1_victim_oh_left_subtree_state_2 = s1_victim_oh_right_subtree_state[1]; // @[package.scala 154:13]
  wire  s1_victim_oh_right_subtree_state_2 = s1_victim_oh_right_subtree_state[0]; // @[Replacement.scala 245:38]
  wire  _s1_victim_oh_T_7 = s1_victim_oh_left_subtree_older_2 ? s1_victim_oh_left_subtree_state_2 :
    s1_victim_oh_right_subtree_state_2; // @[Replacement.scala 250:16]
  wire [1:0] _s1_victim_oh_T_8 = {s1_victim_oh_left_subtree_older_2,_s1_victim_oh_T_7}; // @[Cat.scala 31:58]
  wire [1:0] _s1_victim_oh_T_9 = s1_victim_oh_left_subtree_older ? _s1_victim_oh_T_4 : _s1_victim_oh_T_8; // @[Replacement.scala 250:16]
  wire [2:0] _s1_victim_oh_T_10 = {s1_victim_oh_left_subtree_older,_s1_victim_oh_T_9}; // @[Cat.scala 31:58]
  wire [7:0] _s1_victim_oh_T_11 = 8'h1 << _s1_victim_oh_T_10; // @[OneHot.scala 57:35]
  wire [6:0] _GEN_138 = 5'h1 == s1_req_vsetIdx_1[4:0] ? state_vec_1_1 : state_vec_1_0; // @[Replacement.scala 243:{38,38}]
  wire [6:0] _GEN_139 = 5'h2 == s1_req_vsetIdx_1[4:0] ? state_vec_1_2 : _GEN_138; // @[Replacement.scala 243:{38,38}]
  wire [6:0] _GEN_140 = 5'h3 == s1_req_vsetIdx_1[4:0] ? state_vec_1_3 : _GEN_139; // @[Replacement.scala 243:{38,38}]
  wire [6:0] _GEN_141 = 5'h4 == s1_req_vsetIdx_1[4:0] ? state_vec_1_4 : _GEN_140; // @[Replacement.scala 243:{38,38}]
  wire [6:0] _GEN_142 = 5'h5 == s1_req_vsetIdx_1[4:0] ? state_vec_1_5 : _GEN_141; // @[Replacement.scala 243:{38,38}]
  wire [6:0] _GEN_143 = 5'h6 == s1_req_vsetIdx_1[4:0] ? state_vec_1_6 : _GEN_142; // @[Replacement.scala 243:{38,38}]
  wire [6:0] _GEN_144 = 5'h7 == s1_req_vsetIdx_1[4:0] ? state_vec_1_7 : _GEN_143; // @[Replacement.scala 243:{38,38}]
  wire [6:0] _GEN_145 = 5'h8 == s1_req_vsetIdx_1[4:0] ? state_vec_1_8 : _GEN_144; // @[Replacement.scala 243:{38,38}]
  wire [6:0] _GEN_146 = 5'h9 == s1_req_vsetIdx_1[4:0] ? state_vec_1_9 : _GEN_145; // @[Replacement.scala 243:{38,38}]
  wire [6:0] _GEN_147 = 5'ha == s1_req_vsetIdx_1[4:0] ? state_vec_1_10 : _GEN_146; // @[Replacement.scala 243:{38,38}]
  wire [6:0] _GEN_148 = 5'hb == s1_req_vsetIdx_1[4:0] ? state_vec_1_11 : _GEN_147; // @[Replacement.scala 243:{38,38}]
  wire [6:0] _GEN_149 = 5'hc == s1_req_vsetIdx_1[4:0] ? state_vec_1_12 : _GEN_148; // @[Replacement.scala 243:{38,38}]
  wire [6:0] _GEN_150 = 5'hd == s1_req_vsetIdx_1[4:0] ? state_vec_1_13 : _GEN_149; // @[Replacement.scala 243:{38,38}]
  wire [6:0] _GEN_151 = 5'he == s1_req_vsetIdx_1[4:0] ? state_vec_1_14 : _GEN_150; // @[Replacement.scala 243:{38,38}]
  wire [6:0] _GEN_152 = 5'hf == s1_req_vsetIdx_1[4:0] ? state_vec_1_15 : _GEN_151; // @[Replacement.scala 243:{38,38}]
  wire [6:0] _GEN_153 = 5'h10 == s1_req_vsetIdx_1[4:0] ? state_vec_1_16 : _GEN_152; // @[Replacement.scala 243:{38,38}]
  wire [6:0] _GEN_154 = 5'h11 == s1_req_vsetIdx_1[4:0] ? state_vec_1_17 : _GEN_153; // @[Replacement.scala 243:{38,38}]
  wire [6:0] _GEN_155 = 5'h12 == s1_req_vsetIdx_1[4:0] ? state_vec_1_18 : _GEN_154; // @[Replacement.scala 243:{38,38}]
  wire [6:0] _GEN_156 = 5'h13 == s1_req_vsetIdx_1[4:0] ? state_vec_1_19 : _GEN_155; // @[Replacement.scala 243:{38,38}]
  wire [6:0] _GEN_157 = 5'h14 == s1_req_vsetIdx_1[4:0] ? state_vec_1_20 : _GEN_156; // @[Replacement.scala 243:{38,38}]
  wire [6:0] _GEN_158 = 5'h15 == s1_req_vsetIdx_1[4:0] ? state_vec_1_21 : _GEN_157; // @[Replacement.scala 243:{38,38}]
  wire [6:0] _GEN_159 = 5'h16 == s1_req_vsetIdx_1[4:0] ? state_vec_1_22 : _GEN_158; // @[Replacement.scala 243:{38,38}]
  wire [6:0] _GEN_160 = 5'h17 == s1_req_vsetIdx_1[4:0] ? state_vec_1_23 : _GEN_159; // @[Replacement.scala 243:{38,38}]
  wire [6:0] _GEN_161 = 5'h18 == s1_req_vsetIdx_1[4:0] ? state_vec_1_24 : _GEN_160; // @[Replacement.scala 243:{38,38}]
  wire [6:0] _GEN_162 = 5'h19 == s1_req_vsetIdx_1[4:0] ? state_vec_1_25 : _GEN_161; // @[Replacement.scala 243:{38,38}]
  wire [6:0] _GEN_163 = 5'h1a == s1_req_vsetIdx_1[4:0] ? state_vec_1_26 : _GEN_162; // @[Replacement.scala 243:{38,38}]
  wire [6:0] _GEN_164 = 5'h1b == s1_req_vsetIdx_1[4:0] ? state_vec_1_27 : _GEN_163; // @[Replacement.scala 243:{38,38}]
  wire [6:0] _GEN_165 = 5'h1c == s1_req_vsetIdx_1[4:0] ? state_vec_1_28 : _GEN_164; // @[Replacement.scala 243:{38,38}]
  wire [6:0] _GEN_166 = 5'h1d == s1_req_vsetIdx_1[4:0] ? state_vec_1_29 : _GEN_165; // @[Replacement.scala 243:{38,38}]
  wire [6:0] _GEN_167 = 5'h1e == s1_req_vsetIdx_1[4:0] ? state_vec_1_30 : _GEN_166; // @[Replacement.scala 243:{38,38}]
  wire [6:0] _GEN_168 = 5'h1f == s1_req_vsetIdx_1[4:0] ? state_vec_1_31 : _GEN_167; // @[Replacement.scala 243:{38,38}]
  wire  s1_victim_oh_left_subtree_older_3 = _GEN_168[6]; // @[Replacement.scala 243:38]
  wire [2:0] s1_victim_oh_left_subtree_state_3 = _GEN_168[5:3]; // @[package.scala 154:13]
  wire [2:0] s1_victim_oh_right_subtree_state_3 = _GEN_168[2:0]; // @[Replacement.scala 245:38]
  wire  s1_victim_oh_left_subtree_older_4 = s1_victim_oh_left_subtree_state_3[2]; // @[Replacement.scala 243:38]
  wire  s1_victim_oh_left_subtree_state_4 = s1_victim_oh_left_subtree_state_3[1]; // @[package.scala 154:13]
  wire  s1_victim_oh_right_subtree_state_4 = s1_victim_oh_left_subtree_state_3[0]; // @[Replacement.scala 245:38]
  wire  _s1_victim_oh_T_15 = s1_victim_oh_left_subtree_older_4 ? s1_victim_oh_left_subtree_state_4 :
    s1_victim_oh_right_subtree_state_4; // @[Replacement.scala 250:16]
  wire [1:0] _s1_victim_oh_T_16 = {s1_victim_oh_left_subtree_older_4,_s1_victim_oh_T_15}; // @[Cat.scala 31:58]
  wire  s1_victim_oh_left_subtree_older_5 = s1_victim_oh_right_subtree_state_3[2]; // @[Replacement.scala 243:38]
  wire  s1_victim_oh_left_subtree_state_5 = s1_victim_oh_right_subtree_state_3[1]; // @[package.scala 154:13]
  wire  s1_victim_oh_right_subtree_state_5 = s1_victim_oh_right_subtree_state_3[0]; // @[Replacement.scala 245:38]
  wire  _s1_victim_oh_T_19 = s1_victim_oh_left_subtree_older_5 ? s1_victim_oh_left_subtree_state_5 :
    s1_victim_oh_right_subtree_state_5; // @[Replacement.scala 250:16]
  wire [1:0] _s1_victim_oh_T_20 = {s1_victim_oh_left_subtree_older_5,_s1_victim_oh_T_19}; // @[Cat.scala 31:58]
  wire [1:0] _s1_victim_oh_T_21 = s1_victim_oh_left_subtree_older_3 ? _s1_victim_oh_T_16 : _s1_victim_oh_T_20; // @[Replacement.scala 250:16]
  wire [2:0] _s1_victim_oh_T_22 = {s1_victim_oh_left_subtree_older_3,_s1_victim_oh_T_21}; // @[Cat.scala 31:58]
  wire [7:0] _s1_victim_oh_T_23 = 8'h1 << _s1_victim_oh_T_22; // @[OneHot.scala 57:35]
  reg  s1_victim_oh_REG; // @[ICacheMainPipe.scala 293:166]
  reg [7:0] s1_victim_oh_r0; // @[Reg.scala 16:16]
  reg [7:0] s1_victim_oh_r1; // @[Reg.scala 16:16]
  reg [5:0] s2_req_vsetIdx_0; // @[Reg.scala 16:16]
  wire [4:0] touch_sets_0_0 = s2_req_vsetIdx_0[4:0]; // @[ICacheMainPipe.scala 136:36 671:20]
  wire  touch_ways_0_0_valid = s2_valid & s2_port_hit_0; // @[ICacheMainPipe.scala 672:32]
  wire  set_touch_ways_0_valid = touch_ways_0_0_valid & touch_sets_0_0 == 5'h0; // @[Replacement.scala 315:30]
  wire  touch_ways_0_1_valid = s2_valid & _miss_0_s2_0_T_4; // @[ICacheMainPipe.scala 676:32]
  wire  set_touch_ways_1_valid = touch_ways_0_1_valid & touch_sets_0_0 == 5'h0; // @[Replacement.scala 315:30]
  wire  _T_79 = set_touch_ways_0_valid | set_touch_ways_1_valid; // @[package.scala 72:59]
  reg  s2_tag_match_vec_0_7; // @[Reg.scala 16:16]
  reg  s2_tag_match_vec_0_6; // @[Reg.scala 16:16]
  reg  s2_tag_match_vec_0_5; // @[Reg.scala 16:16]
  reg  s2_tag_match_vec_0_4; // @[Reg.scala 16:16]
  reg  s2_tag_match_vec_0_3; // @[Reg.scala 16:16]
  reg  s2_tag_match_vec_0_2; // @[Reg.scala 16:16]
  reg  s2_tag_match_vec_0_1; // @[Reg.scala 16:16]
  reg  s2_tag_match_vec_0_0; // @[Reg.scala 16:16]
  wire [7:0] _touch_ways_0_0_bits_T = {s2_tag_match_vec_0_7,s2_tag_match_vec_0_6,s2_tag_match_vec_0_5,
    s2_tag_match_vec_0_4,s2_tag_match_vec_0_3,s2_tag_match_vec_0_2,s2_tag_match_vec_0_1,s2_tag_match_vec_0_0}; // @[OneHot.scala 22:45]
  wire [3:0] touch_ways_0_0_bits_hi_1 = _touch_ways_0_0_bits_T[7:4]; // @[OneHot.scala 30:18]
  wire  _touch_ways_0_0_bits_T_1 = |touch_ways_0_0_bits_hi_1; // @[OneHot.scala 32:14]
  wire [3:0] touch_ways_0_0_bits_lo_1 = _touch_ways_0_0_bits_T[3:0]; // @[OneHot.scala 31:18]
  wire [3:0] _touch_ways_0_0_bits_T_2 = touch_ways_0_0_bits_hi_1 | touch_ways_0_0_bits_lo_1; // @[OneHot.scala 32:28]
  wire [1:0] touch_ways_0_0_bits_hi_2 = _touch_ways_0_0_bits_T_2[3:2]; // @[OneHot.scala 30:18]
  wire  _touch_ways_0_0_bits_T_3 = |touch_ways_0_0_bits_hi_2; // @[OneHot.scala 32:14]
  wire [1:0] touch_ways_0_0_bits_lo_2 = _touch_ways_0_0_bits_T_2[1:0]; // @[OneHot.scala 31:18]
  wire [1:0] _touch_ways_0_0_bits_T_4 = touch_ways_0_0_bits_hi_2 | touch_ways_0_0_bits_lo_2; // @[OneHot.scala 32:28]
  wire [2:0] touch_ways_0_0_bits = {_touch_ways_0_0_bits_T_1,_touch_ways_0_0_bits_T_3,_touch_ways_0_0_bits_T_4[1]}; // @[Cat.scala 31:58]
  wire  state_vec_0_set_left_older = ~touch_ways_0_0_bits[2]; // @[Replacement.scala 196:33]
  wire [2:0] state_vec_0_left_subtree_state = state_vec__0[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_0_right_subtree_state = state_vec__0[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_0_set_left_older_1 = ~touch_ways_0_0_bits[1]; // @[Replacement.scala 196:33]
  wire  state_vec_0_left_subtree_state_1 = state_vec_0_left_subtree_state[1]; // @[package.scala 154:13]
  wire  state_vec_0_right_subtree_state_1 = state_vec_0_left_subtree_state[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_0_T_3 = ~touch_ways_0_0_bits[0]; // @[Replacement.scala 218:7]
  wire  _state_vec_0_T_4 = state_vec_0_set_left_older_1 ? state_vec_0_left_subtree_state_1 : _state_vec_0_T_3; // @[Replacement.scala 203:16]
  wire  _state_vec_0_T_8 = state_vec_0_set_left_older_1 ? _state_vec_0_T_3 : state_vec_0_right_subtree_state_1; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_0_T_9 = {state_vec_0_set_left_older_1,_state_vec_0_T_4,_state_vec_0_T_8}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_0_T_10 = state_vec_0_set_left_older ? state_vec_0_left_subtree_state : _state_vec_0_T_9; // @[Replacement.scala 203:16]
  wire  state_vec_0_left_subtree_state_2 = state_vec_0_right_subtree_state[1]; // @[package.scala 154:13]
  wire  state_vec_0_right_subtree_state_2 = state_vec_0_right_subtree_state[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_0_T_15 = state_vec_0_set_left_older_1 ? state_vec_0_left_subtree_state_2 : _state_vec_0_T_3; // @[Replacement.scala 203:16]
  wire  _state_vec_0_T_19 = state_vec_0_set_left_older_1 ? _state_vec_0_T_3 : state_vec_0_right_subtree_state_2; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_0_T_20 = {state_vec_0_set_left_older_1,_state_vec_0_T_15,_state_vec_0_T_19}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_0_T_21 = state_vec_0_set_left_older ? _state_vec_0_T_20 : state_vec_0_right_subtree_state; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_0_T_22 = {state_vec_0_set_left_older,_state_vec_0_T_10,_state_vec_0_T_21}; // @[Cat.scala 31:58]
  wire [6:0] _state_vec_0_T_23 = set_touch_ways_0_valid ? _state_vec_0_T_22 : state_vec__0; // @[Replacement.scala 22:56]
  reg [7:0] s2_waymask_0; // @[Reg.scala 16:16]
  wire [3:0] touch_ways_0_1_bits_hi = s2_waymask_0[7:4]; // @[OneHot.scala 30:18]
  wire  _touch_ways_0_1_bits_T = |touch_ways_0_1_bits_hi; // @[OneHot.scala 32:14]
  wire [3:0] touch_ways_0_1_bits_lo = s2_waymask_0[3:0]; // @[OneHot.scala 31:18]
  wire [3:0] _touch_ways_0_1_bits_T_1 = touch_ways_0_1_bits_hi | touch_ways_0_1_bits_lo; // @[OneHot.scala 32:28]
  wire [1:0] touch_ways_0_1_bits_hi_1 = _touch_ways_0_1_bits_T_1[3:2]; // @[OneHot.scala 30:18]
  wire  _touch_ways_0_1_bits_T_2 = |touch_ways_0_1_bits_hi_1; // @[OneHot.scala 32:14]
  wire [1:0] touch_ways_0_1_bits_lo_1 = _touch_ways_0_1_bits_T_1[1:0]; // @[OneHot.scala 31:18]
  wire [1:0] _touch_ways_0_1_bits_T_3 = touch_ways_0_1_bits_hi_1 | touch_ways_0_1_bits_lo_1; // @[OneHot.scala 32:28]
  wire [2:0] touch_ways_0_1_bits = {_touch_ways_0_1_bits_T,_touch_ways_0_1_bits_T_2,_touch_ways_0_1_bits_T_3[1]}; // @[Cat.scala 31:58]
  wire  state_vec_0_set_left_older_3 = ~touch_ways_0_1_bits[2]; // @[Replacement.scala 196:33]
  wire [2:0] state_vec_0_left_subtree_state_3 = _state_vec_0_T_23[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_0_right_subtree_state_3 = _state_vec_0_T_23[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_0_set_left_older_4 = ~touch_ways_0_1_bits[1]; // @[Replacement.scala 196:33]
  wire  state_vec_0_left_subtree_state_4 = state_vec_0_left_subtree_state_3[1]; // @[package.scala 154:13]
  wire  state_vec_0_right_subtree_state_4 = state_vec_0_left_subtree_state_3[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_0_T_27 = ~touch_ways_0_1_bits[0]; // @[Replacement.scala 218:7]
  wire  _state_vec_0_T_28 = state_vec_0_set_left_older_4 ? state_vec_0_left_subtree_state_4 : _state_vec_0_T_27; // @[Replacement.scala 203:16]
  wire  _state_vec_0_T_32 = state_vec_0_set_left_older_4 ? _state_vec_0_T_27 : state_vec_0_right_subtree_state_4; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_0_T_33 = {state_vec_0_set_left_older_4,_state_vec_0_T_28,_state_vec_0_T_32}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_0_T_34 = state_vec_0_set_left_older_3 ? state_vec_0_left_subtree_state_3 : _state_vec_0_T_33; // @[Replacement.scala 203:16]
  wire  state_vec_0_left_subtree_state_5 = state_vec_0_right_subtree_state_3[1]; // @[package.scala 154:13]
  wire  state_vec_0_right_subtree_state_5 = state_vec_0_right_subtree_state_3[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_0_T_39 = state_vec_0_set_left_older_4 ? state_vec_0_left_subtree_state_5 : _state_vec_0_T_27; // @[Replacement.scala 203:16]
  wire  _state_vec_0_T_43 = state_vec_0_set_left_older_4 ? _state_vec_0_T_27 : state_vec_0_right_subtree_state_5; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_0_T_44 = {state_vec_0_set_left_older_4,_state_vec_0_T_39,_state_vec_0_T_43}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_0_T_45 = state_vec_0_set_left_older_3 ? _state_vec_0_T_44 : state_vec_0_right_subtree_state_3; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_0_T_46 = {state_vec_0_set_left_older_3,_state_vec_0_T_34,_state_vec_0_T_45}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_1_valid = touch_ways_0_0_valid & touch_sets_0_0 == 5'h1; // @[Replacement.scala 315:30]
  wire  set_touch_ways_1_1_valid = touch_ways_0_1_valid & touch_sets_0_0 == 5'h1; // @[Replacement.scala 315:30]
  wire  _T_80 = set_touch_ways_0_1_valid | set_touch_ways_1_1_valid; // @[package.scala 72:59]
  wire [2:0] state_vec_1_left_subtree_state = state_vec__1[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_1_right_subtree_state = state_vec__1[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_1_left_subtree_state_1 = state_vec_1_left_subtree_state[1]; // @[package.scala 154:13]
  wire  state_vec_1_right_subtree_state_1 = state_vec_1_left_subtree_state[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_1_T_4 = state_vec_0_set_left_older_1 ? state_vec_1_left_subtree_state_1 : _state_vec_0_T_3; // @[Replacement.scala 203:16]
  wire  _state_vec_1_T_8 = state_vec_0_set_left_older_1 ? _state_vec_0_T_3 : state_vec_1_right_subtree_state_1; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_1_T_9 = {state_vec_0_set_left_older_1,_state_vec_1_T_4,_state_vec_1_T_8}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_1_T_10 = state_vec_0_set_left_older ? state_vec_1_left_subtree_state : _state_vec_1_T_9; // @[Replacement.scala 203:16]
  wire  state_vec_1_left_subtree_state_2 = state_vec_1_right_subtree_state[1]; // @[package.scala 154:13]
  wire  state_vec_1_right_subtree_state_2 = state_vec_1_right_subtree_state[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_1_T_15 = state_vec_0_set_left_older_1 ? state_vec_1_left_subtree_state_2 : _state_vec_0_T_3; // @[Replacement.scala 203:16]
  wire  _state_vec_1_T_19 = state_vec_0_set_left_older_1 ? _state_vec_0_T_3 : state_vec_1_right_subtree_state_2; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_1_T_20 = {state_vec_0_set_left_older_1,_state_vec_1_T_15,_state_vec_1_T_19}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_1_T_21 = state_vec_0_set_left_older ? _state_vec_1_T_20 : state_vec_1_right_subtree_state; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_1_T_22 = {state_vec_0_set_left_older,_state_vec_1_T_10,_state_vec_1_T_21}; // @[Cat.scala 31:58]
  wire [6:0] _state_vec_1_T_23 = set_touch_ways_0_1_valid ? _state_vec_1_T_22 : state_vec__1; // @[Replacement.scala 22:56]
  wire [2:0] state_vec_1_left_subtree_state_3 = _state_vec_1_T_23[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_1_right_subtree_state_3 = _state_vec_1_T_23[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_1_left_subtree_state_4 = state_vec_1_left_subtree_state_3[1]; // @[package.scala 154:13]
  wire  state_vec_1_right_subtree_state_4 = state_vec_1_left_subtree_state_3[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_1_T_28 = state_vec_0_set_left_older_4 ? state_vec_1_left_subtree_state_4 : _state_vec_0_T_27; // @[Replacement.scala 203:16]
  wire  _state_vec_1_T_32 = state_vec_0_set_left_older_4 ? _state_vec_0_T_27 : state_vec_1_right_subtree_state_4; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_1_T_33 = {state_vec_0_set_left_older_4,_state_vec_1_T_28,_state_vec_1_T_32}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_1_T_34 = state_vec_0_set_left_older_3 ? state_vec_1_left_subtree_state_3 : _state_vec_1_T_33; // @[Replacement.scala 203:16]
  wire  state_vec_1_left_subtree_state_5 = state_vec_1_right_subtree_state_3[1]; // @[package.scala 154:13]
  wire  state_vec_1_right_subtree_state_5 = state_vec_1_right_subtree_state_3[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_1_T_39 = state_vec_0_set_left_older_4 ? state_vec_1_left_subtree_state_5 : _state_vec_0_T_27; // @[Replacement.scala 203:16]
  wire  _state_vec_1_T_43 = state_vec_0_set_left_older_4 ? _state_vec_0_T_27 : state_vec_1_right_subtree_state_5; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_1_T_44 = {state_vec_0_set_left_older_4,_state_vec_1_T_39,_state_vec_1_T_43}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_1_T_45 = state_vec_0_set_left_older_3 ? _state_vec_1_T_44 : state_vec_1_right_subtree_state_3; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_1_T_46 = {state_vec_0_set_left_older_3,_state_vec_1_T_34,_state_vec_1_T_45}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_2_valid = touch_ways_0_0_valid & touch_sets_0_0 == 5'h2; // @[Replacement.scala 315:30]
  wire  set_touch_ways_1_2_valid = touch_ways_0_1_valid & touch_sets_0_0 == 5'h2; // @[Replacement.scala 315:30]
  wire  _T_81 = set_touch_ways_0_2_valid | set_touch_ways_1_2_valid; // @[package.scala 72:59]
  wire [2:0] state_vec_2_left_subtree_state = state_vec__2[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_2_right_subtree_state = state_vec__2[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_2_left_subtree_state_1 = state_vec_2_left_subtree_state[1]; // @[package.scala 154:13]
  wire  state_vec_2_right_subtree_state_1 = state_vec_2_left_subtree_state[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_2_T_4 = state_vec_0_set_left_older_1 ? state_vec_2_left_subtree_state_1 : _state_vec_0_T_3; // @[Replacement.scala 203:16]
  wire  _state_vec_2_T_8 = state_vec_0_set_left_older_1 ? _state_vec_0_T_3 : state_vec_2_right_subtree_state_1; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_2_T_9 = {state_vec_0_set_left_older_1,_state_vec_2_T_4,_state_vec_2_T_8}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_2_T_10 = state_vec_0_set_left_older ? state_vec_2_left_subtree_state : _state_vec_2_T_9; // @[Replacement.scala 203:16]
  wire  state_vec_2_left_subtree_state_2 = state_vec_2_right_subtree_state[1]; // @[package.scala 154:13]
  wire  state_vec_2_right_subtree_state_2 = state_vec_2_right_subtree_state[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_2_T_15 = state_vec_0_set_left_older_1 ? state_vec_2_left_subtree_state_2 : _state_vec_0_T_3; // @[Replacement.scala 203:16]
  wire  _state_vec_2_T_19 = state_vec_0_set_left_older_1 ? _state_vec_0_T_3 : state_vec_2_right_subtree_state_2; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_2_T_20 = {state_vec_0_set_left_older_1,_state_vec_2_T_15,_state_vec_2_T_19}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_2_T_21 = state_vec_0_set_left_older ? _state_vec_2_T_20 : state_vec_2_right_subtree_state; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_2_T_22 = {state_vec_0_set_left_older,_state_vec_2_T_10,_state_vec_2_T_21}; // @[Cat.scala 31:58]
  wire [6:0] _state_vec_2_T_23 = set_touch_ways_0_2_valid ? _state_vec_2_T_22 : state_vec__2; // @[Replacement.scala 22:56]
  wire [2:0] state_vec_2_left_subtree_state_3 = _state_vec_2_T_23[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_2_right_subtree_state_3 = _state_vec_2_T_23[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_2_left_subtree_state_4 = state_vec_2_left_subtree_state_3[1]; // @[package.scala 154:13]
  wire  state_vec_2_right_subtree_state_4 = state_vec_2_left_subtree_state_3[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_2_T_28 = state_vec_0_set_left_older_4 ? state_vec_2_left_subtree_state_4 : _state_vec_0_T_27; // @[Replacement.scala 203:16]
  wire  _state_vec_2_T_32 = state_vec_0_set_left_older_4 ? _state_vec_0_T_27 : state_vec_2_right_subtree_state_4; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_2_T_33 = {state_vec_0_set_left_older_4,_state_vec_2_T_28,_state_vec_2_T_32}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_2_T_34 = state_vec_0_set_left_older_3 ? state_vec_2_left_subtree_state_3 : _state_vec_2_T_33; // @[Replacement.scala 203:16]
  wire  state_vec_2_left_subtree_state_5 = state_vec_2_right_subtree_state_3[1]; // @[package.scala 154:13]
  wire  state_vec_2_right_subtree_state_5 = state_vec_2_right_subtree_state_3[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_2_T_39 = state_vec_0_set_left_older_4 ? state_vec_2_left_subtree_state_5 : _state_vec_0_T_27; // @[Replacement.scala 203:16]
  wire  _state_vec_2_T_43 = state_vec_0_set_left_older_4 ? _state_vec_0_T_27 : state_vec_2_right_subtree_state_5; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_2_T_44 = {state_vec_0_set_left_older_4,_state_vec_2_T_39,_state_vec_2_T_43}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_2_T_45 = state_vec_0_set_left_older_3 ? _state_vec_2_T_44 : state_vec_2_right_subtree_state_3; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_2_T_46 = {state_vec_0_set_left_older_3,_state_vec_2_T_34,_state_vec_2_T_45}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_3_valid = touch_ways_0_0_valid & touch_sets_0_0 == 5'h3; // @[Replacement.scala 315:30]
  wire  set_touch_ways_1_3_valid = touch_ways_0_1_valid & touch_sets_0_0 == 5'h3; // @[Replacement.scala 315:30]
  wire  _T_82 = set_touch_ways_0_3_valid | set_touch_ways_1_3_valid; // @[package.scala 72:59]
  wire [2:0] state_vec_3_left_subtree_state = state_vec__3[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_3_right_subtree_state = state_vec__3[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_3_left_subtree_state_1 = state_vec_3_left_subtree_state[1]; // @[package.scala 154:13]
  wire  state_vec_3_right_subtree_state_1 = state_vec_3_left_subtree_state[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_3_T_4 = state_vec_0_set_left_older_1 ? state_vec_3_left_subtree_state_1 : _state_vec_0_T_3; // @[Replacement.scala 203:16]
  wire  _state_vec_3_T_8 = state_vec_0_set_left_older_1 ? _state_vec_0_T_3 : state_vec_3_right_subtree_state_1; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_3_T_9 = {state_vec_0_set_left_older_1,_state_vec_3_T_4,_state_vec_3_T_8}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_3_T_10 = state_vec_0_set_left_older ? state_vec_3_left_subtree_state : _state_vec_3_T_9; // @[Replacement.scala 203:16]
  wire  state_vec_3_left_subtree_state_2 = state_vec_3_right_subtree_state[1]; // @[package.scala 154:13]
  wire  state_vec_3_right_subtree_state_2 = state_vec_3_right_subtree_state[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_3_T_15 = state_vec_0_set_left_older_1 ? state_vec_3_left_subtree_state_2 : _state_vec_0_T_3; // @[Replacement.scala 203:16]
  wire  _state_vec_3_T_19 = state_vec_0_set_left_older_1 ? _state_vec_0_T_3 : state_vec_3_right_subtree_state_2; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_3_T_20 = {state_vec_0_set_left_older_1,_state_vec_3_T_15,_state_vec_3_T_19}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_3_T_21 = state_vec_0_set_left_older ? _state_vec_3_T_20 : state_vec_3_right_subtree_state; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_3_T_22 = {state_vec_0_set_left_older,_state_vec_3_T_10,_state_vec_3_T_21}; // @[Cat.scala 31:58]
  wire [6:0] _state_vec_3_T_23 = set_touch_ways_0_3_valid ? _state_vec_3_T_22 : state_vec__3; // @[Replacement.scala 22:56]
  wire [2:0] state_vec_3_left_subtree_state_3 = _state_vec_3_T_23[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_3_right_subtree_state_3 = _state_vec_3_T_23[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_3_left_subtree_state_4 = state_vec_3_left_subtree_state_3[1]; // @[package.scala 154:13]
  wire  state_vec_3_right_subtree_state_4 = state_vec_3_left_subtree_state_3[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_3_T_28 = state_vec_0_set_left_older_4 ? state_vec_3_left_subtree_state_4 : _state_vec_0_T_27; // @[Replacement.scala 203:16]
  wire  _state_vec_3_T_32 = state_vec_0_set_left_older_4 ? _state_vec_0_T_27 : state_vec_3_right_subtree_state_4; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_3_T_33 = {state_vec_0_set_left_older_4,_state_vec_3_T_28,_state_vec_3_T_32}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_3_T_34 = state_vec_0_set_left_older_3 ? state_vec_3_left_subtree_state_3 : _state_vec_3_T_33; // @[Replacement.scala 203:16]
  wire  state_vec_3_left_subtree_state_5 = state_vec_3_right_subtree_state_3[1]; // @[package.scala 154:13]
  wire  state_vec_3_right_subtree_state_5 = state_vec_3_right_subtree_state_3[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_3_T_39 = state_vec_0_set_left_older_4 ? state_vec_3_left_subtree_state_5 : _state_vec_0_T_27; // @[Replacement.scala 203:16]
  wire  _state_vec_3_T_43 = state_vec_0_set_left_older_4 ? _state_vec_0_T_27 : state_vec_3_right_subtree_state_5; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_3_T_44 = {state_vec_0_set_left_older_4,_state_vec_3_T_39,_state_vec_3_T_43}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_3_T_45 = state_vec_0_set_left_older_3 ? _state_vec_3_T_44 : state_vec_3_right_subtree_state_3; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_3_T_46 = {state_vec_0_set_left_older_3,_state_vec_3_T_34,_state_vec_3_T_45}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_4_valid = touch_ways_0_0_valid & touch_sets_0_0 == 5'h4; // @[Replacement.scala 315:30]
  wire  set_touch_ways_1_4_valid = touch_ways_0_1_valid & touch_sets_0_0 == 5'h4; // @[Replacement.scala 315:30]
  wire  _T_83 = set_touch_ways_0_4_valid | set_touch_ways_1_4_valid; // @[package.scala 72:59]
  wire [2:0] state_vec_4_left_subtree_state = state_vec__4[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_4_right_subtree_state = state_vec__4[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_4_left_subtree_state_1 = state_vec_4_left_subtree_state[1]; // @[package.scala 154:13]
  wire  state_vec_4_right_subtree_state_1 = state_vec_4_left_subtree_state[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_4_T_4 = state_vec_0_set_left_older_1 ? state_vec_4_left_subtree_state_1 : _state_vec_0_T_3; // @[Replacement.scala 203:16]
  wire  _state_vec_4_T_8 = state_vec_0_set_left_older_1 ? _state_vec_0_T_3 : state_vec_4_right_subtree_state_1; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_4_T_9 = {state_vec_0_set_left_older_1,_state_vec_4_T_4,_state_vec_4_T_8}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_4_T_10 = state_vec_0_set_left_older ? state_vec_4_left_subtree_state : _state_vec_4_T_9; // @[Replacement.scala 203:16]
  wire  state_vec_4_left_subtree_state_2 = state_vec_4_right_subtree_state[1]; // @[package.scala 154:13]
  wire  state_vec_4_right_subtree_state_2 = state_vec_4_right_subtree_state[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_4_T_15 = state_vec_0_set_left_older_1 ? state_vec_4_left_subtree_state_2 : _state_vec_0_T_3; // @[Replacement.scala 203:16]
  wire  _state_vec_4_T_19 = state_vec_0_set_left_older_1 ? _state_vec_0_T_3 : state_vec_4_right_subtree_state_2; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_4_T_20 = {state_vec_0_set_left_older_1,_state_vec_4_T_15,_state_vec_4_T_19}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_4_T_21 = state_vec_0_set_left_older ? _state_vec_4_T_20 : state_vec_4_right_subtree_state; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_4_T_22 = {state_vec_0_set_left_older,_state_vec_4_T_10,_state_vec_4_T_21}; // @[Cat.scala 31:58]
  wire [6:0] _state_vec_4_T_23 = set_touch_ways_0_4_valid ? _state_vec_4_T_22 : state_vec__4; // @[Replacement.scala 22:56]
  wire [2:0] state_vec_4_left_subtree_state_3 = _state_vec_4_T_23[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_4_right_subtree_state_3 = _state_vec_4_T_23[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_4_left_subtree_state_4 = state_vec_4_left_subtree_state_3[1]; // @[package.scala 154:13]
  wire  state_vec_4_right_subtree_state_4 = state_vec_4_left_subtree_state_3[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_4_T_28 = state_vec_0_set_left_older_4 ? state_vec_4_left_subtree_state_4 : _state_vec_0_T_27; // @[Replacement.scala 203:16]
  wire  _state_vec_4_T_32 = state_vec_0_set_left_older_4 ? _state_vec_0_T_27 : state_vec_4_right_subtree_state_4; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_4_T_33 = {state_vec_0_set_left_older_4,_state_vec_4_T_28,_state_vec_4_T_32}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_4_T_34 = state_vec_0_set_left_older_3 ? state_vec_4_left_subtree_state_3 : _state_vec_4_T_33; // @[Replacement.scala 203:16]
  wire  state_vec_4_left_subtree_state_5 = state_vec_4_right_subtree_state_3[1]; // @[package.scala 154:13]
  wire  state_vec_4_right_subtree_state_5 = state_vec_4_right_subtree_state_3[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_4_T_39 = state_vec_0_set_left_older_4 ? state_vec_4_left_subtree_state_5 : _state_vec_0_T_27; // @[Replacement.scala 203:16]
  wire  _state_vec_4_T_43 = state_vec_0_set_left_older_4 ? _state_vec_0_T_27 : state_vec_4_right_subtree_state_5; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_4_T_44 = {state_vec_0_set_left_older_4,_state_vec_4_T_39,_state_vec_4_T_43}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_4_T_45 = state_vec_0_set_left_older_3 ? _state_vec_4_T_44 : state_vec_4_right_subtree_state_3; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_4_T_46 = {state_vec_0_set_left_older_3,_state_vec_4_T_34,_state_vec_4_T_45}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_5_valid = touch_ways_0_0_valid & touch_sets_0_0 == 5'h5; // @[Replacement.scala 315:30]
  wire  set_touch_ways_1_5_valid = touch_ways_0_1_valid & touch_sets_0_0 == 5'h5; // @[Replacement.scala 315:30]
  wire  _T_84 = set_touch_ways_0_5_valid | set_touch_ways_1_5_valid; // @[package.scala 72:59]
  wire [2:0] state_vec_5_left_subtree_state = state_vec__5[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_5_right_subtree_state = state_vec__5[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_5_left_subtree_state_1 = state_vec_5_left_subtree_state[1]; // @[package.scala 154:13]
  wire  state_vec_5_right_subtree_state_1 = state_vec_5_left_subtree_state[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_5_T_4 = state_vec_0_set_left_older_1 ? state_vec_5_left_subtree_state_1 : _state_vec_0_T_3; // @[Replacement.scala 203:16]
  wire  _state_vec_5_T_8 = state_vec_0_set_left_older_1 ? _state_vec_0_T_3 : state_vec_5_right_subtree_state_1; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_5_T_9 = {state_vec_0_set_left_older_1,_state_vec_5_T_4,_state_vec_5_T_8}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_5_T_10 = state_vec_0_set_left_older ? state_vec_5_left_subtree_state : _state_vec_5_T_9; // @[Replacement.scala 203:16]
  wire  state_vec_5_left_subtree_state_2 = state_vec_5_right_subtree_state[1]; // @[package.scala 154:13]
  wire  state_vec_5_right_subtree_state_2 = state_vec_5_right_subtree_state[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_5_T_15 = state_vec_0_set_left_older_1 ? state_vec_5_left_subtree_state_2 : _state_vec_0_T_3; // @[Replacement.scala 203:16]
  wire  _state_vec_5_T_19 = state_vec_0_set_left_older_1 ? _state_vec_0_T_3 : state_vec_5_right_subtree_state_2; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_5_T_20 = {state_vec_0_set_left_older_1,_state_vec_5_T_15,_state_vec_5_T_19}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_5_T_21 = state_vec_0_set_left_older ? _state_vec_5_T_20 : state_vec_5_right_subtree_state; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_5_T_22 = {state_vec_0_set_left_older,_state_vec_5_T_10,_state_vec_5_T_21}; // @[Cat.scala 31:58]
  wire [6:0] _state_vec_5_T_23 = set_touch_ways_0_5_valid ? _state_vec_5_T_22 : state_vec__5; // @[Replacement.scala 22:56]
  wire [2:0] state_vec_5_left_subtree_state_3 = _state_vec_5_T_23[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_5_right_subtree_state_3 = _state_vec_5_T_23[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_5_left_subtree_state_4 = state_vec_5_left_subtree_state_3[1]; // @[package.scala 154:13]
  wire  state_vec_5_right_subtree_state_4 = state_vec_5_left_subtree_state_3[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_5_T_28 = state_vec_0_set_left_older_4 ? state_vec_5_left_subtree_state_4 : _state_vec_0_T_27; // @[Replacement.scala 203:16]
  wire  _state_vec_5_T_32 = state_vec_0_set_left_older_4 ? _state_vec_0_T_27 : state_vec_5_right_subtree_state_4; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_5_T_33 = {state_vec_0_set_left_older_4,_state_vec_5_T_28,_state_vec_5_T_32}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_5_T_34 = state_vec_0_set_left_older_3 ? state_vec_5_left_subtree_state_3 : _state_vec_5_T_33; // @[Replacement.scala 203:16]
  wire  state_vec_5_left_subtree_state_5 = state_vec_5_right_subtree_state_3[1]; // @[package.scala 154:13]
  wire  state_vec_5_right_subtree_state_5 = state_vec_5_right_subtree_state_3[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_5_T_39 = state_vec_0_set_left_older_4 ? state_vec_5_left_subtree_state_5 : _state_vec_0_T_27; // @[Replacement.scala 203:16]
  wire  _state_vec_5_T_43 = state_vec_0_set_left_older_4 ? _state_vec_0_T_27 : state_vec_5_right_subtree_state_5; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_5_T_44 = {state_vec_0_set_left_older_4,_state_vec_5_T_39,_state_vec_5_T_43}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_5_T_45 = state_vec_0_set_left_older_3 ? _state_vec_5_T_44 : state_vec_5_right_subtree_state_3; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_5_T_46 = {state_vec_0_set_left_older_3,_state_vec_5_T_34,_state_vec_5_T_45}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_6_valid = touch_ways_0_0_valid & touch_sets_0_0 == 5'h6; // @[Replacement.scala 315:30]
  wire  set_touch_ways_1_6_valid = touch_ways_0_1_valid & touch_sets_0_0 == 5'h6; // @[Replacement.scala 315:30]
  wire  _T_85 = set_touch_ways_0_6_valid | set_touch_ways_1_6_valid; // @[package.scala 72:59]
  wire [2:0] state_vec_6_left_subtree_state = state_vec__6[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_6_right_subtree_state = state_vec__6[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_6_left_subtree_state_1 = state_vec_6_left_subtree_state[1]; // @[package.scala 154:13]
  wire  state_vec_6_right_subtree_state_1 = state_vec_6_left_subtree_state[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_6_T_4 = state_vec_0_set_left_older_1 ? state_vec_6_left_subtree_state_1 : _state_vec_0_T_3; // @[Replacement.scala 203:16]
  wire  _state_vec_6_T_8 = state_vec_0_set_left_older_1 ? _state_vec_0_T_3 : state_vec_6_right_subtree_state_1; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_6_T_9 = {state_vec_0_set_left_older_1,_state_vec_6_T_4,_state_vec_6_T_8}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_6_T_10 = state_vec_0_set_left_older ? state_vec_6_left_subtree_state : _state_vec_6_T_9; // @[Replacement.scala 203:16]
  wire  state_vec_6_left_subtree_state_2 = state_vec_6_right_subtree_state[1]; // @[package.scala 154:13]
  wire  state_vec_6_right_subtree_state_2 = state_vec_6_right_subtree_state[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_6_T_15 = state_vec_0_set_left_older_1 ? state_vec_6_left_subtree_state_2 : _state_vec_0_T_3; // @[Replacement.scala 203:16]
  wire  _state_vec_6_T_19 = state_vec_0_set_left_older_1 ? _state_vec_0_T_3 : state_vec_6_right_subtree_state_2; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_6_T_20 = {state_vec_0_set_left_older_1,_state_vec_6_T_15,_state_vec_6_T_19}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_6_T_21 = state_vec_0_set_left_older ? _state_vec_6_T_20 : state_vec_6_right_subtree_state; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_6_T_22 = {state_vec_0_set_left_older,_state_vec_6_T_10,_state_vec_6_T_21}; // @[Cat.scala 31:58]
  wire [6:0] _state_vec_6_T_23 = set_touch_ways_0_6_valid ? _state_vec_6_T_22 : state_vec__6; // @[Replacement.scala 22:56]
  wire [2:0] state_vec_6_left_subtree_state_3 = _state_vec_6_T_23[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_6_right_subtree_state_3 = _state_vec_6_T_23[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_6_left_subtree_state_4 = state_vec_6_left_subtree_state_3[1]; // @[package.scala 154:13]
  wire  state_vec_6_right_subtree_state_4 = state_vec_6_left_subtree_state_3[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_6_T_28 = state_vec_0_set_left_older_4 ? state_vec_6_left_subtree_state_4 : _state_vec_0_T_27; // @[Replacement.scala 203:16]
  wire  _state_vec_6_T_32 = state_vec_0_set_left_older_4 ? _state_vec_0_T_27 : state_vec_6_right_subtree_state_4; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_6_T_33 = {state_vec_0_set_left_older_4,_state_vec_6_T_28,_state_vec_6_T_32}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_6_T_34 = state_vec_0_set_left_older_3 ? state_vec_6_left_subtree_state_3 : _state_vec_6_T_33; // @[Replacement.scala 203:16]
  wire  state_vec_6_left_subtree_state_5 = state_vec_6_right_subtree_state_3[1]; // @[package.scala 154:13]
  wire  state_vec_6_right_subtree_state_5 = state_vec_6_right_subtree_state_3[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_6_T_39 = state_vec_0_set_left_older_4 ? state_vec_6_left_subtree_state_5 : _state_vec_0_T_27; // @[Replacement.scala 203:16]
  wire  _state_vec_6_T_43 = state_vec_0_set_left_older_4 ? _state_vec_0_T_27 : state_vec_6_right_subtree_state_5; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_6_T_44 = {state_vec_0_set_left_older_4,_state_vec_6_T_39,_state_vec_6_T_43}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_6_T_45 = state_vec_0_set_left_older_3 ? _state_vec_6_T_44 : state_vec_6_right_subtree_state_3; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_6_T_46 = {state_vec_0_set_left_older_3,_state_vec_6_T_34,_state_vec_6_T_45}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_7_valid = touch_ways_0_0_valid & touch_sets_0_0 == 5'h7; // @[Replacement.scala 315:30]
  wire  set_touch_ways_1_7_valid = touch_ways_0_1_valid & touch_sets_0_0 == 5'h7; // @[Replacement.scala 315:30]
  wire  _T_86 = set_touch_ways_0_7_valid | set_touch_ways_1_7_valid; // @[package.scala 72:59]
  wire [2:0] state_vec_7_left_subtree_state = state_vec__7[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_7_right_subtree_state = state_vec__7[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_7_left_subtree_state_1 = state_vec_7_left_subtree_state[1]; // @[package.scala 154:13]
  wire  state_vec_7_right_subtree_state_1 = state_vec_7_left_subtree_state[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_7_T_4 = state_vec_0_set_left_older_1 ? state_vec_7_left_subtree_state_1 : _state_vec_0_T_3; // @[Replacement.scala 203:16]
  wire  _state_vec_7_T_8 = state_vec_0_set_left_older_1 ? _state_vec_0_T_3 : state_vec_7_right_subtree_state_1; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_7_T_9 = {state_vec_0_set_left_older_1,_state_vec_7_T_4,_state_vec_7_T_8}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_7_T_10 = state_vec_0_set_left_older ? state_vec_7_left_subtree_state : _state_vec_7_T_9; // @[Replacement.scala 203:16]
  wire  state_vec_7_left_subtree_state_2 = state_vec_7_right_subtree_state[1]; // @[package.scala 154:13]
  wire  state_vec_7_right_subtree_state_2 = state_vec_7_right_subtree_state[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_7_T_15 = state_vec_0_set_left_older_1 ? state_vec_7_left_subtree_state_2 : _state_vec_0_T_3; // @[Replacement.scala 203:16]
  wire  _state_vec_7_T_19 = state_vec_0_set_left_older_1 ? _state_vec_0_T_3 : state_vec_7_right_subtree_state_2; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_7_T_20 = {state_vec_0_set_left_older_1,_state_vec_7_T_15,_state_vec_7_T_19}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_7_T_21 = state_vec_0_set_left_older ? _state_vec_7_T_20 : state_vec_7_right_subtree_state; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_7_T_22 = {state_vec_0_set_left_older,_state_vec_7_T_10,_state_vec_7_T_21}; // @[Cat.scala 31:58]
  wire [6:0] _state_vec_7_T_23 = set_touch_ways_0_7_valid ? _state_vec_7_T_22 : state_vec__7; // @[Replacement.scala 22:56]
  wire [2:0] state_vec_7_left_subtree_state_3 = _state_vec_7_T_23[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_7_right_subtree_state_3 = _state_vec_7_T_23[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_7_left_subtree_state_4 = state_vec_7_left_subtree_state_3[1]; // @[package.scala 154:13]
  wire  state_vec_7_right_subtree_state_4 = state_vec_7_left_subtree_state_3[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_7_T_28 = state_vec_0_set_left_older_4 ? state_vec_7_left_subtree_state_4 : _state_vec_0_T_27; // @[Replacement.scala 203:16]
  wire  _state_vec_7_T_32 = state_vec_0_set_left_older_4 ? _state_vec_0_T_27 : state_vec_7_right_subtree_state_4; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_7_T_33 = {state_vec_0_set_left_older_4,_state_vec_7_T_28,_state_vec_7_T_32}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_7_T_34 = state_vec_0_set_left_older_3 ? state_vec_7_left_subtree_state_3 : _state_vec_7_T_33; // @[Replacement.scala 203:16]
  wire  state_vec_7_left_subtree_state_5 = state_vec_7_right_subtree_state_3[1]; // @[package.scala 154:13]
  wire  state_vec_7_right_subtree_state_5 = state_vec_7_right_subtree_state_3[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_7_T_39 = state_vec_0_set_left_older_4 ? state_vec_7_left_subtree_state_5 : _state_vec_0_T_27; // @[Replacement.scala 203:16]
  wire  _state_vec_7_T_43 = state_vec_0_set_left_older_4 ? _state_vec_0_T_27 : state_vec_7_right_subtree_state_5; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_7_T_44 = {state_vec_0_set_left_older_4,_state_vec_7_T_39,_state_vec_7_T_43}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_7_T_45 = state_vec_0_set_left_older_3 ? _state_vec_7_T_44 : state_vec_7_right_subtree_state_3; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_7_T_46 = {state_vec_0_set_left_older_3,_state_vec_7_T_34,_state_vec_7_T_45}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_8_valid = touch_ways_0_0_valid & touch_sets_0_0 == 5'h8; // @[Replacement.scala 315:30]
  wire  set_touch_ways_1_8_valid = touch_ways_0_1_valid & touch_sets_0_0 == 5'h8; // @[Replacement.scala 315:30]
  wire  _T_87 = set_touch_ways_0_8_valid | set_touch_ways_1_8_valid; // @[package.scala 72:59]
  wire [2:0] state_vec_8_left_subtree_state = state_vec__8[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_8_right_subtree_state = state_vec__8[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_8_left_subtree_state_1 = state_vec_8_left_subtree_state[1]; // @[package.scala 154:13]
  wire  state_vec_8_right_subtree_state_1 = state_vec_8_left_subtree_state[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_8_T_4 = state_vec_0_set_left_older_1 ? state_vec_8_left_subtree_state_1 : _state_vec_0_T_3; // @[Replacement.scala 203:16]
  wire  _state_vec_8_T_8 = state_vec_0_set_left_older_1 ? _state_vec_0_T_3 : state_vec_8_right_subtree_state_1; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_8_T_9 = {state_vec_0_set_left_older_1,_state_vec_8_T_4,_state_vec_8_T_8}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_8_T_10 = state_vec_0_set_left_older ? state_vec_8_left_subtree_state : _state_vec_8_T_9; // @[Replacement.scala 203:16]
  wire  state_vec_8_left_subtree_state_2 = state_vec_8_right_subtree_state[1]; // @[package.scala 154:13]
  wire  state_vec_8_right_subtree_state_2 = state_vec_8_right_subtree_state[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_8_T_15 = state_vec_0_set_left_older_1 ? state_vec_8_left_subtree_state_2 : _state_vec_0_T_3; // @[Replacement.scala 203:16]
  wire  _state_vec_8_T_19 = state_vec_0_set_left_older_1 ? _state_vec_0_T_3 : state_vec_8_right_subtree_state_2; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_8_T_20 = {state_vec_0_set_left_older_1,_state_vec_8_T_15,_state_vec_8_T_19}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_8_T_21 = state_vec_0_set_left_older ? _state_vec_8_T_20 : state_vec_8_right_subtree_state; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_8_T_22 = {state_vec_0_set_left_older,_state_vec_8_T_10,_state_vec_8_T_21}; // @[Cat.scala 31:58]
  wire [6:0] _state_vec_8_T_23 = set_touch_ways_0_8_valid ? _state_vec_8_T_22 : state_vec__8; // @[Replacement.scala 22:56]
  wire [2:0] state_vec_8_left_subtree_state_3 = _state_vec_8_T_23[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_8_right_subtree_state_3 = _state_vec_8_T_23[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_8_left_subtree_state_4 = state_vec_8_left_subtree_state_3[1]; // @[package.scala 154:13]
  wire  state_vec_8_right_subtree_state_4 = state_vec_8_left_subtree_state_3[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_8_T_28 = state_vec_0_set_left_older_4 ? state_vec_8_left_subtree_state_4 : _state_vec_0_T_27; // @[Replacement.scala 203:16]
  wire  _state_vec_8_T_32 = state_vec_0_set_left_older_4 ? _state_vec_0_T_27 : state_vec_8_right_subtree_state_4; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_8_T_33 = {state_vec_0_set_left_older_4,_state_vec_8_T_28,_state_vec_8_T_32}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_8_T_34 = state_vec_0_set_left_older_3 ? state_vec_8_left_subtree_state_3 : _state_vec_8_T_33; // @[Replacement.scala 203:16]
  wire  state_vec_8_left_subtree_state_5 = state_vec_8_right_subtree_state_3[1]; // @[package.scala 154:13]
  wire  state_vec_8_right_subtree_state_5 = state_vec_8_right_subtree_state_3[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_8_T_39 = state_vec_0_set_left_older_4 ? state_vec_8_left_subtree_state_5 : _state_vec_0_T_27; // @[Replacement.scala 203:16]
  wire  _state_vec_8_T_43 = state_vec_0_set_left_older_4 ? _state_vec_0_T_27 : state_vec_8_right_subtree_state_5; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_8_T_44 = {state_vec_0_set_left_older_4,_state_vec_8_T_39,_state_vec_8_T_43}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_8_T_45 = state_vec_0_set_left_older_3 ? _state_vec_8_T_44 : state_vec_8_right_subtree_state_3; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_8_T_46 = {state_vec_0_set_left_older_3,_state_vec_8_T_34,_state_vec_8_T_45}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_9_valid = touch_ways_0_0_valid & touch_sets_0_0 == 5'h9; // @[Replacement.scala 315:30]
  wire  set_touch_ways_1_9_valid = touch_ways_0_1_valid & touch_sets_0_0 == 5'h9; // @[Replacement.scala 315:30]
  wire  _T_88 = set_touch_ways_0_9_valid | set_touch_ways_1_9_valid; // @[package.scala 72:59]
  wire [2:0] state_vec_9_left_subtree_state = state_vec__9[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_9_right_subtree_state = state_vec__9[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_9_left_subtree_state_1 = state_vec_9_left_subtree_state[1]; // @[package.scala 154:13]
  wire  state_vec_9_right_subtree_state_1 = state_vec_9_left_subtree_state[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_9_T_4 = state_vec_0_set_left_older_1 ? state_vec_9_left_subtree_state_1 : _state_vec_0_T_3; // @[Replacement.scala 203:16]
  wire  _state_vec_9_T_8 = state_vec_0_set_left_older_1 ? _state_vec_0_T_3 : state_vec_9_right_subtree_state_1; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_9_T_9 = {state_vec_0_set_left_older_1,_state_vec_9_T_4,_state_vec_9_T_8}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_9_T_10 = state_vec_0_set_left_older ? state_vec_9_left_subtree_state : _state_vec_9_T_9; // @[Replacement.scala 203:16]
  wire  state_vec_9_left_subtree_state_2 = state_vec_9_right_subtree_state[1]; // @[package.scala 154:13]
  wire  state_vec_9_right_subtree_state_2 = state_vec_9_right_subtree_state[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_9_T_15 = state_vec_0_set_left_older_1 ? state_vec_9_left_subtree_state_2 : _state_vec_0_T_3; // @[Replacement.scala 203:16]
  wire  _state_vec_9_T_19 = state_vec_0_set_left_older_1 ? _state_vec_0_T_3 : state_vec_9_right_subtree_state_2; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_9_T_20 = {state_vec_0_set_left_older_1,_state_vec_9_T_15,_state_vec_9_T_19}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_9_T_21 = state_vec_0_set_left_older ? _state_vec_9_T_20 : state_vec_9_right_subtree_state; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_9_T_22 = {state_vec_0_set_left_older,_state_vec_9_T_10,_state_vec_9_T_21}; // @[Cat.scala 31:58]
  wire [6:0] _state_vec_9_T_23 = set_touch_ways_0_9_valid ? _state_vec_9_T_22 : state_vec__9; // @[Replacement.scala 22:56]
  wire [2:0] state_vec_9_left_subtree_state_3 = _state_vec_9_T_23[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_9_right_subtree_state_3 = _state_vec_9_T_23[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_9_left_subtree_state_4 = state_vec_9_left_subtree_state_3[1]; // @[package.scala 154:13]
  wire  state_vec_9_right_subtree_state_4 = state_vec_9_left_subtree_state_3[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_9_T_28 = state_vec_0_set_left_older_4 ? state_vec_9_left_subtree_state_4 : _state_vec_0_T_27; // @[Replacement.scala 203:16]
  wire  _state_vec_9_T_32 = state_vec_0_set_left_older_4 ? _state_vec_0_T_27 : state_vec_9_right_subtree_state_4; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_9_T_33 = {state_vec_0_set_left_older_4,_state_vec_9_T_28,_state_vec_9_T_32}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_9_T_34 = state_vec_0_set_left_older_3 ? state_vec_9_left_subtree_state_3 : _state_vec_9_T_33; // @[Replacement.scala 203:16]
  wire  state_vec_9_left_subtree_state_5 = state_vec_9_right_subtree_state_3[1]; // @[package.scala 154:13]
  wire  state_vec_9_right_subtree_state_5 = state_vec_9_right_subtree_state_3[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_9_T_39 = state_vec_0_set_left_older_4 ? state_vec_9_left_subtree_state_5 : _state_vec_0_T_27; // @[Replacement.scala 203:16]
  wire  _state_vec_9_T_43 = state_vec_0_set_left_older_4 ? _state_vec_0_T_27 : state_vec_9_right_subtree_state_5; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_9_T_44 = {state_vec_0_set_left_older_4,_state_vec_9_T_39,_state_vec_9_T_43}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_9_T_45 = state_vec_0_set_left_older_3 ? _state_vec_9_T_44 : state_vec_9_right_subtree_state_3; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_9_T_46 = {state_vec_0_set_left_older_3,_state_vec_9_T_34,_state_vec_9_T_45}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_10_valid = touch_ways_0_0_valid & touch_sets_0_0 == 5'ha; // @[Replacement.scala 315:30]
  wire  set_touch_ways_1_10_valid = touch_ways_0_1_valid & touch_sets_0_0 == 5'ha; // @[Replacement.scala 315:30]
  wire  _T_89 = set_touch_ways_0_10_valid | set_touch_ways_1_10_valid; // @[package.scala 72:59]
  wire [2:0] state_vec_10_left_subtree_state = state_vec__10[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_10_right_subtree_state = state_vec__10[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_10_left_subtree_state_1 = state_vec_10_left_subtree_state[1]; // @[package.scala 154:13]
  wire  state_vec_10_right_subtree_state_1 = state_vec_10_left_subtree_state[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_10_T_4 = state_vec_0_set_left_older_1 ? state_vec_10_left_subtree_state_1 : _state_vec_0_T_3; // @[Replacement.scala 203:16]
  wire  _state_vec_10_T_8 = state_vec_0_set_left_older_1 ? _state_vec_0_T_3 : state_vec_10_right_subtree_state_1; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_10_T_9 = {state_vec_0_set_left_older_1,_state_vec_10_T_4,_state_vec_10_T_8}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_10_T_10 = state_vec_0_set_left_older ? state_vec_10_left_subtree_state : _state_vec_10_T_9; // @[Replacement.scala 203:16]
  wire  state_vec_10_left_subtree_state_2 = state_vec_10_right_subtree_state[1]; // @[package.scala 154:13]
  wire  state_vec_10_right_subtree_state_2 = state_vec_10_right_subtree_state[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_10_T_15 = state_vec_0_set_left_older_1 ? state_vec_10_left_subtree_state_2 : _state_vec_0_T_3; // @[Replacement.scala 203:16]
  wire  _state_vec_10_T_19 = state_vec_0_set_left_older_1 ? _state_vec_0_T_3 : state_vec_10_right_subtree_state_2; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_10_T_20 = {state_vec_0_set_left_older_1,_state_vec_10_T_15,_state_vec_10_T_19}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_10_T_21 = state_vec_0_set_left_older ? _state_vec_10_T_20 : state_vec_10_right_subtree_state; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_10_T_22 = {state_vec_0_set_left_older,_state_vec_10_T_10,_state_vec_10_T_21}; // @[Cat.scala 31:58]
  wire [6:0] _state_vec_10_T_23 = set_touch_ways_0_10_valid ? _state_vec_10_T_22 : state_vec__10; // @[Replacement.scala 22:56]
  wire [2:0] state_vec_10_left_subtree_state_3 = _state_vec_10_T_23[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_10_right_subtree_state_3 = _state_vec_10_T_23[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_10_left_subtree_state_4 = state_vec_10_left_subtree_state_3[1]; // @[package.scala 154:13]
  wire  state_vec_10_right_subtree_state_4 = state_vec_10_left_subtree_state_3[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_10_T_28 = state_vec_0_set_left_older_4 ? state_vec_10_left_subtree_state_4 : _state_vec_0_T_27; // @[Replacement.scala 203:16]
  wire  _state_vec_10_T_32 = state_vec_0_set_left_older_4 ? _state_vec_0_T_27 : state_vec_10_right_subtree_state_4; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_10_T_33 = {state_vec_0_set_left_older_4,_state_vec_10_T_28,_state_vec_10_T_32}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_10_T_34 = state_vec_0_set_left_older_3 ? state_vec_10_left_subtree_state_3 : _state_vec_10_T_33; // @[Replacement.scala 203:16]
  wire  state_vec_10_left_subtree_state_5 = state_vec_10_right_subtree_state_3[1]; // @[package.scala 154:13]
  wire  state_vec_10_right_subtree_state_5 = state_vec_10_right_subtree_state_3[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_10_T_39 = state_vec_0_set_left_older_4 ? state_vec_10_left_subtree_state_5 : _state_vec_0_T_27; // @[Replacement.scala 203:16]
  wire  _state_vec_10_T_43 = state_vec_0_set_left_older_4 ? _state_vec_0_T_27 : state_vec_10_right_subtree_state_5; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_10_T_44 = {state_vec_0_set_left_older_4,_state_vec_10_T_39,_state_vec_10_T_43}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_10_T_45 = state_vec_0_set_left_older_3 ? _state_vec_10_T_44 : state_vec_10_right_subtree_state_3
    ; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_10_T_46 = {state_vec_0_set_left_older_3,_state_vec_10_T_34,_state_vec_10_T_45}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_11_valid = touch_ways_0_0_valid & touch_sets_0_0 == 5'hb; // @[Replacement.scala 315:30]
  wire  set_touch_ways_1_11_valid = touch_ways_0_1_valid & touch_sets_0_0 == 5'hb; // @[Replacement.scala 315:30]
  wire  _T_90 = set_touch_ways_0_11_valid | set_touch_ways_1_11_valid; // @[package.scala 72:59]
  wire [2:0] state_vec_11_left_subtree_state = state_vec__11[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_11_right_subtree_state = state_vec__11[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_11_left_subtree_state_1 = state_vec_11_left_subtree_state[1]; // @[package.scala 154:13]
  wire  state_vec_11_right_subtree_state_1 = state_vec_11_left_subtree_state[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_11_T_4 = state_vec_0_set_left_older_1 ? state_vec_11_left_subtree_state_1 : _state_vec_0_T_3; // @[Replacement.scala 203:16]
  wire  _state_vec_11_T_8 = state_vec_0_set_left_older_1 ? _state_vec_0_T_3 : state_vec_11_right_subtree_state_1; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_11_T_9 = {state_vec_0_set_left_older_1,_state_vec_11_T_4,_state_vec_11_T_8}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_11_T_10 = state_vec_0_set_left_older ? state_vec_11_left_subtree_state : _state_vec_11_T_9; // @[Replacement.scala 203:16]
  wire  state_vec_11_left_subtree_state_2 = state_vec_11_right_subtree_state[1]; // @[package.scala 154:13]
  wire  state_vec_11_right_subtree_state_2 = state_vec_11_right_subtree_state[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_11_T_15 = state_vec_0_set_left_older_1 ? state_vec_11_left_subtree_state_2 : _state_vec_0_T_3; // @[Replacement.scala 203:16]
  wire  _state_vec_11_T_19 = state_vec_0_set_left_older_1 ? _state_vec_0_T_3 : state_vec_11_right_subtree_state_2; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_11_T_20 = {state_vec_0_set_left_older_1,_state_vec_11_T_15,_state_vec_11_T_19}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_11_T_21 = state_vec_0_set_left_older ? _state_vec_11_T_20 : state_vec_11_right_subtree_state; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_11_T_22 = {state_vec_0_set_left_older,_state_vec_11_T_10,_state_vec_11_T_21}; // @[Cat.scala 31:58]
  wire [6:0] _state_vec_11_T_23 = set_touch_ways_0_11_valid ? _state_vec_11_T_22 : state_vec__11; // @[Replacement.scala 22:56]
  wire [2:0] state_vec_11_left_subtree_state_3 = _state_vec_11_T_23[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_11_right_subtree_state_3 = _state_vec_11_T_23[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_11_left_subtree_state_4 = state_vec_11_left_subtree_state_3[1]; // @[package.scala 154:13]
  wire  state_vec_11_right_subtree_state_4 = state_vec_11_left_subtree_state_3[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_11_T_28 = state_vec_0_set_left_older_4 ? state_vec_11_left_subtree_state_4 : _state_vec_0_T_27; // @[Replacement.scala 203:16]
  wire  _state_vec_11_T_32 = state_vec_0_set_left_older_4 ? _state_vec_0_T_27 : state_vec_11_right_subtree_state_4; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_11_T_33 = {state_vec_0_set_left_older_4,_state_vec_11_T_28,_state_vec_11_T_32}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_11_T_34 = state_vec_0_set_left_older_3 ? state_vec_11_left_subtree_state_3 : _state_vec_11_T_33; // @[Replacement.scala 203:16]
  wire  state_vec_11_left_subtree_state_5 = state_vec_11_right_subtree_state_3[1]; // @[package.scala 154:13]
  wire  state_vec_11_right_subtree_state_5 = state_vec_11_right_subtree_state_3[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_11_T_39 = state_vec_0_set_left_older_4 ? state_vec_11_left_subtree_state_5 : _state_vec_0_T_27; // @[Replacement.scala 203:16]
  wire  _state_vec_11_T_43 = state_vec_0_set_left_older_4 ? _state_vec_0_T_27 : state_vec_11_right_subtree_state_5; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_11_T_44 = {state_vec_0_set_left_older_4,_state_vec_11_T_39,_state_vec_11_T_43}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_11_T_45 = state_vec_0_set_left_older_3 ? _state_vec_11_T_44 : state_vec_11_right_subtree_state_3
    ; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_11_T_46 = {state_vec_0_set_left_older_3,_state_vec_11_T_34,_state_vec_11_T_45}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_12_valid = touch_ways_0_0_valid & touch_sets_0_0 == 5'hc; // @[Replacement.scala 315:30]
  wire  set_touch_ways_1_12_valid = touch_ways_0_1_valid & touch_sets_0_0 == 5'hc; // @[Replacement.scala 315:30]
  wire  _T_91 = set_touch_ways_0_12_valid | set_touch_ways_1_12_valid; // @[package.scala 72:59]
  wire [2:0] state_vec_12_left_subtree_state = state_vec__12[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_12_right_subtree_state = state_vec__12[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_12_left_subtree_state_1 = state_vec_12_left_subtree_state[1]; // @[package.scala 154:13]
  wire  state_vec_12_right_subtree_state_1 = state_vec_12_left_subtree_state[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_12_T_4 = state_vec_0_set_left_older_1 ? state_vec_12_left_subtree_state_1 : _state_vec_0_T_3; // @[Replacement.scala 203:16]
  wire  _state_vec_12_T_8 = state_vec_0_set_left_older_1 ? _state_vec_0_T_3 : state_vec_12_right_subtree_state_1; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_12_T_9 = {state_vec_0_set_left_older_1,_state_vec_12_T_4,_state_vec_12_T_8}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_12_T_10 = state_vec_0_set_left_older ? state_vec_12_left_subtree_state : _state_vec_12_T_9; // @[Replacement.scala 203:16]
  wire  state_vec_12_left_subtree_state_2 = state_vec_12_right_subtree_state[1]; // @[package.scala 154:13]
  wire  state_vec_12_right_subtree_state_2 = state_vec_12_right_subtree_state[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_12_T_15 = state_vec_0_set_left_older_1 ? state_vec_12_left_subtree_state_2 : _state_vec_0_T_3; // @[Replacement.scala 203:16]
  wire  _state_vec_12_T_19 = state_vec_0_set_left_older_1 ? _state_vec_0_T_3 : state_vec_12_right_subtree_state_2; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_12_T_20 = {state_vec_0_set_left_older_1,_state_vec_12_T_15,_state_vec_12_T_19}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_12_T_21 = state_vec_0_set_left_older ? _state_vec_12_T_20 : state_vec_12_right_subtree_state; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_12_T_22 = {state_vec_0_set_left_older,_state_vec_12_T_10,_state_vec_12_T_21}; // @[Cat.scala 31:58]
  wire [6:0] _state_vec_12_T_23 = set_touch_ways_0_12_valid ? _state_vec_12_T_22 : state_vec__12; // @[Replacement.scala 22:56]
  wire [2:0] state_vec_12_left_subtree_state_3 = _state_vec_12_T_23[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_12_right_subtree_state_3 = _state_vec_12_T_23[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_12_left_subtree_state_4 = state_vec_12_left_subtree_state_3[1]; // @[package.scala 154:13]
  wire  state_vec_12_right_subtree_state_4 = state_vec_12_left_subtree_state_3[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_12_T_28 = state_vec_0_set_left_older_4 ? state_vec_12_left_subtree_state_4 : _state_vec_0_T_27; // @[Replacement.scala 203:16]
  wire  _state_vec_12_T_32 = state_vec_0_set_left_older_4 ? _state_vec_0_T_27 : state_vec_12_right_subtree_state_4; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_12_T_33 = {state_vec_0_set_left_older_4,_state_vec_12_T_28,_state_vec_12_T_32}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_12_T_34 = state_vec_0_set_left_older_3 ? state_vec_12_left_subtree_state_3 : _state_vec_12_T_33; // @[Replacement.scala 203:16]
  wire  state_vec_12_left_subtree_state_5 = state_vec_12_right_subtree_state_3[1]; // @[package.scala 154:13]
  wire  state_vec_12_right_subtree_state_5 = state_vec_12_right_subtree_state_3[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_12_T_39 = state_vec_0_set_left_older_4 ? state_vec_12_left_subtree_state_5 : _state_vec_0_T_27; // @[Replacement.scala 203:16]
  wire  _state_vec_12_T_43 = state_vec_0_set_left_older_4 ? _state_vec_0_T_27 : state_vec_12_right_subtree_state_5; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_12_T_44 = {state_vec_0_set_left_older_4,_state_vec_12_T_39,_state_vec_12_T_43}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_12_T_45 = state_vec_0_set_left_older_3 ? _state_vec_12_T_44 : state_vec_12_right_subtree_state_3
    ; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_12_T_46 = {state_vec_0_set_left_older_3,_state_vec_12_T_34,_state_vec_12_T_45}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_13_valid = touch_ways_0_0_valid & touch_sets_0_0 == 5'hd; // @[Replacement.scala 315:30]
  wire  set_touch_ways_1_13_valid = touch_ways_0_1_valid & touch_sets_0_0 == 5'hd; // @[Replacement.scala 315:30]
  wire  _T_92 = set_touch_ways_0_13_valid | set_touch_ways_1_13_valid; // @[package.scala 72:59]
  wire [2:0] state_vec_13_left_subtree_state = state_vec__13[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_13_right_subtree_state = state_vec__13[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_13_left_subtree_state_1 = state_vec_13_left_subtree_state[1]; // @[package.scala 154:13]
  wire  state_vec_13_right_subtree_state_1 = state_vec_13_left_subtree_state[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_13_T_4 = state_vec_0_set_left_older_1 ? state_vec_13_left_subtree_state_1 : _state_vec_0_T_3; // @[Replacement.scala 203:16]
  wire  _state_vec_13_T_8 = state_vec_0_set_left_older_1 ? _state_vec_0_T_3 : state_vec_13_right_subtree_state_1; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_13_T_9 = {state_vec_0_set_left_older_1,_state_vec_13_T_4,_state_vec_13_T_8}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_13_T_10 = state_vec_0_set_left_older ? state_vec_13_left_subtree_state : _state_vec_13_T_9; // @[Replacement.scala 203:16]
  wire  state_vec_13_left_subtree_state_2 = state_vec_13_right_subtree_state[1]; // @[package.scala 154:13]
  wire  state_vec_13_right_subtree_state_2 = state_vec_13_right_subtree_state[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_13_T_15 = state_vec_0_set_left_older_1 ? state_vec_13_left_subtree_state_2 : _state_vec_0_T_3; // @[Replacement.scala 203:16]
  wire  _state_vec_13_T_19 = state_vec_0_set_left_older_1 ? _state_vec_0_T_3 : state_vec_13_right_subtree_state_2; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_13_T_20 = {state_vec_0_set_left_older_1,_state_vec_13_T_15,_state_vec_13_T_19}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_13_T_21 = state_vec_0_set_left_older ? _state_vec_13_T_20 : state_vec_13_right_subtree_state; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_13_T_22 = {state_vec_0_set_left_older,_state_vec_13_T_10,_state_vec_13_T_21}; // @[Cat.scala 31:58]
  wire [6:0] _state_vec_13_T_23 = set_touch_ways_0_13_valid ? _state_vec_13_T_22 : state_vec__13; // @[Replacement.scala 22:56]
  wire [2:0] state_vec_13_left_subtree_state_3 = _state_vec_13_T_23[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_13_right_subtree_state_3 = _state_vec_13_T_23[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_13_left_subtree_state_4 = state_vec_13_left_subtree_state_3[1]; // @[package.scala 154:13]
  wire  state_vec_13_right_subtree_state_4 = state_vec_13_left_subtree_state_3[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_13_T_28 = state_vec_0_set_left_older_4 ? state_vec_13_left_subtree_state_4 : _state_vec_0_T_27; // @[Replacement.scala 203:16]
  wire  _state_vec_13_T_32 = state_vec_0_set_left_older_4 ? _state_vec_0_T_27 : state_vec_13_right_subtree_state_4; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_13_T_33 = {state_vec_0_set_left_older_4,_state_vec_13_T_28,_state_vec_13_T_32}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_13_T_34 = state_vec_0_set_left_older_3 ? state_vec_13_left_subtree_state_3 : _state_vec_13_T_33; // @[Replacement.scala 203:16]
  wire  state_vec_13_left_subtree_state_5 = state_vec_13_right_subtree_state_3[1]; // @[package.scala 154:13]
  wire  state_vec_13_right_subtree_state_5 = state_vec_13_right_subtree_state_3[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_13_T_39 = state_vec_0_set_left_older_4 ? state_vec_13_left_subtree_state_5 : _state_vec_0_T_27; // @[Replacement.scala 203:16]
  wire  _state_vec_13_T_43 = state_vec_0_set_left_older_4 ? _state_vec_0_T_27 : state_vec_13_right_subtree_state_5; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_13_T_44 = {state_vec_0_set_left_older_4,_state_vec_13_T_39,_state_vec_13_T_43}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_13_T_45 = state_vec_0_set_left_older_3 ? _state_vec_13_T_44 : state_vec_13_right_subtree_state_3
    ; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_13_T_46 = {state_vec_0_set_left_older_3,_state_vec_13_T_34,_state_vec_13_T_45}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_14_valid = touch_ways_0_0_valid & touch_sets_0_0 == 5'he; // @[Replacement.scala 315:30]
  wire  set_touch_ways_1_14_valid = touch_ways_0_1_valid & touch_sets_0_0 == 5'he; // @[Replacement.scala 315:30]
  wire  _T_93 = set_touch_ways_0_14_valid | set_touch_ways_1_14_valid; // @[package.scala 72:59]
  wire [2:0] state_vec_14_left_subtree_state = state_vec__14[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_14_right_subtree_state = state_vec__14[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_14_left_subtree_state_1 = state_vec_14_left_subtree_state[1]; // @[package.scala 154:13]
  wire  state_vec_14_right_subtree_state_1 = state_vec_14_left_subtree_state[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_14_T_4 = state_vec_0_set_left_older_1 ? state_vec_14_left_subtree_state_1 : _state_vec_0_T_3; // @[Replacement.scala 203:16]
  wire  _state_vec_14_T_8 = state_vec_0_set_left_older_1 ? _state_vec_0_T_3 : state_vec_14_right_subtree_state_1; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_14_T_9 = {state_vec_0_set_left_older_1,_state_vec_14_T_4,_state_vec_14_T_8}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_14_T_10 = state_vec_0_set_left_older ? state_vec_14_left_subtree_state : _state_vec_14_T_9; // @[Replacement.scala 203:16]
  wire  state_vec_14_left_subtree_state_2 = state_vec_14_right_subtree_state[1]; // @[package.scala 154:13]
  wire  state_vec_14_right_subtree_state_2 = state_vec_14_right_subtree_state[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_14_T_15 = state_vec_0_set_left_older_1 ? state_vec_14_left_subtree_state_2 : _state_vec_0_T_3; // @[Replacement.scala 203:16]
  wire  _state_vec_14_T_19 = state_vec_0_set_left_older_1 ? _state_vec_0_T_3 : state_vec_14_right_subtree_state_2; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_14_T_20 = {state_vec_0_set_left_older_1,_state_vec_14_T_15,_state_vec_14_T_19}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_14_T_21 = state_vec_0_set_left_older ? _state_vec_14_T_20 : state_vec_14_right_subtree_state; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_14_T_22 = {state_vec_0_set_left_older,_state_vec_14_T_10,_state_vec_14_T_21}; // @[Cat.scala 31:58]
  wire [6:0] _state_vec_14_T_23 = set_touch_ways_0_14_valid ? _state_vec_14_T_22 : state_vec__14; // @[Replacement.scala 22:56]
  wire [2:0] state_vec_14_left_subtree_state_3 = _state_vec_14_T_23[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_14_right_subtree_state_3 = _state_vec_14_T_23[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_14_left_subtree_state_4 = state_vec_14_left_subtree_state_3[1]; // @[package.scala 154:13]
  wire  state_vec_14_right_subtree_state_4 = state_vec_14_left_subtree_state_3[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_14_T_28 = state_vec_0_set_left_older_4 ? state_vec_14_left_subtree_state_4 : _state_vec_0_T_27; // @[Replacement.scala 203:16]
  wire  _state_vec_14_T_32 = state_vec_0_set_left_older_4 ? _state_vec_0_T_27 : state_vec_14_right_subtree_state_4; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_14_T_33 = {state_vec_0_set_left_older_4,_state_vec_14_T_28,_state_vec_14_T_32}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_14_T_34 = state_vec_0_set_left_older_3 ? state_vec_14_left_subtree_state_3 : _state_vec_14_T_33; // @[Replacement.scala 203:16]
  wire  state_vec_14_left_subtree_state_5 = state_vec_14_right_subtree_state_3[1]; // @[package.scala 154:13]
  wire  state_vec_14_right_subtree_state_5 = state_vec_14_right_subtree_state_3[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_14_T_39 = state_vec_0_set_left_older_4 ? state_vec_14_left_subtree_state_5 : _state_vec_0_T_27; // @[Replacement.scala 203:16]
  wire  _state_vec_14_T_43 = state_vec_0_set_left_older_4 ? _state_vec_0_T_27 : state_vec_14_right_subtree_state_5; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_14_T_44 = {state_vec_0_set_left_older_4,_state_vec_14_T_39,_state_vec_14_T_43}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_14_T_45 = state_vec_0_set_left_older_3 ? _state_vec_14_T_44 : state_vec_14_right_subtree_state_3
    ; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_14_T_46 = {state_vec_0_set_left_older_3,_state_vec_14_T_34,_state_vec_14_T_45}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_15_valid = touch_ways_0_0_valid & touch_sets_0_0 == 5'hf; // @[Replacement.scala 315:30]
  wire  set_touch_ways_1_15_valid = touch_ways_0_1_valid & touch_sets_0_0 == 5'hf; // @[Replacement.scala 315:30]
  wire  _T_94 = set_touch_ways_0_15_valid | set_touch_ways_1_15_valid; // @[package.scala 72:59]
  wire [2:0] state_vec_15_left_subtree_state = state_vec__15[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_15_right_subtree_state = state_vec__15[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_15_left_subtree_state_1 = state_vec_15_left_subtree_state[1]; // @[package.scala 154:13]
  wire  state_vec_15_right_subtree_state_1 = state_vec_15_left_subtree_state[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_15_T_4 = state_vec_0_set_left_older_1 ? state_vec_15_left_subtree_state_1 : _state_vec_0_T_3; // @[Replacement.scala 203:16]
  wire  _state_vec_15_T_8 = state_vec_0_set_left_older_1 ? _state_vec_0_T_3 : state_vec_15_right_subtree_state_1; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_15_T_9 = {state_vec_0_set_left_older_1,_state_vec_15_T_4,_state_vec_15_T_8}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_15_T_10 = state_vec_0_set_left_older ? state_vec_15_left_subtree_state : _state_vec_15_T_9; // @[Replacement.scala 203:16]
  wire  state_vec_15_left_subtree_state_2 = state_vec_15_right_subtree_state[1]; // @[package.scala 154:13]
  wire  state_vec_15_right_subtree_state_2 = state_vec_15_right_subtree_state[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_15_T_15 = state_vec_0_set_left_older_1 ? state_vec_15_left_subtree_state_2 : _state_vec_0_T_3; // @[Replacement.scala 203:16]
  wire  _state_vec_15_T_19 = state_vec_0_set_left_older_1 ? _state_vec_0_T_3 : state_vec_15_right_subtree_state_2; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_15_T_20 = {state_vec_0_set_left_older_1,_state_vec_15_T_15,_state_vec_15_T_19}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_15_T_21 = state_vec_0_set_left_older ? _state_vec_15_T_20 : state_vec_15_right_subtree_state; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_15_T_22 = {state_vec_0_set_left_older,_state_vec_15_T_10,_state_vec_15_T_21}; // @[Cat.scala 31:58]
  wire [6:0] _state_vec_15_T_23 = set_touch_ways_0_15_valid ? _state_vec_15_T_22 : state_vec__15; // @[Replacement.scala 22:56]
  wire [2:0] state_vec_15_left_subtree_state_3 = _state_vec_15_T_23[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_15_right_subtree_state_3 = _state_vec_15_T_23[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_15_left_subtree_state_4 = state_vec_15_left_subtree_state_3[1]; // @[package.scala 154:13]
  wire  state_vec_15_right_subtree_state_4 = state_vec_15_left_subtree_state_3[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_15_T_28 = state_vec_0_set_left_older_4 ? state_vec_15_left_subtree_state_4 : _state_vec_0_T_27; // @[Replacement.scala 203:16]
  wire  _state_vec_15_T_32 = state_vec_0_set_left_older_4 ? _state_vec_0_T_27 : state_vec_15_right_subtree_state_4; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_15_T_33 = {state_vec_0_set_left_older_4,_state_vec_15_T_28,_state_vec_15_T_32}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_15_T_34 = state_vec_0_set_left_older_3 ? state_vec_15_left_subtree_state_3 : _state_vec_15_T_33; // @[Replacement.scala 203:16]
  wire  state_vec_15_left_subtree_state_5 = state_vec_15_right_subtree_state_3[1]; // @[package.scala 154:13]
  wire  state_vec_15_right_subtree_state_5 = state_vec_15_right_subtree_state_3[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_15_T_39 = state_vec_0_set_left_older_4 ? state_vec_15_left_subtree_state_5 : _state_vec_0_T_27; // @[Replacement.scala 203:16]
  wire  _state_vec_15_T_43 = state_vec_0_set_left_older_4 ? _state_vec_0_T_27 : state_vec_15_right_subtree_state_5; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_15_T_44 = {state_vec_0_set_left_older_4,_state_vec_15_T_39,_state_vec_15_T_43}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_15_T_45 = state_vec_0_set_left_older_3 ? _state_vec_15_T_44 : state_vec_15_right_subtree_state_3
    ; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_15_T_46 = {state_vec_0_set_left_older_3,_state_vec_15_T_34,_state_vec_15_T_45}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_16_valid = touch_ways_0_0_valid & touch_sets_0_0 == 5'h10; // @[Replacement.scala 315:30]
  wire  set_touch_ways_1_16_valid = touch_ways_0_1_valid & touch_sets_0_0 == 5'h10; // @[Replacement.scala 315:30]
  wire  _T_95 = set_touch_ways_0_16_valid | set_touch_ways_1_16_valid; // @[package.scala 72:59]
  wire [2:0] state_vec_16_left_subtree_state = state_vec__16[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_16_right_subtree_state = state_vec__16[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_16_left_subtree_state_1 = state_vec_16_left_subtree_state[1]; // @[package.scala 154:13]
  wire  state_vec_16_right_subtree_state_1 = state_vec_16_left_subtree_state[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_16_T_4 = state_vec_0_set_left_older_1 ? state_vec_16_left_subtree_state_1 : _state_vec_0_T_3; // @[Replacement.scala 203:16]
  wire  _state_vec_16_T_8 = state_vec_0_set_left_older_1 ? _state_vec_0_T_3 : state_vec_16_right_subtree_state_1; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_16_T_9 = {state_vec_0_set_left_older_1,_state_vec_16_T_4,_state_vec_16_T_8}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_16_T_10 = state_vec_0_set_left_older ? state_vec_16_left_subtree_state : _state_vec_16_T_9; // @[Replacement.scala 203:16]
  wire  state_vec_16_left_subtree_state_2 = state_vec_16_right_subtree_state[1]; // @[package.scala 154:13]
  wire  state_vec_16_right_subtree_state_2 = state_vec_16_right_subtree_state[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_16_T_15 = state_vec_0_set_left_older_1 ? state_vec_16_left_subtree_state_2 : _state_vec_0_T_3; // @[Replacement.scala 203:16]
  wire  _state_vec_16_T_19 = state_vec_0_set_left_older_1 ? _state_vec_0_T_3 : state_vec_16_right_subtree_state_2; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_16_T_20 = {state_vec_0_set_left_older_1,_state_vec_16_T_15,_state_vec_16_T_19}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_16_T_21 = state_vec_0_set_left_older ? _state_vec_16_T_20 : state_vec_16_right_subtree_state; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_16_T_22 = {state_vec_0_set_left_older,_state_vec_16_T_10,_state_vec_16_T_21}; // @[Cat.scala 31:58]
  wire [6:0] _state_vec_16_T_23 = set_touch_ways_0_16_valid ? _state_vec_16_T_22 : state_vec__16; // @[Replacement.scala 22:56]
  wire [2:0] state_vec_16_left_subtree_state_3 = _state_vec_16_T_23[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_16_right_subtree_state_3 = _state_vec_16_T_23[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_16_left_subtree_state_4 = state_vec_16_left_subtree_state_3[1]; // @[package.scala 154:13]
  wire  state_vec_16_right_subtree_state_4 = state_vec_16_left_subtree_state_3[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_16_T_28 = state_vec_0_set_left_older_4 ? state_vec_16_left_subtree_state_4 : _state_vec_0_T_27; // @[Replacement.scala 203:16]
  wire  _state_vec_16_T_32 = state_vec_0_set_left_older_4 ? _state_vec_0_T_27 : state_vec_16_right_subtree_state_4; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_16_T_33 = {state_vec_0_set_left_older_4,_state_vec_16_T_28,_state_vec_16_T_32}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_16_T_34 = state_vec_0_set_left_older_3 ? state_vec_16_left_subtree_state_3 : _state_vec_16_T_33; // @[Replacement.scala 203:16]
  wire  state_vec_16_left_subtree_state_5 = state_vec_16_right_subtree_state_3[1]; // @[package.scala 154:13]
  wire  state_vec_16_right_subtree_state_5 = state_vec_16_right_subtree_state_3[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_16_T_39 = state_vec_0_set_left_older_4 ? state_vec_16_left_subtree_state_5 : _state_vec_0_T_27; // @[Replacement.scala 203:16]
  wire  _state_vec_16_T_43 = state_vec_0_set_left_older_4 ? _state_vec_0_T_27 : state_vec_16_right_subtree_state_5; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_16_T_44 = {state_vec_0_set_left_older_4,_state_vec_16_T_39,_state_vec_16_T_43}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_16_T_45 = state_vec_0_set_left_older_3 ? _state_vec_16_T_44 : state_vec_16_right_subtree_state_3
    ; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_16_T_46 = {state_vec_0_set_left_older_3,_state_vec_16_T_34,_state_vec_16_T_45}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_17_valid = touch_ways_0_0_valid & touch_sets_0_0 == 5'h11; // @[Replacement.scala 315:30]
  wire  set_touch_ways_1_17_valid = touch_ways_0_1_valid & touch_sets_0_0 == 5'h11; // @[Replacement.scala 315:30]
  wire  _T_96 = set_touch_ways_0_17_valid | set_touch_ways_1_17_valid; // @[package.scala 72:59]
  wire [2:0] state_vec_17_left_subtree_state = state_vec__17[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_17_right_subtree_state = state_vec__17[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_17_left_subtree_state_1 = state_vec_17_left_subtree_state[1]; // @[package.scala 154:13]
  wire  state_vec_17_right_subtree_state_1 = state_vec_17_left_subtree_state[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_17_T_4 = state_vec_0_set_left_older_1 ? state_vec_17_left_subtree_state_1 : _state_vec_0_T_3; // @[Replacement.scala 203:16]
  wire  _state_vec_17_T_8 = state_vec_0_set_left_older_1 ? _state_vec_0_T_3 : state_vec_17_right_subtree_state_1; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_17_T_9 = {state_vec_0_set_left_older_1,_state_vec_17_T_4,_state_vec_17_T_8}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_17_T_10 = state_vec_0_set_left_older ? state_vec_17_left_subtree_state : _state_vec_17_T_9; // @[Replacement.scala 203:16]
  wire  state_vec_17_left_subtree_state_2 = state_vec_17_right_subtree_state[1]; // @[package.scala 154:13]
  wire  state_vec_17_right_subtree_state_2 = state_vec_17_right_subtree_state[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_17_T_15 = state_vec_0_set_left_older_1 ? state_vec_17_left_subtree_state_2 : _state_vec_0_T_3; // @[Replacement.scala 203:16]
  wire  _state_vec_17_T_19 = state_vec_0_set_left_older_1 ? _state_vec_0_T_3 : state_vec_17_right_subtree_state_2; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_17_T_20 = {state_vec_0_set_left_older_1,_state_vec_17_T_15,_state_vec_17_T_19}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_17_T_21 = state_vec_0_set_left_older ? _state_vec_17_T_20 : state_vec_17_right_subtree_state; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_17_T_22 = {state_vec_0_set_left_older,_state_vec_17_T_10,_state_vec_17_T_21}; // @[Cat.scala 31:58]
  wire [6:0] _state_vec_17_T_23 = set_touch_ways_0_17_valid ? _state_vec_17_T_22 : state_vec__17; // @[Replacement.scala 22:56]
  wire [2:0] state_vec_17_left_subtree_state_3 = _state_vec_17_T_23[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_17_right_subtree_state_3 = _state_vec_17_T_23[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_17_left_subtree_state_4 = state_vec_17_left_subtree_state_3[1]; // @[package.scala 154:13]
  wire  state_vec_17_right_subtree_state_4 = state_vec_17_left_subtree_state_3[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_17_T_28 = state_vec_0_set_left_older_4 ? state_vec_17_left_subtree_state_4 : _state_vec_0_T_27; // @[Replacement.scala 203:16]
  wire  _state_vec_17_T_32 = state_vec_0_set_left_older_4 ? _state_vec_0_T_27 : state_vec_17_right_subtree_state_4; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_17_T_33 = {state_vec_0_set_left_older_4,_state_vec_17_T_28,_state_vec_17_T_32}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_17_T_34 = state_vec_0_set_left_older_3 ? state_vec_17_left_subtree_state_3 : _state_vec_17_T_33; // @[Replacement.scala 203:16]
  wire  state_vec_17_left_subtree_state_5 = state_vec_17_right_subtree_state_3[1]; // @[package.scala 154:13]
  wire  state_vec_17_right_subtree_state_5 = state_vec_17_right_subtree_state_3[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_17_T_39 = state_vec_0_set_left_older_4 ? state_vec_17_left_subtree_state_5 : _state_vec_0_T_27; // @[Replacement.scala 203:16]
  wire  _state_vec_17_T_43 = state_vec_0_set_left_older_4 ? _state_vec_0_T_27 : state_vec_17_right_subtree_state_5; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_17_T_44 = {state_vec_0_set_left_older_4,_state_vec_17_T_39,_state_vec_17_T_43}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_17_T_45 = state_vec_0_set_left_older_3 ? _state_vec_17_T_44 : state_vec_17_right_subtree_state_3
    ; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_17_T_46 = {state_vec_0_set_left_older_3,_state_vec_17_T_34,_state_vec_17_T_45}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_18_valid = touch_ways_0_0_valid & touch_sets_0_0 == 5'h12; // @[Replacement.scala 315:30]
  wire  set_touch_ways_1_18_valid = touch_ways_0_1_valid & touch_sets_0_0 == 5'h12; // @[Replacement.scala 315:30]
  wire  _T_97 = set_touch_ways_0_18_valid | set_touch_ways_1_18_valid; // @[package.scala 72:59]
  wire [2:0] state_vec_18_left_subtree_state = state_vec__18[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_18_right_subtree_state = state_vec__18[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_18_left_subtree_state_1 = state_vec_18_left_subtree_state[1]; // @[package.scala 154:13]
  wire  state_vec_18_right_subtree_state_1 = state_vec_18_left_subtree_state[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_18_T_4 = state_vec_0_set_left_older_1 ? state_vec_18_left_subtree_state_1 : _state_vec_0_T_3; // @[Replacement.scala 203:16]
  wire  _state_vec_18_T_8 = state_vec_0_set_left_older_1 ? _state_vec_0_T_3 : state_vec_18_right_subtree_state_1; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_18_T_9 = {state_vec_0_set_left_older_1,_state_vec_18_T_4,_state_vec_18_T_8}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_18_T_10 = state_vec_0_set_left_older ? state_vec_18_left_subtree_state : _state_vec_18_T_9; // @[Replacement.scala 203:16]
  wire  state_vec_18_left_subtree_state_2 = state_vec_18_right_subtree_state[1]; // @[package.scala 154:13]
  wire  state_vec_18_right_subtree_state_2 = state_vec_18_right_subtree_state[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_18_T_15 = state_vec_0_set_left_older_1 ? state_vec_18_left_subtree_state_2 : _state_vec_0_T_3; // @[Replacement.scala 203:16]
  wire  _state_vec_18_T_19 = state_vec_0_set_left_older_1 ? _state_vec_0_T_3 : state_vec_18_right_subtree_state_2; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_18_T_20 = {state_vec_0_set_left_older_1,_state_vec_18_T_15,_state_vec_18_T_19}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_18_T_21 = state_vec_0_set_left_older ? _state_vec_18_T_20 : state_vec_18_right_subtree_state; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_18_T_22 = {state_vec_0_set_left_older,_state_vec_18_T_10,_state_vec_18_T_21}; // @[Cat.scala 31:58]
  wire [6:0] _state_vec_18_T_23 = set_touch_ways_0_18_valid ? _state_vec_18_T_22 : state_vec__18; // @[Replacement.scala 22:56]
  wire [2:0] state_vec_18_left_subtree_state_3 = _state_vec_18_T_23[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_18_right_subtree_state_3 = _state_vec_18_T_23[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_18_left_subtree_state_4 = state_vec_18_left_subtree_state_3[1]; // @[package.scala 154:13]
  wire  state_vec_18_right_subtree_state_4 = state_vec_18_left_subtree_state_3[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_18_T_28 = state_vec_0_set_left_older_4 ? state_vec_18_left_subtree_state_4 : _state_vec_0_T_27; // @[Replacement.scala 203:16]
  wire  _state_vec_18_T_32 = state_vec_0_set_left_older_4 ? _state_vec_0_T_27 : state_vec_18_right_subtree_state_4; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_18_T_33 = {state_vec_0_set_left_older_4,_state_vec_18_T_28,_state_vec_18_T_32}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_18_T_34 = state_vec_0_set_left_older_3 ? state_vec_18_left_subtree_state_3 : _state_vec_18_T_33; // @[Replacement.scala 203:16]
  wire  state_vec_18_left_subtree_state_5 = state_vec_18_right_subtree_state_3[1]; // @[package.scala 154:13]
  wire  state_vec_18_right_subtree_state_5 = state_vec_18_right_subtree_state_3[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_18_T_39 = state_vec_0_set_left_older_4 ? state_vec_18_left_subtree_state_5 : _state_vec_0_T_27; // @[Replacement.scala 203:16]
  wire  _state_vec_18_T_43 = state_vec_0_set_left_older_4 ? _state_vec_0_T_27 : state_vec_18_right_subtree_state_5; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_18_T_44 = {state_vec_0_set_left_older_4,_state_vec_18_T_39,_state_vec_18_T_43}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_18_T_45 = state_vec_0_set_left_older_3 ? _state_vec_18_T_44 : state_vec_18_right_subtree_state_3
    ; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_18_T_46 = {state_vec_0_set_left_older_3,_state_vec_18_T_34,_state_vec_18_T_45}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_19_valid = touch_ways_0_0_valid & touch_sets_0_0 == 5'h13; // @[Replacement.scala 315:30]
  wire  set_touch_ways_1_19_valid = touch_ways_0_1_valid & touch_sets_0_0 == 5'h13; // @[Replacement.scala 315:30]
  wire  _T_98 = set_touch_ways_0_19_valid | set_touch_ways_1_19_valid; // @[package.scala 72:59]
  wire [2:0] state_vec_19_left_subtree_state = state_vec__19[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_19_right_subtree_state = state_vec__19[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_19_left_subtree_state_1 = state_vec_19_left_subtree_state[1]; // @[package.scala 154:13]
  wire  state_vec_19_right_subtree_state_1 = state_vec_19_left_subtree_state[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_19_T_4 = state_vec_0_set_left_older_1 ? state_vec_19_left_subtree_state_1 : _state_vec_0_T_3; // @[Replacement.scala 203:16]
  wire  _state_vec_19_T_8 = state_vec_0_set_left_older_1 ? _state_vec_0_T_3 : state_vec_19_right_subtree_state_1; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_19_T_9 = {state_vec_0_set_left_older_1,_state_vec_19_T_4,_state_vec_19_T_8}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_19_T_10 = state_vec_0_set_left_older ? state_vec_19_left_subtree_state : _state_vec_19_T_9; // @[Replacement.scala 203:16]
  wire  state_vec_19_left_subtree_state_2 = state_vec_19_right_subtree_state[1]; // @[package.scala 154:13]
  wire  state_vec_19_right_subtree_state_2 = state_vec_19_right_subtree_state[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_19_T_15 = state_vec_0_set_left_older_1 ? state_vec_19_left_subtree_state_2 : _state_vec_0_T_3; // @[Replacement.scala 203:16]
  wire  _state_vec_19_T_19 = state_vec_0_set_left_older_1 ? _state_vec_0_T_3 : state_vec_19_right_subtree_state_2; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_19_T_20 = {state_vec_0_set_left_older_1,_state_vec_19_T_15,_state_vec_19_T_19}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_19_T_21 = state_vec_0_set_left_older ? _state_vec_19_T_20 : state_vec_19_right_subtree_state; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_19_T_22 = {state_vec_0_set_left_older,_state_vec_19_T_10,_state_vec_19_T_21}; // @[Cat.scala 31:58]
  wire [6:0] _state_vec_19_T_23 = set_touch_ways_0_19_valid ? _state_vec_19_T_22 : state_vec__19; // @[Replacement.scala 22:56]
  wire [2:0] state_vec_19_left_subtree_state_3 = _state_vec_19_T_23[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_19_right_subtree_state_3 = _state_vec_19_T_23[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_19_left_subtree_state_4 = state_vec_19_left_subtree_state_3[1]; // @[package.scala 154:13]
  wire  state_vec_19_right_subtree_state_4 = state_vec_19_left_subtree_state_3[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_19_T_28 = state_vec_0_set_left_older_4 ? state_vec_19_left_subtree_state_4 : _state_vec_0_T_27; // @[Replacement.scala 203:16]
  wire  _state_vec_19_T_32 = state_vec_0_set_left_older_4 ? _state_vec_0_T_27 : state_vec_19_right_subtree_state_4; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_19_T_33 = {state_vec_0_set_left_older_4,_state_vec_19_T_28,_state_vec_19_T_32}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_19_T_34 = state_vec_0_set_left_older_3 ? state_vec_19_left_subtree_state_3 : _state_vec_19_T_33; // @[Replacement.scala 203:16]
  wire  state_vec_19_left_subtree_state_5 = state_vec_19_right_subtree_state_3[1]; // @[package.scala 154:13]
  wire  state_vec_19_right_subtree_state_5 = state_vec_19_right_subtree_state_3[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_19_T_39 = state_vec_0_set_left_older_4 ? state_vec_19_left_subtree_state_5 : _state_vec_0_T_27; // @[Replacement.scala 203:16]
  wire  _state_vec_19_T_43 = state_vec_0_set_left_older_4 ? _state_vec_0_T_27 : state_vec_19_right_subtree_state_5; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_19_T_44 = {state_vec_0_set_left_older_4,_state_vec_19_T_39,_state_vec_19_T_43}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_19_T_45 = state_vec_0_set_left_older_3 ? _state_vec_19_T_44 : state_vec_19_right_subtree_state_3
    ; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_19_T_46 = {state_vec_0_set_left_older_3,_state_vec_19_T_34,_state_vec_19_T_45}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_20_valid = touch_ways_0_0_valid & touch_sets_0_0 == 5'h14; // @[Replacement.scala 315:30]
  wire  set_touch_ways_1_20_valid = touch_ways_0_1_valid & touch_sets_0_0 == 5'h14; // @[Replacement.scala 315:30]
  wire  _T_99 = set_touch_ways_0_20_valid | set_touch_ways_1_20_valid; // @[package.scala 72:59]
  wire [2:0] state_vec_20_left_subtree_state = state_vec__20[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_20_right_subtree_state = state_vec__20[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_20_left_subtree_state_1 = state_vec_20_left_subtree_state[1]; // @[package.scala 154:13]
  wire  state_vec_20_right_subtree_state_1 = state_vec_20_left_subtree_state[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_20_T_4 = state_vec_0_set_left_older_1 ? state_vec_20_left_subtree_state_1 : _state_vec_0_T_3; // @[Replacement.scala 203:16]
  wire  _state_vec_20_T_8 = state_vec_0_set_left_older_1 ? _state_vec_0_T_3 : state_vec_20_right_subtree_state_1; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_20_T_9 = {state_vec_0_set_left_older_1,_state_vec_20_T_4,_state_vec_20_T_8}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_20_T_10 = state_vec_0_set_left_older ? state_vec_20_left_subtree_state : _state_vec_20_T_9; // @[Replacement.scala 203:16]
  wire  state_vec_20_left_subtree_state_2 = state_vec_20_right_subtree_state[1]; // @[package.scala 154:13]
  wire  state_vec_20_right_subtree_state_2 = state_vec_20_right_subtree_state[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_20_T_15 = state_vec_0_set_left_older_1 ? state_vec_20_left_subtree_state_2 : _state_vec_0_T_3; // @[Replacement.scala 203:16]
  wire  _state_vec_20_T_19 = state_vec_0_set_left_older_1 ? _state_vec_0_T_3 : state_vec_20_right_subtree_state_2; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_20_T_20 = {state_vec_0_set_left_older_1,_state_vec_20_T_15,_state_vec_20_T_19}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_20_T_21 = state_vec_0_set_left_older ? _state_vec_20_T_20 : state_vec_20_right_subtree_state; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_20_T_22 = {state_vec_0_set_left_older,_state_vec_20_T_10,_state_vec_20_T_21}; // @[Cat.scala 31:58]
  wire [6:0] _state_vec_20_T_23 = set_touch_ways_0_20_valid ? _state_vec_20_T_22 : state_vec__20; // @[Replacement.scala 22:56]
  wire [2:0] state_vec_20_left_subtree_state_3 = _state_vec_20_T_23[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_20_right_subtree_state_3 = _state_vec_20_T_23[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_20_left_subtree_state_4 = state_vec_20_left_subtree_state_3[1]; // @[package.scala 154:13]
  wire  state_vec_20_right_subtree_state_4 = state_vec_20_left_subtree_state_3[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_20_T_28 = state_vec_0_set_left_older_4 ? state_vec_20_left_subtree_state_4 : _state_vec_0_T_27; // @[Replacement.scala 203:16]
  wire  _state_vec_20_T_32 = state_vec_0_set_left_older_4 ? _state_vec_0_T_27 : state_vec_20_right_subtree_state_4; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_20_T_33 = {state_vec_0_set_left_older_4,_state_vec_20_T_28,_state_vec_20_T_32}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_20_T_34 = state_vec_0_set_left_older_3 ? state_vec_20_left_subtree_state_3 : _state_vec_20_T_33; // @[Replacement.scala 203:16]
  wire  state_vec_20_left_subtree_state_5 = state_vec_20_right_subtree_state_3[1]; // @[package.scala 154:13]
  wire  state_vec_20_right_subtree_state_5 = state_vec_20_right_subtree_state_3[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_20_T_39 = state_vec_0_set_left_older_4 ? state_vec_20_left_subtree_state_5 : _state_vec_0_T_27; // @[Replacement.scala 203:16]
  wire  _state_vec_20_T_43 = state_vec_0_set_left_older_4 ? _state_vec_0_T_27 : state_vec_20_right_subtree_state_5; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_20_T_44 = {state_vec_0_set_left_older_4,_state_vec_20_T_39,_state_vec_20_T_43}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_20_T_45 = state_vec_0_set_left_older_3 ? _state_vec_20_T_44 : state_vec_20_right_subtree_state_3
    ; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_20_T_46 = {state_vec_0_set_left_older_3,_state_vec_20_T_34,_state_vec_20_T_45}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_21_valid = touch_ways_0_0_valid & touch_sets_0_0 == 5'h15; // @[Replacement.scala 315:30]
  wire  set_touch_ways_1_21_valid = touch_ways_0_1_valid & touch_sets_0_0 == 5'h15; // @[Replacement.scala 315:30]
  wire  _T_100 = set_touch_ways_0_21_valid | set_touch_ways_1_21_valid; // @[package.scala 72:59]
  wire [2:0] state_vec_21_left_subtree_state = state_vec__21[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_21_right_subtree_state = state_vec__21[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_21_left_subtree_state_1 = state_vec_21_left_subtree_state[1]; // @[package.scala 154:13]
  wire  state_vec_21_right_subtree_state_1 = state_vec_21_left_subtree_state[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_21_T_4 = state_vec_0_set_left_older_1 ? state_vec_21_left_subtree_state_1 : _state_vec_0_T_3; // @[Replacement.scala 203:16]
  wire  _state_vec_21_T_8 = state_vec_0_set_left_older_1 ? _state_vec_0_T_3 : state_vec_21_right_subtree_state_1; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_21_T_9 = {state_vec_0_set_left_older_1,_state_vec_21_T_4,_state_vec_21_T_8}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_21_T_10 = state_vec_0_set_left_older ? state_vec_21_left_subtree_state : _state_vec_21_T_9; // @[Replacement.scala 203:16]
  wire  state_vec_21_left_subtree_state_2 = state_vec_21_right_subtree_state[1]; // @[package.scala 154:13]
  wire  state_vec_21_right_subtree_state_2 = state_vec_21_right_subtree_state[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_21_T_15 = state_vec_0_set_left_older_1 ? state_vec_21_left_subtree_state_2 : _state_vec_0_T_3; // @[Replacement.scala 203:16]
  wire  _state_vec_21_T_19 = state_vec_0_set_left_older_1 ? _state_vec_0_T_3 : state_vec_21_right_subtree_state_2; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_21_T_20 = {state_vec_0_set_left_older_1,_state_vec_21_T_15,_state_vec_21_T_19}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_21_T_21 = state_vec_0_set_left_older ? _state_vec_21_T_20 : state_vec_21_right_subtree_state; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_21_T_22 = {state_vec_0_set_left_older,_state_vec_21_T_10,_state_vec_21_T_21}; // @[Cat.scala 31:58]
  wire [6:0] _state_vec_21_T_23 = set_touch_ways_0_21_valid ? _state_vec_21_T_22 : state_vec__21; // @[Replacement.scala 22:56]
  wire [2:0] state_vec_21_left_subtree_state_3 = _state_vec_21_T_23[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_21_right_subtree_state_3 = _state_vec_21_T_23[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_21_left_subtree_state_4 = state_vec_21_left_subtree_state_3[1]; // @[package.scala 154:13]
  wire  state_vec_21_right_subtree_state_4 = state_vec_21_left_subtree_state_3[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_21_T_28 = state_vec_0_set_left_older_4 ? state_vec_21_left_subtree_state_4 : _state_vec_0_T_27; // @[Replacement.scala 203:16]
  wire  _state_vec_21_T_32 = state_vec_0_set_left_older_4 ? _state_vec_0_T_27 : state_vec_21_right_subtree_state_4; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_21_T_33 = {state_vec_0_set_left_older_4,_state_vec_21_T_28,_state_vec_21_T_32}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_21_T_34 = state_vec_0_set_left_older_3 ? state_vec_21_left_subtree_state_3 : _state_vec_21_T_33; // @[Replacement.scala 203:16]
  wire  state_vec_21_left_subtree_state_5 = state_vec_21_right_subtree_state_3[1]; // @[package.scala 154:13]
  wire  state_vec_21_right_subtree_state_5 = state_vec_21_right_subtree_state_3[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_21_T_39 = state_vec_0_set_left_older_4 ? state_vec_21_left_subtree_state_5 : _state_vec_0_T_27; // @[Replacement.scala 203:16]
  wire  _state_vec_21_T_43 = state_vec_0_set_left_older_4 ? _state_vec_0_T_27 : state_vec_21_right_subtree_state_5; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_21_T_44 = {state_vec_0_set_left_older_4,_state_vec_21_T_39,_state_vec_21_T_43}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_21_T_45 = state_vec_0_set_left_older_3 ? _state_vec_21_T_44 : state_vec_21_right_subtree_state_3
    ; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_21_T_46 = {state_vec_0_set_left_older_3,_state_vec_21_T_34,_state_vec_21_T_45}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_22_valid = touch_ways_0_0_valid & touch_sets_0_0 == 5'h16; // @[Replacement.scala 315:30]
  wire  set_touch_ways_1_22_valid = touch_ways_0_1_valid & touch_sets_0_0 == 5'h16; // @[Replacement.scala 315:30]
  wire  _T_101 = set_touch_ways_0_22_valid | set_touch_ways_1_22_valid; // @[package.scala 72:59]
  wire [2:0] state_vec_22_left_subtree_state = state_vec__22[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_22_right_subtree_state = state_vec__22[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_22_left_subtree_state_1 = state_vec_22_left_subtree_state[1]; // @[package.scala 154:13]
  wire  state_vec_22_right_subtree_state_1 = state_vec_22_left_subtree_state[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_22_T_4 = state_vec_0_set_left_older_1 ? state_vec_22_left_subtree_state_1 : _state_vec_0_T_3; // @[Replacement.scala 203:16]
  wire  _state_vec_22_T_8 = state_vec_0_set_left_older_1 ? _state_vec_0_T_3 : state_vec_22_right_subtree_state_1; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_22_T_9 = {state_vec_0_set_left_older_1,_state_vec_22_T_4,_state_vec_22_T_8}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_22_T_10 = state_vec_0_set_left_older ? state_vec_22_left_subtree_state : _state_vec_22_T_9; // @[Replacement.scala 203:16]
  wire  state_vec_22_left_subtree_state_2 = state_vec_22_right_subtree_state[1]; // @[package.scala 154:13]
  wire  state_vec_22_right_subtree_state_2 = state_vec_22_right_subtree_state[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_22_T_15 = state_vec_0_set_left_older_1 ? state_vec_22_left_subtree_state_2 : _state_vec_0_T_3; // @[Replacement.scala 203:16]
  wire  _state_vec_22_T_19 = state_vec_0_set_left_older_1 ? _state_vec_0_T_3 : state_vec_22_right_subtree_state_2; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_22_T_20 = {state_vec_0_set_left_older_1,_state_vec_22_T_15,_state_vec_22_T_19}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_22_T_21 = state_vec_0_set_left_older ? _state_vec_22_T_20 : state_vec_22_right_subtree_state; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_22_T_22 = {state_vec_0_set_left_older,_state_vec_22_T_10,_state_vec_22_T_21}; // @[Cat.scala 31:58]
  wire [6:0] _state_vec_22_T_23 = set_touch_ways_0_22_valid ? _state_vec_22_T_22 : state_vec__22; // @[Replacement.scala 22:56]
  wire [2:0] state_vec_22_left_subtree_state_3 = _state_vec_22_T_23[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_22_right_subtree_state_3 = _state_vec_22_T_23[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_22_left_subtree_state_4 = state_vec_22_left_subtree_state_3[1]; // @[package.scala 154:13]
  wire  state_vec_22_right_subtree_state_4 = state_vec_22_left_subtree_state_3[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_22_T_28 = state_vec_0_set_left_older_4 ? state_vec_22_left_subtree_state_4 : _state_vec_0_T_27; // @[Replacement.scala 203:16]
  wire  _state_vec_22_T_32 = state_vec_0_set_left_older_4 ? _state_vec_0_T_27 : state_vec_22_right_subtree_state_4; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_22_T_33 = {state_vec_0_set_left_older_4,_state_vec_22_T_28,_state_vec_22_T_32}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_22_T_34 = state_vec_0_set_left_older_3 ? state_vec_22_left_subtree_state_3 : _state_vec_22_T_33; // @[Replacement.scala 203:16]
  wire  state_vec_22_left_subtree_state_5 = state_vec_22_right_subtree_state_3[1]; // @[package.scala 154:13]
  wire  state_vec_22_right_subtree_state_5 = state_vec_22_right_subtree_state_3[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_22_T_39 = state_vec_0_set_left_older_4 ? state_vec_22_left_subtree_state_5 : _state_vec_0_T_27; // @[Replacement.scala 203:16]
  wire  _state_vec_22_T_43 = state_vec_0_set_left_older_4 ? _state_vec_0_T_27 : state_vec_22_right_subtree_state_5; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_22_T_44 = {state_vec_0_set_left_older_4,_state_vec_22_T_39,_state_vec_22_T_43}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_22_T_45 = state_vec_0_set_left_older_3 ? _state_vec_22_T_44 : state_vec_22_right_subtree_state_3
    ; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_22_T_46 = {state_vec_0_set_left_older_3,_state_vec_22_T_34,_state_vec_22_T_45}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_23_valid = touch_ways_0_0_valid & touch_sets_0_0 == 5'h17; // @[Replacement.scala 315:30]
  wire  set_touch_ways_1_23_valid = touch_ways_0_1_valid & touch_sets_0_0 == 5'h17; // @[Replacement.scala 315:30]
  wire  _T_102 = set_touch_ways_0_23_valid | set_touch_ways_1_23_valid; // @[package.scala 72:59]
  wire [2:0] state_vec_23_left_subtree_state = state_vec__23[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_23_right_subtree_state = state_vec__23[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_23_left_subtree_state_1 = state_vec_23_left_subtree_state[1]; // @[package.scala 154:13]
  wire  state_vec_23_right_subtree_state_1 = state_vec_23_left_subtree_state[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_23_T_4 = state_vec_0_set_left_older_1 ? state_vec_23_left_subtree_state_1 : _state_vec_0_T_3; // @[Replacement.scala 203:16]
  wire  _state_vec_23_T_8 = state_vec_0_set_left_older_1 ? _state_vec_0_T_3 : state_vec_23_right_subtree_state_1; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_23_T_9 = {state_vec_0_set_left_older_1,_state_vec_23_T_4,_state_vec_23_T_8}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_23_T_10 = state_vec_0_set_left_older ? state_vec_23_left_subtree_state : _state_vec_23_T_9; // @[Replacement.scala 203:16]
  wire  state_vec_23_left_subtree_state_2 = state_vec_23_right_subtree_state[1]; // @[package.scala 154:13]
  wire  state_vec_23_right_subtree_state_2 = state_vec_23_right_subtree_state[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_23_T_15 = state_vec_0_set_left_older_1 ? state_vec_23_left_subtree_state_2 : _state_vec_0_T_3; // @[Replacement.scala 203:16]
  wire  _state_vec_23_T_19 = state_vec_0_set_left_older_1 ? _state_vec_0_T_3 : state_vec_23_right_subtree_state_2; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_23_T_20 = {state_vec_0_set_left_older_1,_state_vec_23_T_15,_state_vec_23_T_19}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_23_T_21 = state_vec_0_set_left_older ? _state_vec_23_T_20 : state_vec_23_right_subtree_state; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_23_T_22 = {state_vec_0_set_left_older,_state_vec_23_T_10,_state_vec_23_T_21}; // @[Cat.scala 31:58]
  wire [6:0] _state_vec_23_T_23 = set_touch_ways_0_23_valid ? _state_vec_23_T_22 : state_vec__23; // @[Replacement.scala 22:56]
  wire [2:0] state_vec_23_left_subtree_state_3 = _state_vec_23_T_23[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_23_right_subtree_state_3 = _state_vec_23_T_23[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_23_left_subtree_state_4 = state_vec_23_left_subtree_state_3[1]; // @[package.scala 154:13]
  wire  state_vec_23_right_subtree_state_4 = state_vec_23_left_subtree_state_3[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_23_T_28 = state_vec_0_set_left_older_4 ? state_vec_23_left_subtree_state_4 : _state_vec_0_T_27; // @[Replacement.scala 203:16]
  wire  _state_vec_23_T_32 = state_vec_0_set_left_older_4 ? _state_vec_0_T_27 : state_vec_23_right_subtree_state_4; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_23_T_33 = {state_vec_0_set_left_older_4,_state_vec_23_T_28,_state_vec_23_T_32}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_23_T_34 = state_vec_0_set_left_older_3 ? state_vec_23_left_subtree_state_3 : _state_vec_23_T_33; // @[Replacement.scala 203:16]
  wire  state_vec_23_left_subtree_state_5 = state_vec_23_right_subtree_state_3[1]; // @[package.scala 154:13]
  wire  state_vec_23_right_subtree_state_5 = state_vec_23_right_subtree_state_3[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_23_T_39 = state_vec_0_set_left_older_4 ? state_vec_23_left_subtree_state_5 : _state_vec_0_T_27; // @[Replacement.scala 203:16]
  wire  _state_vec_23_T_43 = state_vec_0_set_left_older_4 ? _state_vec_0_T_27 : state_vec_23_right_subtree_state_5; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_23_T_44 = {state_vec_0_set_left_older_4,_state_vec_23_T_39,_state_vec_23_T_43}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_23_T_45 = state_vec_0_set_left_older_3 ? _state_vec_23_T_44 : state_vec_23_right_subtree_state_3
    ; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_23_T_46 = {state_vec_0_set_left_older_3,_state_vec_23_T_34,_state_vec_23_T_45}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_24_valid = touch_ways_0_0_valid & touch_sets_0_0 == 5'h18; // @[Replacement.scala 315:30]
  wire  set_touch_ways_1_24_valid = touch_ways_0_1_valid & touch_sets_0_0 == 5'h18; // @[Replacement.scala 315:30]
  wire  _T_103 = set_touch_ways_0_24_valid | set_touch_ways_1_24_valid; // @[package.scala 72:59]
  wire [2:0] state_vec_24_left_subtree_state = state_vec__24[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_24_right_subtree_state = state_vec__24[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_24_left_subtree_state_1 = state_vec_24_left_subtree_state[1]; // @[package.scala 154:13]
  wire  state_vec_24_right_subtree_state_1 = state_vec_24_left_subtree_state[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_24_T_4 = state_vec_0_set_left_older_1 ? state_vec_24_left_subtree_state_1 : _state_vec_0_T_3; // @[Replacement.scala 203:16]
  wire  _state_vec_24_T_8 = state_vec_0_set_left_older_1 ? _state_vec_0_T_3 : state_vec_24_right_subtree_state_1; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_24_T_9 = {state_vec_0_set_left_older_1,_state_vec_24_T_4,_state_vec_24_T_8}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_24_T_10 = state_vec_0_set_left_older ? state_vec_24_left_subtree_state : _state_vec_24_T_9; // @[Replacement.scala 203:16]
  wire  state_vec_24_left_subtree_state_2 = state_vec_24_right_subtree_state[1]; // @[package.scala 154:13]
  wire  state_vec_24_right_subtree_state_2 = state_vec_24_right_subtree_state[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_24_T_15 = state_vec_0_set_left_older_1 ? state_vec_24_left_subtree_state_2 : _state_vec_0_T_3; // @[Replacement.scala 203:16]
  wire  _state_vec_24_T_19 = state_vec_0_set_left_older_1 ? _state_vec_0_T_3 : state_vec_24_right_subtree_state_2; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_24_T_20 = {state_vec_0_set_left_older_1,_state_vec_24_T_15,_state_vec_24_T_19}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_24_T_21 = state_vec_0_set_left_older ? _state_vec_24_T_20 : state_vec_24_right_subtree_state; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_24_T_22 = {state_vec_0_set_left_older,_state_vec_24_T_10,_state_vec_24_T_21}; // @[Cat.scala 31:58]
  wire [6:0] _state_vec_24_T_23 = set_touch_ways_0_24_valid ? _state_vec_24_T_22 : state_vec__24; // @[Replacement.scala 22:56]
  wire [2:0] state_vec_24_left_subtree_state_3 = _state_vec_24_T_23[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_24_right_subtree_state_3 = _state_vec_24_T_23[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_24_left_subtree_state_4 = state_vec_24_left_subtree_state_3[1]; // @[package.scala 154:13]
  wire  state_vec_24_right_subtree_state_4 = state_vec_24_left_subtree_state_3[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_24_T_28 = state_vec_0_set_left_older_4 ? state_vec_24_left_subtree_state_4 : _state_vec_0_T_27; // @[Replacement.scala 203:16]
  wire  _state_vec_24_T_32 = state_vec_0_set_left_older_4 ? _state_vec_0_T_27 : state_vec_24_right_subtree_state_4; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_24_T_33 = {state_vec_0_set_left_older_4,_state_vec_24_T_28,_state_vec_24_T_32}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_24_T_34 = state_vec_0_set_left_older_3 ? state_vec_24_left_subtree_state_3 : _state_vec_24_T_33; // @[Replacement.scala 203:16]
  wire  state_vec_24_left_subtree_state_5 = state_vec_24_right_subtree_state_3[1]; // @[package.scala 154:13]
  wire  state_vec_24_right_subtree_state_5 = state_vec_24_right_subtree_state_3[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_24_T_39 = state_vec_0_set_left_older_4 ? state_vec_24_left_subtree_state_5 : _state_vec_0_T_27; // @[Replacement.scala 203:16]
  wire  _state_vec_24_T_43 = state_vec_0_set_left_older_4 ? _state_vec_0_T_27 : state_vec_24_right_subtree_state_5; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_24_T_44 = {state_vec_0_set_left_older_4,_state_vec_24_T_39,_state_vec_24_T_43}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_24_T_45 = state_vec_0_set_left_older_3 ? _state_vec_24_T_44 : state_vec_24_right_subtree_state_3
    ; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_24_T_46 = {state_vec_0_set_left_older_3,_state_vec_24_T_34,_state_vec_24_T_45}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_25_valid = touch_ways_0_0_valid & touch_sets_0_0 == 5'h19; // @[Replacement.scala 315:30]
  wire  set_touch_ways_1_25_valid = touch_ways_0_1_valid & touch_sets_0_0 == 5'h19; // @[Replacement.scala 315:30]
  wire  _T_104 = set_touch_ways_0_25_valid | set_touch_ways_1_25_valid; // @[package.scala 72:59]
  wire [2:0] state_vec_25_left_subtree_state = state_vec__25[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_25_right_subtree_state = state_vec__25[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_25_left_subtree_state_1 = state_vec_25_left_subtree_state[1]; // @[package.scala 154:13]
  wire  state_vec_25_right_subtree_state_1 = state_vec_25_left_subtree_state[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_25_T_4 = state_vec_0_set_left_older_1 ? state_vec_25_left_subtree_state_1 : _state_vec_0_T_3; // @[Replacement.scala 203:16]
  wire  _state_vec_25_T_8 = state_vec_0_set_left_older_1 ? _state_vec_0_T_3 : state_vec_25_right_subtree_state_1; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_25_T_9 = {state_vec_0_set_left_older_1,_state_vec_25_T_4,_state_vec_25_T_8}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_25_T_10 = state_vec_0_set_left_older ? state_vec_25_left_subtree_state : _state_vec_25_T_9; // @[Replacement.scala 203:16]
  wire  state_vec_25_left_subtree_state_2 = state_vec_25_right_subtree_state[1]; // @[package.scala 154:13]
  wire  state_vec_25_right_subtree_state_2 = state_vec_25_right_subtree_state[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_25_T_15 = state_vec_0_set_left_older_1 ? state_vec_25_left_subtree_state_2 : _state_vec_0_T_3; // @[Replacement.scala 203:16]
  wire  _state_vec_25_T_19 = state_vec_0_set_left_older_1 ? _state_vec_0_T_3 : state_vec_25_right_subtree_state_2; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_25_T_20 = {state_vec_0_set_left_older_1,_state_vec_25_T_15,_state_vec_25_T_19}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_25_T_21 = state_vec_0_set_left_older ? _state_vec_25_T_20 : state_vec_25_right_subtree_state; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_25_T_22 = {state_vec_0_set_left_older,_state_vec_25_T_10,_state_vec_25_T_21}; // @[Cat.scala 31:58]
  wire [6:0] _state_vec_25_T_23 = set_touch_ways_0_25_valid ? _state_vec_25_T_22 : state_vec__25; // @[Replacement.scala 22:56]
  wire [2:0] state_vec_25_left_subtree_state_3 = _state_vec_25_T_23[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_25_right_subtree_state_3 = _state_vec_25_T_23[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_25_left_subtree_state_4 = state_vec_25_left_subtree_state_3[1]; // @[package.scala 154:13]
  wire  state_vec_25_right_subtree_state_4 = state_vec_25_left_subtree_state_3[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_25_T_28 = state_vec_0_set_left_older_4 ? state_vec_25_left_subtree_state_4 : _state_vec_0_T_27; // @[Replacement.scala 203:16]
  wire  _state_vec_25_T_32 = state_vec_0_set_left_older_4 ? _state_vec_0_T_27 : state_vec_25_right_subtree_state_4; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_25_T_33 = {state_vec_0_set_left_older_4,_state_vec_25_T_28,_state_vec_25_T_32}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_25_T_34 = state_vec_0_set_left_older_3 ? state_vec_25_left_subtree_state_3 : _state_vec_25_T_33; // @[Replacement.scala 203:16]
  wire  state_vec_25_left_subtree_state_5 = state_vec_25_right_subtree_state_3[1]; // @[package.scala 154:13]
  wire  state_vec_25_right_subtree_state_5 = state_vec_25_right_subtree_state_3[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_25_T_39 = state_vec_0_set_left_older_4 ? state_vec_25_left_subtree_state_5 : _state_vec_0_T_27; // @[Replacement.scala 203:16]
  wire  _state_vec_25_T_43 = state_vec_0_set_left_older_4 ? _state_vec_0_T_27 : state_vec_25_right_subtree_state_5; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_25_T_44 = {state_vec_0_set_left_older_4,_state_vec_25_T_39,_state_vec_25_T_43}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_25_T_45 = state_vec_0_set_left_older_3 ? _state_vec_25_T_44 : state_vec_25_right_subtree_state_3
    ; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_25_T_46 = {state_vec_0_set_left_older_3,_state_vec_25_T_34,_state_vec_25_T_45}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_26_valid = touch_ways_0_0_valid & touch_sets_0_0 == 5'h1a; // @[Replacement.scala 315:30]
  wire  set_touch_ways_1_26_valid = touch_ways_0_1_valid & touch_sets_0_0 == 5'h1a; // @[Replacement.scala 315:30]
  wire  _T_105 = set_touch_ways_0_26_valid | set_touch_ways_1_26_valid; // @[package.scala 72:59]
  wire [2:0] state_vec_26_left_subtree_state = state_vec__26[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_26_right_subtree_state = state_vec__26[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_26_left_subtree_state_1 = state_vec_26_left_subtree_state[1]; // @[package.scala 154:13]
  wire  state_vec_26_right_subtree_state_1 = state_vec_26_left_subtree_state[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_26_T_4 = state_vec_0_set_left_older_1 ? state_vec_26_left_subtree_state_1 : _state_vec_0_T_3; // @[Replacement.scala 203:16]
  wire  _state_vec_26_T_8 = state_vec_0_set_left_older_1 ? _state_vec_0_T_3 : state_vec_26_right_subtree_state_1; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_26_T_9 = {state_vec_0_set_left_older_1,_state_vec_26_T_4,_state_vec_26_T_8}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_26_T_10 = state_vec_0_set_left_older ? state_vec_26_left_subtree_state : _state_vec_26_T_9; // @[Replacement.scala 203:16]
  wire  state_vec_26_left_subtree_state_2 = state_vec_26_right_subtree_state[1]; // @[package.scala 154:13]
  wire  state_vec_26_right_subtree_state_2 = state_vec_26_right_subtree_state[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_26_T_15 = state_vec_0_set_left_older_1 ? state_vec_26_left_subtree_state_2 : _state_vec_0_T_3; // @[Replacement.scala 203:16]
  wire  _state_vec_26_T_19 = state_vec_0_set_left_older_1 ? _state_vec_0_T_3 : state_vec_26_right_subtree_state_2; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_26_T_20 = {state_vec_0_set_left_older_1,_state_vec_26_T_15,_state_vec_26_T_19}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_26_T_21 = state_vec_0_set_left_older ? _state_vec_26_T_20 : state_vec_26_right_subtree_state; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_26_T_22 = {state_vec_0_set_left_older,_state_vec_26_T_10,_state_vec_26_T_21}; // @[Cat.scala 31:58]
  wire [6:0] _state_vec_26_T_23 = set_touch_ways_0_26_valid ? _state_vec_26_T_22 : state_vec__26; // @[Replacement.scala 22:56]
  wire [2:0] state_vec_26_left_subtree_state_3 = _state_vec_26_T_23[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_26_right_subtree_state_3 = _state_vec_26_T_23[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_26_left_subtree_state_4 = state_vec_26_left_subtree_state_3[1]; // @[package.scala 154:13]
  wire  state_vec_26_right_subtree_state_4 = state_vec_26_left_subtree_state_3[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_26_T_28 = state_vec_0_set_left_older_4 ? state_vec_26_left_subtree_state_4 : _state_vec_0_T_27; // @[Replacement.scala 203:16]
  wire  _state_vec_26_T_32 = state_vec_0_set_left_older_4 ? _state_vec_0_T_27 : state_vec_26_right_subtree_state_4; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_26_T_33 = {state_vec_0_set_left_older_4,_state_vec_26_T_28,_state_vec_26_T_32}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_26_T_34 = state_vec_0_set_left_older_3 ? state_vec_26_left_subtree_state_3 : _state_vec_26_T_33; // @[Replacement.scala 203:16]
  wire  state_vec_26_left_subtree_state_5 = state_vec_26_right_subtree_state_3[1]; // @[package.scala 154:13]
  wire  state_vec_26_right_subtree_state_5 = state_vec_26_right_subtree_state_3[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_26_T_39 = state_vec_0_set_left_older_4 ? state_vec_26_left_subtree_state_5 : _state_vec_0_T_27; // @[Replacement.scala 203:16]
  wire  _state_vec_26_T_43 = state_vec_0_set_left_older_4 ? _state_vec_0_T_27 : state_vec_26_right_subtree_state_5; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_26_T_44 = {state_vec_0_set_left_older_4,_state_vec_26_T_39,_state_vec_26_T_43}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_26_T_45 = state_vec_0_set_left_older_3 ? _state_vec_26_T_44 : state_vec_26_right_subtree_state_3
    ; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_26_T_46 = {state_vec_0_set_left_older_3,_state_vec_26_T_34,_state_vec_26_T_45}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_27_valid = touch_ways_0_0_valid & touch_sets_0_0 == 5'h1b; // @[Replacement.scala 315:30]
  wire  set_touch_ways_1_27_valid = touch_ways_0_1_valid & touch_sets_0_0 == 5'h1b; // @[Replacement.scala 315:30]
  wire  _T_106 = set_touch_ways_0_27_valid | set_touch_ways_1_27_valid; // @[package.scala 72:59]
  wire [2:0] state_vec_27_left_subtree_state = state_vec__27[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_27_right_subtree_state = state_vec__27[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_27_left_subtree_state_1 = state_vec_27_left_subtree_state[1]; // @[package.scala 154:13]
  wire  state_vec_27_right_subtree_state_1 = state_vec_27_left_subtree_state[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_27_T_4 = state_vec_0_set_left_older_1 ? state_vec_27_left_subtree_state_1 : _state_vec_0_T_3; // @[Replacement.scala 203:16]
  wire  _state_vec_27_T_8 = state_vec_0_set_left_older_1 ? _state_vec_0_T_3 : state_vec_27_right_subtree_state_1; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_27_T_9 = {state_vec_0_set_left_older_1,_state_vec_27_T_4,_state_vec_27_T_8}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_27_T_10 = state_vec_0_set_left_older ? state_vec_27_left_subtree_state : _state_vec_27_T_9; // @[Replacement.scala 203:16]
  wire  state_vec_27_left_subtree_state_2 = state_vec_27_right_subtree_state[1]; // @[package.scala 154:13]
  wire  state_vec_27_right_subtree_state_2 = state_vec_27_right_subtree_state[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_27_T_15 = state_vec_0_set_left_older_1 ? state_vec_27_left_subtree_state_2 : _state_vec_0_T_3; // @[Replacement.scala 203:16]
  wire  _state_vec_27_T_19 = state_vec_0_set_left_older_1 ? _state_vec_0_T_3 : state_vec_27_right_subtree_state_2; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_27_T_20 = {state_vec_0_set_left_older_1,_state_vec_27_T_15,_state_vec_27_T_19}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_27_T_21 = state_vec_0_set_left_older ? _state_vec_27_T_20 : state_vec_27_right_subtree_state; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_27_T_22 = {state_vec_0_set_left_older,_state_vec_27_T_10,_state_vec_27_T_21}; // @[Cat.scala 31:58]
  wire [6:0] _state_vec_27_T_23 = set_touch_ways_0_27_valid ? _state_vec_27_T_22 : state_vec__27; // @[Replacement.scala 22:56]
  wire [2:0] state_vec_27_left_subtree_state_3 = _state_vec_27_T_23[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_27_right_subtree_state_3 = _state_vec_27_T_23[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_27_left_subtree_state_4 = state_vec_27_left_subtree_state_3[1]; // @[package.scala 154:13]
  wire  state_vec_27_right_subtree_state_4 = state_vec_27_left_subtree_state_3[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_27_T_28 = state_vec_0_set_left_older_4 ? state_vec_27_left_subtree_state_4 : _state_vec_0_T_27; // @[Replacement.scala 203:16]
  wire  _state_vec_27_T_32 = state_vec_0_set_left_older_4 ? _state_vec_0_T_27 : state_vec_27_right_subtree_state_4; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_27_T_33 = {state_vec_0_set_left_older_4,_state_vec_27_T_28,_state_vec_27_T_32}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_27_T_34 = state_vec_0_set_left_older_3 ? state_vec_27_left_subtree_state_3 : _state_vec_27_T_33; // @[Replacement.scala 203:16]
  wire  state_vec_27_left_subtree_state_5 = state_vec_27_right_subtree_state_3[1]; // @[package.scala 154:13]
  wire  state_vec_27_right_subtree_state_5 = state_vec_27_right_subtree_state_3[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_27_T_39 = state_vec_0_set_left_older_4 ? state_vec_27_left_subtree_state_5 : _state_vec_0_T_27; // @[Replacement.scala 203:16]
  wire  _state_vec_27_T_43 = state_vec_0_set_left_older_4 ? _state_vec_0_T_27 : state_vec_27_right_subtree_state_5; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_27_T_44 = {state_vec_0_set_left_older_4,_state_vec_27_T_39,_state_vec_27_T_43}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_27_T_45 = state_vec_0_set_left_older_3 ? _state_vec_27_T_44 : state_vec_27_right_subtree_state_3
    ; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_27_T_46 = {state_vec_0_set_left_older_3,_state_vec_27_T_34,_state_vec_27_T_45}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_28_valid = touch_ways_0_0_valid & touch_sets_0_0 == 5'h1c; // @[Replacement.scala 315:30]
  wire  set_touch_ways_1_28_valid = touch_ways_0_1_valid & touch_sets_0_0 == 5'h1c; // @[Replacement.scala 315:30]
  wire  _T_107 = set_touch_ways_0_28_valid | set_touch_ways_1_28_valid; // @[package.scala 72:59]
  wire [2:0] state_vec_28_left_subtree_state = state_vec__28[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_28_right_subtree_state = state_vec__28[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_28_left_subtree_state_1 = state_vec_28_left_subtree_state[1]; // @[package.scala 154:13]
  wire  state_vec_28_right_subtree_state_1 = state_vec_28_left_subtree_state[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_28_T_4 = state_vec_0_set_left_older_1 ? state_vec_28_left_subtree_state_1 : _state_vec_0_T_3; // @[Replacement.scala 203:16]
  wire  _state_vec_28_T_8 = state_vec_0_set_left_older_1 ? _state_vec_0_T_3 : state_vec_28_right_subtree_state_1; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_28_T_9 = {state_vec_0_set_left_older_1,_state_vec_28_T_4,_state_vec_28_T_8}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_28_T_10 = state_vec_0_set_left_older ? state_vec_28_left_subtree_state : _state_vec_28_T_9; // @[Replacement.scala 203:16]
  wire  state_vec_28_left_subtree_state_2 = state_vec_28_right_subtree_state[1]; // @[package.scala 154:13]
  wire  state_vec_28_right_subtree_state_2 = state_vec_28_right_subtree_state[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_28_T_15 = state_vec_0_set_left_older_1 ? state_vec_28_left_subtree_state_2 : _state_vec_0_T_3; // @[Replacement.scala 203:16]
  wire  _state_vec_28_T_19 = state_vec_0_set_left_older_1 ? _state_vec_0_T_3 : state_vec_28_right_subtree_state_2; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_28_T_20 = {state_vec_0_set_left_older_1,_state_vec_28_T_15,_state_vec_28_T_19}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_28_T_21 = state_vec_0_set_left_older ? _state_vec_28_T_20 : state_vec_28_right_subtree_state; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_28_T_22 = {state_vec_0_set_left_older,_state_vec_28_T_10,_state_vec_28_T_21}; // @[Cat.scala 31:58]
  wire [6:0] _state_vec_28_T_23 = set_touch_ways_0_28_valid ? _state_vec_28_T_22 : state_vec__28; // @[Replacement.scala 22:56]
  wire [2:0] state_vec_28_left_subtree_state_3 = _state_vec_28_T_23[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_28_right_subtree_state_3 = _state_vec_28_T_23[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_28_left_subtree_state_4 = state_vec_28_left_subtree_state_3[1]; // @[package.scala 154:13]
  wire  state_vec_28_right_subtree_state_4 = state_vec_28_left_subtree_state_3[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_28_T_28 = state_vec_0_set_left_older_4 ? state_vec_28_left_subtree_state_4 : _state_vec_0_T_27; // @[Replacement.scala 203:16]
  wire  _state_vec_28_T_32 = state_vec_0_set_left_older_4 ? _state_vec_0_T_27 : state_vec_28_right_subtree_state_4; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_28_T_33 = {state_vec_0_set_left_older_4,_state_vec_28_T_28,_state_vec_28_T_32}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_28_T_34 = state_vec_0_set_left_older_3 ? state_vec_28_left_subtree_state_3 : _state_vec_28_T_33; // @[Replacement.scala 203:16]
  wire  state_vec_28_left_subtree_state_5 = state_vec_28_right_subtree_state_3[1]; // @[package.scala 154:13]
  wire  state_vec_28_right_subtree_state_5 = state_vec_28_right_subtree_state_3[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_28_T_39 = state_vec_0_set_left_older_4 ? state_vec_28_left_subtree_state_5 : _state_vec_0_T_27; // @[Replacement.scala 203:16]
  wire  _state_vec_28_T_43 = state_vec_0_set_left_older_4 ? _state_vec_0_T_27 : state_vec_28_right_subtree_state_5; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_28_T_44 = {state_vec_0_set_left_older_4,_state_vec_28_T_39,_state_vec_28_T_43}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_28_T_45 = state_vec_0_set_left_older_3 ? _state_vec_28_T_44 : state_vec_28_right_subtree_state_3
    ; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_28_T_46 = {state_vec_0_set_left_older_3,_state_vec_28_T_34,_state_vec_28_T_45}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_29_valid = touch_ways_0_0_valid & touch_sets_0_0 == 5'h1d; // @[Replacement.scala 315:30]
  wire  set_touch_ways_1_29_valid = touch_ways_0_1_valid & touch_sets_0_0 == 5'h1d; // @[Replacement.scala 315:30]
  wire  _T_108 = set_touch_ways_0_29_valid | set_touch_ways_1_29_valid; // @[package.scala 72:59]
  wire [2:0] state_vec_29_left_subtree_state = state_vec__29[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_29_right_subtree_state = state_vec__29[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_29_left_subtree_state_1 = state_vec_29_left_subtree_state[1]; // @[package.scala 154:13]
  wire  state_vec_29_right_subtree_state_1 = state_vec_29_left_subtree_state[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_29_T_4 = state_vec_0_set_left_older_1 ? state_vec_29_left_subtree_state_1 : _state_vec_0_T_3; // @[Replacement.scala 203:16]
  wire  _state_vec_29_T_8 = state_vec_0_set_left_older_1 ? _state_vec_0_T_3 : state_vec_29_right_subtree_state_1; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_29_T_9 = {state_vec_0_set_left_older_1,_state_vec_29_T_4,_state_vec_29_T_8}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_29_T_10 = state_vec_0_set_left_older ? state_vec_29_left_subtree_state : _state_vec_29_T_9; // @[Replacement.scala 203:16]
  wire  state_vec_29_left_subtree_state_2 = state_vec_29_right_subtree_state[1]; // @[package.scala 154:13]
  wire  state_vec_29_right_subtree_state_2 = state_vec_29_right_subtree_state[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_29_T_15 = state_vec_0_set_left_older_1 ? state_vec_29_left_subtree_state_2 : _state_vec_0_T_3; // @[Replacement.scala 203:16]
  wire  _state_vec_29_T_19 = state_vec_0_set_left_older_1 ? _state_vec_0_T_3 : state_vec_29_right_subtree_state_2; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_29_T_20 = {state_vec_0_set_left_older_1,_state_vec_29_T_15,_state_vec_29_T_19}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_29_T_21 = state_vec_0_set_left_older ? _state_vec_29_T_20 : state_vec_29_right_subtree_state; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_29_T_22 = {state_vec_0_set_left_older,_state_vec_29_T_10,_state_vec_29_T_21}; // @[Cat.scala 31:58]
  wire [6:0] _state_vec_29_T_23 = set_touch_ways_0_29_valid ? _state_vec_29_T_22 : state_vec__29; // @[Replacement.scala 22:56]
  wire [2:0] state_vec_29_left_subtree_state_3 = _state_vec_29_T_23[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_29_right_subtree_state_3 = _state_vec_29_T_23[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_29_left_subtree_state_4 = state_vec_29_left_subtree_state_3[1]; // @[package.scala 154:13]
  wire  state_vec_29_right_subtree_state_4 = state_vec_29_left_subtree_state_3[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_29_T_28 = state_vec_0_set_left_older_4 ? state_vec_29_left_subtree_state_4 : _state_vec_0_T_27; // @[Replacement.scala 203:16]
  wire  _state_vec_29_T_32 = state_vec_0_set_left_older_4 ? _state_vec_0_T_27 : state_vec_29_right_subtree_state_4; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_29_T_33 = {state_vec_0_set_left_older_4,_state_vec_29_T_28,_state_vec_29_T_32}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_29_T_34 = state_vec_0_set_left_older_3 ? state_vec_29_left_subtree_state_3 : _state_vec_29_T_33; // @[Replacement.scala 203:16]
  wire  state_vec_29_left_subtree_state_5 = state_vec_29_right_subtree_state_3[1]; // @[package.scala 154:13]
  wire  state_vec_29_right_subtree_state_5 = state_vec_29_right_subtree_state_3[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_29_T_39 = state_vec_0_set_left_older_4 ? state_vec_29_left_subtree_state_5 : _state_vec_0_T_27; // @[Replacement.scala 203:16]
  wire  _state_vec_29_T_43 = state_vec_0_set_left_older_4 ? _state_vec_0_T_27 : state_vec_29_right_subtree_state_5; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_29_T_44 = {state_vec_0_set_left_older_4,_state_vec_29_T_39,_state_vec_29_T_43}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_29_T_45 = state_vec_0_set_left_older_3 ? _state_vec_29_T_44 : state_vec_29_right_subtree_state_3
    ; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_29_T_46 = {state_vec_0_set_left_older_3,_state_vec_29_T_34,_state_vec_29_T_45}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_30_valid = touch_ways_0_0_valid & touch_sets_0_0 == 5'h1e; // @[Replacement.scala 315:30]
  wire  set_touch_ways_1_30_valid = touch_ways_0_1_valid & touch_sets_0_0 == 5'h1e; // @[Replacement.scala 315:30]
  wire  _T_109 = set_touch_ways_0_30_valid | set_touch_ways_1_30_valid; // @[package.scala 72:59]
  wire [2:0] state_vec_30_left_subtree_state = state_vec__30[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_30_right_subtree_state = state_vec__30[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_30_left_subtree_state_1 = state_vec_30_left_subtree_state[1]; // @[package.scala 154:13]
  wire  state_vec_30_right_subtree_state_1 = state_vec_30_left_subtree_state[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_30_T_4 = state_vec_0_set_left_older_1 ? state_vec_30_left_subtree_state_1 : _state_vec_0_T_3; // @[Replacement.scala 203:16]
  wire  _state_vec_30_T_8 = state_vec_0_set_left_older_1 ? _state_vec_0_T_3 : state_vec_30_right_subtree_state_1; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_30_T_9 = {state_vec_0_set_left_older_1,_state_vec_30_T_4,_state_vec_30_T_8}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_30_T_10 = state_vec_0_set_left_older ? state_vec_30_left_subtree_state : _state_vec_30_T_9; // @[Replacement.scala 203:16]
  wire  state_vec_30_left_subtree_state_2 = state_vec_30_right_subtree_state[1]; // @[package.scala 154:13]
  wire  state_vec_30_right_subtree_state_2 = state_vec_30_right_subtree_state[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_30_T_15 = state_vec_0_set_left_older_1 ? state_vec_30_left_subtree_state_2 : _state_vec_0_T_3; // @[Replacement.scala 203:16]
  wire  _state_vec_30_T_19 = state_vec_0_set_left_older_1 ? _state_vec_0_T_3 : state_vec_30_right_subtree_state_2; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_30_T_20 = {state_vec_0_set_left_older_1,_state_vec_30_T_15,_state_vec_30_T_19}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_30_T_21 = state_vec_0_set_left_older ? _state_vec_30_T_20 : state_vec_30_right_subtree_state; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_30_T_22 = {state_vec_0_set_left_older,_state_vec_30_T_10,_state_vec_30_T_21}; // @[Cat.scala 31:58]
  wire [6:0] _state_vec_30_T_23 = set_touch_ways_0_30_valid ? _state_vec_30_T_22 : state_vec__30; // @[Replacement.scala 22:56]
  wire [2:0] state_vec_30_left_subtree_state_3 = _state_vec_30_T_23[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_30_right_subtree_state_3 = _state_vec_30_T_23[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_30_left_subtree_state_4 = state_vec_30_left_subtree_state_3[1]; // @[package.scala 154:13]
  wire  state_vec_30_right_subtree_state_4 = state_vec_30_left_subtree_state_3[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_30_T_28 = state_vec_0_set_left_older_4 ? state_vec_30_left_subtree_state_4 : _state_vec_0_T_27; // @[Replacement.scala 203:16]
  wire  _state_vec_30_T_32 = state_vec_0_set_left_older_4 ? _state_vec_0_T_27 : state_vec_30_right_subtree_state_4; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_30_T_33 = {state_vec_0_set_left_older_4,_state_vec_30_T_28,_state_vec_30_T_32}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_30_T_34 = state_vec_0_set_left_older_3 ? state_vec_30_left_subtree_state_3 : _state_vec_30_T_33; // @[Replacement.scala 203:16]
  wire  state_vec_30_left_subtree_state_5 = state_vec_30_right_subtree_state_3[1]; // @[package.scala 154:13]
  wire  state_vec_30_right_subtree_state_5 = state_vec_30_right_subtree_state_3[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_30_T_39 = state_vec_0_set_left_older_4 ? state_vec_30_left_subtree_state_5 : _state_vec_0_T_27; // @[Replacement.scala 203:16]
  wire  _state_vec_30_T_43 = state_vec_0_set_left_older_4 ? _state_vec_0_T_27 : state_vec_30_right_subtree_state_5; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_30_T_44 = {state_vec_0_set_left_older_4,_state_vec_30_T_39,_state_vec_30_T_43}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_30_T_45 = state_vec_0_set_left_older_3 ? _state_vec_30_T_44 : state_vec_30_right_subtree_state_3
    ; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_30_T_46 = {state_vec_0_set_left_older_3,_state_vec_30_T_34,_state_vec_30_T_45}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_31_valid = touch_ways_0_0_valid & touch_sets_0_0 == 5'h1f; // @[Replacement.scala 315:30]
  wire  set_touch_ways_1_31_valid = touch_ways_0_1_valid & touch_sets_0_0 == 5'h1f; // @[Replacement.scala 315:30]
  wire  _T_110 = set_touch_ways_0_31_valid | set_touch_ways_1_31_valid; // @[package.scala 72:59]
  wire [2:0] state_vec_31_left_subtree_state = state_vec__31[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_31_right_subtree_state = state_vec__31[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_31_left_subtree_state_1 = state_vec_31_left_subtree_state[1]; // @[package.scala 154:13]
  wire  state_vec_31_right_subtree_state_1 = state_vec_31_left_subtree_state[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_31_T_4 = state_vec_0_set_left_older_1 ? state_vec_31_left_subtree_state_1 : _state_vec_0_T_3; // @[Replacement.scala 203:16]
  wire  _state_vec_31_T_8 = state_vec_0_set_left_older_1 ? _state_vec_0_T_3 : state_vec_31_right_subtree_state_1; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_31_T_9 = {state_vec_0_set_left_older_1,_state_vec_31_T_4,_state_vec_31_T_8}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_31_T_10 = state_vec_0_set_left_older ? state_vec_31_left_subtree_state : _state_vec_31_T_9; // @[Replacement.scala 203:16]
  wire  state_vec_31_left_subtree_state_2 = state_vec_31_right_subtree_state[1]; // @[package.scala 154:13]
  wire  state_vec_31_right_subtree_state_2 = state_vec_31_right_subtree_state[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_31_T_15 = state_vec_0_set_left_older_1 ? state_vec_31_left_subtree_state_2 : _state_vec_0_T_3; // @[Replacement.scala 203:16]
  wire  _state_vec_31_T_19 = state_vec_0_set_left_older_1 ? _state_vec_0_T_3 : state_vec_31_right_subtree_state_2; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_31_T_20 = {state_vec_0_set_left_older_1,_state_vec_31_T_15,_state_vec_31_T_19}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_31_T_21 = state_vec_0_set_left_older ? _state_vec_31_T_20 : state_vec_31_right_subtree_state; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_31_T_22 = {state_vec_0_set_left_older,_state_vec_31_T_10,_state_vec_31_T_21}; // @[Cat.scala 31:58]
  wire [6:0] _state_vec_31_T_23 = set_touch_ways_0_31_valid ? _state_vec_31_T_22 : state_vec__31; // @[Replacement.scala 22:56]
  wire [2:0] state_vec_31_left_subtree_state_3 = _state_vec_31_T_23[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_31_right_subtree_state_3 = _state_vec_31_T_23[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_31_left_subtree_state_4 = state_vec_31_left_subtree_state_3[1]; // @[package.scala 154:13]
  wire  state_vec_31_right_subtree_state_4 = state_vec_31_left_subtree_state_3[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_31_T_28 = state_vec_0_set_left_older_4 ? state_vec_31_left_subtree_state_4 : _state_vec_0_T_27; // @[Replacement.scala 203:16]
  wire  _state_vec_31_T_32 = state_vec_0_set_left_older_4 ? _state_vec_0_T_27 : state_vec_31_right_subtree_state_4; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_31_T_33 = {state_vec_0_set_left_older_4,_state_vec_31_T_28,_state_vec_31_T_32}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_31_T_34 = state_vec_0_set_left_older_3 ? state_vec_31_left_subtree_state_3 : _state_vec_31_T_33; // @[Replacement.scala 203:16]
  wire  state_vec_31_left_subtree_state_5 = state_vec_31_right_subtree_state_3[1]; // @[package.scala 154:13]
  wire  state_vec_31_right_subtree_state_5 = state_vec_31_right_subtree_state_3[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_31_T_39 = state_vec_0_set_left_older_4 ? state_vec_31_left_subtree_state_5 : _state_vec_0_T_27; // @[Replacement.scala 203:16]
  wire  _state_vec_31_T_43 = state_vec_0_set_left_older_4 ? _state_vec_0_T_27 : state_vec_31_right_subtree_state_5; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_31_T_44 = {state_vec_0_set_left_older_4,_state_vec_31_T_39,_state_vec_31_T_43}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_31_T_45 = state_vec_0_set_left_older_3 ? _state_vec_31_T_44 : state_vec_31_right_subtree_state_3
    ; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_31_T_46 = {state_vec_0_set_left_older_3,_state_vec_31_T_34,_state_vec_31_T_45}; // @[Cat.scala 31:58]
  reg [5:0] s2_req_vsetIdx_1; // @[Reg.scala 16:16]
  wire [4:0] touch_sets_1_0 = s2_req_vsetIdx_1[4:0]; // @[ICacheMainPipe.scala 136:36 671:20]
  wire  touch_ways_1_0_valid = s2_valid & s2_port_hit_1; // @[ICacheMainPipe.scala 672:32]
  wire  set_touch_ways_0_32_valid = touch_ways_1_0_valid & touch_sets_1_0 == 5'h0; // @[Replacement.scala 315:30]
  wire  touch_ways_1_1_valid = s2_valid & _miss_0_s2_1_T_4; // @[ICacheMainPipe.scala 676:32]
  wire  set_touch_ways_1_32_valid = touch_ways_1_1_valid & touch_sets_1_0 == 5'h0; // @[Replacement.scala 315:30]
  wire  _T_111 = set_touch_ways_0_32_valid | set_touch_ways_1_32_valid; // @[package.scala 72:59]
  reg  s2_tag_match_vec_1_7; // @[Reg.scala 16:16]
  reg  s2_tag_match_vec_1_6; // @[Reg.scala 16:16]
  reg  s2_tag_match_vec_1_5; // @[Reg.scala 16:16]
  reg  s2_tag_match_vec_1_4; // @[Reg.scala 16:16]
  reg  s2_tag_match_vec_1_3; // @[Reg.scala 16:16]
  reg  s2_tag_match_vec_1_2; // @[Reg.scala 16:16]
  reg  s2_tag_match_vec_1_1; // @[Reg.scala 16:16]
  reg  s2_tag_match_vec_1_0; // @[Reg.scala 16:16]
  wire [7:0] _touch_ways_1_0_bits_T = {s2_tag_match_vec_1_7,s2_tag_match_vec_1_6,s2_tag_match_vec_1_5,
    s2_tag_match_vec_1_4,s2_tag_match_vec_1_3,s2_tag_match_vec_1_2,s2_tag_match_vec_1_1,s2_tag_match_vec_1_0}; // @[OneHot.scala 22:45]
  wire [3:0] touch_ways_1_0_bits_hi_1 = _touch_ways_1_0_bits_T[7:4]; // @[OneHot.scala 30:18]
  wire  _touch_ways_1_0_bits_T_1 = |touch_ways_1_0_bits_hi_1; // @[OneHot.scala 32:14]
  wire [3:0] touch_ways_1_0_bits_lo_1 = _touch_ways_1_0_bits_T[3:0]; // @[OneHot.scala 31:18]
  wire [3:0] _touch_ways_1_0_bits_T_2 = touch_ways_1_0_bits_hi_1 | touch_ways_1_0_bits_lo_1; // @[OneHot.scala 32:28]
  wire [1:0] touch_ways_1_0_bits_hi_2 = _touch_ways_1_0_bits_T_2[3:2]; // @[OneHot.scala 30:18]
  wire  _touch_ways_1_0_bits_T_3 = |touch_ways_1_0_bits_hi_2; // @[OneHot.scala 32:14]
  wire [1:0] touch_ways_1_0_bits_lo_2 = _touch_ways_1_0_bits_T_2[1:0]; // @[OneHot.scala 31:18]
  wire [1:0] _touch_ways_1_0_bits_T_4 = touch_ways_1_0_bits_hi_2 | touch_ways_1_0_bits_lo_2; // @[OneHot.scala 32:28]
  wire [2:0] touch_ways_1_0_bits = {_touch_ways_1_0_bits_T_1,_touch_ways_1_0_bits_T_3,_touch_ways_1_0_bits_T_4[1]}; // @[Cat.scala 31:58]
  wire  state_vec_0_set_left_older_6 = ~touch_ways_1_0_bits[2]; // @[Replacement.scala 196:33]
  wire [2:0] state_vec_0_left_subtree_state_6 = state_vec_1_0[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_0_right_subtree_state_6 = state_vec_1_0[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_0_set_left_older_7 = ~touch_ways_1_0_bits[1]; // @[Replacement.scala 196:33]
  wire  state_vec_0_left_subtree_state_7 = state_vec_0_left_subtree_state_6[1]; // @[package.scala 154:13]
  wire  state_vec_0_right_subtree_state_7 = state_vec_0_left_subtree_state_6[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_0_T_51 = ~touch_ways_1_0_bits[0]; // @[Replacement.scala 218:7]
  wire  _state_vec_0_T_52 = state_vec_0_set_left_older_7 ? state_vec_0_left_subtree_state_7 : _state_vec_0_T_51; // @[Replacement.scala 203:16]
  wire  _state_vec_0_T_56 = state_vec_0_set_left_older_7 ? _state_vec_0_T_51 : state_vec_0_right_subtree_state_7; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_0_T_57 = {state_vec_0_set_left_older_7,_state_vec_0_T_52,_state_vec_0_T_56}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_0_T_58 = state_vec_0_set_left_older_6 ? state_vec_0_left_subtree_state_6 : _state_vec_0_T_57; // @[Replacement.scala 203:16]
  wire  state_vec_0_left_subtree_state_8 = state_vec_0_right_subtree_state_6[1]; // @[package.scala 154:13]
  wire  state_vec_0_right_subtree_state_8 = state_vec_0_right_subtree_state_6[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_0_T_63 = state_vec_0_set_left_older_7 ? state_vec_0_left_subtree_state_8 : _state_vec_0_T_51; // @[Replacement.scala 203:16]
  wire  _state_vec_0_T_67 = state_vec_0_set_left_older_7 ? _state_vec_0_T_51 : state_vec_0_right_subtree_state_8; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_0_T_68 = {state_vec_0_set_left_older_7,_state_vec_0_T_63,_state_vec_0_T_67}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_0_T_69 = state_vec_0_set_left_older_6 ? _state_vec_0_T_68 : state_vec_0_right_subtree_state_6; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_0_T_70 = {state_vec_0_set_left_older_6,_state_vec_0_T_58,_state_vec_0_T_69}; // @[Cat.scala 31:58]
  wire [6:0] _state_vec_0_T_71 = set_touch_ways_0_32_valid ? _state_vec_0_T_70 : state_vec_1_0; // @[Replacement.scala 22:56]
  reg [7:0] s2_waymask_1; // @[Reg.scala 16:16]
  wire [3:0] touch_ways_1_1_bits_hi = s2_waymask_1[7:4]; // @[OneHot.scala 30:18]
  wire  _touch_ways_1_1_bits_T = |touch_ways_1_1_bits_hi; // @[OneHot.scala 32:14]
  wire [3:0] touch_ways_1_1_bits_lo = s2_waymask_1[3:0]; // @[OneHot.scala 31:18]
  wire [3:0] _touch_ways_1_1_bits_T_1 = touch_ways_1_1_bits_hi | touch_ways_1_1_bits_lo; // @[OneHot.scala 32:28]
  wire [1:0] touch_ways_1_1_bits_hi_1 = _touch_ways_1_1_bits_T_1[3:2]; // @[OneHot.scala 30:18]
  wire  _touch_ways_1_1_bits_T_2 = |touch_ways_1_1_bits_hi_1; // @[OneHot.scala 32:14]
  wire [1:0] touch_ways_1_1_bits_lo_1 = _touch_ways_1_1_bits_T_1[1:0]; // @[OneHot.scala 31:18]
  wire [1:0] _touch_ways_1_1_bits_T_3 = touch_ways_1_1_bits_hi_1 | touch_ways_1_1_bits_lo_1; // @[OneHot.scala 32:28]
  wire [2:0] touch_ways_1_1_bits = {_touch_ways_1_1_bits_T,_touch_ways_1_1_bits_T_2,_touch_ways_1_1_bits_T_3[1]}; // @[Cat.scala 31:58]
  wire  state_vec_0_set_left_older_9 = ~touch_ways_1_1_bits[2]; // @[Replacement.scala 196:33]
  wire [2:0] state_vec_0_left_subtree_state_9 = _state_vec_0_T_71[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_0_right_subtree_state_9 = _state_vec_0_T_71[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_0_set_left_older_10 = ~touch_ways_1_1_bits[1]; // @[Replacement.scala 196:33]
  wire  state_vec_0_left_subtree_state_10 = state_vec_0_left_subtree_state_9[1]; // @[package.scala 154:13]
  wire  state_vec_0_right_subtree_state_10 = state_vec_0_left_subtree_state_9[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_0_T_75 = ~touch_ways_1_1_bits[0]; // @[Replacement.scala 218:7]
  wire  _state_vec_0_T_76 = state_vec_0_set_left_older_10 ? state_vec_0_left_subtree_state_10 : _state_vec_0_T_75; // @[Replacement.scala 203:16]
  wire  _state_vec_0_T_80 = state_vec_0_set_left_older_10 ? _state_vec_0_T_75 : state_vec_0_right_subtree_state_10; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_0_T_81 = {state_vec_0_set_left_older_10,_state_vec_0_T_76,_state_vec_0_T_80}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_0_T_82 = state_vec_0_set_left_older_9 ? state_vec_0_left_subtree_state_9 : _state_vec_0_T_81; // @[Replacement.scala 203:16]
  wire  state_vec_0_left_subtree_state_11 = state_vec_0_right_subtree_state_9[1]; // @[package.scala 154:13]
  wire  state_vec_0_right_subtree_state_11 = state_vec_0_right_subtree_state_9[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_0_T_87 = state_vec_0_set_left_older_10 ? state_vec_0_left_subtree_state_11 : _state_vec_0_T_75; // @[Replacement.scala 203:16]
  wire  _state_vec_0_T_91 = state_vec_0_set_left_older_10 ? _state_vec_0_T_75 : state_vec_0_right_subtree_state_11; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_0_T_92 = {state_vec_0_set_left_older_10,_state_vec_0_T_87,_state_vec_0_T_91}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_0_T_93 = state_vec_0_set_left_older_9 ? _state_vec_0_T_92 : state_vec_0_right_subtree_state_9; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_0_T_94 = {state_vec_0_set_left_older_9,_state_vec_0_T_82,_state_vec_0_T_93}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_33_valid = touch_ways_1_0_valid & touch_sets_1_0 == 5'h1; // @[Replacement.scala 315:30]
  wire  set_touch_ways_1_33_valid = touch_ways_1_1_valid & touch_sets_1_0 == 5'h1; // @[Replacement.scala 315:30]
  wire  _T_112 = set_touch_ways_0_33_valid | set_touch_ways_1_33_valid; // @[package.scala 72:59]
  wire [2:0] state_vec_1_left_subtree_state_6 = state_vec_1_1[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_1_right_subtree_state_6 = state_vec_1_1[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_1_left_subtree_state_7 = state_vec_1_left_subtree_state_6[1]; // @[package.scala 154:13]
  wire  state_vec_1_right_subtree_state_7 = state_vec_1_left_subtree_state_6[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_1_T_52 = state_vec_0_set_left_older_7 ? state_vec_1_left_subtree_state_7 : _state_vec_0_T_51; // @[Replacement.scala 203:16]
  wire  _state_vec_1_T_56 = state_vec_0_set_left_older_7 ? _state_vec_0_T_51 : state_vec_1_right_subtree_state_7; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_1_T_57 = {state_vec_0_set_left_older_7,_state_vec_1_T_52,_state_vec_1_T_56}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_1_T_58 = state_vec_0_set_left_older_6 ? state_vec_1_left_subtree_state_6 : _state_vec_1_T_57; // @[Replacement.scala 203:16]
  wire  state_vec_1_left_subtree_state_8 = state_vec_1_right_subtree_state_6[1]; // @[package.scala 154:13]
  wire  state_vec_1_right_subtree_state_8 = state_vec_1_right_subtree_state_6[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_1_T_63 = state_vec_0_set_left_older_7 ? state_vec_1_left_subtree_state_8 : _state_vec_0_T_51; // @[Replacement.scala 203:16]
  wire  _state_vec_1_T_67 = state_vec_0_set_left_older_7 ? _state_vec_0_T_51 : state_vec_1_right_subtree_state_8; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_1_T_68 = {state_vec_0_set_left_older_7,_state_vec_1_T_63,_state_vec_1_T_67}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_1_T_69 = state_vec_0_set_left_older_6 ? _state_vec_1_T_68 : state_vec_1_right_subtree_state_6; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_1_T_70 = {state_vec_0_set_left_older_6,_state_vec_1_T_58,_state_vec_1_T_69}; // @[Cat.scala 31:58]
  wire [6:0] _state_vec_1_T_71 = set_touch_ways_0_33_valid ? _state_vec_1_T_70 : state_vec_1_1; // @[Replacement.scala 22:56]
  wire [2:0] state_vec_1_left_subtree_state_9 = _state_vec_1_T_71[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_1_right_subtree_state_9 = _state_vec_1_T_71[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_1_left_subtree_state_10 = state_vec_1_left_subtree_state_9[1]; // @[package.scala 154:13]
  wire  state_vec_1_right_subtree_state_10 = state_vec_1_left_subtree_state_9[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_1_T_76 = state_vec_0_set_left_older_10 ? state_vec_1_left_subtree_state_10 : _state_vec_0_T_75; // @[Replacement.scala 203:16]
  wire  _state_vec_1_T_80 = state_vec_0_set_left_older_10 ? _state_vec_0_T_75 : state_vec_1_right_subtree_state_10; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_1_T_81 = {state_vec_0_set_left_older_10,_state_vec_1_T_76,_state_vec_1_T_80}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_1_T_82 = state_vec_0_set_left_older_9 ? state_vec_1_left_subtree_state_9 : _state_vec_1_T_81; // @[Replacement.scala 203:16]
  wire  state_vec_1_left_subtree_state_11 = state_vec_1_right_subtree_state_9[1]; // @[package.scala 154:13]
  wire  state_vec_1_right_subtree_state_11 = state_vec_1_right_subtree_state_9[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_1_T_87 = state_vec_0_set_left_older_10 ? state_vec_1_left_subtree_state_11 : _state_vec_0_T_75; // @[Replacement.scala 203:16]
  wire  _state_vec_1_T_91 = state_vec_0_set_left_older_10 ? _state_vec_0_T_75 : state_vec_1_right_subtree_state_11; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_1_T_92 = {state_vec_0_set_left_older_10,_state_vec_1_T_87,_state_vec_1_T_91}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_1_T_93 = state_vec_0_set_left_older_9 ? _state_vec_1_T_92 : state_vec_1_right_subtree_state_9; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_1_T_94 = {state_vec_0_set_left_older_9,_state_vec_1_T_82,_state_vec_1_T_93}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_34_valid = touch_ways_1_0_valid & touch_sets_1_0 == 5'h2; // @[Replacement.scala 315:30]
  wire  set_touch_ways_1_34_valid = touch_ways_1_1_valid & touch_sets_1_0 == 5'h2; // @[Replacement.scala 315:30]
  wire  _T_113 = set_touch_ways_0_34_valid | set_touch_ways_1_34_valid; // @[package.scala 72:59]
  wire [2:0] state_vec_2_left_subtree_state_6 = state_vec_1_2[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_2_right_subtree_state_6 = state_vec_1_2[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_2_left_subtree_state_7 = state_vec_2_left_subtree_state_6[1]; // @[package.scala 154:13]
  wire  state_vec_2_right_subtree_state_7 = state_vec_2_left_subtree_state_6[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_2_T_52 = state_vec_0_set_left_older_7 ? state_vec_2_left_subtree_state_7 : _state_vec_0_T_51; // @[Replacement.scala 203:16]
  wire  _state_vec_2_T_56 = state_vec_0_set_left_older_7 ? _state_vec_0_T_51 : state_vec_2_right_subtree_state_7; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_2_T_57 = {state_vec_0_set_left_older_7,_state_vec_2_T_52,_state_vec_2_T_56}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_2_T_58 = state_vec_0_set_left_older_6 ? state_vec_2_left_subtree_state_6 : _state_vec_2_T_57; // @[Replacement.scala 203:16]
  wire  state_vec_2_left_subtree_state_8 = state_vec_2_right_subtree_state_6[1]; // @[package.scala 154:13]
  wire  state_vec_2_right_subtree_state_8 = state_vec_2_right_subtree_state_6[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_2_T_63 = state_vec_0_set_left_older_7 ? state_vec_2_left_subtree_state_8 : _state_vec_0_T_51; // @[Replacement.scala 203:16]
  wire  _state_vec_2_T_67 = state_vec_0_set_left_older_7 ? _state_vec_0_T_51 : state_vec_2_right_subtree_state_8; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_2_T_68 = {state_vec_0_set_left_older_7,_state_vec_2_T_63,_state_vec_2_T_67}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_2_T_69 = state_vec_0_set_left_older_6 ? _state_vec_2_T_68 : state_vec_2_right_subtree_state_6; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_2_T_70 = {state_vec_0_set_left_older_6,_state_vec_2_T_58,_state_vec_2_T_69}; // @[Cat.scala 31:58]
  wire [6:0] _state_vec_2_T_71 = set_touch_ways_0_34_valid ? _state_vec_2_T_70 : state_vec_1_2; // @[Replacement.scala 22:56]
  wire [2:0] state_vec_2_left_subtree_state_9 = _state_vec_2_T_71[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_2_right_subtree_state_9 = _state_vec_2_T_71[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_2_left_subtree_state_10 = state_vec_2_left_subtree_state_9[1]; // @[package.scala 154:13]
  wire  state_vec_2_right_subtree_state_10 = state_vec_2_left_subtree_state_9[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_2_T_76 = state_vec_0_set_left_older_10 ? state_vec_2_left_subtree_state_10 : _state_vec_0_T_75; // @[Replacement.scala 203:16]
  wire  _state_vec_2_T_80 = state_vec_0_set_left_older_10 ? _state_vec_0_T_75 : state_vec_2_right_subtree_state_10; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_2_T_81 = {state_vec_0_set_left_older_10,_state_vec_2_T_76,_state_vec_2_T_80}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_2_T_82 = state_vec_0_set_left_older_9 ? state_vec_2_left_subtree_state_9 : _state_vec_2_T_81; // @[Replacement.scala 203:16]
  wire  state_vec_2_left_subtree_state_11 = state_vec_2_right_subtree_state_9[1]; // @[package.scala 154:13]
  wire  state_vec_2_right_subtree_state_11 = state_vec_2_right_subtree_state_9[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_2_T_87 = state_vec_0_set_left_older_10 ? state_vec_2_left_subtree_state_11 : _state_vec_0_T_75; // @[Replacement.scala 203:16]
  wire  _state_vec_2_T_91 = state_vec_0_set_left_older_10 ? _state_vec_0_T_75 : state_vec_2_right_subtree_state_11; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_2_T_92 = {state_vec_0_set_left_older_10,_state_vec_2_T_87,_state_vec_2_T_91}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_2_T_93 = state_vec_0_set_left_older_9 ? _state_vec_2_T_92 : state_vec_2_right_subtree_state_9; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_2_T_94 = {state_vec_0_set_left_older_9,_state_vec_2_T_82,_state_vec_2_T_93}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_35_valid = touch_ways_1_0_valid & touch_sets_1_0 == 5'h3; // @[Replacement.scala 315:30]
  wire  set_touch_ways_1_35_valid = touch_ways_1_1_valid & touch_sets_1_0 == 5'h3; // @[Replacement.scala 315:30]
  wire  _T_114 = set_touch_ways_0_35_valid | set_touch_ways_1_35_valid; // @[package.scala 72:59]
  wire [2:0] state_vec_3_left_subtree_state_6 = state_vec_1_3[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_3_right_subtree_state_6 = state_vec_1_3[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_3_left_subtree_state_7 = state_vec_3_left_subtree_state_6[1]; // @[package.scala 154:13]
  wire  state_vec_3_right_subtree_state_7 = state_vec_3_left_subtree_state_6[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_3_T_52 = state_vec_0_set_left_older_7 ? state_vec_3_left_subtree_state_7 : _state_vec_0_T_51; // @[Replacement.scala 203:16]
  wire  _state_vec_3_T_56 = state_vec_0_set_left_older_7 ? _state_vec_0_T_51 : state_vec_3_right_subtree_state_7; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_3_T_57 = {state_vec_0_set_left_older_7,_state_vec_3_T_52,_state_vec_3_T_56}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_3_T_58 = state_vec_0_set_left_older_6 ? state_vec_3_left_subtree_state_6 : _state_vec_3_T_57; // @[Replacement.scala 203:16]
  wire  state_vec_3_left_subtree_state_8 = state_vec_3_right_subtree_state_6[1]; // @[package.scala 154:13]
  wire  state_vec_3_right_subtree_state_8 = state_vec_3_right_subtree_state_6[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_3_T_63 = state_vec_0_set_left_older_7 ? state_vec_3_left_subtree_state_8 : _state_vec_0_T_51; // @[Replacement.scala 203:16]
  wire  _state_vec_3_T_67 = state_vec_0_set_left_older_7 ? _state_vec_0_T_51 : state_vec_3_right_subtree_state_8; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_3_T_68 = {state_vec_0_set_left_older_7,_state_vec_3_T_63,_state_vec_3_T_67}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_3_T_69 = state_vec_0_set_left_older_6 ? _state_vec_3_T_68 : state_vec_3_right_subtree_state_6; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_3_T_70 = {state_vec_0_set_left_older_6,_state_vec_3_T_58,_state_vec_3_T_69}; // @[Cat.scala 31:58]
  wire [6:0] _state_vec_3_T_71 = set_touch_ways_0_35_valid ? _state_vec_3_T_70 : state_vec_1_3; // @[Replacement.scala 22:56]
  wire [2:0] state_vec_3_left_subtree_state_9 = _state_vec_3_T_71[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_3_right_subtree_state_9 = _state_vec_3_T_71[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_3_left_subtree_state_10 = state_vec_3_left_subtree_state_9[1]; // @[package.scala 154:13]
  wire  state_vec_3_right_subtree_state_10 = state_vec_3_left_subtree_state_9[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_3_T_76 = state_vec_0_set_left_older_10 ? state_vec_3_left_subtree_state_10 : _state_vec_0_T_75; // @[Replacement.scala 203:16]
  wire  _state_vec_3_T_80 = state_vec_0_set_left_older_10 ? _state_vec_0_T_75 : state_vec_3_right_subtree_state_10; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_3_T_81 = {state_vec_0_set_left_older_10,_state_vec_3_T_76,_state_vec_3_T_80}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_3_T_82 = state_vec_0_set_left_older_9 ? state_vec_3_left_subtree_state_9 : _state_vec_3_T_81; // @[Replacement.scala 203:16]
  wire  state_vec_3_left_subtree_state_11 = state_vec_3_right_subtree_state_9[1]; // @[package.scala 154:13]
  wire  state_vec_3_right_subtree_state_11 = state_vec_3_right_subtree_state_9[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_3_T_87 = state_vec_0_set_left_older_10 ? state_vec_3_left_subtree_state_11 : _state_vec_0_T_75; // @[Replacement.scala 203:16]
  wire  _state_vec_3_T_91 = state_vec_0_set_left_older_10 ? _state_vec_0_T_75 : state_vec_3_right_subtree_state_11; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_3_T_92 = {state_vec_0_set_left_older_10,_state_vec_3_T_87,_state_vec_3_T_91}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_3_T_93 = state_vec_0_set_left_older_9 ? _state_vec_3_T_92 : state_vec_3_right_subtree_state_9; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_3_T_94 = {state_vec_0_set_left_older_9,_state_vec_3_T_82,_state_vec_3_T_93}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_36_valid = touch_ways_1_0_valid & touch_sets_1_0 == 5'h4; // @[Replacement.scala 315:30]
  wire  set_touch_ways_1_36_valid = touch_ways_1_1_valid & touch_sets_1_0 == 5'h4; // @[Replacement.scala 315:30]
  wire  _T_115 = set_touch_ways_0_36_valid | set_touch_ways_1_36_valid; // @[package.scala 72:59]
  wire [2:0] state_vec_4_left_subtree_state_6 = state_vec_1_4[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_4_right_subtree_state_6 = state_vec_1_4[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_4_left_subtree_state_7 = state_vec_4_left_subtree_state_6[1]; // @[package.scala 154:13]
  wire  state_vec_4_right_subtree_state_7 = state_vec_4_left_subtree_state_6[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_4_T_52 = state_vec_0_set_left_older_7 ? state_vec_4_left_subtree_state_7 : _state_vec_0_T_51; // @[Replacement.scala 203:16]
  wire  _state_vec_4_T_56 = state_vec_0_set_left_older_7 ? _state_vec_0_T_51 : state_vec_4_right_subtree_state_7; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_4_T_57 = {state_vec_0_set_left_older_7,_state_vec_4_T_52,_state_vec_4_T_56}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_4_T_58 = state_vec_0_set_left_older_6 ? state_vec_4_left_subtree_state_6 : _state_vec_4_T_57; // @[Replacement.scala 203:16]
  wire  state_vec_4_left_subtree_state_8 = state_vec_4_right_subtree_state_6[1]; // @[package.scala 154:13]
  wire  state_vec_4_right_subtree_state_8 = state_vec_4_right_subtree_state_6[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_4_T_63 = state_vec_0_set_left_older_7 ? state_vec_4_left_subtree_state_8 : _state_vec_0_T_51; // @[Replacement.scala 203:16]
  wire  _state_vec_4_T_67 = state_vec_0_set_left_older_7 ? _state_vec_0_T_51 : state_vec_4_right_subtree_state_8; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_4_T_68 = {state_vec_0_set_left_older_7,_state_vec_4_T_63,_state_vec_4_T_67}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_4_T_69 = state_vec_0_set_left_older_6 ? _state_vec_4_T_68 : state_vec_4_right_subtree_state_6; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_4_T_70 = {state_vec_0_set_left_older_6,_state_vec_4_T_58,_state_vec_4_T_69}; // @[Cat.scala 31:58]
  wire [6:0] _state_vec_4_T_71 = set_touch_ways_0_36_valid ? _state_vec_4_T_70 : state_vec_1_4; // @[Replacement.scala 22:56]
  wire [2:0] state_vec_4_left_subtree_state_9 = _state_vec_4_T_71[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_4_right_subtree_state_9 = _state_vec_4_T_71[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_4_left_subtree_state_10 = state_vec_4_left_subtree_state_9[1]; // @[package.scala 154:13]
  wire  state_vec_4_right_subtree_state_10 = state_vec_4_left_subtree_state_9[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_4_T_76 = state_vec_0_set_left_older_10 ? state_vec_4_left_subtree_state_10 : _state_vec_0_T_75; // @[Replacement.scala 203:16]
  wire  _state_vec_4_T_80 = state_vec_0_set_left_older_10 ? _state_vec_0_T_75 : state_vec_4_right_subtree_state_10; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_4_T_81 = {state_vec_0_set_left_older_10,_state_vec_4_T_76,_state_vec_4_T_80}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_4_T_82 = state_vec_0_set_left_older_9 ? state_vec_4_left_subtree_state_9 : _state_vec_4_T_81; // @[Replacement.scala 203:16]
  wire  state_vec_4_left_subtree_state_11 = state_vec_4_right_subtree_state_9[1]; // @[package.scala 154:13]
  wire  state_vec_4_right_subtree_state_11 = state_vec_4_right_subtree_state_9[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_4_T_87 = state_vec_0_set_left_older_10 ? state_vec_4_left_subtree_state_11 : _state_vec_0_T_75; // @[Replacement.scala 203:16]
  wire  _state_vec_4_T_91 = state_vec_0_set_left_older_10 ? _state_vec_0_T_75 : state_vec_4_right_subtree_state_11; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_4_T_92 = {state_vec_0_set_left_older_10,_state_vec_4_T_87,_state_vec_4_T_91}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_4_T_93 = state_vec_0_set_left_older_9 ? _state_vec_4_T_92 : state_vec_4_right_subtree_state_9; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_4_T_94 = {state_vec_0_set_left_older_9,_state_vec_4_T_82,_state_vec_4_T_93}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_37_valid = touch_ways_1_0_valid & touch_sets_1_0 == 5'h5; // @[Replacement.scala 315:30]
  wire  set_touch_ways_1_37_valid = touch_ways_1_1_valid & touch_sets_1_0 == 5'h5; // @[Replacement.scala 315:30]
  wire  _T_116 = set_touch_ways_0_37_valid | set_touch_ways_1_37_valid; // @[package.scala 72:59]
  wire [2:0] state_vec_5_left_subtree_state_6 = state_vec_1_5[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_5_right_subtree_state_6 = state_vec_1_5[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_5_left_subtree_state_7 = state_vec_5_left_subtree_state_6[1]; // @[package.scala 154:13]
  wire  state_vec_5_right_subtree_state_7 = state_vec_5_left_subtree_state_6[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_5_T_52 = state_vec_0_set_left_older_7 ? state_vec_5_left_subtree_state_7 : _state_vec_0_T_51; // @[Replacement.scala 203:16]
  wire  _state_vec_5_T_56 = state_vec_0_set_left_older_7 ? _state_vec_0_T_51 : state_vec_5_right_subtree_state_7; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_5_T_57 = {state_vec_0_set_left_older_7,_state_vec_5_T_52,_state_vec_5_T_56}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_5_T_58 = state_vec_0_set_left_older_6 ? state_vec_5_left_subtree_state_6 : _state_vec_5_T_57; // @[Replacement.scala 203:16]
  wire  state_vec_5_left_subtree_state_8 = state_vec_5_right_subtree_state_6[1]; // @[package.scala 154:13]
  wire  state_vec_5_right_subtree_state_8 = state_vec_5_right_subtree_state_6[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_5_T_63 = state_vec_0_set_left_older_7 ? state_vec_5_left_subtree_state_8 : _state_vec_0_T_51; // @[Replacement.scala 203:16]
  wire  _state_vec_5_T_67 = state_vec_0_set_left_older_7 ? _state_vec_0_T_51 : state_vec_5_right_subtree_state_8; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_5_T_68 = {state_vec_0_set_left_older_7,_state_vec_5_T_63,_state_vec_5_T_67}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_5_T_69 = state_vec_0_set_left_older_6 ? _state_vec_5_T_68 : state_vec_5_right_subtree_state_6; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_5_T_70 = {state_vec_0_set_left_older_6,_state_vec_5_T_58,_state_vec_5_T_69}; // @[Cat.scala 31:58]
  wire [6:0] _state_vec_5_T_71 = set_touch_ways_0_37_valid ? _state_vec_5_T_70 : state_vec_1_5; // @[Replacement.scala 22:56]
  wire [2:0] state_vec_5_left_subtree_state_9 = _state_vec_5_T_71[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_5_right_subtree_state_9 = _state_vec_5_T_71[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_5_left_subtree_state_10 = state_vec_5_left_subtree_state_9[1]; // @[package.scala 154:13]
  wire  state_vec_5_right_subtree_state_10 = state_vec_5_left_subtree_state_9[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_5_T_76 = state_vec_0_set_left_older_10 ? state_vec_5_left_subtree_state_10 : _state_vec_0_T_75; // @[Replacement.scala 203:16]
  wire  _state_vec_5_T_80 = state_vec_0_set_left_older_10 ? _state_vec_0_T_75 : state_vec_5_right_subtree_state_10; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_5_T_81 = {state_vec_0_set_left_older_10,_state_vec_5_T_76,_state_vec_5_T_80}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_5_T_82 = state_vec_0_set_left_older_9 ? state_vec_5_left_subtree_state_9 : _state_vec_5_T_81; // @[Replacement.scala 203:16]
  wire  state_vec_5_left_subtree_state_11 = state_vec_5_right_subtree_state_9[1]; // @[package.scala 154:13]
  wire  state_vec_5_right_subtree_state_11 = state_vec_5_right_subtree_state_9[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_5_T_87 = state_vec_0_set_left_older_10 ? state_vec_5_left_subtree_state_11 : _state_vec_0_T_75; // @[Replacement.scala 203:16]
  wire  _state_vec_5_T_91 = state_vec_0_set_left_older_10 ? _state_vec_0_T_75 : state_vec_5_right_subtree_state_11; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_5_T_92 = {state_vec_0_set_left_older_10,_state_vec_5_T_87,_state_vec_5_T_91}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_5_T_93 = state_vec_0_set_left_older_9 ? _state_vec_5_T_92 : state_vec_5_right_subtree_state_9; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_5_T_94 = {state_vec_0_set_left_older_9,_state_vec_5_T_82,_state_vec_5_T_93}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_38_valid = touch_ways_1_0_valid & touch_sets_1_0 == 5'h6; // @[Replacement.scala 315:30]
  wire  set_touch_ways_1_38_valid = touch_ways_1_1_valid & touch_sets_1_0 == 5'h6; // @[Replacement.scala 315:30]
  wire  _T_117 = set_touch_ways_0_38_valid | set_touch_ways_1_38_valid; // @[package.scala 72:59]
  wire [2:0] state_vec_6_left_subtree_state_6 = state_vec_1_6[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_6_right_subtree_state_6 = state_vec_1_6[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_6_left_subtree_state_7 = state_vec_6_left_subtree_state_6[1]; // @[package.scala 154:13]
  wire  state_vec_6_right_subtree_state_7 = state_vec_6_left_subtree_state_6[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_6_T_52 = state_vec_0_set_left_older_7 ? state_vec_6_left_subtree_state_7 : _state_vec_0_T_51; // @[Replacement.scala 203:16]
  wire  _state_vec_6_T_56 = state_vec_0_set_left_older_7 ? _state_vec_0_T_51 : state_vec_6_right_subtree_state_7; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_6_T_57 = {state_vec_0_set_left_older_7,_state_vec_6_T_52,_state_vec_6_T_56}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_6_T_58 = state_vec_0_set_left_older_6 ? state_vec_6_left_subtree_state_6 : _state_vec_6_T_57; // @[Replacement.scala 203:16]
  wire  state_vec_6_left_subtree_state_8 = state_vec_6_right_subtree_state_6[1]; // @[package.scala 154:13]
  wire  state_vec_6_right_subtree_state_8 = state_vec_6_right_subtree_state_6[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_6_T_63 = state_vec_0_set_left_older_7 ? state_vec_6_left_subtree_state_8 : _state_vec_0_T_51; // @[Replacement.scala 203:16]
  wire  _state_vec_6_T_67 = state_vec_0_set_left_older_7 ? _state_vec_0_T_51 : state_vec_6_right_subtree_state_8; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_6_T_68 = {state_vec_0_set_left_older_7,_state_vec_6_T_63,_state_vec_6_T_67}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_6_T_69 = state_vec_0_set_left_older_6 ? _state_vec_6_T_68 : state_vec_6_right_subtree_state_6; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_6_T_70 = {state_vec_0_set_left_older_6,_state_vec_6_T_58,_state_vec_6_T_69}; // @[Cat.scala 31:58]
  wire [6:0] _state_vec_6_T_71 = set_touch_ways_0_38_valid ? _state_vec_6_T_70 : state_vec_1_6; // @[Replacement.scala 22:56]
  wire [2:0] state_vec_6_left_subtree_state_9 = _state_vec_6_T_71[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_6_right_subtree_state_9 = _state_vec_6_T_71[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_6_left_subtree_state_10 = state_vec_6_left_subtree_state_9[1]; // @[package.scala 154:13]
  wire  state_vec_6_right_subtree_state_10 = state_vec_6_left_subtree_state_9[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_6_T_76 = state_vec_0_set_left_older_10 ? state_vec_6_left_subtree_state_10 : _state_vec_0_T_75; // @[Replacement.scala 203:16]
  wire  _state_vec_6_T_80 = state_vec_0_set_left_older_10 ? _state_vec_0_T_75 : state_vec_6_right_subtree_state_10; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_6_T_81 = {state_vec_0_set_left_older_10,_state_vec_6_T_76,_state_vec_6_T_80}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_6_T_82 = state_vec_0_set_left_older_9 ? state_vec_6_left_subtree_state_9 : _state_vec_6_T_81; // @[Replacement.scala 203:16]
  wire  state_vec_6_left_subtree_state_11 = state_vec_6_right_subtree_state_9[1]; // @[package.scala 154:13]
  wire  state_vec_6_right_subtree_state_11 = state_vec_6_right_subtree_state_9[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_6_T_87 = state_vec_0_set_left_older_10 ? state_vec_6_left_subtree_state_11 : _state_vec_0_T_75; // @[Replacement.scala 203:16]
  wire  _state_vec_6_T_91 = state_vec_0_set_left_older_10 ? _state_vec_0_T_75 : state_vec_6_right_subtree_state_11; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_6_T_92 = {state_vec_0_set_left_older_10,_state_vec_6_T_87,_state_vec_6_T_91}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_6_T_93 = state_vec_0_set_left_older_9 ? _state_vec_6_T_92 : state_vec_6_right_subtree_state_9; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_6_T_94 = {state_vec_0_set_left_older_9,_state_vec_6_T_82,_state_vec_6_T_93}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_39_valid = touch_ways_1_0_valid & touch_sets_1_0 == 5'h7; // @[Replacement.scala 315:30]
  wire  set_touch_ways_1_39_valid = touch_ways_1_1_valid & touch_sets_1_0 == 5'h7; // @[Replacement.scala 315:30]
  wire  _T_118 = set_touch_ways_0_39_valid | set_touch_ways_1_39_valid; // @[package.scala 72:59]
  wire [2:0] state_vec_7_left_subtree_state_6 = state_vec_1_7[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_7_right_subtree_state_6 = state_vec_1_7[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_7_left_subtree_state_7 = state_vec_7_left_subtree_state_6[1]; // @[package.scala 154:13]
  wire  state_vec_7_right_subtree_state_7 = state_vec_7_left_subtree_state_6[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_7_T_52 = state_vec_0_set_left_older_7 ? state_vec_7_left_subtree_state_7 : _state_vec_0_T_51; // @[Replacement.scala 203:16]
  wire  _state_vec_7_T_56 = state_vec_0_set_left_older_7 ? _state_vec_0_T_51 : state_vec_7_right_subtree_state_7; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_7_T_57 = {state_vec_0_set_left_older_7,_state_vec_7_T_52,_state_vec_7_T_56}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_7_T_58 = state_vec_0_set_left_older_6 ? state_vec_7_left_subtree_state_6 : _state_vec_7_T_57; // @[Replacement.scala 203:16]
  wire  state_vec_7_left_subtree_state_8 = state_vec_7_right_subtree_state_6[1]; // @[package.scala 154:13]
  wire  state_vec_7_right_subtree_state_8 = state_vec_7_right_subtree_state_6[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_7_T_63 = state_vec_0_set_left_older_7 ? state_vec_7_left_subtree_state_8 : _state_vec_0_T_51; // @[Replacement.scala 203:16]
  wire  _state_vec_7_T_67 = state_vec_0_set_left_older_7 ? _state_vec_0_T_51 : state_vec_7_right_subtree_state_8; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_7_T_68 = {state_vec_0_set_left_older_7,_state_vec_7_T_63,_state_vec_7_T_67}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_7_T_69 = state_vec_0_set_left_older_6 ? _state_vec_7_T_68 : state_vec_7_right_subtree_state_6; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_7_T_70 = {state_vec_0_set_left_older_6,_state_vec_7_T_58,_state_vec_7_T_69}; // @[Cat.scala 31:58]
  wire [6:0] _state_vec_7_T_71 = set_touch_ways_0_39_valid ? _state_vec_7_T_70 : state_vec_1_7; // @[Replacement.scala 22:56]
  wire [2:0] state_vec_7_left_subtree_state_9 = _state_vec_7_T_71[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_7_right_subtree_state_9 = _state_vec_7_T_71[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_7_left_subtree_state_10 = state_vec_7_left_subtree_state_9[1]; // @[package.scala 154:13]
  wire  state_vec_7_right_subtree_state_10 = state_vec_7_left_subtree_state_9[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_7_T_76 = state_vec_0_set_left_older_10 ? state_vec_7_left_subtree_state_10 : _state_vec_0_T_75; // @[Replacement.scala 203:16]
  wire  _state_vec_7_T_80 = state_vec_0_set_left_older_10 ? _state_vec_0_T_75 : state_vec_7_right_subtree_state_10; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_7_T_81 = {state_vec_0_set_left_older_10,_state_vec_7_T_76,_state_vec_7_T_80}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_7_T_82 = state_vec_0_set_left_older_9 ? state_vec_7_left_subtree_state_9 : _state_vec_7_T_81; // @[Replacement.scala 203:16]
  wire  state_vec_7_left_subtree_state_11 = state_vec_7_right_subtree_state_9[1]; // @[package.scala 154:13]
  wire  state_vec_7_right_subtree_state_11 = state_vec_7_right_subtree_state_9[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_7_T_87 = state_vec_0_set_left_older_10 ? state_vec_7_left_subtree_state_11 : _state_vec_0_T_75; // @[Replacement.scala 203:16]
  wire  _state_vec_7_T_91 = state_vec_0_set_left_older_10 ? _state_vec_0_T_75 : state_vec_7_right_subtree_state_11; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_7_T_92 = {state_vec_0_set_left_older_10,_state_vec_7_T_87,_state_vec_7_T_91}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_7_T_93 = state_vec_0_set_left_older_9 ? _state_vec_7_T_92 : state_vec_7_right_subtree_state_9; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_7_T_94 = {state_vec_0_set_left_older_9,_state_vec_7_T_82,_state_vec_7_T_93}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_40_valid = touch_ways_1_0_valid & touch_sets_1_0 == 5'h8; // @[Replacement.scala 315:30]
  wire  set_touch_ways_1_40_valid = touch_ways_1_1_valid & touch_sets_1_0 == 5'h8; // @[Replacement.scala 315:30]
  wire  _T_119 = set_touch_ways_0_40_valid | set_touch_ways_1_40_valid; // @[package.scala 72:59]
  wire [2:0] state_vec_8_left_subtree_state_6 = state_vec_1_8[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_8_right_subtree_state_6 = state_vec_1_8[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_8_left_subtree_state_7 = state_vec_8_left_subtree_state_6[1]; // @[package.scala 154:13]
  wire  state_vec_8_right_subtree_state_7 = state_vec_8_left_subtree_state_6[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_8_T_52 = state_vec_0_set_left_older_7 ? state_vec_8_left_subtree_state_7 : _state_vec_0_T_51; // @[Replacement.scala 203:16]
  wire  _state_vec_8_T_56 = state_vec_0_set_left_older_7 ? _state_vec_0_T_51 : state_vec_8_right_subtree_state_7; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_8_T_57 = {state_vec_0_set_left_older_7,_state_vec_8_T_52,_state_vec_8_T_56}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_8_T_58 = state_vec_0_set_left_older_6 ? state_vec_8_left_subtree_state_6 : _state_vec_8_T_57; // @[Replacement.scala 203:16]
  wire  state_vec_8_left_subtree_state_8 = state_vec_8_right_subtree_state_6[1]; // @[package.scala 154:13]
  wire  state_vec_8_right_subtree_state_8 = state_vec_8_right_subtree_state_6[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_8_T_63 = state_vec_0_set_left_older_7 ? state_vec_8_left_subtree_state_8 : _state_vec_0_T_51; // @[Replacement.scala 203:16]
  wire  _state_vec_8_T_67 = state_vec_0_set_left_older_7 ? _state_vec_0_T_51 : state_vec_8_right_subtree_state_8; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_8_T_68 = {state_vec_0_set_left_older_7,_state_vec_8_T_63,_state_vec_8_T_67}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_8_T_69 = state_vec_0_set_left_older_6 ? _state_vec_8_T_68 : state_vec_8_right_subtree_state_6; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_8_T_70 = {state_vec_0_set_left_older_6,_state_vec_8_T_58,_state_vec_8_T_69}; // @[Cat.scala 31:58]
  wire [6:0] _state_vec_8_T_71 = set_touch_ways_0_40_valid ? _state_vec_8_T_70 : state_vec_1_8; // @[Replacement.scala 22:56]
  wire [2:0] state_vec_8_left_subtree_state_9 = _state_vec_8_T_71[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_8_right_subtree_state_9 = _state_vec_8_T_71[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_8_left_subtree_state_10 = state_vec_8_left_subtree_state_9[1]; // @[package.scala 154:13]
  wire  state_vec_8_right_subtree_state_10 = state_vec_8_left_subtree_state_9[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_8_T_76 = state_vec_0_set_left_older_10 ? state_vec_8_left_subtree_state_10 : _state_vec_0_T_75; // @[Replacement.scala 203:16]
  wire  _state_vec_8_T_80 = state_vec_0_set_left_older_10 ? _state_vec_0_T_75 : state_vec_8_right_subtree_state_10; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_8_T_81 = {state_vec_0_set_left_older_10,_state_vec_8_T_76,_state_vec_8_T_80}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_8_T_82 = state_vec_0_set_left_older_9 ? state_vec_8_left_subtree_state_9 : _state_vec_8_T_81; // @[Replacement.scala 203:16]
  wire  state_vec_8_left_subtree_state_11 = state_vec_8_right_subtree_state_9[1]; // @[package.scala 154:13]
  wire  state_vec_8_right_subtree_state_11 = state_vec_8_right_subtree_state_9[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_8_T_87 = state_vec_0_set_left_older_10 ? state_vec_8_left_subtree_state_11 : _state_vec_0_T_75; // @[Replacement.scala 203:16]
  wire  _state_vec_8_T_91 = state_vec_0_set_left_older_10 ? _state_vec_0_T_75 : state_vec_8_right_subtree_state_11; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_8_T_92 = {state_vec_0_set_left_older_10,_state_vec_8_T_87,_state_vec_8_T_91}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_8_T_93 = state_vec_0_set_left_older_9 ? _state_vec_8_T_92 : state_vec_8_right_subtree_state_9; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_8_T_94 = {state_vec_0_set_left_older_9,_state_vec_8_T_82,_state_vec_8_T_93}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_41_valid = touch_ways_1_0_valid & touch_sets_1_0 == 5'h9; // @[Replacement.scala 315:30]
  wire  set_touch_ways_1_41_valid = touch_ways_1_1_valid & touch_sets_1_0 == 5'h9; // @[Replacement.scala 315:30]
  wire  _T_120 = set_touch_ways_0_41_valid | set_touch_ways_1_41_valid; // @[package.scala 72:59]
  wire [2:0] state_vec_9_left_subtree_state_6 = state_vec_1_9[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_9_right_subtree_state_6 = state_vec_1_9[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_9_left_subtree_state_7 = state_vec_9_left_subtree_state_6[1]; // @[package.scala 154:13]
  wire  state_vec_9_right_subtree_state_7 = state_vec_9_left_subtree_state_6[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_9_T_52 = state_vec_0_set_left_older_7 ? state_vec_9_left_subtree_state_7 : _state_vec_0_T_51; // @[Replacement.scala 203:16]
  wire  _state_vec_9_T_56 = state_vec_0_set_left_older_7 ? _state_vec_0_T_51 : state_vec_9_right_subtree_state_7; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_9_T_57 = {state_vec_0_set_left_older_7,_state_vec_9_T_52,_state_vec_9_T_56}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_9_T_58 = state_vec_0_set_left_older_6 ? state_vec_9_left_subtree_state_6 : _state_vec_9_T_57; // @[Replacement.scala 203:16]
  wire  state_vec_9_left_subtree_state_8 = state_vec_9_right_subtree_state_6[1]; // @[package.scala 154:13]
  wire  state_vec_9_right_subtree_state_8 = state_vec_9_right_subtree_state_6[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_9_T_63 = state_vec_0_set_left_older_7 ? state_vec_9_left_subtree_state_8 : _state_vec_0_T_51; // @[Replacement.scala 203:16]
  wire  _state_vec_9_T_67 = state_vec_0_set_left_older_7 ? _state_vec_0_T_51 : state_vec_9_right_subtree_state_8; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_9_T_68 = {state_vec_0_set_left_older_7,_state_vec_9_T_63,_state_vec_9_T_67}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_9_T_69 = state_vec_0_set_left_older_6 ? _state_vec_9_T_68 : state_vec_9_right_subtree_state_6; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_9_T_70 = {state_vec_0_set_left_older_6,_state_vec_9_T_58,_state_vec_9_T_69}; // @[Cat.scala 31:58]
  wire [6:0] _state_vec_9_T_71 = set_touch_ways_0_41_valid ? _state_vec_9_T_70 : state_vec_1_9; // @[Replacement.scala 22:56]
  wire [2:0] state_vec_9_left_subtree_state_9 = _state_vec_9_T_71[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_9_right_subtree_state_9 = _state_vec_9_T_71[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_9_left_subtree_state_10 = state_vec_9_left_subtree_state_9[1]; // @[package.scala 154:13]
  wire  state_vec_9_right_subtree_state_10 = state_vec_9_left_subtree_state_9[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_9_T_76 = state_vec_0_set_left_older_10 ? state_vec_9_left_subtree_state_10 : _state_vec_0_T_75; // @[Replacement.scala 203:16]
  wire  _state_vec_9_T_80 = state_vec_0_set_left_older_10 ? _state_vec_0_T_75 : state_vec_9_right_subtree_state_10; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_9_T_81 = {state_vec_0_set_left_older_10,_state_vec_9_T_76,_state_vec_9_T_80}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_9_T_82 = state_vec_0_set_left_older_9 ? state_vec_9_left_subtree_state_9 : _state_vec_9_T_81; // @[Replacement.scala 203:16]
  wire  state_vec_9_left_subtree_state_11 = state_vec_9_right_subtree_state_9[1]; // @[package.scala 154:13]
  wire  state_vec_9_right_subtree_state_11 = state_vec_9_right_subtree_state_9[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_9_T_87 = state_vec_0_set_left_older_10 ? state_vec_9_left_subtree_state_11 : _state_vec_0_T_75; // @[Replacement.scala 203:16]
  wire  _state_vec_9_T_91 = state_vec_0_set_left_older_10 ? _state_vec_0_T_75 : state_vec_9_right_subtree_state_11; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_9_T_92 = {state_vec_0_set_left_older_10,_state_vec_9_T_87,_state_vec_9_T_91}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_9_T_93 = state_vec_0_set_left_older_9 ? _state_vec_9_T_92 : state_vec_9_right_subtree_state_9; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_9_T_94 = {state_vec_0_set_left_older_9,_state_vec_9_T_82,_state_vec_9_T_93}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_42_valid = touch_ways_1_0_valid & touch_sets_1_0 == 5'ha; // @[Replacement.scala 315:30]
  wire  set_touch_ways_1_42_valid = touch_ways_1_1_valid & touch_sets_1_0 == 5'ha; // @[Replacement.scala 315:30]
  wire  _T_121 = set_touch_ways_0_42_valid | set_touch_ways_1_42_valid; // @[package.scala 72:59]
  wire [2:0] state_vec_10_left_subtree_state_6 = state_vec_1_10[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_10_right_subtree_state_6 = state_vec_1_10[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_10_left_subtree_state_7 = state_vec_10_left_subtree_state_6[1]; // @[package.scala 154:13]
  wire  state_vec_10_right_subtree_state_7 = state_vec_10_left_subtree_state_6[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_10_T_52 = state_vec_0_set_left_older_7 ? state_vec_10_left_subtree_state_7 : _state_vec_0_T_51; // @[Replacement.scala 203:16]
  wire  _state_vec_10_T_56 = state_vec_0_set_left_older_7 ? _state_vec_0_T_51 : state_vec_10_right_subtree_state_7; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_10_T_57 = {state_vec_0_set_left_older_7,_state_vec_10_T_52,_state_vec_10_T_56}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_10_T_58 = state_vec_0_set_left_older_6 ? state_vec_10_left_subtree_state_6 : _state_vec_10_T_57; // @[Replacement.scala 203:16]
  wire  state_vec_10_left_subtree_state_8 = state_vec_10_right_subtree_state_6[1]; // @[package.scala 154:13]
  wire  state_vec_10_right_subtree_state_8 = state_vec_10_right_subtree_state_6[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_10_T_63 = state_vec_0_set_left_older_7 ? state_vec_10_left_subtree_state_8 : _state_vec_0_T_51; // @[Replacement.scala 203:16]
  wire  _state_vec_10_T_67 = state_vec_0_set_left_older_7 ? _state_vec_0_T_51 : state_vec_10_right_subtree_state_8; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_10_T_68 = {state_vec_0_set_left_older_7,_state_vec_10_T_63,_state_vec_10_T_67}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_10_T_69 = state_vec_0_set_left_older_6 ? _state_vec_10_T_68 : state_vec_10_right_subtree_state_6
    ; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_10_T_70 = {state_vec_0_set_left_older_6,_state_vec_10_T_58,_state_vec_10_T_69}; // @[Cat.scala 31:58]
  wire [6:0] _state_vec_10_T_71 = set_touch_ways_0_42_valid ? _state_vec_10_T_70 : state_vec_1_10; // @[Replacement.scala 22:56]
  wire [2:0] state_vec_10_left_subtree_state_9 = _state_vec_10_T_71[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_10_right_subtree_state_9 = _state_vec_10_T_71[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_10_left_subtree_state_10 = state_vec_10_left_subtree_state_9[1]; // @[package.scala 154:13]
  wire  state_vec_10_right_subtree_state_10 = state_vec_10_left_subtree_state_9[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_10_T_76 = state_vec_0_set_left_older_10 ? state_vec_10_left_subtree_state_10 : _state_vec_0_T_75; // @[Replacement.scala 203:16]
  wire  _state_vec_10_T_80 = state_vec_0_set_left_older_10 ? _state_vec_0_T_75 : state_vec_10_right_subtree_state_10; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_10_T_81 = {state_vec_0_set_left_older_10,_state_vec_10_T_76,_state_vec_10_T_80}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_10_T_82 = state_vec_0_set_left_older_9 ? state_vec_10_left_subtree_state_9 : _state_vec_10_T_81; // @[Replacement.scala 203:16]
  wire  state_vec_10_left_subtree_state_11 = state_vec_10_right_subtree_state_9[1]; // @[package.scala 154:13]
  wire  state_vec_10_right_subtree_state_11 = state_vec_10_right_subtree_state_9[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_10_T_87 = state_vec_0_set_left_older_10 ? state_vec_10_left_subtree_state_11 : _state_vec_0_T_75; // @[Replacement.scala 203:16]
  wire  _state_vec_10_T_91 = state_vec_0_set_left_older_10 ? _state_vec_0_T_75 : state_vec_10_right_subtree_state_11; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_10_T_92 = {state_vec_0_set_left_older_10,_state_vec_10_T_87,_state_vec_10_T_91}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_10_T_93 = state_vec_0_set_left_older_9 ? _state_vec_10_T_92 : state_vec_10_right_subtree_state_9
    ; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_10_T_94 = {state_vec_0_set_left_older_9,_state_vec_10_T_82,_state_vec_10_T_93}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_43_valid = touch_ways_1_0_valid & touch_sets_1_0 == 5'hb; // @[Replacement.scala 315:30]
  wire  set_touch_ways_1_43_valid = touch_ways_1_1_valid & touch_sets_1_0 == 5'hb; // @[Replacement.scala 315:30]
  wire  _T_122 = set_touch_ways_0_43_valid | set_touch_ways_1_43_valid; // @[package.scala 72:59]
  wire [2:0] state_vec_11_left_subtree_state_6 = state_vec_1_11[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_11_right_subtree_state_6 = state_vec_1_11[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_11_left_subtree_state_7 = state_vec_11_left_subtree_state_6[1]; // @[package.scala 154:13]
  wire  state_vec_11_right_subtree_state_7 = state_vec_11_left_subtree_state_6[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_11_T_52 = state_vec_0_set_left_older_7 ? state_vec_11_left_subtree_state_7 : _state_vec_0_T_51; // @[Replacement.scala 203:16]
  wire  _state_vec_11_T_56 = state_vec_0_set_left_older_7 ? _state_vec_0_T_51 : state_vec_11_right_subtree_state_7; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_11_T_57 = {state_vec_0_set_left_older_7,_state_vec_11_T_52,_state_vec_11_T_56}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_11_T_58 = state_vec_0_set_left_older_6 ? state_vec_11_left_subtree_state_6 : _state_vec_11_T_57; // @[Replacement.scala 203:16]
  wire  state_vec_11_left_subtree_state_8 = state_vec_11_right_subtree_state_6[1]; // @[package.scala 154:13]
  wire  state_vec_11_right_subtree_state_8 = state_vec_11_right_subtree_state_6[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_11_T_63 = state_vec_0_set_left_older_7 ? state_vec_11_left_subtree_state_8 : _state_vec_0_T_51; // @[Replacement.scala 203:16]
  wire  _state_vec_11_T_67 = state_vec_0_set_left_older_7 ? _state_vec_0_T_51 : state_vec_11_right_subtree_state_8; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_11_T_68 = {state_vec_0_set_left_older_7,_state_vec_11_T_63,_state_vec_11_T_67}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_11_T_69 = state_vec_0_set_left_older_6 ? _state_vec_11_T_68 : state_vec_11_right_subtree_state_6
    ; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_11_T_70 = {state_vec_0_set_left_older_6,_state_vec_11_T_58,_state_vec_11_T_69}; // @[Cat.scala 31:58]
  wire [6:0] _state_vec_11_T_71 = set_touch_ways_0_43_valid ? _state_vec_11_T_70 : state_vec_1_11; // @[Replacement.scala 22:56]
  wire [2:0] state_vec_11_left_subtree_state_9 = _state_vec_11_T_71[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_11_right_subtree_state_9 = _state_vec_11_T_71[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_11_left_subtree_state_10 = state_vec_11_left_subtree_state_9[1]; // @[package.scala 154:13]
  wire  state_vec_11_right_subtree_state_10 = state_vec_11_left_subtree_state_9[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_11_T_76 = state_vec_0_set_left_older_10 ? state_vec_11_left_subtree_state_10 : _state_vec_0_T_75; // @[Replacement.scala 203:16]
  wire  _state_vec_11_T_80 = state_vec_0_set_left_older_10 ? _state_vec_0_T_75 : state_vec_11_right_subtree_state_10; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_11_T_81 = {state_vec_0_set_left_older_10,_state_vec_11_T_76,_state_vec_11_T_80}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_11_T_82 = state_vec_0_set_left_older_9 ? state_vec_11_left_subtree_state_9 : _state_vec_11_T_81; // @[Replacement.scala 203:16]
  wire  state_vec_11_left_subtree_state_11 = state_vec_11_right_subtree_state_9[1]; // @[package.scala 154:13]
  wire  state_vec_11_right_subtree_state_11 = state_vec_11_right_subtree_state_9[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_11_T_87 = state_vec_0_set_left_older_10 ? state_vec_11_left_subtree_state_11 : _state_vec_0_T_75; // @[Replacement.scala 203:16]
  wire  _state_vec_11_T_91 = state_vec_0_set_left_older_10 ? _state_vec_0_T_75 : state_vec_11_right_subtree_state_11; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_11_T_92 = {state_vec_0_set_left_older_10,_state_vec_11_T_87,_state_vec_11_T_91}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_11_T_93 = state_vec_0_set_left_older_9 ? _state_vec_11_T_92 : state_vec_11_right_subtree_state_9
    ; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_11_T_94 = {state_vec_0_set_left_older_9,_state_vec_11_T_82,_state_vec_11_T_93}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_44_valid = touch_ways_1_0_valid & touch_sets_1_0 == 5'hc; // @[Replacement.scala 315:30]
  wire  set_touch_ways_1_44_valid = touch_ways_1_1_valid & touch_sets_1_0 == 5'hc; // @[Replacement.scala 315:30]
  wire  _T_123 = set_touch_ways_0_44_valid | set_touch_ways_1_44_valid; // @[package.scala 72:59]
  wire [2:0] state_vec_12_left_subtree_state_6 = state_vec_1_12[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_12_right_subtree_state_6 = state_vec_1_12[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_12_left_subtree_state_7 = state_vec_12_left_subtree_state_6[1]; // @[package.scala 154:13]
  wire  state_vec_12_right_subtree_state_7 = state_vec_12_left_subtree_state_6[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_12_T_52 = state_vec_0_set_left_older_7 ? state_vec_12_left_subtree_state_7 : _state_vec_0_T_51; // @[Replacement.scala 203:16]
  wire  _state_vec_12_T_56 = state_vec_0_set_left_older_7 ? _state_vec_0_T_51 : state_vec_12_right_subtree_state_7; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_12_T_57 = {state_vec_0_set_left_older_7,_state_vec_12_T_52,_state_vec_12_T_56}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_12_T_58 = state_vec_0_set_left_older_6 ? state_vec_12_left_subtree_state_6 : _state_vec_12_T_57; // @[Replacement.scala 203:16]
  wire  state_vec_12_left_subtree_state_8 = state_vec_12_right_subtree_state_6[1]; // @[package.scala 154:13]
  wire  state_vec_12_right_subtree_state_8 = state_vec_12_right_subtree_state_6[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_12_T_63 = state_vec_0_set_left_older_7 ? state_vec_12_left_subtree_state_8 : _state_vec_0_T_51; // @[Replacement.scala 203:16]
  wire  _state_vec_12_T_67 = state_vec_0_set_left_older_7 ? _state_vec_0_T_51 : state_vec_12_right_subtree_state_8; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_12_T_68 = {state_vec_0_set_left_older_7,_state_vec_12_T_63,_state_vec_12_T_67}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_12_T_69 = state_vec_0_set_left_older_6 ? _state_vec_12_T_68 : state_vec_12_right_subtree_state_6
    ; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_12_T_70 = {state_vec_0_set_left_older_6,_state_vec_12_T_58,_state_vec_12_T_69}; // @[Cat.scala 31:58]
  wire [6:0] _state_vec_12_T_71 = set_touch_ways_0_44_valid ? _state_vec_12_T_70 : state_vec_1_12; // @[Replacement.scala 22:56]
  wire [2:0] state_vec_12_left_subtree_state_9 = _state_vec_12_T_71[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_12_right_subtree_state_9 = _state_vec_12_T_71[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_12_left_subtree_state_10 = state_vec_12_left_subtree_state_9[1]; // @[package.scala 154:13]
  wire  state_vec_12_right_subtree_state_10 = state_vec_12_left_subtree_state_9[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_12_T_76 = state_vec_0_set_left_older_10 ? state_vec_12_left_subtree_state_10 : _state_vec_0_T_75; // @[Replacement.scala 203:16]
  wire  _state_vec_12_T_80 = state_vec_0_set_left_older_10 ? _state_vec_0_T_75 : state_vec_12_right_subtree_state_10; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_12_T_81 = {state_vec_0_set_left_older_10,_state_vec_12_T_76,_state_vec_12_T_80}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_12_T_82 = state_vec_0_set_left_older_9 ? state_vec_12_left_subtree_state_9 : _state_vec_12_T_81; // @[Replacement.scala 203:16]
  wire  state_vec_12_left_subtree_state_11 = state_vec_12_right_subtree_state_9[1]; // @[package.scala 154:13]
  wire  state_vec_12_right_subtree_state_11 = state_vec_12_right_subtree_state_9[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_12_T_87 = state_vec_0_set_left_older_10 ? state_vec_12_left_subtree_state_11 : _state_vec_0_T_75; // @[Replacement.scala 203:16]
  wire  _state_vec_12_T_91 = state_vec_0_set_left_older_10 ? _state_vec_0_T_75 : state_vec_12_right_subtree_state_11; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_12_T_92 = {state_vec_0_set_left_older_10,_state_vec_12_T_87,_state_vec_12_T_91}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_12_T_93 = state_vec_0_set_left_older_9 ? _state_vec_12_T_92 : state_vec_12_right_subtree_state_9
    ; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_12_T_94 = {state_vec_0_set_left_older_9,_state_vec_12_T_82,_state_vec_12_T_93}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_45_valid = touch_ways_1_0_valid & touch_sets_1_0 == 5'hd; // @[Replacement.scala 315:30]
  wire  set_touch_ways_1_45_valid = touch_ways_1_1_valid & touch_sets_1_0 == 5'hd; // @[Replacement.scala 315:30]
  wire  _T_124 = set_touch_ways_0_45_valid | set_touch_ways_1_45_valid; // @[package.scala 72:59]
  wire [2:0] state_vec_13_left_subtree_state_6 = state_vec_1_13[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_13_right_subtree_state_6 = state_vec_1_13[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_13_left_subtree_state_7 = state_vec_13_left_subtree_state_6[1]; // @[package.scala 154:13]
  wire  state_vec_13_right_subtree_state_7 = state_vec_13_left_subtree_state_6[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_13_T_52 = state_vec_0_set_left_older_7 ? state_vec_13_left_subtree_state_7 : _state_vec_0_T_51; // @[Replacement.scala 203:16]
  wire  _state_vec_13_T_56 = state_vec_0_set_left_older_7 ? _state_vec_0_T_51 : state_vec_13_right_subtree_state_7; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_13_T_57 = {state_vec_0_set_left_older_7,_state_vec_13_T_52,_state_vec_13_T_56}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_13_T_58 = state_vec_0_set_left_older_6 ? state_vec_13_left_subtree_state_6 : _state_vec_13_T_57; // @[Replacement.scala 203:16]
  wire  state_vec_13_left_subtree_state_8 = state_vec_13_right_subtree_state_6[1]; // @[package.scala 154:13]
  wire  state_vec_13_right_subtree_state_8 = state_vec_13_right_subtree_state_6[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_13_T_63 = state_vec_0_set_left_older_7 ? state_vec_13_left_subtree_state_8 : _state_vec_0_T_51; // @[Replacement.scala 203:16]
  wire  _state_vec_13_T_67 = state_vec_0_set_left_older_7 ? _state_vec_0_T_51 : state_vec_13_right_subtree_state_8; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_13_T_68 = {state_vec_0_set_left_older_7,_state_vec_13_T_63,_state_vec_13_T_67}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_13_T_69 = state_vec_0_set_left_older_6 ? _state_vec_13_T_68 : state_vec_13_right_subtree_state_6
    ; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_13_T_70 = {state_vec_0_set_left_older_6,_state_vec_13_T_58,_state_vec_13_T_69}; // @[Cat.scala 31:58]
  wire [6:0] _state_vec_13_T_71 = set_touch_ways_0_45_valid ? _state_vec_13_T_70 : state_vec_1_13; // @[Replacement.scala 22:56]
  wire [2:0] state_vec_13_left_subtree_state_9 = _state_vec_13_T_71[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_13_right_subtree_state_9 = _state_vec_13_T_71[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_13_left_subtree_state_10 = state_vec_13_left_subtree_state_9[1]; // @[package.scala 154:13]
  wire  state_vec_13_right_subtree_state_10 = state_vec_13_left_subtree_state_9[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_13_T_76 = state_vec_0_set_left_older_10 ? state_vec_13_left_subtree_state_10 : _state_vec_0_T_75; // @[Replacement.scala 203:16]
  wire  _state_vec_13_T_80 = state_vec_0_set_left_older_10 ? _state_vec_0_T_75 : state_vec_13_right_subtree_state_10; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_13_T_81 = {state_vec_0_set_left_older_10,_state_vec_13_T_76,_state_vec_13_T_80}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_13_T_82 = state_vec_0_set_left_older_9 ? state_vec_13_left_subtree_state_9 : _state_vec_13_T_81; // @[Replacement.scala 203:16]
  wire  state_vec_13_left_subtree_state_11 = state_vec_13_right_subtree_state_9[1]; // @[package.scala 154:13]
  wire  state_vec_13_right_subtree_state_11 = state_vec_13_right_subtree_state_9[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_13_T_87 = state_vec_0_set_left_older_10 ? state_vec_13_left_subtree_state_11 : _state_vec_0_T_75; // @[Replacement.scala 203:16]
  wire  _state_vec_13_T_91 = state_vec_0_set_left_older_10 ? _state_vec_0_T_75 : state_vec_13_right_subtree_state_11; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_13_T_92 = {state_vec_0_set_left_older_10,_state_vec_13_T_87,_state_vec_13_T_91}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_13_T_93 = state_vec_0_set_left_older_9 ? _state_vec_13_T_92 : state_vec_13_right_subtree_state_9
    ; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_13_T_94 = {state_vec_0_set_left_older_9,_state_vec_13_T_82,_state_vec_13_T_93}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_46_valid = touch_ways_1_0_valid & touch_sets_1_0 == 5'he; // @[Replacement.scala 315:30]
  wire  set_touch_ways_1_46_valid = touch_ways_1_1_valid & touch_sets_1_0 == 5'he; // @[Replacement.scala 315:30]
  wire  _T_125 = set_touch_ways_0_46_valid | set_touch_ways_1_46_valid; // @[package.scala 72:59]
  wire [2:0] state_vec_14_left_subtree_state_6 = state_vec_1_14[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_14_right_subtree_state_6 = state_vec_1_14[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_14_left_subtree_state_7 = state_vec_14_left_subtree_state_6[1]; // @[package.scala 154:13]
  wire  state_vec_14_right_subtree_state_7 = state_vec_14_left_subtree_state_6[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_14_T_52 = state_vec_0_set_left_older_7 ? state_vec_14_left_subtree_state_7 : _state_vec_0_T_51; // @[Replacement.scala 203:16]
  wire  _state_vec_14_T_56 = state_vec_0_set_left_older_7 ? _state_vec_0_T_51 : state_vec_14_right_subtree_state_7; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_14_T_57 = {state_vec_0_set_left_older_7,_state_vec_14_T_52,_state_vec_14_T_56}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_14_T_58 = state_vec_0_set_left_older_6 ? state_vec_14_left_subtree_state_6 : _state_vec_14_T_57; // @[Replacement.scala 203:16]
  wire  state_vec_14_left_subtree_state_8 = state_vec_14_right_subtree_state_6[1]; // @[package.scala 154:13]
  wire  state_vec_14_right_subtree_state_8 = state_vec_14_right_subtree_state_6[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_14_T_63 = state_vec_0_set_left_older_7 ? state_vec_14_left_subtree_state_8 : _state_vec_0_T_51; // @[Replacement.scala 203:16]
  wire  _state_vec_14_T_67 = state_vec_0_set_left_older_7 ? _state_vec_0_T_51 : state_vec_14_right_subtree_state_8; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_14_T_68 = {state_vec_0_set_left_older_7,_state_vec_14_T_63,_state_vec_14_T_67}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_14_T_69 = state_vec_0_set_left_older_6 ? _state_vec_14_T_68 : state_vec_14_right_subtree_state_6
    ; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_14_T_70 = {state_vec_0_set_left_older_6,_state_vec_14_T_58,_state_vec_14_T_69}; // @[Cat.scala 31:58]
  wire [6:0] _state_vec_14_T_71 = set_touch_ways_0_46_valid ? _state_vec_14_T_70 : state_vec_1_14; // @[Replacement.scala 22:56]
  wire [2:0] state_vec_14_left_subtree_state_9 = _state_vec_14_T_71[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_14_right_subtree_state_9 = _state_vec_14_T_71[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_14_left_subtree_state_10 = state_vec_14_left_subtree_state_9[1]; // @[package.scala 154:13]
  wire  state_vec_14_right_subtree_state_10 = state_vec_14_left_subtree_state_9[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_14_T_76 = state_vec_0_set_left_older_10 ? state_vec_14_left_subtree_state_10 : _state_vec_0_T_75; // @[Replacement.scala 203:16]
  wire  _state_vec_14_T_80 = state_vec_0_set_left_older_10 ? _state_vec_0_T_75 : state_vec_14_right_subtree_state_10; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_14_T_81 = {state_vec_0_set_left_older_10,_state_vec_14_T_76,_state_vec_14_T_80}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_14_T_82 = state_vec_0_set_left_older_9 ? state_vec_14_left_subtree_state_9 : _state_vec_14_T_81; // @[Replacement.scala 203:16]
  wire  state_vec_14_left_subtree_state_11 = state_vec_14_right_subtree_state_9[1]; // @[package.scala 154:13]
  wire  state_vec_14_right_subtree_state_11 = state_vec_14_right_subtree_state_9[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_14_T_87 = state_vec_0_set_left_older_10 ? state_vec_14_left_subtree_state_11 : _state_vec_0_T_75; // @[Replacement.scala 203:16]
  wire  _state_vec_14_T_91 = state_vec_0_set_left_older_10 ? _state_vec_0_T_75 : state_vec_14_right_subtree_state_11; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_14_T_92 = {state_vec_0_set_left_older_10,_state_vec_14_T_87,_state_vec_14_T_91}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_14_T_93 = state_vec_0_set_left_older_9 ? _state_vec_14_T_92 : state_vec_14_right_subtree_state_9
    ; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_14_T_94 = {state_vec_0_set_left_older_9,_state_vec_14_T_82,_state_vec_14_T_93}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_47_valid = touch_ways_1_0_valid & touch_sets_1_0 == 5'hf; // @[Replacement.scala 315:30]
  wire  set_touch_ways_1_47_valid = touch_ways_1_1_valid & touch_sets_1_0 == 5'hf; // @[Replacement.scala 315:30]
  wire  _T_126 = set_touch_ways_0_47_valid | set_touch_ways_1_47_valid; // @[package.scala 72:59]
  wire [2:0] state_vec_15_left_subtree_state_6 = state_vec_1_15[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_15_right_subtree_state_6 = state_vec_1_15[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_15_left_subtree_state_7 = state_vec_15_left_subtree_state_6[1]; // @[package.scala 154:13]
  wire  state_vec_15_right_subtree_state_7 = state_vec_15_left_subtree_state_6[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_15_T_52 = state_vec_0_set_left_older_7 ? state_vec_15_left_subtree_state_7 : _state_vec_0_T_51; // @[Replacement.scala 203:16]
  wire  _state_vec_15_T_56 = state_vec_0_set_left_older_7 ? _state_vec_0_T_51 : state_vec_15_right_subtree_state_7; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_15_T_57 = {state_vec_0_set_left_older_7,_state_vec_15_T_52,_state_vec_15_T_56}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_15_T_58 = state_vec_0_set_left_older_6 ? state_vec_15_left_subtree_state_6 : _state_vec_15_T_57; // @[Replacement.scala 203:16]
  wire  state_vec_15_left_subtree_state_8 = state_vec_15_right_subtree_state_6[1]; // @[package.scala 154:13]
  wire  state_vec_15_right_subtree_state_8 = state_vec_15_right_subtree_state_6[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_15_T_63 = state_vec_0_set_left_older_7 ? state_vec_15_left_subtree_state_8 : _state_vec_0_T_51; // @[Replacement.scala 203:16]
  wire  _state_vec_15_T_67 = state_vec_0_set_left_older_7 ? _state_vec_0_T_51 : state_vec_15_right_subtree_state_8; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_15_T_68 = {state_vec_0_set_left_older_7,_state_vec_15_T_63,_state_vec_15_T_67}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_15_T_69 = state_vec_0_set_left_older_6 ? _state_vec_15_T_68 : state_vec_15_right_subtree_state_6
    ; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_15_T_70 = {state_vec_0_set_left_older_6,_state_vec_15_T_58,_state_vec_15_T_69}; // @[Cat.scala 31:58]
  wire [6:0] _state_vec_15_T_71 = set_touch_ways_0_47_valid ? _state_vec_15_T_70 : state_vec_1_15; // @[Replacement.scala 22:56]
  wire [2:0] state_vec_15_left_subtree_state_9 = _state_vec_15_T_71[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_15_right_subtree_state_9 = _state_vec_15_T_71[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_15_left_subtree_state_10 = state_vec_15_left_subtree_state_9[1]; // @[package.scala 154:13]
  wire  state_vec_15_right_subtree_state_10 = state_vec_15_left_subtree_state_9[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_15_T_76 = state_vec_0_set_left_older_10 ? state_vec_15_left_subtree_state_10 : _state_vec_0_T_75; // @[Replacement.scala 203:16]
  wire  _state_vec_15_T_80 = state_vec_0_set_left_older_10 ? _state_vec_0_T_75 : state_vec_15_right_subtree_state_10; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_15_T_81 = {state_vec_0_set_left_older_10,_state_vec_15_T_76,_state_vec_15_T_80}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_15_T_82 = state_vec_0_set_left_older_9 ? state_vec_15_left_subtree_state_9 : _state_vec_15_T_81; // @[Replacement.scala 203:16]
  wire  state_vec_15_left_subtree_state_11 = state_vec_15_right_subtree_state_9[1]; // @[package.scala 154:13]
  wire  state_vec_15_right_subtree_state_11 = state_vec_15_right_subtree_state_9[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_15_T_87 = state_vec_0_set_left_older_10 ? state_vec_15_left_subtree_state_11 : _state_vec_0_T_75; // @[Replacement.scala 203:16]
  wire  _state_vec_15_T_91 = state_vec_0_set_left_older_10 ? _state_vec_0_T_75 : state_vec_15_right_subtree_state_11; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_15_T_92 = {state_vec_0_set_left_older_10,_state_vec_15_T_87,_state_vec_15_T_91}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_15_T_93 = state_vec_0_set_left_older_9 ? _state_vec_15_T_92 : state_vec_15_right_subtree_state_9
    ; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_15_T_94 = {state_vec_0_set_left_older_9,_state_vec_15_T_82,_state_vec_15_T_93}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_48_valid = touch_ways_1_0_valid & touch_sets_1_0 == 5'h10; // @[Replacement.scala 315:30]
  wire  set_touch_ways_1_48_valid = touch_ways_1_1_valid & touch_sets_1_0 == 5'h10; // @[Replacement.scala 315:30]
  wire  _T_127 = set_touch_ways_0_48_valid | set_touch_ways_1_48_valid; // @[package.scala 72:59]
  wire [2:0] state_vec_16_left_subtree_state_6 = state_vec_1_16[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_16_right_subtree_state_6 = state_vec_1_16[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_16_left_subtree_state_7 = state_vec_16_left_subtree_state_6[1]; // @[package.scala 154:13]
  wire  state_vec_16_right_subtree_state_7 = state_vec_16_left_subtree_state_6[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_16_T_52 = state_vec_0_set_left_older_7 ? state_vec_16_left_subtree_state_7 : _state_vec_0_T_51; // @[Replacement.scala 203:16]
  wire  _state_vec_16_T_56 = state_vec_0_set_left_older_7 ? _state_vec_0_T_51 : state_vec_16_right_subtree_state_7; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_16_T_57 = {state_vec_0_set_left_older_7,_state_vec_16_T_52,_state_vec_16_T_56}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_16_T_58 = state_vec_0_set_left_older_6 ? state_vec_16_left_subtree_state_6 : _state_vec_16_T_57; // @[Replacement.scala 203:16]
  wire  state_vec_16_left_subtree_state_8 = state_vec_16_right_subtree_state_6[1]; // @[package.scala 154:13]
  wire  state_vec_16_right_subtree_state_8 = state_vec_16_right_subtree_state_6[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_16_T_63 = state_vec_0_set_left_older_7 ? state_vec_16_left_subtree_state_8 : _state_vec_0_T_51; // @[Replacement.scala 203:16]
  wire  _state_vec_16_T_67 = state_vec_0_set_left_older_7 ? _state_vec_0_T_51 : state_vec_16_right_subtree_state_8; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_16_T_68 = {state_vec_0_set_left_older_7,_state_vec_16_T_63,_state_vec_16_T_67}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_16_T_69 = state_vec_0_set_left_older_6 ? _state_vec_16_T_68 : state_vec_16_right_subtree_state_6
    ; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_16_T_70 = {state_vec_0_set_left_older_6,_state_vec_16_T_58,_state_vec_16_T_69}; // @[Cat.scala 31:58]
  wire [6:0] _state_vec_16_T_71 = set_touch_ways_0_48_valid ? _state_vec_16_T_70 : state_vec_1_16; // @[Replacement.scala 22:56]
  wire [2:0] state_vec_16_left_subtree_state_9 = _state_vec_16_T_71[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_16_right_subtree_state_9 = _state_vec_16_T_71[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_16_left_subtree_state_10 = state_vec_16_left_subtree_state_9[1]; // @[package.scala 154:13]
  wire  state_vec_16_right_subtree_state_10 = state_vec_16_left_subtree_state_9[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_16_T_76 = state_vec_0_set_left_older_10 ? state_vec_16_left_subtree_state_10 : _state_vec_0_T_75; // @[Replacement.scala 203:16]
  wire  _state_vec_16_T_80 = state_vec_0_set_left_older_10 ? _state_vec_0_T_75 : state_vec_16_right_subtree_state_10; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_16_T_81 = {state_vec_0_set_left_older_10,_state_vec_16_T_76,_state_vec_16_T_80}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_16_T_82 = state_vec_0_set_left_older_9 ? state_vec_16_left_subtree_state_9 : _state_vec_16_T_81; // @[Replacement.scala 203:16]
  wire  state_vec_16_left_subtree_state_11 = state_vec_16_right_subtree_state_9[1]; // @[package.scala 154:13]
  wire  state_vec_16_right_subtree_state_11 = state_vec_16_right_subtree_state_9[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_16_T_87 = state_vec_0_set_left_older_10 ? state_vec_16_left_subtree_state_11 : _state_vec_0_T_75; // @[Replacement.scala 203:16]
  wire  _state_vec_16_T_91 = state_vec_0_set_left_older_10 ? _state_vec_0_T_75 : state_vec_16_right_subtree_state_11; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_16_T_92 = {state_vec_0_set_left_older_10,_state_vec_16_T_87,_state_vec_16_T_91}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_16_T_93 = state_vec_0_set_left_older_9 ? _state_vec_16_T_92 : state_vec_16_right_subtree_state_9
    ; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_16_T_94 = {state_vec_0_set_left_older_9,_state_vec_16_T_82,_state_vec_16_T_93}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_49_valid = touch_ways_1_0_valid & touch_sets_1_0 == 5'h11; // @[Replacement.scala 315:30]
  wire  set_touch_ways_1_49_valid = touch_ways_1_1_valid & touch_sets_1_0 == 5'h11; // @[Replacement.scala 315:30]
  wire  _T_128 = set_touch_ways_0_49_valid | set_touch_ways_1_49_valid; // @[package.scala 72:59]
  wire [2:0] state_vec_17_left_subtree_state_6 = state_vec_1_17[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_17_right_subtree_state_6 = state_vec_1_17[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_17_left_subtree_state_7 = state_vec_17_left_subtree_state_6[1]; // @[package.scala 154:13]
  wire  state_vec_17_right_subtree_state_7 = state_vec_17_left_subtree_state_6[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_17_T_52 = state_vec_0_set_left_older_7 ? state_vec_17_left_subtree_state_7 : _state_vec_0_T_51; // @[Replacement.scala 203:16]
  wire  _state_vec_17_T_56 = state_vec_0_set_left_older_7 ? _state_vec_0_T_51 : state_vec_17_right_subtree_state_7; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_17_T_57 = {state_vec_0_set_left_older_7,_state_vec_17_T_52,_state_vec_17_T_56}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_17_T_58 = state_vec_0_set_left_older_6 ? state_vec_17_left_subtree_state_6 : _state_vec_17_T_57; // @[Replacement.scala 203:16]
  wire  state_vec_17_left_subtree_state_8 = state_vec_17_right_subtree_state_6[1]; // @[package.scala 154:13]
  wire  state_vec_17_right_subtree_state_8 = state_vec_17_right_subtree_state_6[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_17_T_63 = state_vec_0_set_left_older_7 ? state_vec_17_left_subtree_state_8 : _state_vec_0_T_51; // @[Replacement.scala 203:16]
  wire  _state_vec_17_T_67 = state_vec_0_set_left_older_7 ? _state_vec_0_T_51 : state_vec_17_right_subtree_state_8; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_17_T_68 = {state_vec_0_set_left_older_7,_state_vec_17_T_63,_state_vec_17_T_67}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_17_T_69 = state_vec_0_set_left_older_6 ? _state_vec_17_T_68 : state_vec_17_right_subtree_state_6
    ; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_17_T_70 = {state_vec_0_set_left_older_6,_state_vec_17_T_58,_state_vec_17_T_69}; // @[Cat.scala 31:58]
  wire [6:0] _state_vec_17_T_71 = set_touch_ways_0_49_valid ? _state_vec_17_T_70 : state_vec_1_17; // @[Replacement.scala 22:56]
  wire [2:0] state_vec_17_left_subtree_state_9 = _state_vec_17_T_71[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_17_right_subtree_state_9 = _state_vec_17_T_71[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_17_left_subtree_state_10 = state_vec_17_left_subtree_state_9[1]; // @[package.scala 154:13]
  wire  state_vec_17_right_subtree_state_10 = state_vec_17_left_subtree_state_9[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_17_T_76 = state_vec_0_set_left_older_10 ? state_vec_17_left_subtree_state_10 : _state_vec_0_T_75; // @[Replacement.scala 203:16]
  wire  _state_vec_17_T_80 = state_vec_0_set_left_older_10 ? _state_vec_0_T_75 : state_vec_17_right_subtree_state_10; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_17_T_81 = {state_vec_0_set_left_older_10,_state_vec_17_T_76,_state_vec_17_T_80}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_17_T_82 = state_vec_0_set_left_older_9 ? state_vec_17_left_subtree_state_9 : _state_vec_17_T_81; // @[Replacement.scala 203:16]
  wire  state_vec_17_left_subtree_state_11 = state_vec_17_right_subtree_state_9[1]; // @[package.scala 154:13]
  wire  state_vec_17_right_subtree_state_11 = state_vec_17_right_subtree_state_9[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_17_T_87 = state_vec_0_set_left_older_10 ? state_vec_17_left_subtree_state_11 : _state_vec_0_T_75; // @[Replacement.scala 203:16]
  wire  _state_vec_17_T_91 = state_vec_0_set_left_older_10 ? _state_vec_0_T_75 : state_vec_17_right_subtree_state_11; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_17_T_92 = {state_vec_0_set_left_older_10,_state_vec_17_T_87,_state_vec_17_T_91}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_17_T_93 = state_vec_0_set_left_older_9 ? _state_vec_17_T_92 : state_vec_17_right_subtree_state_9
    ; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_17_T_94 = {state_vec_0_set_left_older_9,_state_vec_17_T_82,_state_vec_17_T_93}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_50_valid = touch_ways_1_0_valid & touch_sets_1_0 == 5'h12; // @[Replacement.scala 315:30]
  wire  set_touch_ways_1_50_valid = touch_ways_1_1_valid & touch_sets_1_0 == 5'h12; // @[Replacement.scala 315:30]
  wire  _T_129 = set_touch_ways_0_50_valid | set_touch_ways_1_50_valid; // @[package.scala 72:59]
  wire [2:0] state_vec_18_left_subtree_state_6 = state_vec_1_18[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_18_right_subtree_state_6 = state_vec_1_18[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_18_left_subtree_state_7 = state_vec_18_left_subtree_state_6[1]; // @[package.scala 154:13]
  wire  state_vec_18_right_subtree_state_7 = state_vec_18_left_subtree_state_6[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_18_T_52 = state_vec_0_set_left_older_7 ? state_vec_18_left_subtree_state_7 : _state_vec_0_T_51; // @[Replacement.scala 203:16]
  wire  _state_vec_18_T_56 = state_vec_0_set_left_older_7 ? _state_vec_0_T_51 : state_vec_18_right_subtree_state_7; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_18_T_57 = {state_vec_0_set_left_older_7,_state_vec_18_T_52,_state_vec_18_T_56}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_18_T_58 = state_vec_0_set_left_older_6 ? state_vec_18_left_subtree_state_6 : _state_vec_18_T_57; // @[Replacement.scala 203:16]
  wire  state_vec_18_left_subtree_state_8 = state_vec_18_right_subtree_state_6[1]; // @[package.scala 154:13]
  wire  state_vec_18_right_subtree_state_8 = state_vec_18_right_subtree_state_6[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_18_T_63 = state_vec_0_set_left_older_7 ? state_vec_18_left_subtree_state_8 : _state_vec_0_T_51; // @[Replacement.scala 203:16]
  wire  _state_vec_18_T_67 = state_vec_0_set_left_older_7 ? _state_vec_0_T_51 : state_vec_18_right_subtree_state_8; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_18_T_68 = {state_vec_0_set_left_older_7,_state_vec_18_T_63,_state_vec_18_T_67}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_18_T_69 = state_vec_0_set_left_older_6 ? _state_vec_18_T_68 : state_vec_18_right_subtree_state_6
    ; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_18_T_70 = {state_vec_0_set_left_older_6,_state_vec_18_T_58,_state_vec_18_T_69}; // @[Cat.scala 31:58]
  wire [6:0] _state_vec_18_T_71 = set_touch_ways_0_50_valid ? _state_vec_18_T_70 : state_vec_1_18; // @[Replacement.scala 22:56]
  wire [2:0] state_vec_18_left_subtree_state_9 = _state_vec_18_T_71[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_18_right_subtree_state_9 = _state_vec_18_T_71[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_18_left_subtree_state_10 = state_vec_18_left_subtree_state_9[1]; // @[package.scala 154:13]
  wire  state_vec_18_right_subtree_state_10 = state_vec_18_left_subtree_state_9[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_18_T_76 = state_vec_0_set_left_older_10 ? state_vec_18_left_subtree_state_10 : _state_vec_0_T_75; // @[Replacement.scala 203:16]
  wire  _state_vec_18_T_80 = state_vec_0_set_left_older_10 ? _state_vec_0_T_75 : state_vec_18_right_subtree_state_10; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_18_T_81 = {state_vec_0_set_left_older_10,_state_vec_18_T_76,_state_vec_18_T_80}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_18_T_82 = state_vec_0_set_left_older_9 ? state_vec_18_left_subtree_state_9 : _state_vec_18_T_81; // @[Replacement.scala 203:16]
  wire  state_vec_18_left_subtree_state_11 = state_vec_18_right_subtree_state_9[1]; // @[package.scala 154:13]
  wire  state_vec_18_right_subtree_state_11 = state_vec_18_right_subtree_state_9[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_18_T_87 = state_vec_0_set_left_older_10 ? state_vec_18_left_subtree_state_11 : _state_vec_0_T_75; // @[Replacement.scala 203:16]
  wire  _state_vec_18_T_91 = state_vec_0_set_left_older_10 ? _state_vec_0_T_75 : state_vec_18_right_subtree_state_11; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_18_T_92 = {state_vec_0_set_left_older_10,_state_vec_18_T_87,_state_vec_18_T_91}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_18_T_93 = state_vec_0_set_left_older_9 ? _state_vec_18_T_92 : state_vec_18_right_subtree_state_9
    ; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_18_T_94 = {state_vec_0_set_left_older_9,_state_vec_18_T_82,_state_vec_18_T_93}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_51_valid = touch_ways_1_0_valid & touch_sets_1_0 == 5'h13; // @[Replacement.scala 315:30]
  wire  set_touch_ways_1_51_valid = touch_ways_1_1_valid & touch_sets_1_0 == 5'h13; // @[Replacement.scala 315:30]
  wire  _T_130 = set_touch_ways_0_51_valid | set_touch_ways_1_51_valid; // @[package.scala 72:59]
  wire [2:0] state_vec_19_left_subtree_state_6 = state_vec_1_19[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_19_right_subtree_state_6 = state_vec_1_19[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_19_left_subtree_state_7 = state_vec_19_left_subtree_state_6[1]; // @[package.scala 154:13]
  wire  state_vec_19_right_subtree_state_7 = state_vec_19_left_subtree_state_6[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_19_T_52 = state_vec_0_set_left_older_7 ? state_vec_19_left_subtree_state_7 : _state_vec_0_T_51; // @[Replacement.scala 203:16]
  wire  _state_vec_19_T_56 = state_vec_0_set_left_older_7 ? _state_vec_0_T_51 : state_vec_19_right_subtree_state_7; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_19_T_57 = {state_vec_0_set_left_older_7,_state_vec_19_T_52,_state_vec_19_T_56}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_19_T_58 = state_vec_0_set_left_older_6 ? state_vec_19_left_subtree_state_6 : _state_vec_19_T_57; // @[Replacement.scala 203:16]
  wire  state_vec_19_left_subtree_state_8 = state_vec_19_right_subtree_state_6[1]; // @[package.scala 154:13]
  wire  state_vec_19_right_subtree_state_8 = state_vec_19_right_subtree_state_6[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_19_T_63 = state_vec_0_set_left_older_7 ? state_vec_19_left_subtree_state_8 : _state_vec_0_T_51; // @[Replacement.scala 203:16]
  wire  _state_vec_19_T_67 = state_vec_0_set_left_older_7 ? _state_vec_0_T_51 : state_vec_19_right_subtree_state_8; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_19_T_68 = {state_vec_0_set_left_older_7,_state_vec_19_T_63,_state_vec_19_T_67}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_19_T_69 = state_vec_0_set_left_older_6 ? _state_vec_19_T_68 : state_vec_19_right_subtree_state_6
    ; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_19_T_70 = {state_vec_0_set_left_older_6,_state_vec_19_T_58,_state_vec_19_T_69}; // @[Cat.scala 31:58]
  wire [6:0] _state_vec_19_T_71 = set_touch_ways_0_51_valid ? _state_vec_19_T_70 : state_vec_1_19; // @[Replacement.scala 22:56]
  wire [2:0] state_vec_19_left_subtree_state_9 = _state_vec_19_T_71[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_19_right_subtree_state_9 = _state_vec_19_T_71[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_19_left_subtree_state_10 = state_vec_19_left_subtree_state_9[1]; // @[package.scala 154:13]
  wire  state_vec_19_right_subtree_state_10 = state_vec_19_left_subtree_state_9[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_19_T_76 = state_vec_0_set_left_older_10 ? state_vec_19_left_subtree_state_10 : _state_vec_0_T_75; // @[Replacement.scala 203:16]
  wire  _state_vec_19_T_80 = state_vec_0_set_left_older_10 ? _state_vec_0_T_75 : state_vec_19_right_subtree_state_10; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_19_T_81 = {state_vec_0_set_left_older_10,_state_vec_19_T_76,_state_vec_19_T_80}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_19_T_82 = state_vec_0_set_left_older_9 ? state_vec_19_left_subtree_state_9 : _state_vec_19_T_81; // @[Replacement.scala 203:16]
  wire  state_vec_19_left_subtree_state_11 = state_vec_19_right_subtree_state_9[1]; // @[package.scala 154:13]
  wire  state_vec_19_right_subtree_state_11 = state_vec_19_right_subtree_state_9[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_19_T_87 = state_vec_0_set_left_older_10 ? state_vec_19_left_subtree_state_11 : _state_vec_0_T_75; // @[Replacement.scala 203:16]
  wire  _state_vec_19_T_91 = state_vec_0_set_left_older_10 ? _state_vec_0_T_75 : state_vec_19_right_subtree_state_11; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_19_T_92 = {state_vec_0_set_left_older_10,_state_vec_19_T_87,_state_vec_19_T_91}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_19_T_93 = state_vec_0_set_left_older_9 ? _state_vec_19_T_92 : state_vec_19_right_subtree_state_9
    ; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_19_T_94 = {state_vec_0_set_left_older_9,_state_vec_19_T_82,_state_vec_19_T_93}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_52_valid = touch_ways_1_0_valid & touch_sets_1_0 == 5'h14; // @[Replacement.scala 315:30]
  wire  set_touch_ways_1_52_valid = touch_ways_1_1_valid & touch_sets_1_0 == 5'h14; // @[Replacement.scala 315:30]
  wire  _T_131 = set_touch_ways_0_52_valid | set_touch_ways_1_52_valid; // @[package.scala 72:59]
  wire [2:0] state_vec_20_left_subtree_state_6 = state_vec_1_20[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_20_right_subtree_state_6 = state_vec_1_20[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_20_left_subtree_state_7 = state_vec_20_left_subtree_state_6[1]; // @[package.scala 154:13]
  wire  state_vec_20_right_subtree_state_7 = state_vec_20_left_subtree_state_6[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_20_T_52 = state_vec_0_set_left_older_7 ? state_vec_20_left_subtree_state_7 : _state_vec_0_T_51; // @[Replacement.scala 203:16]
  wire  _state_vec_20_T_56 = state_vec_0_set_left_older_7 ? _state_vec_0_T_51 : state_vec_20_right_subtree_state_7; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_20_T_57 = {state_vec_0_set_left_older_7,_state_vec_20_T_52,_state_vec_20_T_56}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_20_T_58 = state_vec_0_set_left_older_6 ? state_vec_20_left_subtree_state_6 : _state_vec_20_T_57; // @[Replacement.scala 203:16]
  wire  state_vec_20_left_subtree_state_8 = state_vec_20_right_subtree_state_6[1]; // @[package.scala 154:13]
  wire  state_vec_20_right_subtree_state_8 = state_vec_20_right_subtree_state_6[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_20_T_63 = state_vec_0_set_left_older_7 ? state_vec_20_left_subtree_state_8 : _state_vec_0_T_51; // @[Replacement.scala 203:16]
  wire  _state_vec_20_T_67 = state_vec_0_set_left_older_7 ? _state_vec_0_T_51 : state_vec_20_right_subtree_state_8; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_20_T_68 = {state_vec_0_set_left_older_7,_state_vec_20_T_63,_state_vec_20_T_67}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_20_T_69 = state_vec_0_set_left_older_6 ? _state_vec_20_T_68 : state_vec_20_right_subtree_state_6
    ; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_20_T_70 = {state_vec_0_set_left_older_6,_state_vec_20_T_58,_state_vec_20_T_69}; // @[Cat.scala 31:58]
  wire [6:0] _state_vec_20_T_71 = set_touch_ways_0_52_valid ? _state_vec_20_T_70 : state_vec_1_20; // @[Replacement.scala 22:56]
  wire [2:0] state_vec_20_left_subtree_state_9 = _state_vec_20_T_71[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_20_right_subtree_state_9 = _state_vec_20_T_71[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_20_left_subtree_state_10 = state_vec_20_left_subtree_state_9[1]; // @[package.scala 154:13]
  wire  state_vec_20_right_subtree_state_10 = state_vec_20_left_subtree_state_9[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_20_T_76 = state_vec_0_set_left_older_10 ? state_vec_20_left_subtree_state_10 : _state_vec_0_T_75; // @[Replacement.scala 203:16]
  wire  _state_vec_20_T_80 = state_vec_0_set_left_older_10 ? _state_vec_0_T_75 : state_vec_20_right_subtree_state_10; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_20_T_81 = {state_vec_0_set_left_older_10,_state_vec_20_T_76,_state_vec_20_T_80}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_20_T_82 = state_vec_0_set_left_older_9 ? state_vec_20_left_subtree_state_9 : _state_vec_20_T_81; // @[Replacement.scala 203:16]
  wire  state_vec_20_left_subtree_state_11 = state_vec_20_right_subtree_state_9[1]; // @[package.scala 154:13]
  wire  state_vec_20_right_subtree_state_11 = state_vec_20_right_subtree_state_9[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_20_T_87 = state_vec_0_set_left_older_10 ? state_vec_20_left_subtree_state_11 : _state_vec_0_T_75; // @[Replacement.scala 203:16]
  wire  _state_vec_20_T_91 = state_vec_0_set_left_older_10 ? _state_vec_0_T_75 : state_vec_20_right_subtree_state_11; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_20_T_92 = {state_vec_0_set_left_older_10,_state_vec_20_T_87,_state_vec_20_T_91}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_20_T_93 = state_vec_0_set_left_older_9 ? _state_vec_20_T_92 : state_vec_20_right_subtree_state_9
    ; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_20_T_94 = {state_vec_0_set_left_older_9,_state_vec_20_T_82,_state_vec_20_T_93}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_53_valid = touch_ways_1_0_valid & touch_sets_1_0 == 5'h15; // @[Replacement.scala 315:30]
  wire  set_touch_ways_1_53_valid = touch_ways_1_1_valid & touch_sets_1_0 == 5'h15; // @[Replacement.scala 315:30]
  wire  _T_132 = set_touch_ways_0_53_valid | set_touch_ways_1_53_valid; // @[package.scala 72:59]
  wire [2:0] state_vec_21_left_subtree_state_6 = state_vec_1_21[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_21_right_subtree_state_6 = state_vec_1_21[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_21_left_subtree_state_7 = state_vec_21_left_subtree_state_6[1]; // @[package.scala 154:13]
  wire  state_vec_21_right_subtree_state_7 = state_vec_21_left_subtree_state_6[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_21_T_52 = state_vec_0_set_left_older_7 ? state_vec_21_left_subtree_state_7 : _state_vec_0_T_51; // @[Replacement.scala 203:16]
  wire  _state_vec_21_T_56 = state_vec_0_set_left_older_7 ? _state_vec_0_T_51 : state_vec_21_right_subtree_state_7; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_21_T_57 = {state_vec_0_set_left_older_7,_state_vec_21_T_52,_state_vec_21_T_56}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_21_T_58 = state_vec_0_set_left_older_6 ? state_vec_21_left_subtree_state_6 : _state_vec_21_T_57; // @[Replacement.scala 203:16]
  wire  state_vec_21_left_subtree_state_8 = state_vec_21_right_subtree_state_6[1]; // @[package.scala 154:13]
  wire  state_vec_21_right_subtree_state_8 = state_vec_21_right_subtree_state_6[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_21_T_63 = state_vec_0_set_left_older_7 ? state_vec_21_left_subtree_state_8 : _state_vec_0_T_51; // @[Replacement.scala 203:16]
  wire  _state_vec_21_T_67 = state_vec_0_set_left_older_7 ? _state_vec_0_T_51 : state_vec_21_right_subtree_state_8; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_21_T_68 = {state_vec_0_set_left_older_7,_state_vec_21_T_63,_state_vec_21_T_67}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_21_T_69 = state_vec_0_set_left_older_6 ? _state_vec_21_T_68 : state_vec_21_right_subtree_state_6
    ; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_21_T_70 = {state_vec_0_set_left_older_6,_state_vec_21_T_58,_state_vec_21_T_69}; // @[Cat.scala 31:58]
  wire [6:0] _state_vec_21_T_71 = set_touch_ways_0_53_valid ? _state_vec_21_T_70 : state_vec_1_21; // @[Replacement.scala 22:56]
  wire [2:0] state_vec_21_left_subtree_state_9 = _state_vec_21_T_71[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_21_right_subtree_state_9 = _state_vec_21_T_71[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_21_left_subtree_state_10 = state_vec_21_left_subtree_state_9[1]; // @[package.scala 154:13]
  wire  state_vec_21_right_subtree_state_10 = state_vec_21_left_subtree_state_9[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_21_T_76 = state_vec_0_set_left_older_10 ? state_vec_21_left_subtree_state_10 : _state_vec_0_T_75; // @[Replacement.scala 203:16]
  wire  _state_vec_21_T_80 = state_vec_0_set_left_older_10 ? _state_vec_0_T_75 : state_vec_21_right_subtree_state_10; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_21_T_81 = {state_vec_0_set_left_older_10,_state_vec_21_T_76,_state_vec_21_T_80}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_21_T_82 = state_vec_0_set_left_older_9 ? state_vec_21_left_subtree_state_9 : _state_vec_21_T_81; // @[Replacement.scala 203:16]
  wire  state_vec_21_left_subtree_state_11 = state_vec_21_right_subtree_state_9[1]; // @[package.scala 154:13]
  wire  state_vec_21_right_subtree_state_11 = state_vec_21_right_subtree_state_9[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_21_T_87 = state_vec_0_set_left_older_10 ? state_vec_21_left_subtree_state_11 : _state_vec_0_T_75; // @[Replacement.scala 203:16]
  wire  _state_vec_21_T_91 = state_vec_0_set_left_older_10 ? _state_vec_0_T_75 : state_vec_21_right_subtree_state_11; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_21_T_92 = {state_vec_0_set_left_older_10,_state_vec_21_T_87,_state_vec_21_T_91}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_21_T_93 = state_vec_0_set_left_older_9 ? _state_vec_21_T_92 : state_vec_21_right_subtree_state_9
    ; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_21_T_94 = {state_vec_0_set_left_older_9,_state_vec_21_T_82,_state_vec_21_T_93}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_54_valid = touch_ways_1_0_valid & touch_sets_1_0 == 5'h16; // @[Replacement.scala 315:30]
  wire  set_touch_ways_1_54_valid = touch_ways_1_1_valid & touch_sets_1_0 == 5'h16; // @[Replacement.scala 315:30]
  wire  _T_133 = set_touch_ways_0_54_valid | set_touch_ways_1_54_valid; // @[package.scala 72:59]
  wire [2:0] state_vec_22_left_subtree_state_6 = state_vec_1_22[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_22_right_subtree_state_6 = state_vec_1_22[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_22_left_subtree_state_7 = state_vec_22_left_subtree_state_6[1]; // @[package.scala 154:13]
  wire  state_vec_22_right_subtree_state_7 = state_vec_22_left_subtree_state_6[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_22_T_52 = state_vec_0_set_left_older_7 ? state_vec_22_left_subtree_state_7 : _state_vec_0_T_51; // @[Replacement.scala 203:16]
  wire  _state_vec_22_T_56 = state_vec_0_set_left_older_7 ? _state_vec_0_T_51 : state_vec_22_right_subtree_state_7; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_22_T_57 = {state_vec_0_set_left_older_7,_state_vec_22_T_52,_state_vec_22_T_56}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_22_T_58 = state_vec_0_set_left_older_6 ? state_vec_22_left_subtree_state_6 : _state_vec_22_T_57; // @[Replacement.scala 203:16]
  wire  state_vec_22_left_subtree_state_8 = state_vec_22_right_subtree_state_6[1]; // @[package.scala 154:13]
  wire  state_vec_22_right_subtree_state_8 = state_vec_22_right_subtree_state_6[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_22_T_63 = state_vec_0_set_left_older_7 ? state_vec_22_left_subtree_state_8 : _state_vec_0_T_51; // @[Replacement.scala 203:16]
  wire  _state_vec_22_T_67 = state_vec_0_set_left_older_7 ? _state_vec_0_T_51 : state_vec_22_right_subtree_state_8; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_22_T_68 = {state_vec_0_set_left_older_7,_state_vec_22_T_63,_state_vec_22_T_67}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_22_T_69 = state_vec_0_set_left_older_6 ? _state_vec_22_T_68 : state_vec_22_right_subtree_state_6
    ; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_22_T_70 = {state_vec_0_set_left_older_6,_state_vec_22_T_58,_state_vec_22_T_69}; // @[Cat.scala 31:58]
  wire [6:0] _state_vec_22_T_71 = set_touch_ways_0_54_valid ? _state_vec_22_T_70 : state_vec_1_22; // @[Replacement.scala 22:56]
  wire [2:0] state_vec_22_left_subtree_state_9 = _state_vec_22_T_71[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_22_right_subtree_state_9 = _state_vec_22_T_71[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_22_left_subtree_state_10 = state_vec_22_left_subtree_state_9[1]; // @[package.scala 154:13]
  wire  state_vec_22_right_subtree_state_10 = state_vec_22_left_subtree_state_9[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_22_T_76 = state_vec_0_set_left_older_10 ? state_vec_22_left_subtree_state_10 : _state_vec_0_T_75; // @[Replacement.scala 203:16]
  wire  _state_vec_22_T_80 = state_vec_0_set_left_older_10 ? _state_vec_0_T_75 : state_vec_22_right_subtree_state_10; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_22_T_81 = {state_vec_0_set_left_older_10,_state_vec_22_T_76,_state_vec_22_T_80}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_22_T_82 = state_vec_0_set_left_older_9 ? state_vec_22_left_subtree_state_9 : _state_vec_22_T_81; // @[Replacement.scala 203:16]
  wire  state_vec_22_left_subtree_state_11 = state_vec_22_right_subtree_state_9[1]; // @[package.scala 154:13]
  wire  state_vec_22_right_subtree_state_11 = state_vec_22_right_subtree_state_9[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_22_T_87 = state_vec_0_set_left_older_10 ? state_vec_22_left_subtree_state_11 : _state_vec_0_T_75; // @[Replacement.scala 203:16]
  wire  _state_vec_22_T_91 = state_vec_0_set_left_older_10 ? _state_vec_0_T_75 : state_vec_22_right_subtree_state_11; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_22_T_92 = {state_vec_0_set_left_older_10,_state_vec_22_T_87,_state_vec_22_T_91}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_22_T_93 = state_vec_0_set_left_older_9 ? _state_vec_22_T_92 : state_vec_22_right_subtree_state_9
    ; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_22_T_94 = {state_vec_0_set_left_older_9,_state_vec_22_T_82,_state_vec_22_T_93}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_55_valid = touch_ways_1_0_valid & touch_sets_1_0 == 5'h17; // @[Replacement.scala 315:30]
  wire  set_touch_ways_1_55_valid = touch_ways_1_1_valid & touch_sets_1_0 == 5'h17; // @[Replacement.scala 315:30]
  wire  _T_134 = set_touch_ways_0_55_valid | set_touch_ways_1_55_valid; // @[package.scala 72:59]
  wire [2:0] state_vec_23_left_subtree_state_6 = state_vec_1_23[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_23_right_subtree_state_6 = state_vec_1_23[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_23_left_subtree_state_7 = state_vec_23_left_subtree_state_6[1]; // @[package.scala 154:13]
  wire  state_vec_23_right_subtree_state_7 = state_vec_23_left_subtree_state_6[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_23_T_52 = state_vec_0_set_left_older_7 ? state_vec_23_left_subtree_state_7 : _state_vec_0_T_51; // @[Replacement.scala 203:16]
  wire  _state_vec_23_T_56 = state_vec_0_set_left_older_7 ? _state_vec_0_T_51 : state_vec_23_right_subtree_state_7; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_23_T_57 = {state_vec_0_set_left_older_7,_state_vec_23_T_52,_state_vec_23_T_56}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_23_T_58 = state_vec_0_set_left_older_6 ? state_vec_23_left_subtree_state_6 : _state_vec_23_T_57; // @[Replacement.scala 203:16]
  wire  state_vec_23_left_subtree_state_8 = state_vec_23_right_subtree_state_6[1]; // @[package.scala 154:13]
  wire  state_vec_23_right_subtree_state_8 = state_vec_23_right_subtree_state_6[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_23_T_63 = state_vec_0_set_left_older_7 ? state_vec_23_left_subtree_state_8 : _state_vec_0_T_51; // @[Replacement.scala 203:16]
  wire  _state_vec_23_T_67 = state_vec_0_set_left_older_7 ? _state_vec_0_T_51 : state_vec_23_right_subtree_state_8; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_23_T_68 = {state_vec_0_set_left_older_7,_state_vec_23_T_63,_state_vec_23_T_67}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_23_T_69 = state_vec_0_set_left_older_6 ? _state_vec_23_T_68 : state_vec_23_right_subtree_state_6
    ; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_23_T_70 = {state_vec_0_set_left_older_6,_state_vec_23_T_58,_state_vec_23_T_69}; // @[Cat.scala 31:58]
  wire [6:0] _state_vec_23_T_71 = set_touch_ways_0_55_valid ? _state_vec_23_T_70 : state_vec_1_23; // @[Replacement.scala 22:56]
  wire [2:0] state_vec_23_left_subtree_state_9 = _state_vec_23_T_71[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_23_right_subtree_state_9 = _state_vec_23_T_71[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_23_left_subtree_state_10 = state_vec_23_left_subtree_state_9[1]; // @[package.scala 154:13]
  wire  state_vec_23_right_subtree_state_10 = state_vec_23_left_subtree_state_9[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_23_T_76 = state_vec_0_set_left_older_10 ? state_vec_23_left_subtree_state_10 : _state_vec_0_T_75; // @[Replacement.scala 203:16]
  wire  _state_vec_23_T_80 = state_vec_0_set_left_older_10 ? _state_vec_0_T_75 : state_vec_23_right_subtree_state_10; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_23_T_81 = {state_vec_0_set_left_older_10,_state_vec_23_T_76,_state_vec_23_T_80}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_23_T_82 = state_vec_0_set_left_older_9 ? state_vec_23_left_subtree_state_9 : _state_vec_23_T_81; // @[Replacement.scala 203:16]
  wire  state_vec_23_left_subtree_state_11 = state_vec_23_right_subtree_state_9[1]; // @[package.scala 154:13]
  wire  state_vec_23_right_subtree_state_11 = state_vec_23_right_subtree_state_9[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_23_T_87 = state_vec_0_set_left_older_10 ? state_vec_23_left_subtree_state_11 : _state_vec_0_T_75; // @[Replacement.scala 203:16]
  wire  _state_vec_23_T_91 = state_vec_0_set_left_older_10 ? _state_vec_0_T_75 : state_vec_23_right_subtree_state_11; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_23_T_92 = {state_vec_0_set_left_older_10,_state_vec_23_T_87,_state_vec_23_T_91}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_23_T_93 = state_vec_0_set_left_older_9 ? _state_vec_23_T_92 : state_vec_23_right_subtree_state_9
    ; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_23_T_94 = {state_vec_0_set_left_older_9,_state_vec_23_T_82,_state_vec_23_T_93}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_56_valid = touch_ways_1_0_valid & touch_sets_1_0 == 5'h18; // @[Replacement.scala 315:30]
  wire  set_touch_ways_1_56_valid = touch_ways_1_1_valid & touch_sets_1_0 == 5'h18; // @[Replacement.scala 315:30]
  wire  _T_135 = set_touch_ways_0_56_valid | set_touch_ways_1_56_valid; // @[package.scala 72:59]
  wire [2:0] state_vec_24_left_subtree_state_6 = state_vec_1_24[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_24_right_subtree_state_6 = state_vec_1_24[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_24_left_subtree_state_7 = state_vec_24_left_subtree_state_6[1]; // @[package.scala 154:13]
  wire  state_vec_24_right_subtree_state_7 = state_vec_24_left_subtree_state_6[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_24_T_52 = state_vec_0_set_left_older_7 ? state_vec_24_left_subtree_state_7 : _state_vec_0_T_51; // @[Replacement.scala 203:16]
  wire  _state_vec_24_T_56 = state_vec_0_set_left_older_7 ? _state_vec_0_T_51 : state_vec_24_right_subtree_state_7; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_24_T_57 = {state_vec_0_set_left_older_7,_state_vec_24_T_52,_state_vec_24_T_56}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_24_T_58 = state_vec_0_set_left_older_6 ? state_vec_24_left_subtree_state_6 : _state_vec_24_T_57; // @[Replacement.scala 203:16]
  wire  state_vec_24_left_subtree_state_8 = state_vec_24_right_subtree_state_6[1]; // @[package.scala 154:13]
  wire  state_vec_24_right_subtree_state_8 = state_vec_24_right_subtree_state_6[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_24_T_63 = state_vec_0_set_left_older_7 ? state_vec_24_left_subtree_state_8 : _state_vec_0_T_51; // @[Replacement.scala 203:16]
  wire  _state_vec_24_T_67 = state_vec_0_set_left_older_7 ? _state_vec_0_T_51 : state_vec_24_right_subtree_state_8; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_24_T_68 = {state_vec_0_set_left_older_7,_state_vec_24_T_63,_state_vec_24_T_67}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_24_T_69 = state_vec_0_set_left_older_6 ? _state_vec_24_T_68 : state_vec_24_right_subtree_state_6
    ; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_24_T_70 = {state_vec_0_set_left_older_6,_state_vec_24_T_58,_state_vec_24_T_69}; // @[Cat.scala 31:58]
  wire [6:0] _state_vec_24_T_71 = set_touch_ways_0_56_valid ? _state_vec_24_T_70 : state_vec_1_24; // @[Replacement.scala 22:56]
  wire [2:0] state_vec_24_left_subtree_state_9 = _state_vec_24_T_71[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_24_right_subtree_state_9 = _state_vec_24_T_71[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_24_left_subtree_state_10 = state_vec_24_left_subtree_state_9[1]; // @[package.scala 154:13]
  wire  state_vec_24_right_subtree_state_10 = state_vec_24_left_subtree_state_9[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_24_T_76 = state_vec_0_set_left_older_10 ? state_vec_24_left_subtree_state_10 : _state_vec_0_T_75; // @[Replacement.scala 203:16]
  wire  _state_vec_24_T_80 = state_vec_0_set_left_older_10 ? _state_vec_0_T_75 : state_vec_24_right_subtree_state_10; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_24_T_81 = {state_vec_0_set_left_older_10,_state_vec_24_T_76,_state_vec_24_T_80}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_24_T_82 = state_vec_0_set_left_older_9 ? state_vec_24_left_subtree_state_9 : _state_vec_24_T_81; // @[Replacement.scala 203:16]
  wire  state_vec_24_left_subtree_state_11 = state_vec_24_right_subtree_state_9[1]; // @[package.scala 154:13]
  wire  state_vec_24_right_subtree_state_11 = state_vec_24_right_subtree_state_9[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_24_T_87 = state_vec_0_set_left_older_10 ? state_vec_24_left_subtree_state_11 : _state_vec_0_T_75; // @[Replacement.scala 203:16]
  wire  _state_vec_24_T_91 = state_vec_0_set_left_older_10 ? _state_vec_0_T_75 : state_vec_24_right_subtree_state_11; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_24_T_92 = {state_vec_0_set_left_older_10,_state_vec_24_T_87,_state_vec_24_T_91}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_24_T_93 = state_vec_0_set_left_older_9 ? _state_vec_24_T_92 : state_vec_24_right_subtree_state_9
    ; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_24_T_94 = {state_vec_0_set_left_older_9,_state_vec_24_T_82,_state_vec_24_T_93}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_57_valid = touch_ways_1_0_valid & touch_sets_1_0 == 5'h19; // @[Replacement.scala 315:30]
  wire  set_touch_ways_1_57_valid = touch_ways_1_1_valid & touch_sets_1_0 == 5'h19; // @[Replacement.scala 315:30]
  wire  _T_136 = set_touch_ways_0_57_valid | set_touch_ways_1_57_valid; // @[package.scala 72:59]
  wire [2:0] state_vec_25_left_subtree_state_6 = state_vec_1_25[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_25_right_subtree_state_6 = state_vec_1_25[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_25_left_subtree_state_7 = state_vec_25_left_subtree_state_6[1]; // @[package.scala 154:13]
  wire  state_vec_25_right_subtree_state_7 = state_vec_25_left_subtree_state_6[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_25_T_52 = state_vec_0_set_left_older_7 ? state_vec_25_left_subtree_state_7 : _state_vec_0_T_51; // @[Replacement.scala 203:16]
  wire  _state_vec_25_T_56 = state_vec_0_set_left_older_7 ? _state_vec_0_T_51 : state_vec_25_right_subtree_state_7; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_25_T_57 = {state_vec_0_set_left_older_7,_state_vec_25_T_52,_state_vec_25_T_56}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_25_T_58 = state_vec_0_set_left_older_6 ? state_vec_25_left_subtree_state_6 : _state_vec_25_T_57; // @[Replacement.scala 203:16]
  wire  state_vec_25_left_subtree_state_8 = state_vec_25_right_subtree_state_6[1]; // @[package.scala 154:13]
  wire  state_vec_25_right_subtree_state_8 = state_vec_25_right_subtree_state_6[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_25_T_63 = state_vec_0_set_left_older_7 ? state_vec_25_left_subtree_state_8 : _state_vec_0_T_51; // @[Replacement.scala 203:16]
  wire  _state_vec_25_T_67 = state_vec_0_set_left_older_7 ? _state_vec_0_T_51 : state_vec_25_right_subtree_state_8; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_25_T_68 = {state_vec_0_set_left_older_7,_state_vec_25_T_63,_state_vec_25_T_67}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_25_T_69 = state_vec_0_set_left_older_6 ? _state_vec_25_T_68 : state_vec_25_right_subtree_state_6
    ; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_25_T_70 = {state_vec_0_set_left_older_6,_state_vec_25_T_58,_state_vec_25_T_69}; // @[Cat.scala 31:58]
  wire [6:0] _state_vec_25_T_71 = set_touch_ways_0_57_valid ? _state_vec_25_T_70 : state_vec_1_25; // @[Replacement.scala 22:56]
  wire [2:0] state_vec_25_left_subtree_state_9 = _state_vec_25_T_71[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_25_right_subtree_state_9 = _state_vec_25_T_71[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_25_left_subtree_state_10 = state_vec_25_left_subtree_state_9[1]; // @[package.scala 154:13]
  wire  state_vec_25_right_subtree_state_10 = state_vec_25_left_subtree_state_9[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_25_T_76 = state_vec_0_set_left_older_10 ? state_vec_25_left_subtree_state_10 : _state_vec_0_T_75; // @[Replacement.scala 203:16]
  wire  _state_vec_25_T_80 = state_vec_0_set_left_older_10 ? _state_vec_0_T_75 : state_vec_25_right_subtree_state_10; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_25_T_81 = {state_vec_0_set_left_older_10,_state_vec_25_T_76,_state_vec_25_T_80}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_25_T_82 = state_vec_0_set_left_older_9 ? state_vec_25_left_subtree_state_9 : _state_vec_25_T_81; // @[Replacement.scala 203:16]
  wire  state_vec_25_left_subtree_state_11 = state_vec_25_right_subtree_state_9[1]; // @[package.scala 154:13]
  wire  state_vec_25_right_subtree_state_11 = state_vec_25_right_subtree_state_9[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_25_T_87 = state_vec_0_set_left_older_10 ? state_vec_25_left_subtree_state_11 : _state_vec_0_T_75; // @[Replacement.scala 203:16]
  wire  _state_vec_25_T_91 = state_vec_0_set_left_older_10 ? _state_vec_0_T_75 : state_vec_25_right_subtree_state_11; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_25_T_92 = {state_vec_0_set_left_older_10,_state_vec_25_T_87,_state_vec_25_T_91}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_25_T_93 = state_vec_0_set_left_older_9 ? _state_vec_25_T_92 : state_vec_25_right_subtree_state_9
    ; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_25_T_94 = {state_vec_0_set_left_older_9,_state_vec_25_T_82,_state_vec_25_T_93}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_58_valid = touch_ways_1_0_valid & touch_sets_1_0 == 5'h1a; // @[Replacement.scala 315:30]
  wire  set_touch_ways_1_58_valid = touch_ways_1_1_valid & touch_sets_1_0 == 5'h1a; // @[Replacement.scala 315:30]
  wire  _T_137 = set_touch_ways_0_58_valid | set_touch_ways_1_58_valid; // @[package.scala 72:59]
  wire [2:0] state_vec_26_left_subtree_state_6 = state_vec_1_26[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_26_right_subtree_state_6 = state_vec_1_26[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_26_left_subtree_state_7 = state_vec_26_left_subtree_state_6[1]; // @[package.scala 154:13]
  wire  state_vec_26_right_subtree_state_7 = state_vec_26_left_subtree_state_6[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_26_T_52 = state_vec_0_set_left_older_7 ? state_vec_26_left_subtree_state_7 : _state_vec_0_T_51; // @[Replacement.scala 203:16]
  wire  _state_vec_26_T_56 = state_vec_0_set_left_older_7 ? _state_vec_0_T_51 : state_vec_26_right_subtree_state_7; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_26_T_57 = {state_vec_0_set_left_older_7,_state_vec_26_T_52,_state_vec_26_T_56}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_26_T_58 = state_vec_0_set_left_older_6 ? state_vec_26_left_subtree_state_6 : _state_vec_26_T_57; // @[Replacement.scala 203:16]
  wire  state_vec_26_left_subtree_state_8 = state_vec_26_right_subtree_state_6[1]; // @[package.scala 154:13]
  wire  state_vec_26_right_subtree_state_8 = state_vec_26_right_subtree_state_6[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_26_T_63 = state_vec_0_set_left_older_7 ? state_vec_26_left_subtree_state_8 : _state_vec_0_T_51; // @[Replacement.scala 203:16]
  wire  _state_vec_26_T_67 = state_vec_0_set_left_older_7 ? _state_vec_0_T_51 : state_vec_26_right_subtree_state_8; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_26_T_68 = {state_vec_0_set_left_older_7,_state_vec_26_T_63,_state_vec_26_T_67}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_26_T_69 = state_vec_0_set_left_older_6 ? _state_vec_26_T_68 : state_vec_26_right_subtree_state_6
    ; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_26_T_70 = {state_vec_0_set_left_older_6,_state_vec_26_T_58,_state_vec_26_T_69}; // @[Cat.scala 31:58]
  wire [6:0] _state_vec_26_T_71 = set_touch_ways_0_58_valid ? _state_vec_26_T_70 : state_vec_1_26; // @[Replacement.scala 22:56]
  wire [2:0] state_vec_26_left_subtree_state_9 = _state_vec_26_T_71[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_26_right_subtree_state_9 = _state_vec_26_T_71[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_26_left_subtree_state_10 = state_vec_26_left_subtree_state_9[1]; // @[package.scala 154:13]
  wire  state_vec_26_right_subtree_state_10 = state_vec_26_left_subtree_state_9[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_26_T_76 = state_vec_0_set_left_older_10 ? state_vec_26_left_subtree_state_10 : _state_vec_0_T_75; // @[Replacement.scala 203:16]
  wire  _state_vec_26_T_80 = state_vec_0_set_left_older_10 ? _state_vec_0_T_75 : state_vec_26_right_subtree_state_10; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_26_T_81 = {state_vec_0_set_left_older_10,_state_vec_26_T_76,_state_vec_26_T_80}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_26_T_82 = state_vec_0_set_left_older_9 ? state_vec_26_left_subtree_state_9 : _state_vec_26_T_81; // @[Replacement.scala 203:16]
  wire  state_vec_26_left_subtree_state_11 = state_vec_26_right_subtree_state_9[1]; // @[package.scala 154:13]
  wire  state_vec_26_right_subtree_state_11 = state_vec_26_right_subtree_state_9[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_26_T_87 = state_vec_0_set_left_older_10 ? state_vec_26_left_subtree_state_11 : _state_vec_0_T_75; // @[Replacement.scala 203:16]
  wire  _state_vec_26_T_91 = state_vec_0_set_left_older_10 ? _state_vec_0_T_75 : state_vec_26_right_subtree_state_11; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_26_T_92 = {state_vec_0_set_left_older_10,_state_vec_26_T_87,_state_vec_26_T_91}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_26_T_93 = state_vec_0_set_left_older_9 ? _state_vec_26_T_92 : state_vec_26_right_subtree_state_9
    ; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_26_T_94 = {state_vec_0_set_left_older_9,_state_vec_26_T_82,_state_vec_26_T_93}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_59_valid = touch_ways_1_0_valid & touch_sets_1_0 == 5'h1b; // @[Replacement.scala 315:30]
  wire  set_touch_ways_1_59_valid = touch_ways_1_1_valid & touch_sets_1_0 == 5'h1b; // @[Replacement.scala 315:30]
  wire  _T_138 = set_touch_ways_0_59_valid | set_touch_ways_1_59_valid; // @[package.scala 72:59]
  wire [2:0] state_vec_27_left_subtree_state_6 = state_vec_1_27[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_27_right_subtree_state_6 = state_vec_1_27[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_27_left_subtree_state_7 = state_vec_27_left_subtree_state_6[1]; // @[package.scala 154:13]
  wire  state_vec_27_right_subtree_state_7 = state_vec_27_left_subtree_state_6[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_27_T_52 = state_vec_0_set_left_older_7 ? state_vec_27_left_subtree_state_7 : _state_vec_0_T_51; // @[Replacement.scala 203:16]
  wire  _state_vec_27_T_56 = state_vec_0_set_left_older_7 ? _state_vec_0_T_51 : state_vec_27_right_subtree_state_7; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_27_T_57 = {state_vec_0_set_left_older_7,_state_vec_27_T_52,_state_vec_27_T_56}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_27_T_58 = state_vec_0_set_left_older_6 ? state_vec_27_left_subtree_state_6 : _state_vec_27_T_57; // @[Replacement.scala 203:16]
  wire  state_vec_27_left_subtree_state_8 = state_vec_27_right_subtree_state_6[1]; // @[package.scala 154:13]
  wire  state_vec_27_right_subtree_state_8 = state_vec_27_right_subtree_state_6[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_27_T_63 = state_vec_0_set_left_older_7 ? state_vec_27_left_subtree_state_8 : _state_vec_0_T_51; // @[Replacement.scala 203:16]
  wire  _state_vec_27_T_67 = state_vec_0_set_left_older_7 ? _state_vec_0_T_51 : state_vec_27_right_subtree_state_8; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_27_T_68 = {state_vec_0_set_left_older_7,_state_vec_27_T_63,_state_vec_27_T_67}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_27_T_69 = state_vec_0_set_left_older_6 ? _state_vec_27_T_68 : state_vec_27_right_subtree_state_6
    ; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_27_T_70 = {state_vec_0_set_left_older_6,_state_vec_27_T_58,_state_vec_27_T_69}; // @[Cat.scala 31:58]
  wire [6:0] _state_vec_27_T_71 = set_touch_ways_0_59_valid ? _state_vec_27_T_70 : state_vec_1_27; // @[Replacement.scala 22:56]
  wire [2:0] state_vec_27_left_subtree_state_9 = _state_vec_27_T_71[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_27_right_subtree_state_9 = _state_vec_27_T_71[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_27_left_subtree_state_10 = state_vec_27_left_subtree_state_9[1]; // @[package.scala 154:13]
  wire  state_vec_27_right_subtree_state_10 = state_vec_27_left_subtree_state_9[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_27_T_76 = state_vec_0_set_left_older_10 ? state_vec_27_left_subtree_state_10 : _state_vec_0_T_75; // @[Replacement.scala 203:16]
  wire  _state_vec_27_T_80 = state_vec_0_set_left_older_10 ? _state_vec_0_T_75 : state_vec_27_right_subtree_state_10; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_27_T_81 = {state_vec_0_set_left_older_10,_state_vec_27_T_76,_state_vec_27_T_80}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_27_T_82 = state_vec_0_set_left_older_9 ? state_vec_27_left_subtree_state_9 : _state_vec_27_T_81; // @[Replacement.scala 203:16]
  wire  state_vec_27_left_subtree_state_11 = state_vec_27_right_subtree_state_9[1]; // @[package.scala 154:13]
  wire  state_vec_27_right_subtree_state_11 = state_vec_27_right_subtree_state_9[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_27_T_87 = state_vec_0_set_left_older_10 ? state_vec_27_left_subtree_state_11 : _state_vec_0_T_75; // @[Replacement.scala 203:16]
  wire  _state_vec_27_T_91 = state_vec_0_set_left_older_10 ? _state_vec_0_T_75 : state_vec_27_right_subtree_state_11; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_27_T_92 = {state_vec_0_set_left_older_10,_state_vec_27_T_87,_state_vec_27_T_91}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_27_T_93 = state_vec_0_set_left_older_9 ? _state_vec_27_T_92 : state_vec_27_right_subtree_state_9
    ; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_27_T_94 = {state_vec_0_set_left_older_9,_state_vec_27_T_82,_state_vec_27_T_93}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_60_valid = touch_ways_1_0_valid & touch_sets_1_0 == 5'h1c; // @[Replacement.scala 315:30]
  wire  set_touch_ways_1_60_valid = touch_ways_1_1_valid & touch_sets_1_0 == 5'h1c; // @[Replacement.scala 315:30]
  wire  _T_139 = set_touch_ways_0_60_valid | set_touch_ways_1_60_valid; // @[package.scala 72:59]
  wire [2:0] state_vec_28_left_subtree_state_6 = state_vec_1_28[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_28_right_subtree_state_6 = state_vec_1_28[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_28_left_subtree_state_7 = state_vec_28_left_subtree_state_6[1]; // @[package.scala 154:13]
  wire  state_vec_28_right_subtree_state_7 = state_vec_28_left_subtree_state_6[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_28_T_52 = state_vec_0_set_left_older_7 ? state_vec_28_left_subtree_state_7 : _state_vec_0_T_51; // @[Replacement.scala 203:16]
  wire  _state_vec_28_T_56 = state_vec_0_set_left_older_7 ? _state_vec_0_T_51 : state_vec_28_right_subtree_state_7; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_28_T_57 = {state_vec_0_set_left_older_7,_state_vec_28_T_52,_state_vec_28_T_56}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_28_T_58 = state_vec_0_set_left_older_6 ? state_vec_28_left_subtree_state_6 : _state_vec_28_T_57; // @[Replacement.scala 203:16]
  wire  state_vec_28_left_subtree_state_8 = state_vec_28_right_subtree_state_6[1]; // @[package.scala 154:13]
  wire  state_vec_28_right_subtree_state_8 = state_vec_28_right_subtree_state_6[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_28_T_63 = state_vec_0_set_left_older_7 ? state_vec_28_left_subtree_state_8 : _state_vec_0_T_51; // @[Replacement.scala 203:16]
  wire  _state_vec_28_T_67 = state_vec_0_set_left_older_7 ? _state_vec_0_T_51 : state_vec_28_right_subtree_state_8; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_28_T_68 = {state_vec_0_set_left_older_7,_state_vec_28_T_63,_state_vec_28_T_67}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_28_T_69 = state_vec_0_set_left_older_6 ? _state_vec_28_T_68 : state_vec_28_right_subtree_state_6
    ; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_28_T_70 = {state_vec_0_set_left_older_6,_state_vec_28_T_58,_state_vec_28_T_69}; // @[Cat.scala 31:58]
  wire [6:0] _state_vec_28_T_71 = set_touch_ways_0_60_valid ? _state_vec_28_T_70 : state_vec_1_28; // @[Replacement.scala 22:56]
  wire [2:0] state_vec_28_left_subtree_state_9 = _state_vec_28_T_71[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_28_right_subtree_state_9 = _state_vec_28_T_71[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_28_left_subtree_state_10 = state_vec_28_left_subtree_state_9[1]; // @[package.scala 154:13]
  wire  state_vec_28_right_subtree_state_10 = state_vec_28_left_subtree_state_9[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_28_T_76 = state_vec_0_set_left_older_10 ? state_vec_28_left_subtree_state_10 : _state_vec_0_T_75; // @[Replacement.scala 203:16]
  wire  _state_vec_28_T_80 = state_vec_0_set_left_older_10 ? _state_vec_0_T_75 : state_vec_28_right_subtree_state_10; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_28_T_81 = {state_vec_0_set_left_older_10,_state_vec_28_T_76,_state_vec_28_T_80}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_28_T_82 = state_vec_0_set_left_older_9 ? state_vec_28_left_subtree_state_9 : _state_vec_28_T_81; // @[Replacement.scala 203:16]
  wire  state_vec_28_left_subtree_state_11 = state_vec_28_right_subtree_state_9[1]; // @[package.scala 154:13]
  wire  state_vec_28_right_subtree_state_11 = state_vec_28_right_subtree_state_9[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_28_T_87 = state_vec_0_set_left_older_10 ? state_vec_28_left_subtree_state_11 : _state_vec_0_T_75; // @[Replacement.scala 203:16]
  wire  _state_vec_28_T_91 = state_vec_0_set_left_older_10 ? _state_vec_0_T_75 : state_vec_28_right_subtree_state_11; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_28_T_92 = {state_vec_0_set_left_older_10,_state_vec_28_T_87,_state_vec_28_T_91}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_28_T_93 = state_vec_0_set_left_older_9 ? _state_vec_28_T_92 : state_vec_28_right_subtree_state_9
    ; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_28_T_94 = {state_vec_0_set_left_older_9,_state_vec_28_T_82,_state_vec_28_T_93}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_61_valid = touch_ways_1_0_valid & touch_sets_1_0 == 5'h1d; // @[Replacement.scala 315:30]
  wire  set_touch_ways_1_61_valid = touch_ways_1_1_valid & touch_sets_1_0 == 5'h1d; // @[Replacement.scala 315:30]
  wire  _T_140 = set_touch_ways_0_61_valid | set_touch_ways_1_61_valid; // @[package.scala 72:59]
  wire [2:0] state_vec_29_left_subtree_state_6 = state_vec_1_29[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_29_right_subtree_state_6 = state_vec_1_29[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_29_left_subtree_state_7 = state_vec_29_left_subtree_state_6[1]; // @[package.scala 154:13]
  wire  state_vec_29_right_subtree_state_7 = state_vec_29_left_subtree_state_6[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_29_T_52 = state_vec_0_set_left_older_7 ? state_vec_29_left_subtree_state_7 : _state_vec_0_T_51; // @[Replacement.scala 203:16]
  wire  _state_vec_29_T_56 = state_vec_0_set_left_older_7 ? _state_vec_0_T_51 : state_vec_29_right_subtree_state_7; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_29_T_57 = {state_vec_0_set_left_older_7,_state_vec_29_T_52,_state_vec_29_T_56}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_29_T_58 = state_vec_0_set_left_older_6 ? state_vec_29_left_subtree_state_6 : _state_vec_29_T_57; // @[Replacement.scala 203:16]
  wire  state_vec_29_left_subtree_state_8 = state_vec_29_right_subtree_state_6[1]; // @[package.scala 154:13]
  wire  state_vec_29_right_subtree_state_8 = state_vec_29_right_subtree_state_6[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_29_T_63 = state_vec_0_set_left_older_7 ? state_vec_29_left_subtree_state_8 : _state_vec_0_T_51; // @[Replacement.scala 203:16]
  wire  _state_vec_29_T_67 = state_vec_0_set_left_older_7 ? _state_vec_0_T_51 : state_vec_29_right_subtree_state_8; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_29_T_68 = {state_vec_0_set_left_older_7,_state_vec_29_T_63,_state_vec_29_T_67}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_29_T_69 = state_vec_0_set_left_older_6 ? _state_vec_29_T_68 : state_vec_29_right_subtree_state_6
    ; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_29_T_70 = {state_vec_0_set_left_older_6,_state_vec_29_T_58,_state_vec_29_T_69}; // @[Cat.scala 31:58]
  wire [6:0] _state_vec_29_T_71 = set_touch_ways_0_61_valid ? _state_vec_29_T_70 : state_vec_1_29; // @[Replacement.scala 22:56]
  wire [2:0] state_vec_29_left_subtree_state_9 = _state_vec_29_T_71[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_29_right_subtree_state_9 = _state_vec_29_T_71[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_29_left_subtree_state_10 = state_vec_29_left_subtree_state_9[1]; // @[package.scala 154:13]
  wire  state_vec_29_right_subtree_state_10 = state_vec_29_left_subtree_state_9[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_29_T_76 = state_vec_0_set_left_older_10 ? state_vec_29_left_subtree_state_10 : _state_vec_0_T_75; // @[Replacement.scala 203:16]
  wire  _state_vec_29_T_80 = state_vec_0_set_left_older_10 ? _state_vec_0_T_75 : state_vec_29_right_subtree_state_10; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_29_T_81 = {state_vec_0_set_left_older_10,_state_vec_29_T_76,_state_vec_29_T_80}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_29_T_82 = state_vec_0_set_left_older_9 ? state_vec_29_left_subtree_state_9 : _state_vec_29_T_81; // @[Replacement.scala 203:16]
  wire  state_vec_29_left_subtree_state_11 = state_vec_29_right_subtree_state_9[1]; // @[package.scala 154:13]
  wire  state_vec_29_right_subtree_state_11 = state_vec_29_right_subtree_state_9[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_29_T_87 = state_vec_0_set_left_older_10 ? state_vec_29_left_subtree_state_11 : _state_vec_0_T_75; // @[Replacement.scala 203:16]
  wire  _state_vec_29_T_91 = state_vec_0_set_left_older_10 ? _state_vec_0_T_75 : state_vec_29_right_subtree_state_11; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_29_T_92 = {state_vec_0_set_left_older_10,_state_vec_29_T_87,_state_vec_29_T_91}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_29_T_93 = state_vec_0_set_left_older_9 ? _state_vec_29_T_92 : state_vec_29_right_subtree_state_9
    ; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_29_T_94 = {state_vec_0_set_left_older_9,_state_vec_29_T_82,_state_vec_29_T_93}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_62_valid = touch_ways_1_0_valid & touch_sets_1_0 == 5'h1e; // @[Replacement.scala 315:30]
  wire  set_touch_ways_1_62_valid = touch_ways_1_1_valid & touch_sets_1_0 == 5'h1e; // @[Replacement.scala 315:30]
  wire  _T_141 = set_touch_ways_0_62_valid | set_touch_ways_1_62_valid; // @[package.scala 72:59]
  wire [2:0] state_vec_30_left_subtree_state_6 = state_vec_1_30[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_30_right_subtree_state_6 = state_vec_1_30[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_30_left_subtree_state_7 = state_vec_30_left_subtree_state_6[1]; // @[package.scala 154:13]
  wire  state_vec_30_right_subtree_state_7 = state_vec_30_left_subtree_state_6[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_30_T_52 = state_vec_0_set_left_older_7 ? state_vec_30_left_subtree_state_7 : _state_vec_0_T_51; // @[Replacement.scala 203:16]
  wire  _state_vec_30_T_56 = state_vec_0_set_left_older_7 ? _state_vec_0_T_51 : state_vec_30_right_subtree_state_7; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_30_T_57 = {state_vec_0_set_left_older_7,_state_vec_30_T_52,_state_vec_30_T_56}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_30_T_58 = state_vec_0_set_left_older_6 ? state_vec_30_left_subtree_state_6 : _state_vec_30_T_57; // @[Replacement.scala 203:16]
  wire  state_vec_30_left_subtree_state_8 = state_vec_30_right_subtree_state_6[1]; // @[package.scala 154:13]
  wire  state_vec_30_right_subtree_state_8 = state_vec_30_right_subtree_state_6[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_30_T_63 = state_vec_0_set_left_older_7 ? state_vec_30_left_subtree_state_8 : _state_vec_0_T_51; // @[Replacement.scala 203:16]
  wire  _state_vec_30_T_67 = state_vec_0_set_left_older_7 ? _state_vec_0_T_51 : state_vec_30_right_subtree_state_8; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_30_T_68 = {state_vec_0_set_left_older_7,_state_vec_30_T_63,_state_vec_30_T_67}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_30_T_69 = state_vec_0_set_left_older_6 ? _state_vec_30_T_68 : state_vec_30_right_subtree_state_6
    ; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_30_T_70 = {state_vec_0_set_left_older_6,_state_vec_30_T_58,_state_vec_30_T_69}; // @[Cat.scala 31:58]
  wire [6:0] _state_vec_30_T_71 = set_touch_ways_0_62_valid ? _state_vec_30_T_70 : state_vec_1_30; // @[Replacement.scala 22:56]
  wire [2:0] state_vec_30_left_subtree_state_9 = _state_vec_30_T_71[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_30_right_subtree_state_9 = _state_vec_30_T_71[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_30_left_subtree_state_10 = state_vec_30_left_subtree_state_9[1]; // @[package.scala 154:13]
  wire  state_vec_30_right_subtree_state_10 = state_vec_30_left_subtree_state_9[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_30_T_76 = state_vec_0_set_left_older_10 ? state_vec_30_left_subtree_state_10 : _state_vec_0_T_75; // @[Replacement.scala 203:16]
  wire  _state_vec_30_T_80 = state_vec_0_set_left_older_10 ? _state_vec_0_T_75 : state_vec_30_right_subtree_state_10; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_30_T_81 = {state_vec_0_set_left_older_10,_state_vec_30_T_76,_state_vec_30_T_80}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_30_T_82 = state_vec_0_set_left_older_9 ? state_vec_30_left_subtree_state_9 : _state_vec_30_T_81; // @[Replacement.scala 203:16]
  wire  state_vec_30_left_subtree_state_11 = state_vec_30_right_subtree_state_9[1]; // @[package.scala 154:13]
  wire  state_vec_30_right_subtree_state_11 = state_vec_30_right_subtree_state_9[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_30_T_87 = state_vec_0_set_left_older_10 ? state_vec_30_left_subtree_state_11 : _state_vec_0_T_75; // @[Replacement.scala 203:16]
  wire  _state_vec_30_T_91 = state_vec_0_set_left_older_10 ? _state_vec_0_T_75 : state_vec_30_right_subtree_state_11; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_30_T_92 = {state_vec_0_set_left_older_10,_state_vec_30_T_87,_state_vec_30_T_91}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_30_T_93 = state_vec_0_set_left_older_9 ? _state_vec_30_T_92 : state_vec_30_right_subtree_state_9
    ; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_30_T_94 = {state_vec_0_set_left_older_9,_state_vec_30_T_82,_state_vec_30_T_93}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_63_valid = touch_ways_1_0_valid & touch_sets_1_0 == 5'h1f; // @[Replacement.scala 315:30]
  wire  set_touch_ways_1_63_valid = touch_ways_1_1_valid & touch_sets_1_0 == 5'h1f; // @[Replacement.scala 315:30]
  wire  _T_142 = set_touch_ways_0_63_valid | set_touch_ways_1_63_valid; // @[package.scala 72:59]
  wire [2:0] state_vec_31_left_subtree_state_6 = state_vec_1_31[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_31_right_subtree_state_6 = state_vec_1_31[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_31_left_subtree_state_7 = state_vec_31_left_subtree_state_6[1]; // @[package.scala 154:13]
  wire  state_vec_31_right_subtree_state_7 = state_vec_31_left_subtree_state_6[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_31_T_52 = state_vec_0_set_left_older_7 ? state_vec_31_left_subtree_state_7 : _state_vec_0_T_51; // @[Replacement.scala 203:16]
  wire  _state_vec_31_T_56 = state_vec_0_set_left_older_7 ? _state_vec_0_T_51 : state_vec_31_right_subtree_state_7; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_31_T_57 = {state_vec_0_set_left_older_7,_state_vec_31_T_52,_state_vec_31_T_56}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_31_T_58 = state_vec_0_set_left_older_6 ? state_vec_31_left_subtree_state_6 : _state_vec_31_T_57; // @[Replacement.scala 203:16]
  wire  state_vec_31_left_subtree_state_8 = state_vec_31_right_subtree_state_6[1]; // @[package.scala 154:13]
  wire  state_vec_31_right_subtree_state_8 = state_vec_31_right_subtree_state_6[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_31_T_63 = state_vec_0_set_left_older_7 ? state_vec_31_left_subtree_state_8 : _state_vec_0_T_51; // @[Replacement.scala 203:16]
  wire  _state_vec_31_T_67 = state_vec_0_set_left_older_7 ? _state_vec_0_T_51 : state_vec_31_right_subtree_state_8; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_31_T_68 = {state_vec_0_set_left_older_7,_state_vec_31_T_63,_state_vec_31_T_67}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_31_T_69 = state_vec_0_set_left_older_6 ? _state_vec_31_T_68 : state_vec_31_right_subtree_state_6
    ; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_31_T_70 = {state_vec_0_set_left_older_6,_state_vec_31_T_58,_state_vec_31_T_69}; // @[Cat.scala 31:58]
  wire [6:0] _state_vec_31_T_71 = set_touch_ways_0_63_valid ? _state_vec_31_T_70 : state_vec_1_31; // @[Replacement.scala 22:56]
  wire [2:0] state_vec_31_left_subtree_state_9 = _state_vec_31_T_71[5:3]; // @[package.scala 154:13]
  wire [2:0] state_vec_31_right_subtree_state_9 = _state_vec_31_T_71[2:0]; // @[Replacement.scala 198:38]
  wire  state_vec_31_left_subtree_state_10 = state_vec_31_left_subtree_state_9[1]; // @[package.scala 154:13]
  wire  state_vec_31_right_subtree_state_10 = state_vec_31_left_subtree_state_9[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_31_T_76 = state_vec_0_set_left_older_10 ? state_vec_31_left_subtree_state_10 : _state_vec_0_T_75; // @[Replacement.scala 203:16]
  wire  _state_vec_31_T_80 = state_vec_0_set_left_older_10 ? _state_vec_0_T_75 : state_vec_31_right_subtree_state_10; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_31_T_81 = {state_vec_0_set_left_older_10,_state_vec_31_T_76,_state_vec_31_T_80}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_31_T_82 = state_vec_0_set_left_older_9 ? state_vec_31_left_subtree_state_9 : _state_vec_31_T_81; // @[Replacement.scala 203:16]
  wire  state_vec_31_left_subtree_state_11 = state_vec_31_right_subtree_state_9[1]; // @[package.scala 154:13]
  wire  state_vec_31_right_subtree_state_11 = state_vec_31_right_subtree_state_9[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_31_T_87 = state_vec_0_set_left_older_10 ? state_vec_31_left_subtree_state_11 : _state_vec_0_T_75; // @[Replacement.scala 203:16]
  wire  _state_vec_31_T_91 = state_vec_0_set_left_older_10 ? _state_vec_0_T_75 : state_vec_31_right_subtree_state_11; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_31_T_92 = {state_vec_0_set_left_older_10,_state_vec_31_T_87,_state_vec_31_T_91}; // @[Cat.scala 31:58]
  wire [2:0] _state_vec_31_T_93 = state_vec_0_set_left_older_9 ? _state_vec_31_T_92 : state_vec_31_right_subtree_state_9
    ; // @[Replacement.scala 206:16]
  wire [6:0] _state_vec_31_T_94 = {state_vec_0_set_left_older_9,_state_vec_31_T_82,_state_vec_31_T_93}; // @[Cat.scala 31:58]
  wire  _GEN_235 = _s2_ready_T_2 ? 1'h0 : s2_valid; // @[ICache.scala 101:{43,51} 98:25]
  reg [35:0] s2_req_paddr_0; // @[Reg.scala 16:16]
  reg [35:0] s2_req_paddr_1; // @[Reg.scala 16:16]
  reg [38:0] s2_req_vaddr_0; // @[Reg.scala 16:16]
  reg [38:0] s2_req_vaddr_1; // @[Reg.scala 16:16]
  reg  s2_meta_errors_0_0; // @[Reg.scala 16:16]
  reg  s2_meta_errors_0_1; // @[Reg.scala 16:16]
  reg  s2_meta_errors_0_2; // @[Reg.scala 16:16]
  reg  s2_meta_errors_0_3; // @[Reg.scala 16:16]
  reg  s2_meta_errors_0_4; // @[Reg.scala 16:16]
  reg  s2_meta_errors_0_5; // @[Reg.scala 16:16]
  reg  s2_meta_errors_0_6; // @[Reg.scala 16:16]
  reg  s2_meta_errors_0_7; // @[Reg.scala 16:16]
  reg  s2_meta_errors_1_0; // @[Reg.scala 16:16]
  reg  s2_meta_errors_1_1; // @[Reg.scala 16:16]
  reg  s2_meta_errors_1_2; // @[Reg.scala 16:16]
  reg  s2_meta_errors_1_3; // @[Reg.scala 16:16]
  reg  s2_meta_errors_1_4; // @[Reg.scala 16:16]
  reg  s2_meta_errors_1_5; // @[Reg.scala 16:16]
  reg  s2_meta_errors_1_6; // @[Reg.scala 16:16]
  reg  s2_meta_errors_1_7; // @[Reg.scala 16:16]
  reg [31:0] s2_data_errorBits_0_0; // @[Reg.scala 16:16]
  reg [31:0] s2_data_errorBits_0_1; // @[Reg.scala 16:16]
  reg [31:0] s2_data_errorBits_0_2; // @[Reg.scala 16:16]
  reg [31:0] s2_data_errorBits_0_3; // @[Reg.scala 16:16]
  reg [31:0] s2_data_errorBits_0_4; // @[Reg.scala 16:16]
  reg [31:0] s2_data_errorBits_0_5; // @[Reg.scala 16:16]
  reg [31:0] s2_data_errorBits_0_6; // @[Reg.scala 16:16]
  reg [31:0] s2_data_errorBits_0_7; // @[Reg.scala 16:16]
  reg [31:0] s2_data_errorBits_1_0; // @[Reg.scala 16:16]
  reg [31:0] s2_data_errorBits_1_1; // @[Reg.scala 16:16]
  reg [31:0] s2_data_errorBits_1_2; // @[Reg.scala 16:16]
  reg [31:0] s2_data_errorBits_1_3; // @[Reg.scala 16:16]
  reg [31:0] s2_data_errorBits_1_4; // @[Reg.scala 16:16]
  reg [31:0] s2_data_errorBits_1_5; // @[Reg.scala 16:16]
  reg [31:0] s2_data_errorBits_1_6; // @[Reg.scala 16:16]
  reg [31:0] s2_data_errorBits_1_7; // @[Reg.scala 16:16]
  reg [511:0] s2_data_cacheline_0_0; // @[Reg.scala 16:16]
  reg [511:0] s2_data_cacheline_0_1; // @[Reg.scala 16:16]
  reg [511:0] s2_data_cacheline_0_2; // @[Reg.scala 16:16]
  reg [511:0] s2_data_cacheline_0_3; // @[Reg.scala 16:16]
  reg [511:0] s2_data_cacheline_0_4; // @[Reg.scala 16:16]
  reg [511:0] s2_data_cacheline_0_5; // @[Reg.scala 16:16]
  reg [511:0] s2_data_cacheline_0_6; // @[Reg.scala 16:16]
  reg [511:0] s2_data_cacheline_0_7; // @[Reg.scala 16:16]
  reg [511:0] s2_data_cacheline_1_0; // @[Reg.scala 16:16]
  reg [511:0] s2_data_cacheline_1_1; // @[Reg.scala 16:16]
  reg [511:0] s2_data_cacheline_1_2; // @[Reg.scala 16:16]
  reg [511:0] s2_data_cacheline_1_3; // @[Reg.scala 16:16]
  reg [511:0] s2_data_cacheline_1_4; // @[Reg.scala 16:16]
  reg [511:0] s2_data_cacheline_1_5; // @[Reg.scala 16:16]
  reg [511:0] s2_data_cacheline_1_6; // @[Reg.scala 16:16]
  reg [511:0] s2_data_cacheline_1_7; // @[Reg.scala 16:16]
  wire [4095:0] _read_datas_T = {s2_data_cacheline_0_7,s2_data_cacheline_0_6,s2_data_cacheline_0_5,s2_data_cacheline_0_4
    ,s2_data_cacheline_0_3,s2_data_cacheline_0_2,s2_data_cacheline_0_1,s2_data_cacheline_0_0}; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__0_0 = _read_datas_T[15:0]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__0_1 = _read_datas_T[31:16]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__0_2 = _read_datas_T[47:32]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__0_3 = _read_datas_T[63:48]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__0_4 = _read_datas_T[79:64]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__0_5 = _read_datas_T[95:80]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__0_6 = _read_datas_T[111:96]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__0_7 = _read_datas_T[127:112]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__0_8 = _read_datas_T[143:128]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__0_9 = _read_datas_T[159:144]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__0_10 = _read_datas_T[175:160]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__0_11 = _read_datas_T[191:176]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__0_12 = _read_datas_T[207:192]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__0_13 = _read_datas_T[223:208]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__0_14 = _read_datas_T[239:224]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__0_15 = _read_datas_T[255:240]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__0_16 = _read_datas_T[271:256]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__0_17 = _read_datas_T[287:272]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__0_18 = _read_datas_T[303:288]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__0_19 = _read_datas_T[319:304]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__0_20 = _read_datas_T[335:320]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__0_21 = _read_datas_T[351:336]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__0_22 = _read_datas_T[367:352]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__0_23 = _read_datas_T[383:368]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__0_24 = _read_datas_T[399:384]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__0_25 = _read_datas_T[415:400]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__0_26 = _read_datas_T[431:416]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__0_27 = _read_datas_T[447:432]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__0_28 = _read_datas_T[463:448]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__0_29 = _read_datas_T[479:464]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__0_30 = _read_datas_T[495:480]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__0_31 = _read_datas_T[511:496]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__1_0 = _read_datas_T[527:512]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__1_1 = _read_datas_T[543:528]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__1_2 = _read_datas_T[559:544]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__1_3 = _read_datas_T[575:560]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__1_4 = _read_datas_T[591:576]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__1_5 = _read_datas_T[607:592]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__1_6 = _read_datas_T[623:608]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__1_7 = _read_datas_T[639:624]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__1_8 = _read_datas_T[655:640]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__1_9 = _read_datas_T[671:656]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__1_10 = _read_datas_T[687:672]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__1_11 = _read_datas_T[703:688]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__1_12 = _read_datas_T[719:704]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__1_13 = _read_datas_T[735:720]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__1_14 = _read_datas_T[751:736]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__1_15 = _read_datas_T[767:752]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__1_16 = _read_datas_T[783:768]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__1_17 = _read_datas_T[799:784]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__1_18 = _read_datas_T[815:800]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__1_19 = _read_datas_T[831:816]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__1_20 = _read_datas_T[847:832]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__1_21 = _read_datas_T[863:848]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__1_22 = _read_datas_T[879:864]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__1_23 = _read_datas_T[895:880]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__1_24 = _read_datas_T[911:896]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__1_25 = _read_datas_T[927:912]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__1_26 = _read_datas_T[943:928]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__1_27 = _read_datas_T[959:944]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__1_28 = _read_datas_T[975:960]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__1_29 = _read_datas_T[991:976]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__1_30 = _read_datas_T[1007:992]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__1_31 = _read_datas_T[1023:1008]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__2_0 = _read_datas_T[1039:1024]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__2_1 = _read_datas_T[1055:1040]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__2_2 = _read_datas_T[1071:1056]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__2_3 = _read_datas_T[1087:1072]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__2_4 = _read_datas_T[1103:1088]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__2_5 = _read_datas_T[1119:1104]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__2_6 = _read_datas_T[1135:1120]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__2_7 = _read_datas_T[1151:1136]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__2_8 = _read_datas_T[1167:1152]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__2_9 = _read_datas_T[1183:1168]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__2_10 = _read_datas_T[1199:1184]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__2_11 = _read_datas_T[1215:1200]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__2_12 = _read_datas_T[1231:1216]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__2_13 = _read_datas_T[1247:1232]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__2_14 = _read_datas_T[1263:1248]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__2_15 = _read_datas_T[1279:1264]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__2_16 = _read_datas_T[1295:1280]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__2_17 = _read_datas_T[1311:1296]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__2_18 = _read_datas_T[1327:1312]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__2_19 = _read_datas_T[1343:1328]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__2_20 = _read_datas_T[1359:1344]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__2_21 = _read_datas_T[1375:1360]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__2_22 = _read_datas_T[1391:1376]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__2_23 = _read_datas_T[1407:1392]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__2_24 = _read_datas_T[1423:1408]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__2_25 = _read_datas_T[1439:1424]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__2_26 = _read_datas_T[1455:1440]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__2_27 = _read_datas_T[1471:1456]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__2_28 = _read_datas_T[1487:1472]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__2_29 = _read_datas_T[1503:1488]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__2_30 = _read_datas_T[1519:1504]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__2_31 = _read_datas_T[1535:1520]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__3_0 = _read_datas_T[1551:1536]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__3_1 = _read_datas_T[1567:1552]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__3_2 = _read_datas_T[1583:1568]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__3_3 = _read_datas_T[1599:1584]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__3_4 = _read_datas_T[1615:1600]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__3_5 = _read_datas_T[1631:1616]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__3_6 = _read_datas_T[1647:1632]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__3_7 = _read_datas_T[1663:1648]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__3_8 = _read_datas_T[1679:1664]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__3_9 = _read_datas_T[1695:1680]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__3_10 = _read_datas_T[1711:1696]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__3_11 = _read_datas_T[1727:1712]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__3_12 = _read_datas_T[1743:1728]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__3_13 = _read_datas_T[1759:1744]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__3_14 = _read_datas_T[1775:1760]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__3_15 = _read_datas_T[1791:1776]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__3_16 = _read_datas_T[1807:1792]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__3_17 = _read_datas_T[1823:1808]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__3_18 = _read_datas_T[1839:1824]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__3_19 = _read_datas_T[1855:1840]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__3_20 = _read_datas_T[1871:1856]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__3_21 = _read_datas_T[1887:1872]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__3_22 = _read_datas_T[1903:1888]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__3_23 = _read_datas_T[1919:1904]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__3_24 = _read_datas_T[1935:1920]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__3_25 = _read_datas_T[1951:1936]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__3_26 = _read_datas_T[1967:1952]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__3_27 = _read_datas_T[1983:1968]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__3_28 = _read_datas_T[1999:1984]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__3_29 = _read_datas_T[2015:2000]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__3_30 = _read_datas_T[2031:2016]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__3_31 = _read_datas_T[2047:2032]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__4_0 = _read_datas_T[2063:2048]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__4_1 = _read_datas_T[2079:2064]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__4_2 = _read_datas_T[2095:2080]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__4_3 = _read_datas_T[2111:2096]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__4_4 = _read_datas_T[2127:2112]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__4_5 = _read_datas_T[2143:2128]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__4_6 = _read_datas_T[2159:2144]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__4_7 = _read_datas_T[2175:2160]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__4_8 = _read_datas_T[2191:2176]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__4_9 = _read_datas_T[2207:2192]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__4_10 = _read_datas_T[2223:2208]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__4_11 = _read_datas_T[2239:2224]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__4_12 = _read_datas_T[2255:2240]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__4_13 = _read_datas_T[2271:2256]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__4_14 = _read_datas_T[2287:2272]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__4_15 = _read_datas_T[2303:2288]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__4_16 = _read_datas_T[2319:2304]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__4_17 = _read_datas_T[2335:2320]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__4_18 = _read_datas_T[2351:2336]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__4_19 = _read_datas_T[2367:2352]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__4_20 = _read_datas_T[2383:2368]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__4_21 = _read_datas_T[2399:2384]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__4_22 = _read_datas_T[2415:2400]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__4_23 = _read_datas_T[2431:2416]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__4_24 = _read_datas_T[2447:2432]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__4_25 = _read_datas_T[2463:2448]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__4_26 = _read_datas_T[2479:2464]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__4_27 = _read_datas_T[2495:2480]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__4_28 = _read_datas_T[2511:2496]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__4_29 = _read_datas_T[2527:2512]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__4_30 = _read_datas_T[2543:2528]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__4_31 = _read_datas_T[2559:2544]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__5_0 = _read_datas_T[2575:2560]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__5_1 = _read_datas_T[2591:2576]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__5_2 = _read_datas_T[2607:2592]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__5_3 = _read_datas_T[2623:2608]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__5_4 = _read_datas_T[2639:2624]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__5_5 = _read_datas_T[2655:2640]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__5_6 = _read_datas_T[2671:2656]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__5_7 = _read_datas_T[2687:2672]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__5_8 = _read_datas_T[2703:2688]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__5_9 = _read_datas_T[2719:2704]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__5_10 = _read_datas_T[2735:2720]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__5_11 = _read_datas_T[2751:2736]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__5_12 = _read_datas_T[2767:2752]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__5_13 = _read_datas_T[2783:2768]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__5_14 = _read_datas_T[2799:2784]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__5_15 = _read_datas_T[2815:2800]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__5_16 = _read_datas_T[2831:2816]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__5_17 = _read_datas_T[2847:2832]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__5_18 = _read_datas_T[2863:2848]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__5_19 = _read_datas_T[2879:2864]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__5_20 = _read_datas_T[2895:2880]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__5_21 = _read_datas_T[2911:2896]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__5_22 = _read_datas_T[2927:2912]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__5_23 = _read_datas_T[2943:2928]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__5_24 = _read_datas_T[2959:2944]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__5_25 = _read_datas_T[2975:2960]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__5_26 = _read_datas_T[2991:2976]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__5_27 = _read_datas_T[3007:2992]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__5_28 = _read_datas_T[3023:3008]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__5_29 = _read_datas_T[3039:3024]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__5_30 = _read_datas_T[3055:3040]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__5_31 = _read_datas_T[3071:3056]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__6_0 = _read_datas_T[3087:3072]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__6_1 = _read_datas_T[3103:3088]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__6_2 = _read_datas_T[3119:3104]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__6_3 = _read_datas_T[3135:3120]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__6_4 = _read_datas_T[3151:3136]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__6_5 = _read_datas_T[3167:3152]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__6_6 = _read_datas_T[3183:3168]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__6_7 = _read_datas_T[3199:3184]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__6_8 = _read_datas_T[3215:3200]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__6_9 = _read_datas_T[3231:3216]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__6_10 = _read_datas_T[3247:3232]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__6_11 = _read_datas_T[3263:3248]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__6_12 = _read_datas_T[3279:3264]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__6_13 = _read_datas_T[3295:3280]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__6_14 = _read_datas_T[3311:3296]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__6_15 = _read_datas_T[3327:3312]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__6_16 = _read_datas_T[3343:3328]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__6_17 = _read_datas_T[3359:3344]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__6_18 = _read_datas_T[3375:3360]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__6_19 = _read_datas_T[3391:3376]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__6_20 = _read_datas_T[3407:3392]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__6_21 = _read_datas_T[3423:3408]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__6_22 = _read_datas_T[3439:3424]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__6_23 = _read_datas_T[3455:3440]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__6_24 = _read_datas_T[3471:3456]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__6_25 = _read_datas_T[3487:3472]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__6_26 = _read_datas_T[3503:3488]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__6_27 = _read_datas_T[3519:3504]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__6_28 = _read_datas_T[3535:3520]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__6_29 = _read_datas_T[3551:3536]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__6_30 = _read_datas_T[3567:3552]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__6_31 = _read_datas_T[3583:3568]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__7_0 = _read_datas_T[3599:3584]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__7_1 = _read_datas_T[3615:3600]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__7_2 = _read_datas_T[3631:3616]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__7_3 = _read_datas_T[3647:3632]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__7_4 = _read_datas_T[3663:3648]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__7_5 = _read_datas_T[3679:3664]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__7_6 = _read_datas_T[3695:3680]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__7_7 = _read_datas_T[3711:3696]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__7_8 = _read_datas_T[3727:3712]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__7_9 = _read_datas_T[3743:3728]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__7_10 = _read_datas_T[3759:3744]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__7_11 = _read_datas_T[3775:3760]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__7_12 = _read_datas_T[3791:3776]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__7_13 = _read_datas_T[3807:3792]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__7_14 = _read_datas_T[3823:3808]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__7_15 = _read_datas_T[3839:3824]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__7_16 = _read_datas_T[3855:3840]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__7_17 = _read_datas_T[3871:3856]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__7_18 = _read_datas_T[3887:3872]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__7_19 = _read_datas_T[3903:3888]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__7_20 = _read_datas_T[3919:3904]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__7_21 = _read_datas_T[3935:3920]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__7_22 = _read_datas_T[3951:3936]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__7_23 = _read_datas_T[3967:3952]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__7_24 = _read_datas_T[3983:3968]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__7_25 = _read_datas_T[3999:3984]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__7_26 = _read_datas_T[4015:4000]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__7_27 = _read_datas_T[4031:4016]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__7_28 = _read_datas_T[4047:4032]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__7_29 = _read_datas_T[4063:4048]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__7_30 = _read_datas_T[4079:4064]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas__7_31 = _read_datas_T[4095:4080]; // @[ICacheMainPipe.scala 369:51]
  wire [255:0] _read_codes_T = {s2_data_errorBits_0_7,s2_data_errorBits_0_6,s2_data_errorBits_0_5,s2_data_errorBits_0_4,
    s2_data_errorBits_0_3,s2_data_errorBits_0_2,s2_data_errorBits_0_1,s2_data_errorBits_0_0}; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__0_0 = _read_codes_T[0]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__0_1 = _read_codes_T[1]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__0_2 = _read_codes_T[2]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__0_3 = _read_codes_T[3]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__0_4 = _read_codes_T[4]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__0_5 = _read_codes_T[5]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__0_6 = _read_codes_T[6]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__0_7 = _read_codes_T[7]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__0_8 = _read_codes_T[8]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__0_9 = _read_codes_T[9]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__0_10 = _read_codes_T[10]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__0_11 = _read_codes_T[11]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__0_12 = _read_codes_T[12]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__0_13 = _read_codes_T[13]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__0_14 = _read_codes_T[14]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__0_15 = _read_codes_T[15]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__0_16 = _read_codes_T[16]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__0_17 = _read_codes_T[17]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__0_18 = _read_codes_T[18]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__0_19 = _read_codes_T[19]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__0_20 = _read_codes_T[20]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__0_21 = _read_codes_T[21]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__0_22 = _read_codes_T[22]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__0_23 = _read_codes_T[23]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__0_24 = _read_codes_T[24]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__0_25 = _read_codes_T[25]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__0_26 = _read_codes_T[26]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__0_27 = _read_codes_T[27]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__0_28 = _read_codes_T[28]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__0_29 = _read_codes_T[29]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__0_30 = _read_codes_T[30]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__0_31 = _read_codes_T[31]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__1_0 = _read_codes_T[32]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__1_1 = _read_codes_T[33]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__1_2 = _read_codes_T[34]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__1_3 = _read_codes_T[35]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__1_4 = _read_codes_T[36]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__1_5 = _read_codes_T[37]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__1_6 = _read_codes_T[38]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__1_7 = _read_codes_T[39]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__1_8 = _read_codes_T[40]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__1_9 = _read_codes_T[41]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__1_10 = _read_codes_T[42]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__1_11 = _read_codes_T[43]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__1_12 = _read_codes_T[44]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__1_13 = _read_codes_T[45]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__1_14 = _read_codes_T[46]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__1_15 = _read_codes_T[47]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__1_16 = _read_codes_T[48]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__1_17 = _read_codes_T[49]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__1_18 = _read_codes_T[50]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__1_19 = _read_codes_T[51]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__1_20 = _read_codes_T[52]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__1_21 = _read_codes_T[53]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__1_22 = _read_codes_T[54]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__1_23 = _read_codes_T[55]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__1_24 = _read_codes_T[56]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__1_25 = _read_codes_T[57]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__1_26 = _read_codes_T[58]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__1_27 = _read_codes_T[59]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__1_28 = _read_codes_T[60]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__1_29 = _read_codes_T[61]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__1_30 = _read_codes_T[62]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__1_31 = _read_codes_T[63]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__2_0 = _read_codes_T[64]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__2_1 = _read_codes_T[65]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__2_2 = _read_codes_T[66]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__2_3 = _read_codes_T[67]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__2_4 = _read_codes_T[68]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__2_5 = _read_codes_T[69]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__2_6 = _read_codes_T[70]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__2_7 = _read_codes_T[71]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__2_8 = _read_codes_T[72]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__2_9 = _read_codes_T[73]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__2_10 = _read_codes_T[74]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__2_11 = _read_codes_T[75]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__2_12 = _read_codes_T[76]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__2_13 = _read_codes_T[77]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__2_14 = _read_codes_T[78]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__2_15 = _read_codes_T[79]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__2_16 = _read_codes_T[80]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__2_17 = _read_codes_T[81]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__2_18 = _read_codes_T[82]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__2_19 = _read_codes_T[83]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__2_20 = _read_codes_T[84]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__2_21 = _read_codes_T[85]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__2_22 = _read_codes_T[86]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__2_23 = _read_codes_T[87]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__2_24 = _read_codes_T[88]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__2_25 = _read_codes_T[89]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__2_26 = _read_codes_T[90]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__2_27 = _read_codes_T[91]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__2_28 = _read_codes_T[92]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__2_29 = _read_codes_T[93]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__2_30 = _read_codes_T[94]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__2_31 = _read_codes_T[95]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__3_0 = _read_codes_T[96]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__3_1 = _read_codes_T[97]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__3_2 = _read_codes_T[98]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__3_3 = _read_codes_T[99]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__3_4 = _read_codes_T[100]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__3_5 = _read_codes_T[101]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__3_6 = _read_codes_T[102]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__3_7 = _read_codes_T[103]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__3_8 = _read_codes_T[104]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__3_9 = _read_codes_T[105]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__3_10 = _read_codes_T[106]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__3_11 = _read_codes_T[107]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__3_12 = _read_codes_T[108]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__3_13 = _read_codes_T[109]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__3_14 = _read_codes_T[110]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__3_15 = _read_codes_T[111]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__3_16 = _read_codes_T[112]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__3_17 = _read_codes_T[113]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__3_18 = _read_codes_T[114]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__3_19 = _read_codes_T[115]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__3_20 = _read_codes_T[116]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__3_21 = _read_codes_T[117]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__3_22 = _read_codes_T[118]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__3_23 = _read_codes_T[119]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__3_24 = _read_codes_T[120]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__3_25 = _read_codes_T[121]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__3_26 = _read_codes_T[122]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__3_27 = _read_codes_T[123]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__3_28 = _read_codes_T[124]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__3_29 = _read_codes_T[125]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__3_30 = _read_codes_T[126]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__3_31 = _read_codes_T[127]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__4_0 = _read_codes_T[128]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__4_1 = _read_codes_T[129]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__4_2 = _read_codes_T[130]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__4_3 = _read_codes_T[131]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__4_4 = _read_codes_T[132]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__4_5 = _read_codes_T[133]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__4_6 = _read_codes_T[134]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__4_7 = _read_codes_T[135]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__4_8 = _read_codes_T[136]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__4_9 = _read_codes_T[137]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__4_10 = _read_codes_T[138]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__4_11 = _read_codes_T[139]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__4_12 = _read_codes_T[140]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__4_13 = _read_codes_T[141]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__4_14 = _read_codes_T[142]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__4_15 = _read_codes_T[143]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__4_16 = _read_codes_T[144]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__4_17 = _read_codes_T[145]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__4_18 = _read_codes_T[146]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__4_19 = _read_codes_T[147]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__4_20 = _read_codes_T[148]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__4_21 = _read_codes_T[149]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__4_22 = _read_codes_T[150]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__4_23 = _read_codes_T[151]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__4_24 = _read_codes_T[152]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__4_25 = _read_codes_T[153]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__4_26 = _read_codes_T[154]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__4_27 = _read_codes_T[155]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__4_28 = _read_codes_T[156]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__4_29 = _read_codes_T[157]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__4_30 = _read_codes_T[158]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__4_31 = _read_codes_T[159]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__5_0 = _read_codes_T[160]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__5_1 = _read_codes_T[161]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__5_2 = _read_codes_T[162]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__5_3 = _read_codes_T[163]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__5_4 = _read_codes_T[164]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__5_5 = _read_codes_T[165]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__5_6 = _read_codes_T[166]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__5_7 = _read_codes_T[167]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__5_8 = _read_codes_T[168]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__5_9 = _read_codes_T[169]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__5_10 = _read_codes_T[170]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__5_11 = _read_codes_T[171]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__5_12 = _read_codes_T[172]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__5_13 = _read_codes_T[173]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__5_14 = _read_codes_T[174]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__5_15 = _read_codes_T[175]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__5_16 = _read_codes_T[176]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__5_17 = _read_codes_T[177]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__5_18 = _read_codes_T[178]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__5_19 = _read_codes_T[179]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__5_20 = _read_codes_T[180]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__5_21 = _read_codes_T[181]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__5_22 = _read_codes_T[182]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__5_23 = _read_codes_T[183]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__5_24 = _read_codes_T[184]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__5_25 = _read_codes_T[185]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__5_26 = _read_codes_T[186]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__5_27 = _read_codes_T[187]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__5_28 = _read_codes_T[188]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__5_29 = _read_codes_T[189]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__5_30 = _read_codes_T[190]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__5_31 = _read_codes_T[191]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__6_0 = _read_codes_T[192]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__6_1 = _read_codes_T[193]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__6_2 = _read_codes_T[194]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__6_3 = _read_codes_T[195]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__6_4 = _read_codes_T[196]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__6_5 = _read_codes_T[197]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__6_6 = _read_codes_T[198]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__6_7 = _read_codes_T[199]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__6_8 = _read_codes_T[200]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__6_9 = _read_codes_T[201]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__6_10 = _read_codes_T[202]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__6_11 = _read_codes_T[203]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__6_12 = _read_codes_T[204]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__6_13 = _read_codes_T[205]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__6_14 = _read_codes_T[206]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__6_15 = _read_codes_T[207]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__6_16 = _read_codes_T[208]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__6_17 = _read_codes_T[209]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__6_18 = _read_codes_T[210]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__6_19 = _read_codes_T[211]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__6_20 = _read_codes_T[212]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__6_21 = _read_codes_T[213]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__6_22 = _read_codes_T[214]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__6_23 = _read_codes_T[215]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__6_24 = _read_codes_T[216]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__6_25 = _read_codes_T[217]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__6_26 = _read_codes_T[218]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__6_27 = _read_codes_T[219]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__6_28 = _read_codes_T[220]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__6_29 = _read_codes_T[221]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__6_30 = _read_codes_T[222]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__6_31 = _read_codes_T[223]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__7_0 = _read_codes_T[224]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__7_1 = _read_codes_T[225]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__7_2 = _read_codes_T[226]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__7_3 = _read_codes_T[227]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__7_4 = _read_codes_T[228]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__7_5 = _read_codes_T[229]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__7_6 = _read_codes_T[230]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__7_7 = _read_codes_T[231]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__7_8 = _read_codes_T[232]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__7_9 = _read_codes_T[233]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__7_10 = _read_codes_T[234]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__7_11 = _read_codes_T[235]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__7_12 = _read_codes_T[236]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__7_13 = _read_codes_T[237]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__7_14 = _read_codes_T[238]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__7_15 = _read_codes_T[239]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__7_16 = _read_codes_T[240]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__7_17 = _read_codes_T[241]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__7_18 = _read_codes_T[242]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__7_19 = _read_codes_T[243]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__7_20 = _read_codes_T[244]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__7_21 = _read_codes_T[245]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__7_22 = _read_codes_T[246]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__7_23 = _read_codes_T[247]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__7_24 = _read_codes_T[248]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__7_25 = _read_codes_T[249]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__7_26 = _read_codes_T[250]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__7_27 = _read_codes_T[251]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__7_28 = _read_codes_T[252]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__7_29 = _read_codes_T[253]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__7_30 = _read_codes_T[254]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes__7_31 = _read_codes_T[255]; // @[ICacheMainPipe.scala 370:51]
  wire [16:0] data_full_wayBits__0_0 = {read_codes__0_0,read_datas__0_0}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__0_1 = {read_codes__0_1,read_datas__0_1}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__0_2 = {read_codes__0_2,read_datas__0_2}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__0_3 = {read_codes__0_3,read_datas__0_3}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__0_4 = {read_codes__0_4,read_datas__0_4}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__0_5 = {read_codes__0_5,read_datas__0_5}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__0_6 = {read_codes__0_6,read_datas__0_6}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__0_7 = {read_codes__0_7,read_datas__0_7}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__0_8 = {read_codes__0_8,read_datas__0_8}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__0_9 = {read_codes__0_9,read_datas__0_9}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__0_10 = {read_codes__0_10,read_datas__0_10}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__0_11 = {read_codes__0_11,read_datas__0_11}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__0_12 = {read_codes__0_12,read_datas__0_12}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__0_13 = {read_codes__0_13,read_datas__0_13}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__0_14 = {read_codes__0_14,read_datas__0_14}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__0_15 = {read_codes__0_15,read_datas__0_15}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__0_16 = {read_codes__0_16,read_datas__0_16}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__0_17 = {read_codes__0_17,read_datas__0_17}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__0_18 = {read_codes__0_18,read_datas__0_18}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__0_19 = {read_codes__0_19,read_datas__0_19}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__0_20 = {read_codes__0_20,read_datas__0_20}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__0_21 = {read_codes__0_21,read_datas__0_21}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__0_22 = {read_codes__0_22,read_datas__0_22}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__0_23 = {read_codes__0_23,read_datas__0_23}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__0_24 = {read_codes__0_24,read_datas__0_24}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__0_25 = {read_codes__0_25,read_datas__0_25}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__0_26 = {read_codes__0_26,read_datas__0_26}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__0_27 = {read_codes__0_27,read_datas__0_27}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__0_28 = {read_codes__0_28,read_datas__0_28}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__0_29 = {read_codes__0_29,read_datas__0_29}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__0_30 = {read_codes__0_30,read_datas__0_30}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__0_31 = {read_codes__0_31,read_datas__0_31}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__1_0 = {read_codes__1_0,read_datas__1_0}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__1_1 = {read_codes__1_1,read_datas__1_1}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__1_2 = {read_codes__1_2,read_datas__1_2}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__1_3 = {read_codes__1_3,read_datas__1_3}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__1_4 = {read_codes__1_4,read_datas__1_4}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__1_5 = {read_codes__1_5,read_datas__1_5}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__1_6 = {read_codes__1_6,read_datas__1_6}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__1_7 = {read_codes__1_7,read_datas__1_7}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__1_8 = {read_codes__1_8,read_datas__1_8}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__1_9 = {read_codes__1_9,read_datas__1_9}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__1_10 = {read_codes__1_10,read_datas__1_10}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__1_11 = {read_codes__1_11,read_datas__1_11}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__1_12 = {read_codes__1_12,read_datas__1_12}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__1_13 = {read_codes__1_13,read_datas__1_13}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__1_14 = {read_codes__1_14,read_datas__1_14}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__1_15 = {read_codes__1_15,read_datas__1_15}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__1_16 = {read_codes__1_16,read_datas__1_16}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__1_17 = {read_codes__1_17,read_datas__1_17}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__1_18 = {read_codes__1_18,read_datas__1_18}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__1_19 = {read_codes__1_19,read_datas__1_19}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__1_20 = {read_codes__1_20,read_datas__1_20}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__1_21 = {read_codes__1_21,read_datas__1_21}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__1_22 = {read_codes__1_22,read_datas__1_22}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__1_23 = {read_codes__1_23,read_datas__1_23}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__1_24 = {read_codes__1_24,read_datas__1_24}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__1_25 = {read_codes__1_25,read_datas__1_25}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__1_26 = {read_codes__1_26,read_datas__1_26}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__1_27 = {read_codes__1_27,read_datas__1_27}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__1_28 = {read_codes__1_28,read_datas__1_28}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__1_29 = {read_codes__1_29,read_datas__1_29}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__1_30 = {read_codes__1_30,read_datas__1_30}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__1_31 = {read_codes__1_31,read_datas__1_31}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__2_0 = {read_codes__2_0,read_datas__2_0}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__2_1 = {read_codes__2_1,read_datas__2_1}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__2_2 = {read_codes__2_2,read_datas__2_2}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__2_3 = {read_codes__2_3,read_datas__2_3}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__2_4 = {read_codes__2_4,read_datas__2_4}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__2_5 = {read_codes__2_5,read_datas__2_5}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__2_6 = {read_codes__2_6,read_datas__2_6}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__2_7 = {read_codes__2_7,read_datas__2_7}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__2_8 = {read_codes__2_8,read_datas__2_8}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__2_9 = {read_codes__2_9,read_datas__2_9}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__2_10 = {read_codes__2_10,read_datas__2_10}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__2_11 = {read_codes__2_11,read_datas__2_11}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__2_12 = {read_codes__2_12,read_datas__2_12}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__2_13 = {read_codes__2_13,read_datas__2_13}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__2_14 = {read_codes__2_14,read_datas__2_14}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__2_15 = {read_codes__2_15,read_datas__2_15}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__2_16 = {read_codes__2_16,read_datas__2_16}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__2_17 = {read_codes__2_17,read_datas__2_17}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__2_18 = {read_codes__2_18,read_datas__2_18}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__2_19 = {read_codes__2_19,read_datas__2_19}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__2_20 = {read_codes__2_20,read_datas__2_20}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__2_21 = {read_codes__2_21,read_datas__2_21}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__2_22 = {read_codes__2_22,read_datas__2_22}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__2_23 = {read_codes__2_23,read_datas__2_23}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__2_24 = {read_codes__2_24,read_datas__2_24}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__2_25 = {read_codes__2_25,read_datas__2_25}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__2_26 = {read_codes__2_26,read_datas__2_26}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__2_27 = {read_codes__2_27,read_datas__2_27}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__2_28 = {read_codes__2_28,read_datas__2_28}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__2_29 = {read_codes__2_29,read_datas__2_29}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__2_30 = {read_codes__2_30,read_datas__2_30}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__2_31 = {read_codes__2_31,read_datas__2_31}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__3_0 = {read_codes__3_0,read_datas__3_0}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__3_1 = {read_codes__3_1,read_datas__3_1}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__3_2 = {read_codes__3_2,read_datas__3_2}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__3_3 = {read_codes__3_3,read_datas__3_3}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__3_4 = {read_codes__3_4,read_datas__3_4}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__3_5 = {read_codes__3_5,read_datas__3_5}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__3_6 = {read_codes__3_6,read_datas__3_6}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__3_7 = {read_codes__3_7,read_datas__3_7}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__3_8 = {read_codes__3_8,read_datas__3_8}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__3_9 = {read_codes__3_9,read_datas__3_9}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__3_10 = {read_codes__3_10,read_datas__3_10}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__3_11 = {read_codes__3_11,read_datas__3_11}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__3_12 = {read_codes__3_12,read_datas__3_12}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__3_13 = {read_codes__3_13,read_datas__3_13}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__3_14 = {read_codes__3_14,read_datas__3_14}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__3_15 = {read_codes__3_15,read_datas__3_15}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__3_16 = {read_codes__3_16,read_datas__3_16}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__3_17 = {read_codes__3_17,read_datas__3_17}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__3_18 = {read_codes__3_18,read_datas__3_18}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__3_19 = {read_codes__3_19,read_datas__3_19}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__3_20 = {read_codes__3_20,read_datas__3_20}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__3_21 = {read_codes__3_21,read_datas__3_21}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__3_22 = {read_codes__3_22,read_datas__3_22}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__3_23 = {read_codes__3_23,read_datas__3_23}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__3_24 = {read_codes__3_24,read_datas__3_24}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__3_25 = {read_codes__3_25,read_datas__3_25}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__3_26 = {read_codes__3_26,read_datas__3_26}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__3_27 = {read_codes__3_27,read_datas__3_27}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__3_28 = {read_codes__3_28,read_datas__3_28}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__3_29 = {read_codes__3_29,read_datas__3_29}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__3_30 = {read_codes__3_30,read_datas__3_30}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__3_31 = {read_codes__3_31,read_datas__3_31}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__4_0 = {read_codes__4_0,read_datas__4_0}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__4_1 = {read_codes__4_1,read_datas__4_1}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__4_2 = {read_codes__4_2,read_datas__4_2}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__4_3 = {read_codes__4_3,read_datas__4_3}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__4_4 = {read_codes__4_4,read_datas__4_4}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__4_5 = {read_codes__4_5,read_datas__4_5}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__4_6 = {read_codes__4_6,read_datas__4_6}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__4_7 = {read_codes__4_7,read_datas__4_7}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__4_8 = {read_codes__4_8,read_datas__4_8}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__4_9 = {read_codes__4_9,read_datas__4_9}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__4_10 = {read_codes__4_10,read_datas__4_10}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__4_11 = {read_codes__4_11,read_datas__4_11}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__4_12 = {read_codes__4_12,read_datas__4_12}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__4_13 = {read_codes__4_13,read_datas__4_13}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__4_14 = {read_codes__4_14,read_datas__4_14}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__4_15 = {read_codes__4_15,read_datas__4_15}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__4_16 = {read_codes__4_16,read_datas__4_16}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__4_17 = {read_codes__4_17,read_datas__4_17}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__4_18 = {read_codes__4_18,read_datas__4_18}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__4_19 = {read_codes__4_19,read_datas__4_19}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__4_20 = {read_codes__4_20,read_datas__4_20}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__4_21 = {read_codes__4_21,read_datas__4_21}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__4_22 = {read_codes__4_22,read_datas__4_22}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__4_23 = {read_codes__4_23,read_datas__4_23}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__4_24 = {read_codes__4_24,read_datas__4_24}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__4_25 = {read_codes__4_25,read_datas__4_25}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__4_26 = {read_codes__4_26,read_datas__4_26}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__4_27 = {read_codes__4_27,read_datas__4_27}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__4_28 = {read_codes__4_28,read_datas__4_28}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__4_29 = {read_codes__4_29,read_datas__4_29}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__4_30 = {read_codes__4_30,read_datas__4_30}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__4_31 = {read_codes__4_31,read_datas__4_31}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__5_0 = {read_codes__5_0,read_datas__5_0}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__5_1 = {read_codes__5_1,read_datas__5_1}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__5_2 = {read_codes__5_2,read_datas__5_2}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__5_3 = {read_codes__5_3,read_datas__5_3}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__5_4 = {read_codes__5_4,read_datas__5_4}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__5_5 = {read_codes__5_5,read_datas__5_5}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__5_6 = {read_codes__5_6,read_datas__5_6}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__5_7 = {read_codes__5_7,read_datas__5_7}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__5_8 = {read_codes__5_8,read_datas__5_8}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__5_9 = {read_codes__5_9,read_datas__5_9}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__5_10 = {read_codes__5_10,read_datas__5_10}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__5_11 = {read_codes__5_11,read_datas__5_11}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__5_12 = {read_codes__5_12,read_datas__5_12}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__5_13 = {read_codes__5_13,read_datas__5_13}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__5_14 = {read_codes__5_14,read_datas__5_14}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__5_15 = {read_codes__5_15,read_datas__5_15}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__5_16 = {read_codes__5_16,read_datas__5_16}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__5_17 = {read_codes__5_17,read_datas__5_17}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__5_18 = {read_codes__5_18,read_datas__5_18}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__5_19 = {read_codes__5_19,read_datas__5_19}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__5_20 = {read_codes__5_20,read_datas__5_20}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__5_21 = {read_codes__5_21,read_datas__5_21}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__5_22 = {read_codes__5_22,read_datas__5_22}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__5_23 = {read_codes__5_23,read_datas__5_23}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__5_24 = {read_codes__5_24,read_datas__5_24}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__5_25 = {read_codes__5_25,read_datas__5_25}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__5_26 = {read_codes__5_26,read_datas__5_26}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__5_27 = {read_codes__5_27,read_datas__5_27}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__5_28 = {read_codes__5_28,read_datas__5_28}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__5_29 = {read_codes__5_29,read_datas__5_29}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__5_30 = {read_codes__5_30,read_datas__5_30}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__5_31 = {read_codes__5_31,read_datas__5_31}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__6_0 = {read_codes__6_0,read_datas__6_0}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__6_1 = {read_codes__6_1,read_datas__6_1}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__6_2 = {read_codes__6_2,read_datas__6_2}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__6_3 = {read_codes__6_3,read_datas__6_3}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__6_4 = {read_codes__6_4,read_datas__6_4}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__6_5 = {read_codes__6_5,read_datas__6_5}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__6_6 = {read_codes__6_6,read_datas__6_6}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__6_7 = {read_codes__6_7,read_datas__6_7}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__6_8 = {read_codes__6_8,read_datas__6_8}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__6_9 = {read_codes__6_9,read_datas__6_9}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__6_10 = {read_codes__6_10,read_datas__6_10}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__6_11 = {read_codes__6_11,read_datas__6_11}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__6_12 = {read_codes__6_12,read_datas__6_12}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__6_13 = {read_codes__6_13,read_datas__6_13}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__6_14 = {read_codes__6_14,read_datas__6_14}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__6_15 = {read_codes__6_15,read_datas__6_15}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__6_16 = {read_codes__6_16,read_datas__6_16}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__6_17 = {read_codes__6_17,read_datas__6_17}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__6_18 = {read_codes__6_18,read_datas__6_18}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__6_19 = {read_codes__6_19,read_datas__6_19}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__6_20 = {read_codes__6_20,read_datas__6_20}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__6_21 = {read_codes__6_21,read_datas__6_21}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__6_22 = {read_codes__6_22,read_datas__6_22}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__6_23 = {read_codes__6_23,read_datas__6_23}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__6_24 = {read_codes__6_24,read_datas__6_24}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__6_25 = {read_codes__6_25,read_datas__6_25}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__6_26 = {read_codes__6_26,read_datas__6_26}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__6_27 = {read_codes__6_27,read_datas__6_27}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__6_28 = {read_codes__6_28,read_datas__6_28}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__6_29 = {read_codes__6_29,read_datas__6_29}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__6_30 = {read_codes__6_30,read_datas__6_30}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__6_31 = {read_codes__6_31,read_datas__6_31}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__7_0 = {read_codes__7_0,read_datas__7_0}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__7_1 = {read_codes__7_1,read_datas__7_1}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__7_2 = {read_codes__7_2,read_datas__7_2}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__7_3 = {read_codes__7_3,read_datas__7_3}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__7_4 = {read_codes__7_4,read_datas__7_4}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__7_5 = {read_codes__7_5,read_datas__7_5}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__7_6 = {read_codes__7_6,read_datas__7_6}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__7_7 = {read_codes__7_7,read_datas__7_7}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__7_8 = {read_codes__7_8,read_datas__7_8}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__7_9 = {read_codes__7_9,read_datas__7_9}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__7_10 = {read_codes__7_10,read_datas__7_10}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__7_11 = {read_codes__7_11,read_datas__7_11}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__7_12 = {read_codes__7_12,read_datas__7_12}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__7_13 = {read_codes__7_13,read_datas__7_13}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__7_14 = {read_codes__7_14,read_datas__7_14}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__7_15 = {read_codes__7_15,read_datas__7_15}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__7_16 = {read_codes__7_16,read_datas__7_16}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__7_17 = {read_codes__7_17,read_datas__7_17}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__7_18 = {read_codes__7_18,read_datas__7_18}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__7_19 = {read_codes__7_19,read_datas__7_19}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__7_20 = {read_codes__7_20,read_datas__7_20}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__7_21 = {read_codes__7_21,read_datas__7_21}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__7_22 = {read_codes__7_22,read_datas__7_22}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__7_23 = {read_codes__7_23,read_datas__7_23}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__7_24 = {read_codes__7_24,read_datas__7_24}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__7_25 = {read_codes__7_25,read_datas__7_25}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__7_26 = {read_codes__7_26,read_datas__7_26}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__7_27 = {read_codes__7_27,read_datas__7_27}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__7_28 = {read_codes__7_28,read_datas__7_28}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__7_29 = {read_codes__7_29,read_datas__7_29}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__7_30 = {read_codes__7_30,read_datas__7_30}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits__7_31 = {read_codes__7_31,read_datas__7_31}; // @[Cat.scala 31:58]
  reg  s2_data_errors_0_0_REG; // @[ICacheMainPipe.scala 379:48]
  reg  s2_data_errors_0_0_REG_1; // @[ICacheMainPipe.scala 379:40]
  reg  s2_data_errors_0_0_REG_2_0; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_0_REG_2_1; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_0_REG_2_2; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_0_REG_2_3; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_0_REG_2_4; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_0_REG_2_5; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_0_REG_2_6; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_0_REG_2_7; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_0_REG_2_8; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_0_REG_2_9; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_0_REG_2_10; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_0_REG_2_11; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_0_REG_2_12; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_0_REG_2_13; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_0_REG_2_14; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_0_REG_2_15; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_0_REG_2_16; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_0_REG_2_17; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_0_REG_2_18; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_0_REG_2_19; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_0_REG_2_20; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_0_REG_2_21; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_0_REG_2_22; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_0_REG_2_23; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_0_REG_2_24; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_0_REG_2_25; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_0_REG_2_26; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_0_REG_2_27; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_0_REG_2_28; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_0_REG_2_29; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_0_REG_2_30; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_0_REG_2_31; // @[ICacheMainPipe.scala 379:69]
  wire  _s2_data_errors_0_0_T_29 = s2_data_errors_0_0_REG_2_0 | s2_data_errors_0_0_REG_2_1 | s2_data_errors_0_0_REG_2_2
     | s2_data_errors_0_0_REG_2_3 | s2_data_errors_0_0_REG_2_4 | s2_data_errors_0_0_REG_2_5 | s2_data_errors_0_0_REG_2_6
     | s2_data_errors_0_0_REG_2_7 | s2_data_errors_0_0_REG_2_8 | s2_data_errors_0_0_REG_2_9 |
    s2_data_errors_0_0_REG_2_10 | s2_data_errors_0_0_REG_2_11 | s2_data_errors_0_0_REG_2_12 |
    s2_data_errors_0_0_REG_2_13 | s2_data_errors_0_0_REG_2_14 | s2_data_errors_0_0_REG_2_15 |
    s2_data_errors_0_0_REG_2_16 | s2_data_errors_0_0_REG_2_17 | s2_data_errors_0_0_REG_2_18 |
    s2_data_errors_0_0_REG_2_19 | s2_data_errors_0_0_REG_2_20 | s2_data_errors_0_0_REG_2_21 |
    s2_data_errors_0_0_REG_2_22 | s2_data_errors_0_0_REG_2_23 | s2_data_errors_0_0_REG_2_24 |
    s2_data_errors_0_0_REG_2_25 | s2_data_errors_0_0_REG_2_26 | s2_data_errors_0_0_REG_2_27 |
    s2_data_errors_0_0_REG_2_28 | s2_data_errors_0_0_REG_2_29 | s2_data_errors_0_0_REG_2_30; // @[ICacheMainPipe.scala 379:101]
  wire  s2_data_errors_0_0 = s2_data_errors_0_0_REG_1 & (_s2_data_errors_0_0_T_29 | s2_data_errors_0_0_REG_2_31); // @[ICacheMainPipe.scala 379:59]
  reg  s2_data_errors_0_1_REG; // @[ICacheMainPipe.scala 379:48]
  reg  s2_data_errors_0_1_REG_1; // @[ICacheMainPipe.scala 379:40]
  reg  s2_data_errors_0_1_REG_2_0; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_1_REG_2_1; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_1_REG_2_2; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_1_REG_2_3; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_1_REG_2_4; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_1_REG_2_5; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_1_REG_2_6; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_1_REG_2_7; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_1_REG_2_8; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_1_REG_2_9; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_1_REG_2_10; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_1_REG_2_11; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_1_REG_2_12; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_1_REG_2_13; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_1_REG_2_14; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_1_REG_2_15; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_1_REG_2_16; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_1_REG_2_17; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_1_REG_2_18; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_1_REG_2_19; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_1_REG_2_20; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_1_REG_2_21; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_1_REG_2_22; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_1_REG_2_23; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_1_REG_2_24; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_1_REG_2_25; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_1_REG_2_26; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_1_REG_2_27; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_1_REG_2_28; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_1_REG_2_29; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_1_REG_2_30; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_1_REG_2_31; // @[ICacheMainPipe.scala 379:69]
  wire  _s2_data_errors_0_1_T_29 = s2_data_errors_0_1_REG_2_0 | s2_data_errors_0_1_REG_2_1 | s2_data_errors_0_1_REG_2_2
     | s2_data_errors_0_1_REG_2_3 | s2_data_errors_0_1_REG_2_4 | s2_data_errors_0_1_REG_2_5 | s2_data_errors_0_1_REG_2_6
     | s2_data_errors_0_1_REG_2_7 | s2_data_errors_0_1_REG_2_8 | s2_data_errors_0_1_REG_2_9 |
    s2_data_errors_0_1_REG_2_10 | s2_data_errors_0_1_REG_2_11 | s2_data_errors_0_1_REG_2_12 |
    s2_data_errors_0_1_REG_2_13 | s2_data_errors_0_1_REG_2_14 | s2_data_errors_0_1_REG_2_15 |
    s2_data_errors_0_1_REG_2_16 | s2_data_errors_0_1_REG_2_17 | s2_data_errors_0_1_REG_2_18 |
    s2_data_errors_0_1_REG_2_19 | s2_data_errors_0_1_REG_2_20 | s2_data_errors_0_1_REG_2_21 |
    s2_data_errors_0_1_REG_2_22 | s2_data_errors_0_1_REG_2_23 | s2_data_errors_0_1_REG_2_24 |
    s2_data_errors_0_1_REG_2_25 | s2_data_errors_0_1_REG_2_26 | s2_data_errors_0_1_REG_2_27 |
    s2_data_errors_0_1_REG_2_28 | s2_data_errors_0_1_REG_2_29 | s2_data_errors_0_1_REG_2_30; // @[ICacheMainPipe.scala 379:101]
  wire  s2_data_errors_0_1 = s2_data_errors_0_1_REG_1 & (_s2_data_errors_0_1_T_29 | s2_data_errors_0_1_REG_2_31); // @[ICacheMainPipe.scala 379:59]
  reg  s2_data_errors_0_2_REG; // @[ICacheMainPipe.scala 379:48]
  reg  s2_data_errors_0_2_REG_1; // @[ICacheMainPipe.scala 379:40]
  reg  s2_data_errors_0_2_REG_2_0; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_2_REG_2_1; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_2_REG_2_2; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_2_REG_2_3; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_2_REG_2_4; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_2_REG_2_5; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_2_REG_2_6; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_2_REG_2_7; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_2_REG_2_8; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_2_REG_2_9; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_2_REG_2_10; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_2_REG_2_11; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_2_REG_2_12; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_2_REG_2_13; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_2_REG_2_14; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_2_REG_2_15; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_2_REG_2_16; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_2_REG_2_17; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_2_REG_2_18; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_2_REG_2_19; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_2_REG_2_20; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_2_REG_2_21; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_2_REG_2_22; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_2_REG_2_23; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_2_REG_2_24; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_2_REG_2_25; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_2_REG_2_26; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_2_REG_2_27; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_2_REG_2_28; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_2_REG_2_29; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_2_REG_2_30; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_2_REG_2_31; // @[ICacheMainPipe.scala 379:69]
  wire  _s2_data_errors_0_2_T_29 = s2_data_errors_0_2_REG_2_0 | s2_data_errors_0_2_REG_2_1 | s2_data_errors_0_2_REG_2_2
     | s2_data_errors_0_2_REG_2_3 | s2_data_errors_0_2_REG_2_4 | s2_data_errors_0_2_REG_2_5 | s2_data_errors_0_2_REG_2_6
     | s2_data_errors_0_2_REG_2_7 | s2_data_errors_0_2_REG_2_8 | s2_data_errors_0_2_REG_2_9 |
    s2_data_errors_0_2_REG_2_10 | s2_data_errors_0_2_REG_2_11 | s2_data_errors_0_2_REG_2_12 |
    s2_data_errors_0_2_REG_2_13 | s2_data_errors_0_2_REG_2_14 | s2_data_errors_0_2_REG_2_15 |
    s2_data_errors_0_2_REG_2_16 | s2_data_errors_0_2_REG_2_17 | s2_data_errors_0_2_REG_2_18 |
    s2_data_errors_0_2_REG_2_19 | s2_data_errors_0_2_REG_2_20 | s2_data_errors_0_2_REG_2_21 |
    s2_data_errors_0_2_REG_2_22 | s2_data_errors_0_2_REG_2_23 | s2_data_errors_0_2_REG_2_24 |
    s2_data_errors_0_2_REG_2_25 | s2_data_errors_0_2_REG_2_26 | s2_data_errors_0_2_REG_2_27 |
    s2_data_errors_0_2_REG_2_28 | s2_data_errors_0_2_REG_2_29 | s2_data_errors_0_2_REG_2_30; // @[ICacheMainPipe.scala 379:101]
  wire  s2_data_errors_0_2 = s2_data_errors_0_2_REG_1 & (_s2_data_errors_0_2_T_29 | s2_data_errors_0_2_REG_2_31); // @[ICacheMainPipe.scala 379:59]
  reg  s2_data_errors_0_3_REG; // @[ICacheMainPipe.scala 379:48]
  reg  s2_data_errors_0_3_REG_1; // @[ICacheMainPipe.scala 379:40]
  reg  s2_data_errors_0_3_REG_2_0; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_3_REG_2_1; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_3_REG_2_2; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_3_REG_2_3; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_3_REG_2_4; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_3_REG_2_5; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_3_REG_2_6; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_3_REG_2_7; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_3_REG_2_8; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_3_REG_2_9; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_3_REG_2_10; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_3_REG_2_11; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_3_REG_2_12; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_3_REG_2_13; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_3_REG_2_14; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_3_REG_2_15; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_3_REG_2_16; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_3_REG_2_17; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_3_REG_2_18; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_3_REG_2_19; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_3_REG_2_20; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_3_REG_2_21; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_3_REG_2_22; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_3_REG_2_23; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_3_REG_2_24; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_3_REG_2_25; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_3_REG_2_26; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_3_REG_2_27; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_3_REG_2_28; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_3_REG_2_29; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_3_REG_2_30; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_3_REG_2_31; // @[ICacheMainPipe.scala 379:69]
  wire  _s2_data_errors_0_3_T_29 = s2_data_errors_0_3_REG_2_0 | s2_data_errors_0_3_REG_2_1 | s2_data_errors_0_3_REG_2_2
     | s2_data_errors_0_3_REG_2_3 | s2_data_errors_0_3_REG_2_4 | s2_data_errors_0_3_REG_2_5 | s2_data_errors_0_3_REG_2_6
     | s2_data_errors_0_3_REG_2_7 | s2_data_errors_0_3_REG_2_8 | s2_data_errors_0_3_REG_2_9 |
    s2_data_errors_0_3_REG_2_10 | s2_data_errors_0_3_REG_2_11 | s2_data_errors_0_3_REG_2_12 |
    s2_data_errors_0_3_REG_2_13 | s2_data_errors_0_3_REG_2_14 | s2_data_errors_0_3_REG_2_15 |
    s2_data_errors_0_3_REG_2_16 | s2_data_errors_0_3_REG_2_17 | s2_data_errors_0_3_REG_2_18 |
    s2_data_errors_0_3_REG_2_19 | s2_data_errors_0_3_REG_2_20 | s2_data_errors_0_3_REG_2_21 |
    s2_data_errors_0_3_REG_2_22 | s2_data_errors_0_3_REG_2_23 | s2_data_errors_0_3_REG_2_24 |
    s2_data_errors_0_3_REG_2_25 | s2_data_errors_0_3_REG_2_26 | s2_data_errors_0_3_REG_2_27 |
    s2_data_errors_0_3_REG_2_28 | s2_data_errors_0_3_REG_2_29 | s2_data_errors_0_3_REG_2_30; // @[ICacheMainPipe.scala 379:101]
  wire  s2_data_errors_0_3 = s2_data_errors_0_3_REG_1 & (_s2_data_errors_0_3_T_29 | s2_data_errors_0_3_REG_2_31); // @[ICacheMainPipe.scala 379:59]
  reg  s2_data_errors_0_4_REG; // @[ICacheMainPipe.scala 379:48]
  reg  s2_data_errors_0_4_REG_1; // @[ICacheMainPipe.scala 379:40]
  reg  s2_data_errors_0_4_REG_2_0; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_4_REG_2_1; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_4_REG_2_2; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_4_REG_2_3; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_4_REG_2_4; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_4_REG_2_5; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_4_REG_2_6; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_4_REG_2_7; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_4_REG_2_8; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_4_REG_2_9; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_4_REG_2_10; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_4_REG_2_11; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_4_REG_2_12; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_4_REG_2_13; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_4_REG_2_14; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_4_REG_2_15; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_4_REG_2_16; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_4_REG_2_17; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_4_REG_2_18; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_4_REG_2_19; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_4_REG_2_20; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_4_REG_2_21; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_4_REG_2_22; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_4_REG_2_23; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_4_REG_2_24; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_4_REG_2_25; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_4_REG_2_26; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_4_REG_2_27; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_4_REG_2_28; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_4_REG_2_29; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_4_REG_2_30; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_4_REG_2_31; // @[ICacheMainPipe.scala 379:69]
  wire  _s2_data_errors_0_4_T_29 = s2_data_errors_0_4_REG_2_0 | s2_data_errors_0_4_REG_2_1 | s2_data_errors_0_4_REG_2_2
     | s2_data_errors_0_4_REG_2_3 | s2_data_errors_0_4_REG_2_4 | s2_data_errors_0_4_REG_2_5 | s2_data_errors_0_4_REG_2_6
     | s2_data_errors_0_4_REG_2_7 | s2_data_errors_0_4_REG_2_8 | s2_data_errors_0_4_REG_2_9 |
    s2_data_errors_0_4_REG_2_10 | s2_data_errors_0_4_REG_2_11 | s2_data_errors_0_4_REG_2_12 |
    s2_data_errors_0_4_REG_2_13 | s2_data_errors_0_4_REG_2_14 | s2_data_errors_0_4_REG_2_15 |
    s2_data_errors_0_4_REG_2_16 | s2_data_errors_0_4_REG_2_17 | s2_data_errors_0_4_REG_2_18 |
    s2_data_errors_0_4_REG_2_19 | s2_data_errors_0_4_REG_2_20 | s2_data_errors_0_4_REG_2_21 |
    s2_data_errors_0_4_REG_2_22 | s2_data_errors_0_4_REG_2_23 | s2_data_errors_0_4_REG_2_24 |
    s2_data_errors_0_4_REG_2_25 | s2_data_errors_0_4_REG_2_26 | s2_data_errors_0_4_REG_2_27 |
    s2_data_errors_0_4_REG_2_28 | s2_data_errors_0_4_REG_2_29 | s2_data_errors_0_4_REG_2_30; // @[ICacheMainPipe.scala 379:101]
  wire  s2_data_errors_0_4 = s2_data_errors_0_4_REG_1 & (_s2_data_errors_0_4_T_29 | s2_data_errors_0_4_REG_2_31); // @[ICacheMainPipe.scala 379:59]
  reg  s2_data_errors_0_5_REG; // @[ICacheMainPipe.scala 379:48]
  reg  s2_data_errors_0_5_REG_1; // @[ICacheMainPipe.scala 379:40]
  reg  s2_data_errors_0_5_REG_2_0; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_5_REG_2_1; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_5_REG_2_2; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_5_REG_2_3; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_5_REG_2_4; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_5_REG_2_5; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_5_REG_2_6; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_5_REG_2_7; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_5_REG_2_8; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_5_REG_2_9; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_5_REG_2_10; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_5_REG_2_11; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_5_REG_2_12; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_5_REG_2_13; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_5_REG_2_14; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_5_REG_2_15; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_5_REG_2_16; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_5_REG_2_17; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_5_REG_2_18; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_5_REG_2_19; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_5_REG_2_20; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_5_REG_2_21; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_5_REG_2_22; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_5_REG_2_23; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_5_REG_2_24; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_5_REG_2_25; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_5_REG_2_26; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_5_REG_2_27; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_5_REG_2_28; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_5_REG_2_29; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_5_REG_2_30; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_5_REG_2_31; // @[ICacheMainPipe.scala 379:69]
  wire  _s2_data_errors_0_5_T_29 = s2_data_errors_0_5_REG_2_0 | s2_data_errors_0_5_REG_2_1 | s2_data_errors_0_5_REG_2_2
     | s2_data_errors_0_5_REG_2_3 | s2_data_errors_0_5_REG_2_4 | s2_data_errors_0_5_REG_2_5 | s2_data_errors_0_5_REG_2_6
     | s2_data_errors_0_5_REG_2_7 | s2_data_errors_0_5_REG_2_8 | s2_data_errors_0_5_REG_2_9 |
    s2_data_errors_0_5_REG_2_10 | s2_data_errors_0_5_REG_2_11 | s2_data_errors_0_5_REG_2_12 |
    s2_data_errors_0_5_REG_2_13 | s2_data_errors_0_5_REG_2_14 | s2_data_errors_0_5_REG_2_15 |
    s2_data_errors_0_5_REG_2_16 | s2_data_errors_0_5_REG_2_17 | s2_data_errors_0_5_REG_2_18 |
    s2_data_errors_0_5_REG_2_19 | s2_data_errors_0_5_REG_2_20 | s2_data_errors_0_5_REG_2_21 |
    s2_data_errors_0_5_REG_2_22 | s2_data_errors_0_5_REG_2_23 | s2_data_errors_0_5_REG_2_24 |
    s2_data_errors_0_5_REG_2_25 | s2_data_errors_0_5_REG_2_26 | s2_data_errors_0_5_REG_2_27 |
    s2_data_errors_0_5_REG_2_28 | s2_data_errors_0_5_REG_2_29 | s2_data_errors_0_5_REG_2_30; // @[ICacheMainPipe.scala 379:101]
  wire  s2_data_errors_0_5 = s2_data_errors_0_5_REG_1 & (_s2_data_errors_0_5_T_29 | s2_data_errors_0_5_REG_2_31); // @[ICacheMainPipe.scala 379:59]
  reg  s2_data_errors_0_6_REG; // @[ICacheMainPipe.scala 379:48]
  reg  s2_data_errors_0_6_REG_1; // @[ICacheMainPipe.scala 379:40]
  reg  s2_data_errors_0_6_REG_2_0; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_6_REG_2_1; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_6_REG_2_2; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_6_REG_2_3; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_6_REG_2_4; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_6_REG_2_5; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_6_REG_2_6; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_6_REG_2_7; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_6_REG_2_8; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_6_REG_2_9; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_6_REG_2_10; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_6_REG_2_11; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_6_REG_2_12; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_6_REG_2_13; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_6_REG_2_14; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_6_REG_2_15; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_6_REG_2_16; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_6_REG_2_17; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_6_REG_2_18; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_6_REG_2_19; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_6_REG_2_20; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_6_REG_2_21; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_6_REG_2_22; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_6_REG_2_23; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_6_REG_2_24; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_6_REG_2_25; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_6_REG_2_26; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_6_REG_2_27; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_6_REG_2_28; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_6_REG_2_29; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_6_REG_2_30; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_6_REG_2_31; // @[ICacheMainPipe.scala 379:69]
  wire  _s2_data_errors_0_6_T_29 = s2_data_errors_0_6_REG_2_0 | s2_data_errors_0_6_REG_2_1 | s2_data_errors_0_6_REG_2_2
     | s2_data_errors_0_6_REG_2_3 | s2_data_errors_0_6_REG_2_4 | s2_data_errors_0_6_REG_2_5 | s2_data_errors_0_6_REG_2_6
     | s2_data_errors_0_6_REG_2_7 | s2_data_errors_0_6_REG_2_8 | s2_data_errors_0_6_REG_2_9 |
    s2_data_errors_0_6_REG_2_10 | s2_data_errors_0_6_REG_2_11 | s2_data_errors_0_6_REG_2_12 |
    s2_data_errors_0_6_REG_2_13 | s2_data_errors_0_6_REG_2_14 | s2_data_errors_0_6_REG_2_15 |
    s2_data_errors_0_6_REG_2_16 | s2_data_errors_0_6_REG_2_17 | s2_data_errors_0_6_REG_2_18 |
    s2_data_errors_0_6_REG_2_19 | s2_data_errors_0_6_REG_2_20 | s2_data_errors_0_6_REG_2_21 |
    s2_data_errors_0_6_REG_2_22 | s2_data_errors_0_6_REG_2_23 | s2_data_errors_0_6_REG_2_24 |
    s2_data_errors_0_6_REG_2_25 | s2_data_errors_0_6_REG_2_26 | s2_data_errors_0_6_REG_2_27 |
    s2_data_errors_0_6_REG_2_28 | s2_data_errors_0_6_REG_2_29 | s2_data_errors_0_6_REG_2_30; // @[ICacheMainPipe.scala 379:101]
  wire  s2_data_errors_0_6 = s2_data_errors_0_6_REG_1 & (_s2_data_errors_0_6_T_29 | s2_data_errors_0_6_REG_2_31); // @[ICacheMainPipe.scala 379:59]
  reg  s2_data_errors_0_7_REG; // @[ICacheMainPipe.scala 379:48]
  reg  s2_data_errors_0_7_REG_1; // @[ICacheMainPipe.scala 379:40]
  reg  s2_data_errors_0_7_REG_2_0; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_7_REG_2_1; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_7_REG_2_2; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_7_REG_2_3; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_7_REG_2_4; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_7_REG_2_5; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_7_REG_2_6; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_7_REG_2_7; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_7_REG_2_8; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_7_REG_2_9; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_7_REG_2_10; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_7_REG_2_11; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_7_REG_2_12; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_7_REG_2_13; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_7_REG_2_14; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_7_REG_2_15; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_7_REG_2_16; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_7_REG_2_17; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_7_REG_2_18; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_7_REG_2_19; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_7_REG_2_20; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_7_REG_2_21; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_7_REG_2_22; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_7_REG_2_23; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_7_REG_2_24; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_7_REG_2_25; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_7_REG_2_26; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_7_REG_2_27; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_7_REG_2_28; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_7_REG_2_29; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_7_REG_2_30; // @[ICacheMainPipe.scala 379:69]
  reg  s2_data_errors_0_7_REG_2_31; // @[ICacheMainPipe.scala 379:69]
  wire  _s2_data_errors_0_7_T_29 = s2_data_errors_0_7_REG_2_0 | s2_data_errors_0_7_REG_2_1 | s2_data_errors_0_7_REG_2_2
     | s2_data_errors_0_7_REG_2_3 | s2_data_errors_0_7_REG_2_4 | s2_data_errors_0_7_REG_2_5 | s2_data_errors_0_7_REG_2_6
     | s2_data_errors_0_7_REG_2_7 | s2_data_errors_0_7_REG_2_8 | s2_data_errors_0_7_REG_2_9 |
    s2_data_errors_0_7_REG_2_10 | s2_data_errors_0_7_REG_2_11 | s2_data_errors_0_7_REG_2_12 |
    s2_data_errors_0_7_REG_2_13 | s2_data_errors_0_7_REG_2_14 | s2_data_errors_0_7_REG_2_15 |
    s2_data_errors_0_7_REG_2_16 | s2_data_errors_0_7_REG_2_17 | s2_data_errors_0_7_REG_2_18 |
    s2_data_errors_0_7_REG_2_19 | s2_data_errors_0_7_REG_2_20 | s2_data_errors_0_7_REG_2_21 |
    s2_data_errors_0_7_REG_2_22 | s2_data_errors_0_7_REG_2_23 | s2_data_errors_0_7_REG_2_24 |
    s2_data_errors_0_7_REG_2_25 | s2_data_errors_0_7_REG_2_26 | s2_data_errors_0_7_REG_2_27 |
    s2_data_errors_0_7_REG_2_28 | s2_data_errors_0_7_REG_2_29 | s2_data_errors_0_7_REG_2_30; // @[ICacheMainPipe.scala 379:101]
  wire  s2_data_errors_0_7 = s2_data_errors_0_7_REG_1 & (_s2_data_errors_0_7_T_29 | s2_data_errors_0_7_REG_2_31); // @[ICacheMainPipe.scala 379:59]
  wire [4095:0] _read_datas_T_257 = {s2_data_cacheline_1_7,s2_data_cacheline_1_6,s2_data_cacheline_1_5,
    s2_data_cacheline_1_4,s2_data_cacheline_1_3,s2_data_cacheline_1_2,s2_data_cacheline_1_1,s2_data_cacheline_1_0}; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_0_0 = _read_datas_T_257[15:0]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_0_1 = _read_datas_T_257[31:16]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_0_2 = _read_datas_T_257[47:32]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_0_3 = _read_datas_T_257[63:48]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_0_4 = _read_datas_T_257[79:64]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_0_5 = _read_datas_T_257[95:80]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_0_6 = _read_datas_T_257[111:96]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_0_7 = _read_datas_T_257[127:112]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_0_8 = _read_datas_T_257[143:128]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_0_9 = _read_datas_T_257[159:144]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_0_10 = _read_datas_T_257[175:160]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_0_11 = _read_datas_T_257[191:176]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_0_12 = _read_datas_T_257[207:192]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_0_13 = _read_datas_T_257[223:208]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_0_14 = _read_datas_T_257[239:224]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_0_15 = _read_datas_T_257[255:240]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_0_16 = _read_datas_T_257[271:256]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_0_17 = _read_datas_T_257[287:272]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_0_18 = _read_datas_T_257[303:288]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_0_19 = _read_datas_T_257[319:304]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_0_20 = _read_datas_T_257[335:320]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_0_21 = _read_datas_T_257[351:336]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_0_22 = _read_datas_T_257[367:352]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_0_23 = _read_datas_T_257[383:368]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_0_24 = _read_datas_T_257[399:384]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_0_25 = _read_datas_T_257[415:400]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_0_26 = _read_datas_T_257[431:416]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_0_27 = _read_datas_T_257[447:432]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_0_28 = _read_datas_T_257[463:448]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_0_29 = _read_datas_T_257[479:464]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_0_30 = _read_datas_T_257[495:480]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_0_31 = _read_datas_T_257[511:496]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_1_0 = _read_datas_T_257[527:512]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_1_1 = _read_datas_T_257[543:528]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_1_2 = _read_datas_T_257[559:544]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_1_3 = _read_datas_T_257[575:560]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_1_4 = _read_datas_T_257[591:576]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_1_5 = _read_datas_T_257[607:592]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_1_6 = _read_datas_T_257[623:608]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_1_7 = _read_datas_T_257[639:624]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_1_8 = _read_datas_T_257[655:640]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_1_9 = _read_datas_T_257[671:656]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_1_10 = _read_datas_T_257[687:672]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_1_11 = _read_datas_T_257[703:688]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_1_12 = _read_datas_T_257[719:704]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_1_13 = _read_datas_T_257[735:720]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_1_14 = _read_datas_T_257[751:736]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_1_15 = _read_datas_T_257[767:752]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_1_16 = _read_datas_T_257[783:768]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_1_17 = _read_datas_T_257[799:784]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_1_18 = _read_datas_T_257[815:800]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_1_19 = _read_datas_T_257[831:816]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_1_20 = _read_datas_T_257[847:832]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_1_21 = _read_datas_T_257[863:848]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_1_22 = _read_datas_T_257[879:864]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_1_23 = _read_datas_T_257[895:880]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_1_24 = _read_datas_T_257[911:896]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_1_25 = _read_datas_T_257[927:912]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_1_26 = _read_datas_T_257[943:928]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_1_27 = _read_datas_T_257[959:944]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_1_28 = _read_datas_T_257[975:960]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_1_29 = _read_datas_T_257[991:976]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_1_30 = _read_datas_T_257[1007:992]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_1_31 = _read_datas_T_257[1023:1008]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_2_0 = _read_datas_T_257[1039:1024]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_2_1 = _read_datas_T_257[1055:1040]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_2_2 = _read_datas_T_257[1071:1056]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_2_3 = _read_datas_T_257[1087:1072]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_2_4 = _read_datas_T_257[1103:1088]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_2_5 = _read_datas_T_257[1119:1104]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_2_6 = _read_datas_T_257[1135:1120]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_2_7 = _read_datas_T_257[1151:1136]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_2_8 = _read_datas_T_257[1167:1152]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_2_9 = _read_datas_T_257[1183:1168]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_2_10 = _read_datas_T_257[1199:1184]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_2_11 = _read_datas_T_257[1215:1200]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_2_12 = _read_datas_T_257[1231:1216]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_2_13 = _read_datas_T_257[1247:1232]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_2_14 = _read_datas_T_257[1263:1248]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_2_15 = _read_datas_T_257[1279:1264]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_2_16 = _read_datas_T_257[1295:1280]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_2_17 = _read_datas_T_257[1311:1296]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_2_18 = _read_datas_T_257[1327:1312]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_2_19 = _read_datas_T_257[1343:1328]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_2_20 = _read_datas_T_257[1359:1344]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_2_21 = _read_datas_T_257[1375:1360]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_2_22 = _read_datas_T_257[1391:1376]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_2_23 = _read_datas_T_257[1407:1392]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_2_24 = _read_datas_T_257[1423:1408]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_2_25 = _read_datas_T_257[1439:1424]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_2_26 = _read_datas_T_257[1455:1440]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_2_27 = _read_datas_T_257[1471:1456]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_2_28 = _read_datas_T_257[1487:1472]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_2_29 = _read_datas_T_257[1503:1488]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_2_30 = _read_datas_T_257[1519:1504]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_2_31 = _read_datas_T_257[1535:1520]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_3_0 = _read_datas_T_257[1551:1536]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_3_1 = _read_datas_T_257[1567:1552]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_3_2 = _read_datas_T_257[1583:1568]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_3_3 = _read_datas_T_257[1599:1584]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_3_4 = _read_datas_T_257[1615:1600]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_3_5 = _read_datas_T_257[1631:1616]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_3_6 = _read_datas_T_257[1647:1632]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_3_7 = _read_datas_T_257[1663:1648]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_3_8 = _read_datas_T_257[1679:1664]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_3_9 = _read_datas_T_257[1695:1680]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_3_10 = _read_datas_T_257[1711:1696]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_3_11 = _read_datas_T_257[1727:1712]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_3_12 = _read_datas_T_257[1743:1728]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_3_13 = _read_datas_T_257[1759:1744]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_3_14 = _read_datas_T_257[1775:1760]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_3_15 = _read_datas_T_257[1791:1776]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_3_16 = _read_datas_T_257[1807:1792]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_3_17 = _read_datas_T_257[1823:1808]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_3_18 = _read_datas_T_257[1839:1824]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_3_19 = _read_datas_T_257[1855:1840]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_3_20 = _read_datas_T_257[1871:1856]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_3_21 = _read_datas_T_257[1887:1872]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_3_22 = _read_datas_T_257[1903:1888]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_3_23 = _read_datas_T_257[1919:1904]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_3_24 = _read_datas_T_257[1935:1920]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_3_25 = _read_datas_T_257[1951:1936]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_3_26 = _read_datas_T_257[1967:1952]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_3_27 = _read_datas_T_257[1983:1968]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_3_28 = _read_datas_T_257[1999:1984]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_3_29 = _read_datas_T_257[2015:2000]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_3_30 = _read_datas_T_257[2031:2016]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_3_31 = _read_datas_T_257[2047:2032]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_4_0 = _read_datas_T_257[2063:2048]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_4_1 = _read_datas_T_257[2079:2064]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_4_2 = _read_datas_T_257[2095:2080]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_4_3 = _read_datas_T_257[2111:2096]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_4_4 = _read_datas_T_257[2127:2112]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_4_5 = _read_datas_T_257[2143:2128]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_4_6 = _read_datas_T_257[2159:2144]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_4_7 = _read_datas_T_257[2175:2160]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_4_8 = _read_datas_T_257[2191:2176]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_4_9 = _read_datas_T_257[2207:2192]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_4_10 = _read_datas_T_257[2223:2208]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_4_11 = _read_datas_T_257[2239:2224]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_4_12 = _read_datas_T_257[2255:2240]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_4_13 = _read_datas_T_257[2271:2256]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_4_14 = _read_datas_T_257[2287:2272]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_4_15 = _read_datas_T_257[2303:2288]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_4_16 = _read_datas_T_257[2319:2304]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_4_17 = _read_datas_T_257[2335:2320]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_4_18 = _read_datas_T_257[2351:2336]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_4_19 = _read_datas_T_257[2367:2352]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_4_20 = _read_datas_T_257[2383:2368]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_4_21 = _read_datas_T_257[2399:2384]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_4_22 = _read_datas_T_257[2415:2400]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_4_23 = _read_datas_T_257[2431:2416]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_4_24 = _read_datas_T_257[2447:2432]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_4_25 = _read_datas_T_257[2463:2448]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_4_26 = _read_datas_T_257[2479:2464]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_4_27 = _read_datas_T_257[2495:2480]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_4_28 = _read_datas_T_257[2511:2496]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_4_29 = _read_datas_T_257[2527:2512]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_4_30 = _read_datas_T_257[2543:2528]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_4_31 = _read_datas_T_257[2559:2544]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_5_0 = _read_datas_T_257[2575:2560]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_5_1 = _read_datas_T_257[2591:2576]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_5_2 = _read_datas_T_257[2607:2592]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_5_3 = _read_datas_T_257[2623:2608]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_5_4 = _read_datas_T_257[2639:2624]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_5_5 = _read_datas_T_257[2655:2640]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_5_6 = _read_datas_T_257[2671:2656]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_5_7 = _read_datas_T_257[2687:2672]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_5_8 = _read_datas_T_257[2703:2688]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_5_9 = _read_datas_T_257[2719:2704]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_5_10 = _read_datas_T_257[2735:2720]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_5_11 = _read_datas_T_257[2751:2736]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_5_12 = _read_datas_T_257[2767:2752]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_5_13 = _read_datas_T_257[2783:2768]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_5_14 = _read_datas_T_257[2799:2784]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_5_15 = _read_datas_T_257[2815:2800]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_5_16 = _read_datas_T_257[2831:2816]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_5_17 = _read_datas_T_257[2847:2832]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_5_18 = _read_datas_T_257[2863:2848]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_5_19 = _read_datas_T_257[2879:2864]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_5_20 = _read_datas_T_257[2895:2880]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_5_21 = _read_datas_T_257[2911:2896]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_5_22 = _read_datas_T_257[2927:2912]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_5_23 = _read_datas_T_257[2943:2928]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_5_24 = _read_datas_T_257[2959:2944]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_5_25 = _read_datas_T_257[2975:2960]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_5_26 = _read_datas_T_257[2991:2976]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_5_27 = _read_datas_T_257[3007:2992]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_5_28 = _read_datas_T_257[3023:3008]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_5_29 = _read_datas_T_257[3039:3024]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_5_30 = _read_datas_T_257[3055:3040]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_5_31 = _read_datas_T_257[3071:3056]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_6_0 = _read_datas_T_257[3087:3072]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_6_1 = _read_datas_T_257[3103:3088]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_6_2 = _read_datas_T_257[3119:3104]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_6_3 = _read_datas_T_257[3135:3120]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_6_4 = _read_datas_T_257[3151:3136]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_6_5 = _read_datas_T_257[3167:3152]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_6_6 = _read_datas_T_257[3183:3168]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_6_7 = _read_datas_T_257[3199:3184]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_6_8 = _read_datas_T_257[3215:3200]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_6_9 = _read_datas_T_257[3231:3216]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_6_10 = _read_datas_T_257[3247:3232]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_6_11 = _read_datas_T_257[3263:3248]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_6_12 = _read_datas_T_257[3279:3264]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_6_13 = _read_datas_T_257[3295:3280]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_6_14 = _read_datas_T_257[3311:3296]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_6_15 = _read_datas_T_257[3327:3312]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_6_16 = _read_datas_T_257[3343:3328]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_6_17 = _read_datas_T_257[3359:3344]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_6_18 = _read_datas_T_257[3375:3360]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_6_19 = _read_datas_T_257[3391:3376]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_6_20 = _read_datas_T_257[3407:3392]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_6_21 = _read_datas_T_257[3423:3408]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_6_22 = _read_datas_T_257[3439:3424]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_6_23 = _read_datas_T_257[3455:3440]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_6_24 = _read_datas_T_257[3471:3456]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_6_25 = _read_datas_T_257[3487:3472]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_6_26 = _read_datas_T_257[3503:3488]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_6_27 = _read_datas_T_257[3519:3504]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_6_28 = _read_datas_T_257[3535:3520]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_6_29 = _read_datas_T_257[3551:3536]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_6_30 = _read_datas_T_257[3567:3552]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_6_31 = _read_datas_T_257[3583:3568]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_7_0 = _read_datas_T_257[3599:3584]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_7_1 = _read_datas_T_257[3615:3600]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_7_2 = _read_datas_T_257[3631:3616]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_7_3 = _read_datas_T_257[3647:3632]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_7_4 = _read_datas_T_257[3663:3648]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_7_5 = _read_datas_T_257[3679:3664]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_7_6 = _read_datas_T_257[3695:3680]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_7_7 = _read_datas_T_257[3711:3696]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_7_8 = _read_datas_T_257[3727:3712]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_7_9 = _read_datas_T_257[3743:3728]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_7_10 = _read_datas_T_257[3759:3744]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_7_11 = _read_datas_T_257[3775:3760]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_7_12 = _read_datas_T_257[3791:3776]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_7_13 = _read_datas_T_257[3807:3792]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_7_14 = _read_datas_T_257[3823:3808]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_7_15 = _read_datas_T_257[3839:3824]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_7_16 = _read_datas_T_257[3855:3840]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_7_17 = _read_datas_T_257[3871:3856]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_7_18 = _read_datas_T_257[3887:3872]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_7_19 = _read_datas_T_257[3903:3888]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_7_20 = _read_datas_T_257[3919:3904]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_7_21 = _read_datas_T_257[3935:3920]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_7_22 = _read_datas_T_257[3951:3936]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_7_23 = _read_datas_T_257[3967:3952]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_7_24 = _read_datas_T_257[3983:3968]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_7_25 = _read_datas_T_257[3999:3984]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_7_26 = _read_datas_T_257[4015:4000]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_7_27 = _read_datas_T_257[4031:4016]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_7_28 = _read_datas_T_257[4047:4032]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_7_29 = _read_datas_T_257[4063:4048]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_7_30 = _read_datas_T_257[4079:4064]; // @[ICacheMainPipe.scala 369:51]
  wire [15:0] read_datas_1_7_31 = _read_datas_T_257[4095:4080]; // @[ICacheMainPipe.scala 369:51]
  wire [255:0] _read_codes_T_257 = {s2_data_errorBits_1_7,s2_data_errorBits_1_6,s2_data_errorBits_1_5,
    s2_data_errorBits_1_4,s2_data_errorBits_1_3,s2_data_errorBits_1_2,s2_data_errorBits_1_1,s2_data_errorBits_1_0}; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_0_0 = _read_codes_T_257[0]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_0_1 = _read_codes_T_257[1]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_0_2 = _read_codes_T_257[2]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_0_3 = _read_codes_T_257[3]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_0_4 = _read_codes_T_257[4]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_0_5 = _read_codes_T_257[5]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_0_6 = _read_codes_T_257[6]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_0_7 = _read_codes_T_257[7]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_0_8 = _read_codes_T_257[8]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_0_9 = _read_codes_T_257[9]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_0_10 = _read_codes_T_257[10]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_0_11 = _read_codes_T_257[11]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_0_12 = _read_codes_T_257[12]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_0_13 = _read_codes_T_257[13]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_0_14 = _read_codes_T_257[14]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_0_15 = _read_codes_T_257[15]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_0_16 = _read_codes_T_257[16]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_0_17 = _read_codes_T_257[17]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_0_18 = _read_codes_T_257[18]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_0_19 = _read_codes_T_257[19]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_0_20 = _read_codes_T_257[20]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_0_21 = _read_codes_T_257[21]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_0_22 = _read_codes_T_257[22]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_0_23 = _read_codes_T_257[23]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_0_24 = _read_codes_T_257[24]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_0_25 = _read_codes_T_257[25]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_0_26 = _read_codes_T_257[26]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_0_27 = _read_codes_T_257[27]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_0_28 = _read_codes_T_257[28]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_0_29 = _read_codes_T_257[29]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_0_30 = _read_codes_T_257[30]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_0_31 = _read_codes_T_257[31]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_1_0 = _read_codes_T_257[32]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_1_1 = _read_codes_T_257[33]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_1_2 = _read_codes_T_257[34]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_1_3 = _read_codes_T_257[35]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_1_4 = _read_codes_T_257[36]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_1_5 = _read_codes_T_257[37]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_1_6 = _read_codes_T_257[38]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_1_7 = _read_codes_T_257[39]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_1_8 = _read_codes_T_257[40]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_1_9 = _read_codes_T_257[41]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_1_10 = _read_codes_T_257[42]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_1_11 = _read_codes_T_257[43]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_1_12 = _read_codes_T_257[44]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_1_13 = _read_codes_T_257[45]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_1_14 = _read_codes_T_257[46]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_1_15 = _read_codes_T_257[47]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_1_16 = _read_codes_T_257[48]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_1_17 = _read_codes_T_257[49]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_1_18 = _read_codes_T_257[50]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_1_19 = _read_codes_T_257[51]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_1_20 = _read_codes_T_257[52]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_1_21 = _read_codes_T_257[53]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_1_22 = _read_codes_T_257[54]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_1_23 = _read_codes_T_257[55]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_1_24 = _read_codes_T_257[56]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_1_25 = _read_codes_T_257[57]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_1_26 = _read_codes_T_257[58]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_1_27 = _read_codes_T_257[59]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_1_28 = _read_codes_T_257[60]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_1_29 = _read_codes_T_257[61]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_1_30 = _read_codes_T_257[62]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_1_31 = _read_codes_T_257[63]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_2_0 = _read_codes_T_257[64]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_2_1 = _read_codes_T_257[65]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_2_2 = _read_codes_T_257[66]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_2_3 = _read_codes_T_257[67]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_2_4 = _read_codes_T_257[68]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_2_5 = _read_codes_T_257[69]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_2_6 = _read_codes_T_257[70]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_2_7 = _read_codes_T_257[71]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_2_8 = _read_codes_T_257[72]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_2_9 = _read_codes_T_257[73]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_2_10 = _read_codes_T_257[74]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_2_11 = _read_codes_T_257[75]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_2_12 = _read_codes_T_257[76]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_2_13 = _read_codes_T_257[77]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_2_14 = _read_codes_T_257[78]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_2_15 = _read_codes_T_257[79]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_2_16 = _read_codes_T_257[80]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_2_17 = _read_codes_T_257[81]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_2_18 = _read_codes_T_257[82]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_2_19 = _read_codes_T_257[83]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_2_20 = _read_codes_T_257[84]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_2_21 = _read_codes_T_257[85]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_2_22 = _read_codes_T_257[86]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_2_23 = _read_codes_T_257[87]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_2_24 = _read_codes_T_257[88]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_2_25 = _read_codes_T_257[89]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_2_26 = _read_codes_T_257[90]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_2_27 = _read_codes_T_257[91]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_2_28 = _read_codes_T_257[92]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_2_29 = _read_codes_T_257[93]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_2_30 = _read_codes_T_257[94]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_2_31 = _read_codes_T_257[95]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_3_0 = _read_codes_T_257[96]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_3_1 = _read_codes_T_257[97]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_3_2 = _read_codes_T_257[98]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_3_3 = _read_codes_T_257[99]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_3_4 = _read_codes_T_257[100]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_3_5 = _read_codes_T_257[101]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_3_6 = _read_codes_T_257[102]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_3_7 = _read_codes_T_257[103]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_3_8 = _read_codes_T_257[104]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_3_9 = _read_codes_T_257[105]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_3_10 = _read_codes_T_257[106]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_3_11 = _read_codes_T_257[107]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_3_12 = _read_codes_T_257[108]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_3_13 = _read_codes_T_257[109]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_3_14 = _read_codes_T_257[110]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_3_15 = _read_codes_T_257[111]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_3_16 = _read_codes_T_257[112]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_3_17 = _read_codes_T_257[113]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_3_18 = _read_codes_T_257[114]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_3_19 = _read_codes_T_257[115]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_3_20 = _read_codes_T_257[116]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_3_21 = _read_codes_T_257[117]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_3_22 = _read_codes_T_257[118]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_3_23 = _read_codes_T_257[119]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_3_24 = _read_codes_T_257[120]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_3_25 = _read_codes_T_257[121]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_3_26 = _read_codes_T_257[122]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_3_27 = _read_codes_T_257[123]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_3_28 = _read_codes_T_257[124]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_3_29 = _read_codes_T_257[125]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_3_30 = _read_codes_T_257[126]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_3_31 = _read_codes_T_257[127]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_4_0 = _read_codes_T_257[128]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_4_1 = _read_codes_T_257[129]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_4_2 = _read_codes_T_257[130]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_4_3 = _read_codes_T_257[131]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_4_4 = _read_codes_T_257[132]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_4_5 = _read_codes_T_257[133]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_4_6 = _read_codes_T_257[134]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_4_7 = _read_codes_T_257[135]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_4_8 = _read_codes_T_257[136]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_4_9 = _read_codes_T_257[137]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_4_10 = _read_codes_T_257[138]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_4_11 = _read_codes_T_257[139]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_4_12 = _read_codes_T_257[140]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_4_13 = _read_codes_T_257[141]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_4_14 = _read_codes_T_257[142]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_4_15 = _read_codes_T_257[143]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_4_16 = _read_codes_T_257[144]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_4_17 = _read_codes_T_257[145]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_4_18 = _read_codes_T_257[146]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_4_19 = _read_codes_T_257[147]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_4_20 = _read_codes_T_257[148]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_4_21 = _read_codes_T_257[149]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_4_22 = _read_codes_T_257[150]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_4_23 = _read_codes_T_257[151]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_4_24 = _read_codes_T_257[152]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_4_25 = _read_codes_T_257[153]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_4_26 = _read_codes_T_257[154]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_4_27 = _read_codes_T_257[155]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_4_28 = _read_codes_T_257[156]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_4_29 = _read_codes_T_257[157]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_4_30 = _read_codes_T_257[158]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_4_31 = _read_codes_T_257[159]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_5_0 = _read_codes_T_257[160]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_5_1 = _read_codes_T_257[161]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_5_2 = _read_codes_T_257[162]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_5_3 = _read_codes_T_257[163]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_5_4 = _read_codes_T_257[164]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_5_5 = _read_codes_T_257[165]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_5_6 = _read_codes_T_257[166]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_5_7 = _read_codes_T_257[167]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_5_8 = _read_codes_T_257[168]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_5_9 = _read_codes_T_257[169]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_5_10 = _read_codes_T_257[170]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_5_11 = _read_codes_T_257[171]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_5_12 = _read_codes_T_257[172]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_5_13 = _read_codes_T_257[173]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_5_14 = _read_codes_T_257[174]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_5_15 = _read_codes_T_257[175]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_5_16 = _read_codes_T_257[176]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_5_17 = _read_codes_T_257[177]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_5_18 = _read_codes_T_257[178]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_5_19 = _read_codes_T_257[179]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_5_20 = _read_codes_T_257[180]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_5_21 = _read_codes_T_257[181]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_5_22 = _read_codes_T_257[182]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_5_23 = _read_codes_T_257[183]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_5_24 = _read_codes_T_257[184]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_5_25 = _read_codes_T_257[185]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_5_26 = _read_codes_T_257[186]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_5_27 = _read_codes_T_257[187]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_5_28 = _read_codes_T_257[188]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_5_29 = _read_codes_T_257[189]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_5_30 = _read_codes_T_257[190]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_5_31 = _read_codes_T_257[191]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_6_0 = _read_codes_T_257[192]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_6_1 = _read_codes_T_257[193]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_6_2 = _read_codes_T_257[194]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_6_3 = _read_codes_T_257[195]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_6_4 = _read_codes_T_257[196]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_6_5 = _read_codes_T_257[197]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_6_6 = _read_codes_T_257[198]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_6_7 = _read_codes_T_257[199]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_6_8 = _read_codes_T_257[200]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_6_9 = _read_codes_T_257[201]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_6_10 = _read_codes_T_257[202]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_6_11 = _read_codes_T_257[203]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_6_12 = _read_codes_T_257[204]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_6_13 = _read_codes_T_257[205]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_6_14 = _read_codes_T_257[206]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_6_15 = _read_codes_T_257[207]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_6_16 = _read_codes_T_257[208]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_6_17 = _read_codes_T_257[209]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_6_18 = _read_codes_T_257[210]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_6_19 = _read_codes_T_257[211]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_6_20 = _read_codes_T_257[212]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_6_21 = _read_codes_T_257[213]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_6_22 = _read_codes_T_257[214]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_6_23 = _read_codes_T_257[215]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_6_24 = _read_codes_T_257[216]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_6_25 = _read_codes_T_257[217]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_6_26 = _read_codes_T_257[218]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_6_27 = _read_codes_T_257[219]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_6_28 = _read_codes_T_257[220]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_6_29 = _read_codes_T_257[221]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_6_30 = _read_codes_T_257[222]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_6_31 = _read_codes_T_257[223]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_7_0 = _read_codes_T_257[224]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_7_1 = _read_codes_T_257[225]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_7_2 = _read_codes_T_257[226]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_7_3 = _read_codes_T_257[227]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_7_4 = _read_codes_T_257[228]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_7_5 = _read_codes_T_257[229]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_7_6 = _read_codes_T_257[230]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_7_7 = _read_codes_T_257[231]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_7_8 = _read_codes_T_257[232]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_7_9 = _read_codes_T_257[233]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_7_10 = _read_codes_T_257[234]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_7_11 = _read_codes_T_257[235]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_7_12 = _read_codes_T_257[236]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_7_13 = _read_codes_T_257[237]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_7_14 = _read_codes_T_257[238]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_7_15 = _read_codes_T_257[239]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_7_16 = _read_codes_T_257[240]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_7_17 = _read_codes_T_257[241]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_7_18 = _read_codes_T_257[242]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_7_19 = _read_codes_T_257[243]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_7_20 = _read_codes_T_257[244]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_7_21 = _read_codes_T_257[245]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_7_22 = _read_codes_T_257[246]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_7_23 = _read_codes_T_257[247]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_7_24 = _read_codes_T_257[248]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_7_25 = _read_codes_T_257[249]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_7_26 = _read_codes_T_257[250]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_7_27 = _read_codes_T_257[251]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_7_28 = _read_codes_T_257[252]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_7_29 = _read_codes_T_257[253]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_7_30 = _read_codes_T_257[254]; // @[ICacheMainPipe.scala 370:51]
  wire  read_codes_1_7_31 = _read_codes_T_257[255]; // @[ICacheMainPipe.scala 370:51]
  wire [16:0] data_full_wayBits_1_0_0 = {read_codes_1_0_0,read_datas_1_0_0}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_0_1 = {read_codes_1_0_1,read_datas_1_0_1}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_0_2 = {read_codes_1_0_2,read_datas_1_0_2}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_0_3 = {read_codes_1_0_3,read_datas_1_0_3}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_0_4 = {read_codes_1_0_4,read_datas_1_0_4}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_0_5 = {read_codes_1_0_5,read_datas_1_0_5}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_0_6 = {read_codes_1_0_6,read_datas_1_0_6}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_0_7 = {read_codes_1_0_7,read_datas_1_0_7}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_0_8 = {read_codes_1_0_8,read_datas_1_0_8}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_0_9 = {read_codes_1_0_9,read_datas_1_0_9}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_0_10 = {read_codes_1_0_10,read_datas_1_0_10}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_0_11 = {read_codes_1_0_11,read_datas_1_0_11}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_0_12 = {read_codes_1_0_12,read_datas_1_0_12}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_0_13 = {read_codes_1_0_13,read_datas_1_0_13}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_0_14 = {read_codes_1_0_14,read_datas_1_0_14}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_0_15 = {read_codes_1_0_15,read_datas_1_0_15}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_0_16 = {read_codes_1_0_16,read_datas_1_0_16}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_0_17 = {read_codes_1_0_17,read_datas_1_0_17}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_0_18 = {read_codes_1_0_18,read_datas_1_0_18}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_0_19 = {read_codes_1_0_19,read_datas_1_0_19}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_0_20 = {read_codes_1_0_20,read_datas_1_0_20}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_0_21 = {read_codes_1_0_21,read_datas_1_0_21}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_0_22 = {read_codes_1_0_22,read_datas_1_0_22}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_0_23 = {read_codes_1_0_23,read_datas_1_0_23}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_0_24 = {read_codes_1_0_24,read_datas_1_0_24}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_0_25 = {read_codes_1_0_25,read_datas_1_0_25}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_0_26 = {read_codes_1_0_26,read_datas_1_0_26}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_0_27 = {read_codes_1_0_27,read_datas_1_0_27}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_0_28 = {read_codes_1_0_28,read_datas_1_0_28}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_0_29 = {read_codes_1_0_29,read_datas_1_0_29}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_0_30 = {read_codes_1_0_30,read_datas_1_0_30}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_0_31 = {read_codes_1_0_31,read_datas_1_0_31}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_1_0 = {read_codes_1_1_0,read_datas_1_1_0}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_1_1 = {read_codes_1_1_1,read_datas_1_1_1}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_1_2 = {read_codes_1_1_2,read_datas_1_1_2}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_1_3 = {read_codes_1_1_3,read_datas_1_1_3}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_1_4 = {read_codes_1_1_4,read_datas_1_1_4}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_1_5 = {read_codes_1_1_5,read_datas_1_1_5}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_1_6 = {read_codes_1_1_6,read_datas_1_1_6}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_1_7 = {read_codes_1_1_7,read_datas_1_1_7}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_1_8 = {read_codes_1_1_8,read_datas_1_1_8}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_1_9 = {read_codes_1_1_9,read_datas_1_1_9}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_1_10 = {read_codes_1_1_10,read_datas_1_1_10}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_1_11 = {read_codes_1_1_11,read_datas_1_1_11}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_1_12 = {read_codes_1_1_12,read_datas_1_1_12}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_1_13 = {read_codes_1_1_13,read_datas_1_1_13}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_1_14 = {read_codes_1_1_14,read_datas_1_1_14}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_1_15 = {read_codes_1_1_15,read_datas_1_1_15}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_1_16 = {read_codes_1_1_16,read_datas_1_1_16}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_1_17 = {read_codes_1_1_17,read_datas_1_1_17}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_1_18 = {read_codes_1_1_18,read_datas_1_1_18}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_1_19 = {read_codes_1_1_19,read_datas_1_1_19}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_1_20 = {read_codes_1_1_20,read_datas_1_1_20}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_1_21 = {read_codes_1_1_21,read_datas_1_1_21}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_1_22 = {read_codes_1_1_22,read_datas_1_1_22}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_1_23 = {read_codes_1_1_23,read_datas_1_1_23}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_1_24 = {read_codes_1_1_24,read_datas_1_1_24}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_1_25 = {read_codes_1_1_25,read_datas_1_1_25}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_1_26 = {read_codes_1_1_26,read_datas_1_1_26}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_1_27 = {read_codes_1_1_27,read_datas_1_1_27}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_1_28 = {read_codes_1_1_28,read_datas_1_1_28}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_1_29 = {read_codes_1_1_29,read_datas_1_1_29}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_1_30 = {read_codes_1_1_30,read_datas_1_1_30}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_1_31 = {read_codes_1_1_31,read_datas_1_1_31}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_2_0 = {read_codes_1_2_0,read_datas_1_2_0}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_2_1 = {read_codes_1_2_1,read_datas_1_2_1}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_2_2 = {read_codes_1_2_2,read_datas_1_2_2}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_2_3 = {read_codes_1_2_3,read_datas_1_2_3}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_2_4 = {read_codes_1_2_4,read_datas_1_2_4}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_2_5 = {read_codes_1_2_5,read_datas_1_2_5}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_2_6 = {read_codes_1_2_6,read_datas_1_2_6}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_2_7 = {read_codes_1_2_7,read_datas_1_2_7}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_2_8 = {read_codes_1_2_8,read_datas_1_2_8}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_2_9 = {read_codes_1_2_9,read_datas_1_2_9}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_2_10 = {read_codes_1_2_10,read_datas_1_2_10}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_2_11 = {read_codes_1_2_11,read_datas_1_2_11}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_2_12 = {read_codes_1_2_12,read_datas_1_2_12}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_2_13 = {read_codes_1_2_13,read_datas_1_2_13}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_2_14 = {read_codes_1_2_14,read_datas_1_2_14}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_2_15 = {read_codes_1_2_15,read_datas_1_2_15}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_2_16 = {read_codes_1_2_16,read_datas_1_2_16}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_2_17 = {read_codes_1_2_17,read_datas_1_2_17}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_2_18 = {read_codes_1_2_18,read_datas_1_2_18}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_2_19 = {read_codes_1_2_19,read_datas_1_2_19}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_2_20 = {read_codes_1_2_20,read_datas_1_2_20}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_2_21 = {read_codes_1_2_21,read_datas_1_2_21}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_2_22 = {read_codes_1_2_22,read_datas_1_2_22}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_2_23 = {read_codes_1_2_23,read_datas_1_2_23}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_2_24 = {read_codes_1_2_24,read_datas_1_2_24}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_2_25 = {read_codes_1_2_25,read_datas_1_2_25}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_2_26 = {read_codes_1_2_26,read_datas_1_2_26}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_2_27 = {read_codes_1_2_27,read_datas_1_2_27}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_2_28 = {read_codes_1_2_28,read_datas_1_2_28}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_2_29 = {read_codes_1_2_29,read_datas_1_2_29}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_2_30 = {read_codes_1_2_30,read_datas_1_2_30}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_2_31 = {read_codes_1_2_31,read_datas_1_2_31}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_3_0 = {read_codes_1_3_0,read_datas_1_3_0}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_3_1 = {read_codes_1_3_1,read_datas_1_3_1}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_3_2 = {read_codes_1_3_2,read_datas_1_3_2}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_3_3 = {read_codes_1_3_3,read_datas_1_3_3}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_3_4 = {read_codes_1_3_4,read_datas_1_3_4}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_3_5 = {read_codes_1_3_5,read_datas_1_3_5}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_3_6 = {read_codes_1_3_6,read_datas_1_3_6}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_3_7 = {read_codes_1_3_7,read_datas_1_3_7}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_3_8 = {read_codes_1_3_8,read_datas_1_3_8}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_3_9 = {read_codes_1_3_9,read_datas_1_3_9}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_3_10 = {read_codes_1_3_10,read_datas_1_3_10}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_3_11 = {read_codes_1_3_11,read_datas_1_3_11}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_3_12 = {read_codes_1_3_12,read_datas_1_3_12}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_3_13 = {read_codes_1_3_13,read_datas_1_3_13}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_3_14 = {read_codes_1_3_14,read_datas_1_3_14}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_3_15 = {read_codes_1_3_15,read_datas_1_3_15}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_3_16 = {read_codes_1_3_16,read_datas_1_3_16}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_3_17 = {read_codes_1_3_17,read_datas_1_3_17}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_3_18 = {read_codes_1_3_18,read_datas_1_3_18}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_3_19 = {read_codes_1_3_19,read_datas_1_3_19}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_3_20 = {read_codes_1_3_20,read_datas_1_3_20}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_3_21 = {read_codes_1_3_21,read_datas_1_3_21}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_3_22 = {read_codes_1_3_22,read_datas_1_3_22}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_3_23 = {read_codes_1_3_23,read_datas_1_3_23}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_3_24 = {read_codes_1_3_24,read_datas_1_3_24}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_3_25 = {read_codes_1_3_25,read_datas_1_3_25}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_3_26 = {read_codes_1_3_26,read_datas_1_3_26}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_3_27 = {read_codes_1_3_27,read_datas_1_3_27}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_3_28 = {read_codes_1_3_28,read_datas_1_3_28}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_3_29 = {read_codes_1_3_29,read_datas_1_3_29}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_3_30 = {read_codes_1_3_30,read_datas_1_3_30}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_3_31 = {read_codes_1_3_31,read_datas_1_3_31}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_4_0 = {read_codes_1_4_0,read_datas_1_4_0}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_4_1 = {read_codes_1_4_1,read_datas_1_4_1}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_4_2 = {read_codes_1_4_2,read_datas_1_4_2}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_4_3 = {read_codes_1_4_3,read_datas_1_4_3}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_4_4 = {read_codes_1_4_4,read_datas_1_4_4}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_4_5 = {read_codes_1_4_5,read_datas_1_4_5}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_4_6 = {read_codes_1_4_6,read_datas_1_4_6}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_4_7 = {read_codes_1_4_7,read_datas_1_4_7}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_4_8 = {read_codes_1_4_8,read_datas_1_4_8}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_4_9 = {read_codes_1_4_9,read_datas_1_4_9}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_4_10 = {read_codes_1_4_10,read_datas_1_4_10}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_4_11 = {read_codes_1_4_11,read_datas_1_4_11}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_4_12 = {read_codes_1_4_12,read_datas_1_4_12}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_4_13 = {read_codes_1_4_13,read_datas_1_4_13}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_4_14 = {read_codes_1_4_14,read_datas_1_4_14}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_4_15 = {read_codes_1_4_15,read_datas_1_4_15}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_4_16 = {read_codes_1_4_16,read_datas_1_4_16}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_4_17 = {read_codes_1_4_17,read_datas_1_4_17}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_4_18 = {read_codes_1_4_18,read_datas_1_4_18}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_4_19 = {read_codes_1_4_19,read_datas_1_4_19}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_4_20 = {read_codes_1_4_20,read_datas_1_4_20}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_4_21 = {read_codes_1_4_21,read_datas_1_4_21}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_4_22 = {read_codes_1_4_22,read_datas_1_4_22}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_4_23 = {read_codes_1_4_23,read_datas_1_4_23}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_4_24 = {read_codes_1_4_24,read_datas_1_4_24}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_4_25 = {read_codes_1_4_25,read_datas_1_4_25}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_4_26 = {read_codes_1_4_26,read_datas_1_4_26}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_4_27 = {read_codes_1_4_27,read_datas_1_4_27}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_4_28 = {read_codes_1_4_28,read_datas_1_4_28}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_4_29 = {read_codes_1_4_29,read_datas_1_4_29}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_4_30 = {read_codes_1_4_30,read_datas_1_4_30}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_4_31 = {read_codes_1_4_31,read_datas_1_4_31}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_5_0 = {read_codes_1_5_0,read_datas_1_5_0}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_5_1 = {read_codes_1_5_1,read_datas_1_5_1}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_5_2 = {read_codes_1_5_2,read_datas_1_5_2}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_5_3 = {read_codes_1_5_3,read_datas_1_5_3}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_5_4 = {read_codes_1_5_4,read_datas_1_5_4}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_5_5 = {read_codes_1_5_5,read_datas_1_5_5}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_5_6 = {read_codes_1_5_6,read_datas_1_5_6}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_5_7 = {read_codes_1_5_7,read_datas_1_5_7}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_5_8 = {read_codes_1_5_8,read_datas_1_5_8}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_5_9 = {read_codes_1_5_9,read_datas_1_5_9}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_5_10 = {read_codes_1_5_10,read_datas_1_5_10}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_5_11 = {read_codes_1_5_11,read_datas_1_5_11}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_5_12 = {read_codes_1_5_12,read_datas_1_5_12}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_5_13 = {read_codes_1_5_13,read_datas_1_5_13}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_5_14 = {read_codes_1_5_14,read_datas_1_5_14}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_5_15 = {read_codes_1_5_15,read_datas_1_5_15}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_5_16 = {read_codes_1_5_16,read_datas_1_5_16}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_5_17 = {read_codes_1_5_17,read_datas_1_5_17}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_5_18 = {read_codes_1_5_18,read_datas_1_5_18}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_5_19 = {read_codes_1_5_19,read_datas_1_5_19}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_5_20 = {read_codes_1_5_20,read_datas_1_5_20}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_5_21 = {read_codes_1_5_21,read_datas_1_5_21}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_5_22 = {read_codes_1_5_22,read_datas_1_5_22}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_5_23 = {read_codes_1_5_23,read_datas_1_5_23}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_5_24 = {read_codes_1_5_24,read_datas_1_5_24}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_5_25 = {read_codes_1_5_25,read_datas_1_5_25}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_5_26 = {read_codes_1_5_26,read_datas_1_5_26}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_5_27 = {read_codes_1_5_27,read_datas_1_5_27}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_5_28 = {read_codes_1_5_28,read_datas_1_5_28}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_5_29 = {read_codes_1_5_29,read_datas_1_5_29}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_5_30 = {read_codes_1_5_30,read_datas_1_5_30}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_5_31 = {read_codes_1_5_31,read_datas_1_5_31}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_6_0 = {read_codes_1_6_0,read_datas_1_6_0}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_6_1 = {read_codes_1_6_1,read_datas_1_6_1}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_6_2 = {read_codes_1_6_2,read_datas_1_6_2}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_6_3 = {read_codes_1_6_3,read_datas_1_6_3}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_6_4 = {read_codes_1_6_4,read_datas_1_6_4}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_6_5 = {read_codes_1_6_5,read_datas_1_6_5}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_6_6 = {read_codes_1_6_6,read_datas_1_6_6}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_6_7 = {read_codes_1_6_7,read_datas_1_6_7}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_6_8 = {read_codes_1_6_8,read_datas_1_6_8}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_6_9 = {read_codes_1_6_9,read_datas_1_6_9}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_6_10 = {read_codes_1_6_10,read_datas_1_6_10}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_6_11 = {read_codes_1_6_11,read_datas_1_6_11}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_6_12 = {read_codes_1_6_12,read_datas_1_6_12}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_6_13 = {read_codes_1_6_13,read_datas_1_6_13}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_6_14 = {read_codes_1_6_14,read_datas_1_6_14}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_6_15 = {read_codes_1_6_15,read_datas_1_6_15}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_6_16 = {read_codes_1_6_16,read_datas_1_6_16}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_6_17 = {read_codes_1_6_17,read_datas_1_6_17}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_6_18 = {read_codes_1_6_18,read_datas_1_6_18}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_6_19 = {read_codes_1_6_19,read_datas_1_6_19}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_6_20 = {read_codes_1_6_20,read_datas_1_6_20}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_6_21 = {read_codes_1_6_21,read_datas_1_6_21}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_6_22 = {read_codes_1_6_22,read_datas_1_6_22}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_6_23 = {read_codes_1_6_23,read_datas_1_6_23}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_6_24 = {read_codes_1_6_24,read_datas_1_6_24}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_6_25 = {read_codes_1_6_25,read_datas_1_6_25}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_6_26 = {read_codes_1_6_26,read_datas_1_6_26}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_6_27 = {read_codes_1_6_27,read_datas_1_6_27}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_6_28 = {read_codes_1_6_28,read_datas_1_6_28}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_6_29 = {read_codes_1_6_29,read_datas_1_6_29}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_6_30 = {read_codes_1_6_30,read_datas_1_6_30}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_6_31 = {read_codes_1_6_31,read_datas_1_6_31}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_7_0 = {read_codes_1_7_0,read_datas_1_7_0}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_7_1 = {read_codes_1_7_1,read_datas_1_7_1}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_7_2 = {read_codes_1_7_2,read_datas_1_7_2}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_7_3 = {read_codes_1_7_3,read_datas_1_7_3}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_7_4 = {read_codes_1_7_4,read_datas_1_7_4}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_7_5 = {read_codes_1_7_5,read_datas_1_7_5}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_7_6 = {read_codes_1_7_6,read_datas_1_7_6}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_7_7 = {read_codes_1_7_7,read_datas_1_7_7}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_7_8 = {read_codes_1_7_8,read_datas_1_7_8}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_7_9 = {read_codes_1_7_9,read_datas_1_7_9}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_7_10 = {read_codes_1_7_10,read_datas_1_7_10}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_7_11 = {read_codes_1_7_11,read_datas_1_7_11}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_7_12 = {read_codes_1_7_12,read_datas_1_7_12}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_7_13 = {read_codes_1_7_13,read_datas_1_7_13}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_7_14 = {read_codes_1_7_14,read_datas_1_7_14}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_7_15 = {read_codes_1_7_15,read_datas_1_7_15}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_7_16 = {read_codes_1_7_16,read_datas_1_7_16}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_7_17 = {read_codes_1_7_17,read_datas_1_7_17}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_7_18 = {read_codes_1_7_18,read_datas_1_7_18}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_7_19 = {read_codes_1_7_19,read_datas_1_7_19}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_7_20 = {read_codes_1_7_20,read_datas_1_7_20}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_7_21 = {read_codes_1_7_21,read_datas_1_7_21}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_7_22 = {read_codes_1_7_22,read_datas_1_7_22}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_7_23 = {read_codes_1_7_23,read_datas_1_7_23}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_7_24 = {read_codes_1_7_24,read_datas_1_7_24}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_7_25 = {read_codes_1_7_25,read_datas_1_7_25}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_7_26 = {read_codes_1_7_26,read_datas_1_7_26}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_7_27 = {read_codes_1_7_27,read_datas_1_7_27}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_7_28 = {read_codes_1_7_28,read_datas_1_7_28}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_7_29 = {read_codes_1_7_29,read_datas_1_7_29}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_7_30 = {read_codes_1_7_30,read_datas_1_7_30}; // @[Cat.scala 31:58]
  wire [16:0] data_full_wayBits_1_7_31 = {read_codes_1_7_31,read_datas_1_7_31}; // @[Cat.scala 31:58]
  reg  s2_data_errors_1_0_REG; // @[ICacheMainPipe.scala 383:48]
  reg  s2_data_errors_1_0_REG_1; // @[ICacheMainPipe.scala 383:40]
  reg  s2_data_errors_1_0_REG_2; // @[ICacheMainPipe.scala 383:77]
  reg  s2_data_errors_1_0_REG_3; // @[ICacheMainPipe.scala 383:69]
  reg  s2_data_errors_1_0_REG_4_0; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_0_REG_4_1; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_0_REG_4_2; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_0_REG_4_3; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_0_REG_4_4; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_0_REG_4_5; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_0_REG_4_6; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_0_REG_4_7; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_0_REG_4_8; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_0_REG_4_9; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_0_REG_4_10; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_0_REG_4_11; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_0_REG_4_12; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_0_REG_4_13; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_0_REG_4_14; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_0_REG_4_15; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_0_REG_4_16; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_0_REG_4_17; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_0_REG_4_18; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_0_REG_4_19; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_0_REG_4_20; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_0_REG_4_21; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_0_REG_4_22; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_0_REG_4_23; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_0_REG_4_24; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_0_REG_4_25; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_0_REG_4_26; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_0_REG_4_27; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_0_REG_4_28; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_0_REG_4_29; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_0_REG_4_30; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_0_REG_4_31; // @[ICacheMainPipe.scala 383:105]
  wire  _s2_data_errors_1_0_T_30 = s2_data_errors_1_0_REG_4_0 | s2_data_errors_1_0_REG_4_1 | s2_data_errors_1_0_REG_4_2
     | s2_data_errors_1_0_REG_4_3 | s2_data_errors_1_0_REG_4_4 | s2_data_errors_1_0_REG_4_5 | s2_data_errors_1_0_REG_4_6
     | s2_data_errors_1_0_REG_4_7 | s2_data_errors_1_0_REG_4_8 | s2_data_errors_1_0_REG_4_9 |
    s2_data_errors_1_0_REG_4_10 | s2_data_errors_1_0_REG_4_11 | s2_data_errors_1_0_REG_4_12 |
    s2_data_errors_1_0_REG_4_13 | s2_data_errors_1_0_REG_4_14 | s2_data_errors_1_0_REG_4_15 |
    s2_data_errors_1_0_REG_4_16 | s2_data_errors_1_0_REG_4_17 | s2_data_errors_1_0_REG_4_18 |
    s2_data_errors_1_0_REG_4_19 | s2_data_errors_1_0_REG_4_20 | s2_data_errors_1_0_REG_4_21 |
    s2_data_errors_1_0_REG_4_22 | s2_data_errors_1_0_REG_4_23 | s2_data_errors_1_0_REG_4_24 |
    s2_data_errors_1_0_REG_4_25 | s2_data_errors_1_0_REG_4_26 | s2_data_errors_1_0_REG_4_27 |
    s2_data_errors_1_0_REG_4_28 | s2_data_errors_1_0_REG_4_29 | s2_data_errors_1_0_REG_4_30; // @[ICacheMainPipe.scala 383:137]
  wire  s2_data_errors_1_0 = s2_data_errors_1_0_REG_1 & s2_data_errors_1_0_REG_3 & (_s2_data_errors_1_0_T_30 |
    s2_data_errors_1_0_REG_4_31); // @[ICacheMainPipe.scala 383:95]
  reg  s2_data_errors_1_1_REG; // @[ICacheMainPipe.scala 383:48]
  reg  s2_data_errors_1_1_REG_1; // @[ICacheMainPipe.scala 383:40]
  reg  s2_data_errors_1_1_REG_2; // @[ICacheMainPipe.scala 383:77]
  reg  s2_data_errors_1_1_REG_3; // @[ICacheMainPipe.scala 383:69]
  reg  s2_data_errors_1_1_REG_4_0; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_1_REG_4_1; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_1_REG_4_2; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_1_REG_4_3; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_1_REG_4_4; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_1_REG_4_5; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_1_REG_4_6; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_1_REG_4_7; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_1_REG_4_8; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_1_REG_4_9; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_1_REG_4_10; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_1_REG_4_11; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_1_REG_4_12; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_1_REG_4_13; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_1_REG_4_14; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_1_REG_4_15; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_1_REG_4_16; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_1_REG_4_17; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_1_REG_4_18; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_1_REG_4_19; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_1_REG_4_20; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_1_REG_4_21; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_1_REG_4_22; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_1_REG_4_23; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_1_REG_4_24; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_1_REG_4_25; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_1_REG_4_26; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_1_REG_4_27; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_1_REG_4_28; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_1_REG_4_29; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_1_REG_4_30; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_1_REG_4_31; // @[ICacheMainPipe.scala 383:105]
  wire  _s2_data_errors_1_1_T_30 = s2_data_errors_1_1_REG_4_0 | s2_data_errors_1_1_REG_4_1 | s2_data_errors_1_1_REG_4_2
     | s2_data_errors_1_1_REG_4_3 | s2_data_errors_1_1_REG_4_4 | s2_data_errors_1_1_REG_4_5 | s2_data_errors_1_1_REG_4_6
     | s2_data_errors_1_1_REG_4_7 | s2_data_errors_1_1_REG_4_8 | s2_data_errors_1_1_REG_4_9 |
    s2_data_errors_1_1_REG_4_10 | s2_data_errors_1_1_REG_4_11 | s2_data_errors_1_1_REG_4_12 |
    s2_data_errors_1_1_REG_4_13 | s2_data_errors_1_1_REG_4_14 | s2_data_errors_1_1_REG_4_15 |
    s2_data_errors_1_1_REG_4_16 | s2_data_errors_1_1_REG_4_17 | s2_data_errors_1_1_REG_4_18 |
    s2_data_errors_1_1_REG_4_19 | s2_data_errors_1_1_REG_4_20 | s2_data_errors_1_1_REG_4_21 |
    s2_data_errors_1_1_REG_4_22 | s2_data_errors_1_1_REG_4_23 | s2_data_errors_1_1_REG_4_24 |
    s2_data_errors_1_1_REG_4_25 | s2_data_errors_1_1_REG_4_26 | s2_data_errors_1_1_REG_4_27 |
    s2_data_errors_1_1_REG_4_28 | s2_data_errors_1_1_REG_4_29 | s2_data_errors_1_1_REG_4_30; // @[ICacheMainPipe.scala 383:137]
  wire  s2_data_errors_1_1 = s2_data_errors_1_1_REG_1 & s2_data_errors_1_1_REG_3 & (_s2_data_errors_1_1_T_30 |
    s2_data_errors_1_1_REG_4_31); // @[ICacheMainPipe.scala 383:95]
  reg  s2_data_errors_1_2_REG; // @[ICacheMainPipe.scala 383:48]
  reg  s2_data_errors_1_2_REG_1; // @[ICacheMainPipe.scala 383:40]
  reg  s2_data_errors_1_2_REG_2; // @[ICacheMainPipe.scala 383:77]
  reg  s2_data_errors_1_2_REG_3; // @[ICacheMainPipe.scala 383:69]
  reg  s2_data_errors_1_2_REG_4_0; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_2_REG_4_1; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_2_REG_4_2; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_2_REG_4_3; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_2_REG_4_4; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_2_REG_4_5; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_2_REG_4_6; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_2_REG_4_7; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_2_REG_4_8; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_2_REG_4_9; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_2_REG_4_10; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_2_REG_4_11; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_2_REG_4_12; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_2_REG_4_13; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_2_REG_4_14; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_2_REG_4_15; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_2_REG_4_16; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_2_REG_4_17; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_2_REG_4_18; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_2_REG_4_19; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_2_REG_4_20; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_2_REG_4_21; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_2_REG_4_22; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_2_REG_4_23; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_2_REG_4_24; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_2_REG_4_25; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_2_REG_4_26; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_2_REG_4_27; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_2_REG_4_28; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_2_REG_4_29; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_2_REG_4_30; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_2_REG_4_31; // @[ICacheMainPipe.scala 383:105]
  wire  _s2_data_errors_1_2_T_30 = s2_data_errors_1_2_REG_4_0 | s2_data_errors_1_2_REG_4_1 | s2_data_errors_1_2_REG_4_2
     | s2_data_errors_1_2_REG_4_3 | s2_data_errors_1_2_REG_4_4 | s2_data_errors_1_2_REG_4_5 | s2_data_errors_1_2_REG_4_6
     | s2_data_errors_1_2_REG_4_7 | s2_data_errors_1_2_REG_4_8 | s2_data_errors_1_2_REG_4_9 |
    s2_data_errors_1_2_REG_4_10 | s2_data_errors_1_2_REG_4_11 | s2_data_errors_1_2_REG_4_12 |
    s2_data_errors_1_2_REG_4_13 | s2_data_errors_1_2_REG_4_14 | s2_data_errors_1_2_REG_4_15 |
    s2_data_errors_1_2_REG_4_16 | s2_data_errors_1_2_REG_4_17 | s2_data_errors_1_2_REG_4_18 |
    s2_data_errors_1_2_REG_4_19 | s2_data_errors_1_2_REG_4_20 | s2_data_errors_1_2_REG_4_21 |
    s2_data_errors_1_2_REG_4_22 | s2_data_errors_1_2_REG_4_23 | s2_data_errors_1_2_REG_4_24 |
    s2_data_errors_1_2_REG_4_25 | s2_data_errors_1_2_REG_4_26 | s2_data_errors_1_2_REG_4_27 |
    s2_data_errors_1_2_REG_4_28 | s2_data_errors_1_2_REG_4_29 | s2_data_errors_1_2_REG_4_30; // @[ICacheMainPipe.scala 383:137]
  wire  s2_data_errors_1_2 = s2_data_errors_1_2_REG_1 & s2_data_errors_1_2_REG_3 & (_s2_data_errors_1_2_T_30 |
    s2_data_errors_1_2_REG_4_31); // @[ICacheMainPipe.scala 383:95]
  reg  s2_data_errors_1_3_REG; // @[ICacheMainPipe.scala 383:48]
  reg  s2_data_errors_1_3_REG_1; // @[ICacheMainPipe.scala 383:40]
  reg  s2_data_errors_1_3_REG_2; // @[ICacheMainPipe.scala 383:77]
  reg  s2_data_errors_1_3_REG_3; // @[ICacheMainPipe.scala 383:69]
  reg  s2_data_errors_1_3_REG_4_0; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_3_REG_4_1; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_3_REG_4_2; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_3_REG_4_3; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_3_REG_4_4; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_3_REG_4_5; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_3_REG_4_6; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_3_REG_4_7; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_3_REG_4_8; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_3_REG_4_9; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_3_REG_4_10; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_3_REG_4_11; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_3_REG_4_12; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_3_REG_4_13; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_3_REG_4_14; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_3_REG_4_15; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_3_REG_4_16; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_3_REG_4_17; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_3_REG_4_18; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_3_REG_4_19; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_3_REG_4_20; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_3_REG_4_21; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_3_REG_4_22; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_3_REG_4_23; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_3_REG_4_24; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_3_REG_4_25; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_3_REG_4_26; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_3_REG_4_27; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_3_REG_4_28; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_3_REG_4_29; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_3_REG_4_30; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_3_REG_4_31; // @[ICacheMainPipe.scala 383:105]
  wire  _s2_data_errors_1_3_T_30 = s2_data_errors_1_3_REG_4_0 | s2_data_errors_1_3_REG_4_1 | s2_data_errors_1_3_REG_4_2
     | s2_data_errors_1_3_REG_4_3 | s2_data_errors_1_3_REG_4_4 | s2_data_errors_1_3_REG_4_5 | s2_data_errors_1_3_REG_4_6
     | s2_data_errors_1_3_REG_4_7 | s2_data_errors_1_3_REG_4_8 | s2_data_errors_1_3_REG_4_9 |
    s2_data_errors_1_3_REG_4_10 | s2_data_errors_1_3_REG_4_11 | s2_data_errors_1_3_REG_4_12 |
    s2_data_errors_1_3_REG_4_13 | s2_data_errors_1_3_REG_4_14 | s2_data_errors_1_3_REG_4_15 |
    s2_data_errors_1_3_REG_4_16 | s2_data_errors_1_3_REG_4_17 | s2_data_errors_1_3_REG_4_18 |
    s2_data_errors_1_3_REG_4_19 | s2_data_errors_1_3_REG_4_20 | s2_data_errors_1_3_REG_4_21 |
    s2_data_errors_1_3_REG_4_22 | s2_data_errors_1_3_REG_4_23 | s2_data_errors_1_3_REG_4_24 |
    s2_data_errors_1_3_REG_4_25 | s2_data_errors_1_3_REG_4_26 | s2_data_errors_1_3_REG_4_27 |
    s2_data_errors_1_3_REG_4_28 | s2_data_errors_1_3_REG_4_29 | s2_data_errors_1_3_REG_4_30; // @[ICacheMainPipe.scala 383:137]
  wire  s2_data_errors_1_3 = s2_data_errors_1_3_REG_1 & s2_data_errors_1_3_REG_3 & (_s2_data_errors_1_3_T_30 |
    s2_data_errors_1_3_REG_4_31); // @[ICacheMainPipe.scala 383:95]
  reg  s2_data_errors_1_4_REG; // @[ICacheMainPipe.scala 383:48]
  reg  s2_data_errors_1_4_REG_1; // @[ICacheMainPipe.scala 383:40]
  reg  s2_data_errors_1_4_REG_2; // @[ICacheMainPipe.scala 383:77]
  reg  s2_data_errors_1_4_REG_3; // @[ICacheMainPipe.scala 383:69]
  reg  s2_data_errors_1_4_REG_4_0; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_4_REG_4_1; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_4_REG_4_2; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_4_REG_4_3; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_4_REG_4_4; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_4_REG_4_5; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_4_REG_4_6; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_4_REG_4_7; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_4_REG_4_8; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_4_REG_4_9; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_4_REG_4_10; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_4_REG_4_11; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_4_REG_4_12; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_4_REG_4_13; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_4_REG_4_14; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_4_REG_4_15; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_4_REG_4_16; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_4_REG_4_17; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_4_REG_4_18; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_4_REG_4_19; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_4_REG_4_20; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_4_REG_4_21; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_4_REG_4_22; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_4_REG_4_23; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_4_REG_4_24; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_4_REG_4_25; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_4_REG_4_26; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_4_REG_4_27; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_4_REG_4_28; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_4_REG_4_29; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_4_REG_4_30; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_4_REG_4_31; // @[ICacheMainPipe.scala 383:105]
  wire  _s2_data_errors_1_4_T_30 = s2_data_errors_1_4_REG_4_0 | s2_data_errors_1_4_REG_4_1 | s2_data_errors_1_4_REG_4_2
     | s2_data_errors_1_4_REG_4_3 | s2_data_errors_1_4_REG_4_4 | s2_data_errors_1_4_REG_4_5 | s2_data_errors_1_4_REG_4_6
     | s2_data_errors_1_4_REG_4_7 | s2_data_errors_1_4_REG_4_8 | s2_data_errors_1_4_REG_4_9 |
    s2_data_errors_1_4_REG_4_10 | s2_data_errors_1_4_REG_4_11 | s2_data_errors_1_4_REG_4_12 |
    s2_data_errors_1_4_REG_4_13 | s2_data_errors_1_4_REG_4_14 | s2_data_errors_1_4_REG_4_15 |
    s2_data_errors_1_4_REG_4_16 | s2_data_errors_1_4_REG_4_17 | s2_data_errors_1_4_REG_4_18 |
    s2_data_errors_1_4_REG_4_19 | s2_data_errors_1_4_REG_4_20 | s2_data_errors_1_4_REG_4_21 |
    s2_data_errors_1_4_REG_4_22 | s2_data_errors_1_4_REG_4_23 | s2_data_errors_1_4_REG_4_24 |
    s2_data_errors_1_4_REG_4_25 | s2_data_errors_1_4_REG_4_26 | s2_data_errors_1_4_REG_4_27 |
    s2_data_errors_1_4_REG_4_28 | s2_data_errors_1_4_REG_4_29 | s2_data_errors_1_4_REG_4_30; // @[ICacheMainPipe.scala 383:137]
  wire  s2_data_errors_1_4 = s2_data_errors_1_4_REG_1 & s2_data_errors_1_4_REG_3 & (_s2_data_errors_1_4_T_30 |
    s2_data_errors_1_4_REG_4_31); // @[ICacheMainPipe.scala 383:95]
  reg  s2_data_errors_1_5_REG; // @[ICacheMainPipe.scala 383:48]
  reg  s2_data_errors_1_5_REG_1; // @[ICacheMainPipe.scala 383:40]
  reg  s2_data_errors_1_5_REG_2; // @[ICacheMainPipe.scala 383:77]
  reg  s2_data_errors_1_5_REG_3; // @[ICacheMainPipe.scala 383:69]
  reg  s2_data_errors_1_5_REG_4_0; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_5_REG_4_1; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_5_REG_4_2; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_5_REG_4_3; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_5_REG_4_4; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_5_REG_4_5; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_5_REG_4_6; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_5_REG_4_7; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_5_REG_4_8; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_5_REG_4_9; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_5_REG_4_10; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_5_REG_4_11; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_5_REG_4_12; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_5_REG_4_13; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_5_REG_4_14; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_5_REG_4_15; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_5_REG_4_16; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_5_REG_4_17; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_5_REG_4_18; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_5_REG_4_19; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_5_REG_4_20; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_5_REG_4_21; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_5_REG_4_22; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_5_REG_4_23; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_5_REG_4_24; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_5_REG_4_25; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_5_REG_4_26; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_5_REG_4_27; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_5_REG_4_28; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_5_REG_4_29; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_5_REG_4_30; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_5_REG_4_31; // @[ICacheMainPipe.scala 383:105]
  wire  _s2_data_errors_1_5_T_30 = s2_data_errors_1_5_REG_4_0 | s2_data_errors_1_5_REG_4_1 | s2_data_errors_1_5_REG_4_2
     | s2_data_errors_1_5_REG_4_3 | s2_data_errors_1_5_REG_4_4 | s2_data_errors_1_5_REG_4_5 | s2_data_errors_1_5_REG_4_6
     | s2_data_errors_1_5_REG_4_7 | s2_data_errors_1_5_REG_4_8 | s2_data_errors_1_5_REG_4_9 |
    s2_data_errors_1_5_REG_4_10 | s2_data_errors_1_5_REG_4_11 | s2_data_errors_1_5_REG_4_12 |
    s2_data_errors_1_5_REG_4_13 | s2_data_errors_1_5_REG_4_14 | s2_data_errors_1_5_REG_4_15 |
    s2_data_errors_1_5_REG_4_16 | s2_data_errors_1_5_REG_4_17 | s2_data_errors_1_5_REG_4_18 |
    s2_data_errors_1_5_REG_4_19 | s2_data_errors_1_5_REG_4_20 | s2_data_errors_1_5_REG_4_21 |
    s2_data_errors_1_5_REG_4_22 | s2_data_errors_1_5_REG_4_23 | s2_data_errors_1_5_REG_4_24 |
    s2_data_errors_1_5_REG_4_25 | s2_data_errors_1_5_REG_4_26 | s2_data_errors_1_5_REG_4_27 |
    s2_data_errors_1_5_REG_4_28 | s2_data_errors_1_5_REG_4_29 | s2_data_errors_1_5_REG_4_30; // @[ICacheMainPipe.scala 383:137]
  wire  s2_data_errors_1_5 = s2_data_errors_1_5_REG_1 & s2_data_errors_1_5_REG_3 & (_s2_data_errors_1_5_T_30 |
    s2_data_errors_1_5_REG_4_31); // @[ICacheMainPipe.scala 383:95]
  reg  s2_data_errors_1_6_REG; // @[ICacheMainPipe.scala 383:48]
  reg  s2_data_errors_1_6_REG_1; // @[ICacheMainPipe.scala 383:40]
  reg  s2_data_errors_1_6_REG_2; // @[ICacheMainPipe.scala 383:77]
  reg  s2_data_errors_1_6_REG_3; // @[ICacheMainPipe.scala 383:69]
  reg  s2_data_errors_1_6_REG_4_0; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_6_REG_4_1; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_6_REG_4_2; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_6_REG_4_3; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_6_REG_4_4; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_6_REG_4_5; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_6_REG_4_6; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_6_REG_4_7; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_6_REG_4_8; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_6_REG_4_9; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_6_REG_4_10; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_6_REG_4_11; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_6_REG_4_12; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_6_REG_4_13; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_6_REG_4_14; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_6_REG_4_15; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_6_REG_4_16; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_6_REG_4_17; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_6_REG_4_18; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_6_REG_4_19; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_6_REG_4_20; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_6_REG_4_21; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_6_REG_4_22; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_6_REG_4_23; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_6_REG_4_24; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_6_REG_4_25; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_6_REG_4_26; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_6_REG_4_27; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_6_REG_4_28; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_6_REG_4_29; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_6_REG_4_30; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_6_REG_4_31; // @[ICacheMainPipe.scala 383:105]
  wire  _s2_data_errors_1_6_T_30 = s2_data_errors_1_6_REG_4_0 | s2_data_errors_1_6_REG_4_1 | s2_data_errors_1_6_REG_4_2
     | s2_data_errors_1_6_REG_4_3 | s2_data_errors_1_6_REG_4_4 | s2_data_errors_1_6_REG_4_5 | s2_data_errors_1_6_REG_4_6
     | s2_data_errors_1_6_REG_4_7 | s2_data_errors_1_6_REG_4_8 | s2_data_errors_1_6_REG_4_9 |
    s2_data_errors_1_6_REG_4_10 | s2_data_errors_1_6_REG_4_11 | s2_data_errors_1_6_REG_4_12 |
    s2_data_errors_1_6_REG_4_13 | s2_data_errors_1_6_REG_4_14 | s2_data_errors_1_6_REG_4_15 |
    s2_data_errors_1_6_REG_4_16 | s2_data_errors_1_6_REG_4_17 | s2_data_errors_1_6_REG_4_18 |
    s2_data_errors_1_6_REG_4_19 | s2_data_errors_1_6_REG_4_20 | s2_data_errors_1_6_REG_4_21 |
    s2_data_errors_1_6_REG_4_22 | s2_data_errors_1_6_REG_4_23 | s2_data_errors_1_6_REG_4_24 |
    s2_data_errors_1_6_REG_4_25 | s2_data_errors_1_6_REG_4_26 | s2_data_errors_1_6_REG_4_27 |
    s2_data_errors_1_6_REG_4_28 | s2_data_errors_1_6_REG_4_29 | s2_data_errors_1_6_REG_4_30; // @[ICacheMainPipe.scala 383:137]
  wire  s2_data_errors_1_6 = s2_data_errors_1_6_REG_1 & s2_data_errors_1_6_REG_3 & (_s2_data_errors_1_6_T_30 |
    s2_data_errors_1_6_REG_4_31); // @[ICacheMainPipe.scala 383:95]
  reg  s2_data_errors_1_7_REG; // @[ICacheMainPipe.scala 383:48]
  reg  s2_data_errors_1_7_REG_1; // @[ICacheMainPipe.scala 383:40]
  reg  s2_data_errors_1_7_REG_2; // @[ICacheMainPipe.scala 383:77]
  reg  s2_data_errors_1_7_REG_3; // @[ICacheMainPipe.scala 383:69]
  reg  s2_data_errors_1_7_REG_4_0; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_7_REG_4_1; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_7_REG_4_2; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_7_REG_4_3; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_7_REG_4_4; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_7_REG_4_5; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_7_REG_4_6; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_7_REG_4_7; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_7_REG_4_8; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_7_REG_4_9; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_7_REG_4_10; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_7_REG_4_11; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_7_REG_4_12; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_7_REG_4_13; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_7_REG_4_14; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_7_REG_4_15; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_7_REG_4_16; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_7_REG_4_17; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_7_REG_4_18; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_7_REG_4_19; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_7_REG_4_20; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_7_REG_4_21; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_7_REG_4_22; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_7_REG_4_23; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_7_REG_4_24; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_7_REG_4_25; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_7_REG_4_26; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_7_REG_4_27; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_7_REG_4_28; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_7_REG_4_29; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_7_REG_4_30; // @[ICacheMainPipe.scala 383:105]
  reg  s2_data_errors_1_7_REG_4_31; // @[ICacheMainPipe.scala 383:105]
  wire  _s2_data_errors_1_7_T_30 = s2_data_errors_1_7_REG_4_0 | s2_data_errors_1_7_REG_4_1 | s2_data_errors_1_7_REG_4_2
     | s2_data_errors_1_7_REG_4_3 | s2_data_errors_1_7_REG_4_4 | s2_data_errors_1_7_REG_4_5 | s2_data_errors_1_7_REG_4_6
     | s2_data_errors_1_7_REG_4_7 | s2_data_errors_1_7_REG_4_8 | s2_data_errors_1_7_REG_4_9 |
    s2_data_errors_1_7_REG_4_10 | s2_data_errors_1_7_REG_4_11 | s2_data_errors_1_7_REG_4_12 |
    s2_data_errors_1_7_REG_4_13 | s2_data_errors_1_7_REG_4_14 | s2_data_errors_1_7_REG_4_15 |
    s2_data_errors_1_7_REG_4_16 | s2_data_errors_1_7_REG_4_17 | s2_data_errors_1_7_REG_4_18 |
    s2_data_errors_1_7_REG_4_19 | s2_data_errors_1_7_REG_4_20 | s2_data_errors_1_7_REG_4_21 |
    s2_data_errors_1_7_REG_4_22 | s2_data_errors_1_7_REG_4_23 | s2_data_errors_1_7_REG_4_24 |
    s2_data_errors_1_7_REG_4_25 | s2_data_errors_1_7_REG_4_26 | s2_data_errors_1_7_REG_4_27 |
    s2_data_errors_1_7_REG_4_28 | s2_data_errors_1_7_REG_4_29 | s2_data_errors_1_7_REG_4_30; // @[ICacheMainPipe.scala 383:137]
  wire  s2_data_errors_1_7 = s2_data_errors_1_7_REG_1 & s2_data_errors_1_7_REG_3 & (_s2_data_errors_1_7_T_30 |
    s2_data_errors_1_7_REG_4_31); // @[ICacheMainPipe.scala 383:95]
  wire  s2_parity_data_error_0 = (s2_data_errors_0_0 | s2_data_errors_0_1 | s2_data_errors_0_2 | s2_data_errors_0_3 |
    s2_data_errors_0_4 | s2_data_errors_0_5 | s2_data_errors_0_6 | s2_data_errors_0_7) & io_csr_parity_enable; // @[ICacheMainPipe.scala 389:100]
  wire  s2_parity_data_error_1 = (s2_data_errors_1_0 | s2_data_errors_1_1 | s2_data_errors_1_2 | s2_data_errors_1_3 |
    s2_data_errors_1_4 | s2_data_errors_1_5 | s2_data_errors_1_6 | s2_data_errors_1_7) & io_csr_parity_enable; // @[ICacheMainPipe.scala 389:100]
  reg  s2_parity_error_REG; // @[ICacheMainPipe.scala 390:76]
  wire  s2_parity_error_0 = s2_parity_error_REG | s2_parity_data_error_0; // @[ICacheMainPipe.scala 390:102]
  reg  s2_parity_error_REG_1; // @[ICacheMainPipe.scala 390:76]
  wire  s2_parity_error_1 = s2_parity_error_REG_1 | s2_parity_data_error_1; // @[ICacheMainPipe.scala 390:102]
  reg  io_errors_0_valid_REG; // @[ICacheMainPipe.scala 393:83]
  reg  io_errors_0_valid_REG_1; // @[ICacheMainPipe.scala 393:75]
  reg  io_errors_0_valid_REG_2; // @[ICacheMainPipe.scala 393:45]
  reg  io_errors_0_report_to_beu_REG; // @[ICacheMainPipe.scala 394:83]
  reg  io_errors_0_report_to_beu_REG_1; // @[ICacheMainPipe.scala 394:75]
  reg  io_errors_0_report_to_beu_REG_2; // @[ICacheMainPipe.scala 394:45]
  reg [35:0] io_errors_0_paddr_REG; // @[ICacheMainPipe.scala 395:53]
  reg [35:0] io_errors_0_paddr_REG_1; // @[ICacheMainPipe.scala 395:45]
  reg  io_errors_0_source_tag_REG; // @[ICacheMainPipe.scala 397:53]
  reg  io_errors_0_source_tag_REG_1; // @[ICacheMainPipe.scala 397:45]
  reg  io_errors_0_source_data_REG; // @[ICacheMainPipe.scala 398:45]
  reg  io_errors_1_valid_REG; // @[ICacheMainPipe.scala 393:83]
  reg  io_errors_1_valid_REG_1; // @[ICacheMainPipe.scala 393:75]
  reg  io_errors_1_valid_REG_2; // @[ICacheMainPipe.scala 393:45]
  reg  io_errors_1_report_to_beu_REG; // @[ICacheMainPipe.scala 394:83]
  reg  io_errors_1_report_to_beu_REG_1; // @[ICacheMainPipe.scala 394:75]
  reg  io_errors_1_report_to_beu_REG_2; // @[ICacheMainPipe.scala 394:45]
  reg [35:0] io_errors_1_paddr_REG; // @[ICacheMainPipe.scala 395:53]
  reg [35:0] io_errors_1_paddr_REG_1; // @[ICacheMainPipe.scala 395:45]
  reg  io_errors_1_source_tag_REG; // @[ICacheMainPipe.scala 397:53]
  reg  io_errors_1_source_tag_REG_1; // @[ICacheMainPipe.scala 397:45]
  reg  io_errors_1_source_data_REG; // @[ICacheMainPipe.scala 398:45]
  wire  _s2_tlb_need_back_T = tlb_need_back_valid & s1_fire; // @[ICacheMainPipe.scala 408:91]
  reg  s2_tlb_need_back_valid; // @[Hold.scala 40:24]
  wire  _GEN_321 = _s2_ready_T_2 ? 1'h0 : s2_tlb_need_back_valid; // @[Hold.scala 41:20 40:24 41:28]
  wire  _s2_tlb_need_back_T_1 = tlb_need_back_valid_1 & s1_fire; // @[ICacheMainPipe.scala 408:91]
  reg  s2_tlb_need_back_valid_1; // @[Hold.scala 40:24]
  wire  _GEN_324 = _s2_ready_T_2 ? 1'h0 : s2_tlb_need_back_valid_1; // @[Hold.scala 41:20 40:24 41:28]
  wire  pmpExcpAF_0 = io_pmp_0_resp_instr & s2_tlb_need_back_valid; // @[ICacheMainPipe.scala 410:37]
  wire  pmpExcpAF_1 = io_pmp_1_resp_instr & s2_double_line & s2_tlb_need_back_valid_1; // @[ICacheMainPipe.scala 411:55]
  reg  s2_except_pmp_af_REG; // @[ICacheMainPipe.scala 417:63]
  reg  s2_except_pmp_af_r0; // @[Reg.scala 16:16]
  reg  s2_except_pmp_af_r1; // @[Reg.scala 16:16]
  wire  _GEN_331 = s2_except_pmp_af_REG ? pmpExcpAF_0 : s2_except_pmp_af_r0; // @[Reg.scala 16:16 17:{18,22}]
  wire  _GEN_332 = s2_except_pmp_af_REG ? pmpExcpAF_1 : s2_except_pmp_af_r1; // @[Reg.scala 16:16 17:{18,22}]
  wire  s2_has_except = s2_valid & (s2_except_tlb_af_0 | s2_except_tlb_af_1 | (s2_except_pf_0 | s2_except_pf_1)); // @[ICacheMainPipe.scala 421:32]
  wire  _s2_mmio_T_5 = io_pmp_0_resp_mmio & ~s2_except_tlb_af_0 & ~_GEN_331 & ~s2_except_pf_0; // @[ICacheMainPipe.scala 423:105]
  reg  s2_mmio_REG; // @[ICacheMainPipe.scala 423:133]
  reg  s2_mmio_r; // @[Reg.scala 16:16]
  wire  _GEN_333 = s2_mmio_REG ? _s2_mmio_T_5 : s2_mmio_r; // @[Reg.scala 16:16 17:{18,22}]
  wire  s2_mmio = _GEN_333 & s2_valid; // @[ICacheMainPipe.scala 423:153]
  reg [5:0] missSlot_0_m_vSetIdx; // @[ICacheMainPipe.scala 447:40]
  reg [23:0] missSlot_0_m_pTag; // @[ICacheMainPipe.scala 447:40]
  reg [511:0] missSlot_0_m_data; // @[ICacheMainPipe.scala 447:40]
  reg  missSlot_0_m_corrupt; // @[ICacheMainPipe.scala 447:40]
  reg [5:0] missSlot_1_m_vSetIdx; // @[ICacheMainPipe.scala 447:40]
  reg [23:0] missSlot_1_m_pTag; // @[ICacheMainPipe.scala 447:40]
  reg [511:0] missSlot_1_m_data; // @[ICacheMainPipe.scala 447:40]
  reg  missSlot_1_m_corrupt; // @[ICacheMainPipe.scala 447:40]
  wire  cacheline_0_miss = _miss_0_s2_0_T_4 & ~sec_meet_0_miss; // @[ICacheMainPipe.scala 461:42]
  wire  cacheline_1_miss = _miss_0_s2_1_T_4 & ~sec_meet_1_miss; // @[ICacheMainPipe.scala 464:42]
  reg  only_0_miss_REG; // @[ICacheMainPipe.scala 466:34]
  wire  _only_0_miss_T_3 = ~s2_has_except; // @[ICacheMainPipe.scala 466:86]
  wire  _only_0_miss_T_5 = ~s2_mmio; // @[ICacheMainPipe.scala 466:104]
  wire  only_0_miss = only_0_miss_REG & cacheline_0_miss & _s2_fixed_hit_T_4 & ~s2_has_except & ~s2_mmio; // @[ICacheMainPipe.scala 466:101]
  reg  only_0_hit_REG; // @[ICacheMainPipe.scala 467:34]
  wire  only_0_hit = only_0_hit_REG & s2_fixed_hit_vec_0 & _s2_fixed_hit_T_4 & _only_0_miss_T_5; // @[ICacheMainPipe.scala 467:83]
  reg  hit_0_hit_1_REG; // @[ICacheMainPipe.scala 468:34]
  wire  hit_0_hit_1 = hit_0_hit_1_REG & s2_fixed_hit_vec_0 & s2_fixed_hit_vec_1 & s2_double_line & _only_0_miss_T_5; // @[ICacheMainPipe.scala 468:102]
  reg  hit_0_miss_1_REG; // @[ICacheMainPipe.scala 469:34]
  wire  hit_0_miss_1 = hit_0_miss_1_REG & s2_fixed_hit_vec_0 & cacheline_1_miss & s2_double_line & _only_0_miss_T_3 &
    _only_0_miss_T_5; // @[ICacheMainPipe.scala 469:121]
  reg  miss_0_hit_1_REG; // @[ICacheMainPipe.scala 470:34]
  wire  miss_0_hit_1 = miss_0_hit_1_REG & cacheline_0_miss & s2_fixed_hit_vec_1 & s2_double_line & _only_0_miss_T_3 &
    _only_0_miss_T_5; // @[ICacheMainPipe.scala 470:120]
  reg  miss_0_miss_1_REG; // @[ICacheMainPipe.scala 471:34]
  wire  miss_0_miss_1 = miss_0_miss_1_REG & cacheline_0_miss & cacheline_1_miss & s2_double_line & _only_0_miss_T_3 &
    _only_0_miss_T_5; // @[ICacheMainPipe.scala 471:121]
  reg  miss_0_except_1_REG; // @[ICacheMainPipe.scala 474:34]
  wire  miss_0_except_1 = miss_0_except_1_REG & s2_double_line & _hit_0_except_1_T_1 & s2_except_1 & cacheline_0_miss; // @[ICacheMainPipe.scala 474:97]
  reg  miss_0_hit_1_latch_bit; // @[ICacheMainPipe.scala 478:22]
  wire  _miss_0_hit_1_latch_T = ~_s2_ready_T_2; // @[ICacheMainPipe.scala 480:24]
  wire  _GEN_334 = _s2_ready_T_2 ? 1'h0 : miss_0_hit_1_latch_bit; // @[ICacheMainPipe.scala 478:22 481:{35,41}]
  wire  miss_0_hit_1_latch = miss_0_hit_1_latch_bit | miss_0_hit_1; // @[ICacheMainPipe.scala 482:9]
  reg  miss_0_miss_1_latch_bit; // @[ICacheMainPipe.scala 478:22]
  wire  _GEN_337 = _s2_ready_T_2 ? 1'h0 : miss_0_miss_1_latch_bit; // @[ICacheMainPipe.scala 478:22 481:{35,41}]
  wire  miss_0_miss_1_latch = miss_0_miss_1_latch_bit | miss_0_miss_1; // @[ICacheMainPipe.scala 482:9]
  reg  only_0_miss_latch_bit; // @[ICacheMainPipe.scala 478:22]
  wire  _GEN_340 = _s2_ready_T_2 ? 1'h0 : only_0_miss_latch_bit; // @[ICacheMainPipe.scala 478:22 481:{35,41}]
  wire  only_0_miss_latch = only_0_miss_latch_bit | only_0_miss; // @[ICacheMainPipe.scala 482:9]
  reg  hit_0_miss_1_latch_bit; // @[ICacheMainPipe.scala 478:22]
  wire  _GEN_343 = _s2_ready_T_2 ? 1'h0 : hit_0_miss_1_latch_bit; // @[ICacheMainPipe.scala 478:22 481:{35,41}]
  wire  hit_0_miss_1_latch = hit_0_miss_1_latch_bit | hit_0_miss_1; // @[ICacheMainPipe.scala 482:9]
  reg  miss_0_except_1_latch_bit; // @[ICacheMainPipe.scala 478:22]
  wire  _GEN_346 = _s2_ready_T_2 ? 1'h0 : miss_0_except_1_latch_bit; // @[ICacheMainPipe.scala 478:22 481:{35,41}]
  wire  miss_0_except_1_latch = miss_0_except_1_latch_bit | miss_0_except_1; // @[ICacheMainPipe.scala 482:9]
  wire  _GEN_349 = _s2_ready_T_2 ? 1'h0 : except_0_latch_bit; // @[ICacheMainPipe.scala 478:22 481:{35,41}]
  wire  _GEN_352 = _s2_ready_T_2 ? 1'h0 : hit_0_except_1_latch_bit; // @[ICacheMainPipe.scala 478:22 481:{35,41}]
  reg  only_0_hit_latch_bit; // @[ICacheMainPipe.scala 478:22]
  wire  _GEN_355 = _s2_ready_T_2 ? 1'h0 : only_0_hit_latch_bit; // @[ICacheMainPipe.scala 478:22 481:{35,41}]
  wire  only_0_hit_latch = only_0_hit_latch_bit | only_0_hit; // @[ICacheMainPipe.scala 482:9]
  reg  hit_0_hit_1_latch_bit; // @[ICacheMainPipe.scala 478:22]
  wire  _GEN_358 = _s2_ready_T_2 ? 1'h0 : hit_0_hit_1_latch_bit; // @[ICacheMainPipe.scala 478:22 481:{35,41}]
  wire  hit_0_hit_1_latch = hit_0_hit_1_latch_bit | hit_0_hit_1; // @[ICacheMainPipe.scala 482:9]
  wire  _GEN_361 = _s2_ready_T_2 ? 1'h0 : miss_0_s2_0_latch_bit; // @[ICacheMainPipe.scala 478:22 481:{35,41}]
  wire  _GEN_364 = _s2_ready_T_2 ? 1'h0 : miss_0_s2_1_latch_bit; // @[ICacheMainPipe.scala 478:22 481:{35,41}]
  wire  _GEN_367 = _s2_ready_T_2 ? 1'h0 : miss_1_s2_0_latch_bit; // @[ICacheMainPipe.scala 478:22 481:{35,41}]
  wire  _GEN_370 = _s2_ready_T_2 ? 1'h0 : miss_1_s2_1_latch_bit; // @[ICacheMainPipe.scala 478:22 481:{35,41}]
  wire  slot_0_solve = miss_0_s2_0_latch | miss_0_s2_1_latch; // @[ICacheMainPipe.scala 522:38]
  wire  slot_1_solve = miss_1_s2_0_latch | miss_1_s2_1_latch; // @[ICacheMainPipe.scala 523:38]
  wire  _reservedRefillData_0_T = miss_0_s2_0 | miss_0_s2_1; // @[ICacheMainPipe.scala 530:90]
  reg [511:0] reservedRefillData_0_r; // @[Reg.scala 16:16]
  wire [511:0] _GEN_373 = _reservedRefillData_0_T ? missSlot_0_m_data : reservedRefillData_0_r; // @[Reg.scala 16:16 17:{18,22}]
  wire  _reservedRefillData_1_T = miss_1_s2_0 | miss_1_s2_1; // @[ICacheMainPipe.scala 531:90]
  reg [511:0] reservedRefillData_1_r; // @[Reg.scala 16:16]
  wire [511:0] _GEN_374 = _reservedRefillData_1_T ? missSlot_1_m_data : reservedRefillData_1_r; // @[Reg.scala 16:16 17:{18,22}]
  wire  only_pmp_af_0 = _GEN_331 & cacheline_0_miss & _hit_0_except_1_T_1 & s2_valid; // @[ICacheMainPipe.scala 537:78]
  wire  only_pmp_af_1 = _GEN_332 & cacheline_1_miss & ~s2_except_1 & s2_valid & s2_double_line; // @[ICacheMainPipe.scala 538:90]
  wire [3:0] _wait_state_T = io_mshr_0_toMSHR_ready ? 4'h1 : 4'h0; // @[ICacheMainPipe.scala 548:27]
  wire  _T_524 = only_0_miss_latch | miss_0_hit_1_latch; // @[ICacheMainPipe.scala 549:38]
  wire [3:0] _wait_state_T_2 = io_mshr_1_toMSHR_ready ? 4'h1 : 4'h0; // @[ICacheMainPipe.scala 552:27]
  wire [3:0] _wait_state_T_4 = io_mshr_0_toMSHR_ready & io_mshr_1_toMSHR_ready ? 4'h1 : 4'h0; // @[ICacheMainPipe.scala 554:26]
  wire [3:0] _GEN_375 = miss_0_miss_1_latch ? _wait_state_T_4 : wait_state; // @[ICacheMainPipe.scala 553:40 554:20 435:27]
  wire [3:0] _GEN_376 = hit_0_miss_1_latch ? _wait_state_T_2 : _GEN_375; // @[ICacheMainPipe.scala 551:37 552:20]
  wire  _T_527 = miss_0_except_1_latch | only_0_miss_latch; // @[ICacheMainPipe.scala 563:34]
  wire [3:0] _GEN_380 = miss_0_miss_1_latch ? 4'h3 : wait_state; // @[ICacheMainPipe.scala 565:40 566:20 435:27]
  wire [3:0] _GEN_382 = hit_0_miss_1_latch & io_mshr_1_fromMSHR_valid ? 4'h7 : wait_state; // @[ICacheMainPipe.scala 573:60 574:20 435:27]
  wire [3:0] _GEN_383 = (_T_527 | miss_0_hit_1_latch) & io_mshr_0_fromMSHR_valid ? 4'h7 : _GEN_382; // @[ICacheMainPipe.scala 571:101 572:20]
  wire [3:0] _GEN_384 = io_mshr_0_fromMSHR_valid & ~io_mshr_1_fromMSHR_valid ? 4'h5 : wait_state; // @[ICacheMainPipe.scala 583:60 584:20 435:27]
  wire [3:0] _GEN_385 = ~io_mshr_0_fromMSHR_valid & io_mshr_1_fromMSHR_valid ? 4'h4 : _GEN_384; // @[ICacheMainPipe.scala 581:62 582:20]
  wire [3:0] _GEN_386 = io_mshr_0_fromMSHR_valid & io_mshr_1_fromMSHR_valid ? 4'h7 : _GEN_385; // @[ICacheMainPipe.scala 579:53 580:20]
  wire [3:0] _GEN_387 = io_mshr_0_fromMSHR_valid ? 4'h7 : wait_state; // @[ICacheMainPipe.scala 589:31 590:20 435:27]
  wire [3:0] _GEN_388 = io_mshr_1_fromMSHR_valid ? 4'h7 : wait_state; // @[ICacheMainPipe.scala 595:31 596:20 435:27]
  wire [3:0] _GEN_389 = _s2_ready_T_2 ? 4'h0 : wait_state; // @[ICacheMainPipe.scala 435:27 600:{36,48}]
  wire [3:0] _GEN_390 = 4'h7 == wait_state ? _GEN_389 : wait_state; // @[ICacheMainPipe.scala 540:21 435:27]
  wire [3:0] _GEN_391 = 4'h5 == wait_state ? _GEN_388 : _GEN_390; // @[ICacheMainPipe.scala 540:21]
  wire [3:0] _GEN_392 = 4'h4 == wait_state ? _GEN_387 : _GEN_391; // @[ICacheMainPipe.scala 540:21]
  wire [3:0] _GEN_393 = 4'h3 == wait_state ? _GEN_386 : _GEN_392; // @[ICacheMainPipe.scala 540:21]
  wire  _io_mshr_0_toMSHR_valid_T_3 = wait_state == 4'h1; // @[ICacheMainPipe.scala 609:141]
  wire  _T_544 = io_mshr_0_toMSHR_ready & io_mshr_0_toMSHR_valid; // @[Decoupled.scala 50:35]
  wire [2:0] _GEN_398 = _T_544 & _s2_miss_available_T ? 3'h1 : missStateQueue_0; // @[ICacheMainPipe.scala 616:62 617:29 449:31]
  wire [2:0] _GEN_401 = io_mshr_0_fromMSHR_valid & missStateQueue_0 == 3'h1 ? 3'h2 : _GEN_398; // @[ICacheMainPipe.scala 622:63 623:33]
  wire [2:0] _GEN_404 = _s2_ready_T_2 & missStateQueue_0 == 3'h2 ? 3'h4 : _GEN_401; // @[ICacheMainPipe.scala 629:54 630:29]
  wire  _T_553 = ~slot_0_solve; // @[ICacheMainPipe.scala 636:43]
  wire [2:0] _GEN_405 = slot_0_solve & _miss_0_hit_1_latch_T & s2_valid | s2_valid & _T_553 & _miss_0_hit_1_latch_T ? 3'h5
     : _GEN_404; // @[ICacheMainPipe.scala 640:103 641:31]
  wire  _T_564 = missStateQueue_0 == 3'h5; // @[ICacheMainPipe.scala 645:28]
  wire  _T_568 = io_mshr_1_toMSHR_ready & io_mshr_1_toMSHR_valid; // @[Decoupled.scala 50:35]
  wire [2:0] _GEN_412 = _T_568 & _s2_miss_available_T_3 ? 3'h1 : missStateQueue_1; // @[ICacheMainPipe.scala 616:62 617:29 449:31]
  wire [2:0] _GEN_415 = io_mshr_1_fromMSHR_valid & missStateQueue_1 == 3'h1 ? 3'h2 : _GEN_412; // @[ICacheMainPipe.scala 622:63 623:33]
  wire [2:0] _GEN_418 = _s2_ready_T_2 & missStateQueue_1 == 3'h2 ? 3'h4 : _GEN_415; // @[ICacheMainPipe.scala 629:54 630:29]
  wire  _T_577 = ~slot_1_solve; // @[ICacheMainPipe.scala 636:43]
  wire [2:0] _GEN_419 = slot_1_solve & _miss_0_hit_1_latch_T & s2_valid | s2_valid & _T_577 & _miss_0_hit_1_latch_T ? 3'h5
     : _GEN_418; // @[ICacheMainPipe.scala 640:103 641:31]
  wire  _T_588 = missStateQueue_1 == 3'h5; // @[ICacheMainPipe.scala 645:28]
  wire  _GEN_426 = missSwitchBit & s2_fetch_finish ? 1'h0 : missSwitchBit; // @[ICacheMainPipe.scala 659:47 660:19 133:30]
  wire [511:0] _s2_hit_datas_port_hit_data_T_9 = _touch_ways_0_0_bits_T[0] ? s2_data_cacheline_0_0 : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _s2_hit_datas_port_hit_data_T_10 = _touch_ways_0_0_bits_T[1] ? s2_data_cacheline_0_1 : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _s2_hit_datas_port_hit_data_T_11 = _touch_ways_0_0_bits_T[2] ? s2_data_cacheline_0_2 : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _s2_hit_datas_port_hit_data_T_12 = _touch_ways_0_0_bits_T[3] ? s2_data_cacheline_0_3 : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _s2_hit_datas_port_hit_data_T_13 = _touch_ways_0_0_bits_T[4] ? s2_data_cacheline_0_4 : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _s2_hit_datas_port_hit_data_T_14 = _touch_ways_0_0_bits_T[5] ? s2_data_cacheline_0_5 : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _s2_hit_datas_port_hit_data_T_15 = _touch_ways_0_0_bits_T[6] ? s2_data_cacheline_0_6 : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _s2_hit_datas_port_hit_data_T_16 = _touch_ways_0_0_bits_T[7] ? s2_data_cacheline_0_7 : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _s2_hit_datas_port_hit_data_T_17 = _s2_hit_datas_port_hit_data_T_9 | _s2_hit_datas_port_hit_data_T_10; // @[Mux.scala 27:73]
  wire [511:0] _s2_hit_datas_port_hit_data_T_18 = _s2_hit_datas_port_hit_data_T_17 | _s2_hit_datas_port_hit_data_T_11; // @[Mux.scala 27:73]
  wire [511:0] _s2_hit_datas_port_hit_data_T_19 = _s2_hit_datas_port_hit_data_T_18 | _s2_hit_datas_port_hit_data_T_12; // @[Mux.scala 27:73]
  wire [511:0] _s2_hit_datas_port_hit_data_T_20 = _s2_hit_datas_port_hit_data_T_19 | _s2_hit_datas_port_hit_data_T_13; // @[Mux.scala 27:73]
  wire [511:0] _s2_hit_datas_port_hit_data_T_21 = _s2_hit_datas_port_hit_data_T_20 | _s2_hit_datas_port_hit_data_T_14; // @[Mux.scala 27:73]
  wire [511:0] _s2_hit_datas_port_hit_data_T_22 = _s2_hit_datas_port_hit_data_T_21 | _s2_hit_datas_port_hit_data_T_15; // @[Mux.scala 27:73]
  wire [511:0] _s2_hit_datas_port_hit_data_T_33 = _touch_ways_1_0_bits_T[0] ? s2_data_cacheline_1_0 : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _s2_hit_datas_port_hit_data_T_34 = _touch_ways_1_0_bits_T[1] ? s2_data_cacheline_1_1 : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _s2_hit_datas_port_hit_data_T_35 = _touch_ways_1_0_bits_T[2] ? s2_data_cacheline_1_2 : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _s2_hit_datas_port_hit_data_T_36 = _touch_ways_1_0_bits_T[3] ? s2_data_cacheline_1_3 : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _s2_hit_datas_port_hit_data_T_37 = _touch_ways_1_0_bits_T[4] ? s2_data_cacheline_1_4 : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _s2_hit_datas_port_hit_data_T_38 = _touch_ways_1_0_bits_T[5] ? s2_data_cacheline_1_5 : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _s2_hit_datas_port_hit_data_T_39 = _touch_ways_1_0_bits_T[6] ? s2_data_cacheline_1_6 : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _s2_hit_datas_port_hit_data_T_40 = _touch_ways_1_0_bits_T[7] ? s2_data_cacheline_1_7 : 512'h0; // @[Mux.scala 27:73]
  wire [511:0] _s2_hit_datas_port_hit_data_T_41 = _s2_hit_datas_port_hit_data_T_33 | _s2_hit_datas_port_hit_data_T_34; // @[Mux.scala 27:73]
  wire [511:0] _s2_hit_datas_port_hit_data_T_42 = _s2_hit_datas_port_hit_data_T_41 | _s2_hit_datas_port_hit_data_T_35; // @[Mux.scala 27:73]
  wire [511:0] _s2_hit_datas_port_hit_data_T_43 = _s2_hit_datas_port_hit_data_T_42 | _s2_hit_datas_port_hit_data_T_36; // @[Mux.scala 27:73]
  wire [511:0] _s2_hit_datas_port_hit_data_T_44 = _s2_hit_datas_port_hit_data_T_43 | _s2_hit_datas_port_hit_data_T_37; // @[Mux.scala 27:73]
  wire [511:0] _s2_hit_datas_port_hit_data_T_45 = _s2_hit_datas_port_hit_data_T_44 | _s2_hit_datas_port_hit_data_T_38; // @[Mux.scala 27:73]
  wire [511:0] _s2_hit_datas_port_hit_data_T_46 = _s2_hit_datas_port_hit_data_T_45 | _s2_hit_datas_port_hit_data_T_39; // @[Mux.scala 27:73]
  wire [511:0] _s2_register_datas_0_T = miss_1_s2_0_latch ? _GEN_374 : missSlot_0_m_data; // @[ICacheMainPipe.scala 691:72]
  wire [511:0] _s2_register_datas_1_T = miss_1_s2_1_latch ? _GEN_374 : missSlot_1_m_data; // @[ICacheMainPipe.scala 692:72]
  reg  REG_8; // @[ICacheMainPipe.scala 710:17]
  reg [35:0] io_errors_0_paddr_REG_2; // @[ICacheMainPipe.scala 713:47]
  reg  REG_9; // @[ICacheMainPipe.scala 710:17]
  reg [35:0] io_errors_1_paddr_REG_2; // @[ICacheMainPipe.scala 713:47]
  assign io_metaArray_toIMeta_valid = io_fetch_req_valid & _io_dataArray_toIData_valid_T; // @[ICacheMainPipe.scala 181:42]
  assign io_metaArray_toIMeta_bits_isDoubleLine = io_fetch_req_bits_readValid_0 &
    io_fetch_req_bits_pcMemRead_0_startAddr[5]; // @[ICacheMainPipe.scala 152:84]
  assign io_metaArray_toIMeta_bits_vSetIdx_0 = io_fetch_req_bits_pcMemRead_0_startAddr[11:6]; // @[L1Cache.scala 81:33]
  assign io_metaArray_toIMeta_bits_vSetIdx_1 = io_fetch_req_bits_pcMemRead_0_nextlineStart[11:6]; // @[L1Cache.scala 81:33]
  assign io_dataArray_toIData_valid = io_fetch_req_bits_readValid_3 & ~missSwitchBit; // @[ICacheMainPipe.scala 176:63]
  assign io_dataArray_toIData_bits_0_isDoubleLine = io_fetch_req_bits_readValid_0 &
    io_fetch_req_bits_pcMemRead_0_startAddr[5]; // @[ICacheMainPipe.scala 152:84]
  assign io_dataArray_toIData_bits_0_vSetIdx_0 = io_fetch_req_bits_pcMemRead_0_startAddr[11:6]; // @[L1Cache.scala 81:33]
  assign io_dataArray_toIData_bits_0_vSetIdx_1 = io_fetch_req_bits_pcMemRead_0_nextlineStart[11:6]; // @[L1Cache.scala 81:33]
  assign io_dataArray_toIData_bits_1_isDoubleLine = io_fetch_req_bits_readValid_1 &
    io_fetch_req_bits_pcMemRead_1_startAddr[5]; // @[ICacheMainPipe.scala 152:84]
  assign io_dataArray_toIData_bits_1_vSetIdx_0 = io_fetch_req_bits_pcMemRead_1_startAddr[11:6]; // @[L1Cache.scala 81:33]
  assign io_dataArray_toIData_bits_1_vSetIdx_1 = io_fetch_req_bits_pcMemRead_1_nextlineStart[11:6]; // @[L1Cache.scala 81:33]
  assign io_dataArray_toIData_bits_2_isDoubleLine = io_fetch_req_bits_readValid_2 &
    io_fetch_req_bits_pcMemRead_2_startAddr[5]; // @[ICacheMainPipe.scala 152:84]
  assign io_dataArray_toIData_bits_2_vSetIdx_0 = io_fetch_req_bits_pcMemRead_2_startAddr[11:6]; // @[L1Cache.scala 81:33]
  assign io_dataArray_toIData_bits_2_vSetIdx_1 = io_fetch_req_bits_pcMemRead_2_nextlineStart[11:6]; // @[L1Cache.scala 81:33]
  assign io_dataArray_toIData_bits_3_isDoubleLine = io_fetch_req_bits_readValid_3 &
    io_fetch_req_bits_pcMemRead_3_startAddr[5]; // @[ICacheMainPipe.scala 152:84]
  assign io_dataArray_toIData_bits_3_vSetIdx_0 = io_fetch_req_bits_pcMemRead_3_startAddr[11:6]; // @[L1Cache.scala 81:33]
  assign io_dataArray_toIData_bits_3_vSetIdx_1 = io_fetch_req_bits_pcMemRead_3_nextlineStart[11:6]; // @[L1Cache.scala 81:33]
  assign io_mshr_0_toMSHR_valid = (_T_524 | miss_0_miss_1_latch | miss_0_except_1_latch) & wait_state == 4'h1 &
    _only_0_miss_T_5; // @[ICacheMainPipe.scala 609:162]
  assign io_mshr_0_toMSHR_bits_paddr = s2_req_paddr_0; // @[ICacheMainPipe.scala 610:29]
  assign io_mshr_0_toMSHR_bits_vaddr = s2_req_vaddr_0; // @[ICacheMainPipe.scala 611:29]
  assign io_mshr_0_toMSHR_bits_waymask = s2_waymask_0; // @[ICacheMainPipe.scala 612:29]
  assign io_mshr_1_toMSHR_valid = (hit_0_miss_1_latch | miss_0_miss_1_latch) & _io_mshr_0_toMSHR_valid_T_3 &
    _only_0_miss_T_5; // @[ICacheMainPipe.scala 608:116]
  assign io_mshr_1_toMSHR_bits_paddr = s2_req_paddr_1; // @[ICacheMainPipe.scala 610:29]
  assign io_mshr_1_toMSHR_bits_vaddr = s2_req_vaddr_1; // @[ICacheMainPipe.scala 611:29]
  assign io_mshr_1_toMSHR_bits_waymask = s2_waymask_1; // @[ICacheMainPipe.scala 612:29]
  assign io_errors_0_source_tag = REG_8 ? 1'h0 : io_errors_0_source_tag_REG_1; // @[ICacheMainPipe.scala 397:35 710:52 714:37]
  assign io_errors_0_source_data = REG_8 ? 1'h0 : io_errors_0_source_data_REG; // @[ICacheMainPipe.scala 398:35 710:52 715:37]
  assign io_errors_0_source_l2 = REG_8; // @[ICacheMainPipe.scala 399:35 710:52 716:37]
  assign io_errors_0_paddr = REG_8 ? io_errors_0_paddr_REG_2 : io_errors_0_paddr_REG_1; // @[ICacheMainPipe.scala 395:35 710:52 713:37]
  assign io_errors_0_report_to_beu = REG_8 ? 1'h0 : io_errors_0_report_to_beu_REG_2; // @[ICacheMainPipe.scala 394:35 710:52 712:37]
  assign io_errors_0_valid = REG_8 | io_errors_0_valid_REG_2; // @[ICacheMainPipe.scala 393:35 710:52 711:37]
  assign io_errors_1_source_tag = REG_9 ? 1'h0 : io_errors_1_source_tag_REG_1; // @[ICacheMainPipe.scala 397:35 710:52 714:37]
  assign io_errors_1_source_data = REG_9 ? 1'h0 : io_errors_1_source_data_REG; // @[ICacheMainPipe.scala 398:35 710:52 715:37]
  assign io_errors_1_source_l2 = REG_9; // @[ICacheMainPipe.scala 399:35 710:52 716:37]
  assign io_errors_1_paddr = REG_9 ? io_errors_1_paddr_REG_2 : io_errors_1_paddr_REG_1; // @[ICacheMainPipe.scala 395:35 710:52 713:37]
  assign io_errors_1_report_to_beu = REG_9 ? 1'h0 : io_errors_1_report_to_beu_REG_2; // @[ICacheMainPipe.scala 394:35 710:52 712:37]
  assign io_errors_1_valid = REG_9 | io_errors_1_valid_REG_2; // @[ICacheMainPipe.scala 393:35 710:52 711:37]
  assign io_fetch_req_ready = itlb_can_go & icache_can_go & pipe_can_go; // @[ICacheMainPipe.scala 214:53]
  assign io_fetch_resp_0_valid = _s2_ready_T & _s2_ready_T_1; // @[ICacheMainPipe.scala 338:48]
  assign io_fetch_resp_0_bits_vaddr = s2_req_vaddr_0; // @[ICacheMainPipe.scala 705:29]
  assign io_fetch_resp_0_bits_registerData = miss_0_s2_0_latch ? _GEN_373 : _s2_register_datas_0_T; // @[ICacheMainPipe.scala 691:27]
  assign io_fetch_resp_0_bits_sramData = _s2_hit_datas_port_hit_data_T_22 | _s2_hit_datas_port_hit_data_T_16; // @[Mux.scala 27:73]
  assign io_fetch_resp_0_bits_select = s2_port_hit_0; // @[ICacheMainPipe.scala 703:29]
  assign io_fetch_resp_0_bits_paddr = s2_req_paddr_0; // @[ICacheMainPipe.scala 704:29]
  assign io_fetch_resp_0_bits_tlbExcp_pageFault = s2_except_pf_0; // @[ICacheMainPipe.scala 706:41]
  assign io_fetch_resp_0_bits_tlbExcp_accessFault = s2_except_tlb_af_0 | missSlot_0_m_corrupt | _GEN_331; // @[ICacheMainPipe.scala 707:89]
  assign io_fetch_resp_0_bits_tlbExcp_mmio = _GEN_333 & s2_valid; // @[ICacheMainPipe.scala 423:153]
  assign io_fetch_resp_1_valid = _s2_ready_T_2 & s2_double_line; // @[ICacheMainPipe.scala 699:50]
  assign io_fetch_resp_1_bits_vaddr = s2_req_vaddr_1; // @[ICacheMainPipe.scala 705:29]
  assign io_fetch_resp_1_bits_registerData = miss_0_s2_1_latch ? _GEN_373 : _s2_register_datas_1_T; // @[ICacheMainPipe.scala 692:27]
  assign io_fetch_resp_1_bits_sramData = _s2_hit_datas_port_hit_data_T_46 | _s2_hit_datas_port_hit_data_T_40; // @[Mux.scala 27:73]
  assign io_fetch_resp_1_bits_select = s2_port_hit_1; // @[ICacheMainPipe.scala 703:29]
  assign io_fetch_resp_1_bits_tlbExcp_pageFault = s2_except_pf_1; // @[ICacheMainPipe.scala 706:41]
  assign io_fetch_resp_1_bits_tlbExcp_accessFault = s2_except_tlb_af_1 | missSlot_1_m_corrupt | _GEN_332; // @[ICacheMainPipe.scala 707:89]
  assign io_pmp_0_req_bits_addr = s2_req_paddr_0; // @[ICacheMainPipe.scala 428:21]
  assign io_pmp_1_req_bits_addr = s2_req_paddr_1; // @[ICacheMainPipe.scala 428:21]
  assign io_itlb_0_req_valid = io_fetch_req_valid; // @[ICacheMainPipe.scala 186:27]
  assign io_itlb_0_req_bits_vaddr = io_fetch_req_bits_pcMemRead_4_startAddr; // @[ICacheMainPipe.scala 149:{65,65}]
  assign io_itlb_0_req_bits_kill = ~icache_can_go | ~pipe_can_go; // @[ICacheMainPipe.scala 217:55]
  assign io_itlb_0_resp_ready = tlb_ready_recv_REG | s1_valid & ~tlb_already_recv_0; // @[ICacheMainPipe.scala 244:88]
  assign io_itlb_1_req_valid = io_fetch_req_valid & ftq_req_to_itlb_doubleline; // @[ICacheMainPipe.scala 191:39]
  assign io_itlb_1_req_bits_vaddr = io_fetch_req_bits_pcMemRead_4_nextlineStart; // @[ICacheMainPipe.scala 149:{65,65}]
  assign io_itlb_1_req_bits_kill = ~icache_can_go | ~pipe_can_go; // @[ICacheMainPipe.scala 217:55]
  assign io_itlb_1_resp_ready = tlb_ready_recv_REG_1 | s1_valid & ~tlb_already_recv_1; // @[ICacheMainPipe.scala 244:88]
  assign io_perfInfo_only_0_hit = only_0_hit_latch_bit | only_0_hit; // @[ICacheMainPipe.scala 482:9]
  assign io_perfInfo_only_0_miss = only_0_miss_latch_bit | only_0_miss; // @[ICacheMainPipe.scala 482:9]
  assign io_perfInfo_hit_0_hit_1 = hit_0_hit_1_latch_bit | hit_0_hit_1; // @[ICacheMainPipe.scala 482:9]
  assign io_perfInfo_hit_0_miss_1 = hit_0_miss_1_latch_bit | hit_0_miss_1; // @[ICacheMainPipe.scala 482:9]
  assign io_perfInfo_miss_0_hit_1 = miss_0_hit_1_latch_bit | miss_0_hit_1; // @[ICacheMainPipe.scala 482:9]
  assign io_perfInfo_miss_0_miss_1 = miss_0_miss_1_latch_bit | miss_0_miss_1; // @[ICacheMainPipe.scala 482:9]
  assign io_perfInfo_hit_0_except_1 = hit_0_except_1_latch_bit | hit_0_except_1; // @[ICacheMainPipe.scala 482:9]
  assign io_perfInfo_miss_0_except_1 = miss_0_except_1_latch_bit | miss_0_except_1; // @[ICacheMainPipe.scala 482:9]
  assign io_perfInfo_except_0 = except_0_latch_bit | except_0; // @[ICacheMainPipe.scala 482:9]
  assign io_perfInfo_bank_hit_1 = miss_0_hit_1_latch | hit_0_hit_1_latch; // @[ICacheMainPipe.scala 730:51]
  assign io_perfInfo_hit = hit_0_hit_1_latch | only_0_hit_latch | hit_0_except_1_latch | except_0_latch; // @[ICacheMainPipe.scala 731:94]
  always @(posedge clock) begin
    if (s1_fire) begin // @[Reg.scala 17:18]
      s2_port_hit_0 <= s1_port_hit_0; // @[Reg.scala 17:22]
    end
    miss_0_s2_0_REG <= s1_valid & tlbRespAllValid & s2_ready; // @[ICacheMainPipe.scala 270:43]
    miss_0_s2_0_REG_1 <= missSlot_0_m_vSetIdx == s1_req_vsetIdx_0; // @[ICacheMainPipe.scala 505:41]
    miss_0_s2_0_REG_2 <= missSlot_0_m_pTag == s1_req_ptags_0; // @[ICacheMainPipe.scala 506:39]
    miss_1_s2_0_REG <= s1_valid & tlbRespAllValid & s2_ready; // @[ICacheMainPipe.scala 270:43]
    miss_1_s2_0_REG_1 <= missSlot_1_m_vSetIdx == s1_req_vsetIdx_0; // @[ICacheMainPipe.scala 505:41]
    miss_1_s2_0_REG_2 <= missSlot_1_m_pTag == s1_req_ptags_0; // @[ICacheMainPipe.scala 506:39]
    if (s1_fire) begin // @[Reg.scala 17:18]
      s2_port_hit_1 <= s1_port_hit_1; // @[Reg.scala 17:22]
    end
    miss_0_s2_1_REG <= s1_valid & tlbRespAllValid & s2_ready; // @[ICacheMainPipe.scala 270:43]
    miss_0_s2_1_REG_1 <= missSlot_0_m_vSetIdx == s1_req_vsetIdx_1; // @[ICacheMainPipe.scala 505:41]
    miss_0_s2_1_REG_2 <= missSlot_0_m_pTag == s1_req_ptags_1; // @[ICacheMainPipe.scala 506:39]
    miss_1_s2_1_REG <= s1_valid & tlbRespAllValid & s2_ready; // @[ICacheMainPipe.scala 270:43]
    miss_1_s2_1_REG_1 <= missSlot_1_m_vSetIdx == s1_req_vsetIdx_1; // @[ICacheMainPipe.scala 505:41]
    miss_1_s2_1_REG_2 <= missSlot_1_m_pTag == s1_req_ptags_1; // @[ICacheMainPipe.scala 506:39]
    if (s1_fire) begin // @[Reg.scala 17:18]
      s2_double_line <= s1_double_line; // @[Reg.scala 17:22]
    end
    hit_0_except_1_REG <= s1_valid & tlbRespAllValid & s2_ready; // @[ICacheMainPipe.scala 270:43]
    if (s1_fire) begin // @[Reg.scala 17:18]
      s2_except_pf_0 <= tlbExcpPF_0; // @[Reg.scala 17:22]
    end
    if (s1_fire) begin // @[Reg.scala 17:18]
      s2_except_tlb_af_0 <= tlbExcpAF_0; // @[Reg.scala 17:22]
    end
    if (s1_fire) begin // @[Reg.scala 17:18]
      s2_except_pf_1 <= tlbExcpPF_1; // @[Reg.scala 17:22]
    end
    if (s1_fire) begin // @[Reg.scala 17:18]
      s2_except_tlb_af_1 <= tlbExcpAF_1; // @[Reg.scala 17:22]
    end
    except_0_REG <= s1_valid & tlbRespAllValid & s2_ready; // @[ICacheMainPipe.scala 270:43]
    if (s0_fetch_fire) begin // @[Reg.scala 17:18]
      s1_req_vaddr_0 <= io_fetch_req_bits_pcMemRead_0_startAddr; // @[Reg.scala 17:22]
    end
    if (s0_fetch_fire) begin // @[Reg.scala 17:18]
      s1_req_vaddr_1 <= io_fetch_req_bits_pcMemRead_0_nextlineStart; // @[Reg.scala 17:22]
    end
    if (s0_fetch_fire) begin // @[Reg.scala 17:18]
      s1_req_vsetIdx_0 <= ftq_req_to_data_vset_idx_0_0; // @[Reg.scala 17:22]
    end
    if (s0_fetch_fire) begin // @[Reg.scala 17:18]
      s1_req_vsetIdx_1 <= ftq_req_to_data_vset_idx_0_1; // @[Reg.scala 17:22]
    end
    if (s0_fetch_fire) begin // @[Reg.scala 17:18]
      s1_double_line <= ftq_req_to_data_doubleline_0; // @[Reg.scala 17:22]
    end
    if (tlb_back_0) begin // @[Reg.scala 17:18]
      tlbRespPAddr_r <= io_itlb_0_resp_bits_paddr_0; // @[Reg.scala 17:22]
    end
    if (tlb_back_1) begin // @[Reg.scala 17:18]
      tlbRespPAddr_r1 <= io_itlb_1_resp_bits_paddr_0; // @[Reg.scala 17:22]
    end
    if (tlb_back_0) begin // @[Reg.scala 17:18]
      tlbExcpPF_r <= io_itlb_0_resp_bits_excp_0_pf_instr; // @[Reg.scala 17:22]
    end
    if (tlb_back_1) begin // @[Reg.scala 17:18]
      tlbExcpPF_r1 <= io_itlb_1_resp_bits_excp_0_pf_instr; // @[Reg.scala 17:22]
    end
    if (tlb_back_0) begin // @[Reg.scala 17:18]
      tlbExcpAF_r <= io_itlb_0_resp_bits_excp_0_af_instr; // @[Reg.scala 17:22]
    end
    if (tlb_back_1) begin // @[Reg.scala 17:18]
      tlbExcpAF_r1 <= io_itlb_1_resp_bits_excp_0_af_instr; // @[Reg.scala 17:22]
    end
    s1_meta_ptags_REG <= io_fetch_req_valid & s0_can_go; // @[ICacheMainPipe.scala 215:33]
    if (s1_meta_ptags_REG) begin // @[Reg.scala 17:18]
      s1_meta_ptags_r0_0 <= io_metaArray_fromIMeta_metaData_0_0_tag; // @[Reg.scala 17:22]
    end
    if (s1_meta_ptags_REG) begin // @[Reg.scala 17:18]
      s1_meta_ptags_r0_1 <= io_metaArray_fromIMeta_metaData_0_1_tag; // @[Reg.scala 17:22]
    end
    if (s1_meta_ptags_REG) begin // @[Reg.scala 17:18]
      s1_meta_ptags_r0_2 <= io_metaArray_fromIMeta_metaData_0_2_tag; // @[Reg.scala 17:22]
    end
    if (s1_meta_ptags_REG) begin // @[Reg.scala 17:18]
      s1_meta_ptags_r0_3 <= io_metaArray_fromIMeta_metaData_0_3_tag; // @[Reg.scala 17:22]
    end
    if (s1_meta_ptags_REG) begin // @[Reg.scala 17:18]
      s1_meta_ptags_r0_4 <= io_metaArray_fromIMeta_metaData_0_4_tag; // @[Reg.scala 17:22]
    end
    if (s1_meta_ptags_REG) begin // @[Reg.scala 17:18]
      s1_meta_ptags_r0_5 <= io_metaArray_fromIMeta_metaData_0_5_tag; // @[Reg.scala 17:22]
    end
    if (s1_meta_ptags_REG) begin // @[Reg.scala 17:18]
      s1_meta_ptags_r0_6 <= io_metaArray_fromIMeta_metaData_0_6_tag; // @[Reg.scala 17:22]
    end
    if (s1_meta_ptags_REG) begin // @[Reg.scala 17:18]
      s1_meta_ptags_r0_7 <= io_metaArray_fromIMeta_metaData_0_7_tag; // @[Reg.scala 17:22]
    end
    if (s1_meta_ptags_REG) begin // @[Reg.scala 17:18]
      s1_meta_ptags_r1_0 <= io_metaArray_fromIMeta_metaData_1_0_tag; // @[Reg.scala 17:22]
    end
    if (s1_meta_ptags_REG) begin // @[Reg.scala 17:18]
      s1_meta_ptags_r1_1 <= io_metaArray_fromIMeta_metaData_1_1_tag; // @[Reg.scala 17:22]
    end
    if (s1_meta_ptags_REG) begin // @[Reg.scala 17:18]
      s1_meta_ptags_r1_2 <= io_metaArray_fromIMeta_metaData_1_2_tag; // @[Reg.scala 17:22]
    end
    if (s1_meta_ptags_REG) begin // @[Reg.scala 17:18]
      s1_meta_ptags_r1_3 <= io_metaArray_fromIMeta_metaData_1_3_tag; // @[Reg.scala 17:22]
    end
    if (s1_meta_ptags_REG) begin // @[Reg.scala 17:18]
      s1_meta_ptags_r1_4 <= io_metaArray_fromIMeta_metaData_1_4_tag; // @[Reg.scala 17:22]
    end
    if (s1_meta_ptags_REG) begin // @[Reg.scala 17:18]
      s1_meta_ptags_r1_5 <= io_metaArray_fromIMeta_metaData_1_5_tag; // @[Reg.scala 17:22]
    end
    if (s1_meta_ptags_REG) begin // @[Reg.scala 17:18]
      s1_meta_ptags_r1_6 <= io_metaArray_fromIMeta_metaData_1_6_tag; // @[Reg.scala 17:22]
    end
    if (s1_meta_ptags_REG) begin // @[Reg.scala 17:18]
      s1_meta_ptags_r1_7 <= io_metaArray_fromIMeta_metaData_1_7_tag; // @[Reg.scala 17:22]
    end
    s1_meta_cohs_REG <= io_fetch_req_valid & s0_can_go; // @[ICacheMainPipe.scala 215:33]
    if (s1_meta_cohs_REG) begin // @[Reg.scala 17:18]
      s1_meta_cohs_r0_0_state <= io_metaArray_fromIMeta_metaData_0_0_coh_state; // @[Reg.scala 17:22]
    end
    if (s1_meta_cohs_REG) begin // @[Reg.scala 17:18]
      s1_meta_cohs_r0_1_state <= io_metaArray_fromIMeta_metaData_0_1_coh_state; // @[Reg.scala 17:22]
    end
    if (s1_meta_cohs_REG) begin // @[Reg.scala 17:18]
      s1_meta_cohs_r0_2_state <= io_metaArray_fromIMeta_metaData_0_2_coh_state; // @[Reg.scala 17:22]
    end
    if (s1_meta_cohs_REG) begin // @[Reg.scala 17:18]
      s1_meta_cohs_r0_3_state <= io_metaArray_fromIMeta_metaData_0_3_coh_state; // @[Reg.scala 17:22]
    end
    if (s1_meta_cohs_REG) begin // @[Reg.scala 17:18]
      s1_meta_cohs_r0_4_state <= io_metaArray_fromIMeta_metaData_0_4_coh_state; // @[Reg.scala 17:22]
    end
    if (s1_meta_cohs_REG) begin // @[Reg.scala 17:18]
      s1_meta_cohs_r0_5_state <= io_metaArray_fromIMeta_metaData_0_5_coh_state; // @[Reg.scala 17:22]
    end
    if (s1_meta_cohs_REG) begin // @[Reg.scala 17:18]
      s1_meta_cohs_r0_6_state <= io_metaArray_fromIMeta_metaData_0_6_coh_state; // @[Reg.scala 17:22]
    end
    if (s1_meta_cohs_REG) begin // @[Reg.scala 17:18]
      s1_meta_cohs_r0_7_state <= io_metaArray_fromIMeta_metaData_0_7_coh_state; // @[Reg.scala 17:22]
    end
    if (s1_meta_cohs_REG) begin // @[Reg.scala 17:18]
      s1_meta_cohs_r1_0_state <= io_metaArray_fromIMeta_metaData_1_0_coh_state; // @[Reg.scala 17:22]
    end
    if (s1_meta_cohs_REG) begin // @[Reg.scala 17:18]
      s1_meta_cohs_r1_1_state <= io_metaArray_fromIMeta_metaData_1_1_coh_state; // @[Reg.scala 17:22]
    end
    if (s1_meta_cohs_REG) begin // @[Reg.scala 17:18]
      s1_meta_cohs_r1_2_state <= io_metaArray_fromIMeta_metaData_1_2_coh_state; // @[Reg.scala 17:22]
    end
    if (s1_meta_cohs_REG) begin // @[Reg.scala 17:18]
      s1_meta_cohs_r1_3_state <= io_metaArray_fromIMeta_metaData_1_3_coh_state; // @[Reg.scala 17:22]
    end
    if (s1_meta_cohs_REG) begin // @[Reg.scala 17:18]
      s1_meta_cohs_r1_4_state <= io_metaArray_fromIMeta_metaData_1_4_coh_state; // @[Reg.scala 17:22]
    end
    if (s1_meta_cohs_REG) begin // @[Reg.scala 17:18]
      s1_meta_cohs_r1_5_state <= io_metaArray_fromIMeta_metaData_1_5_coh_state; // @[Reg.scala 17:22]
    end
    if (s1_meta_cohs_REG) begin // @[Reg.scala 17:18]
      s1_meta_cohs_r1_6_state <= io_metaArray_fromIMeta_metaData_1_6_coh_state; // @[Reg.scala 17:22]
    end
    if (s1_meta_cohs_REG) begin // @[Reg.scala 17:18]
      s1_meta_cohs_r1_7_state <= io_metaArray_fromIMeta_metaData_1_7_coh_state; // @[Reg.scala 17:22]
    end
    s1_meta_errors_REG <= io_fetch_req_valid & s0_can_go; // @[ICacheMainPipe.scala 215:33]
    if (s1_meta_errors_REG) begin // @[Reg.scala 17:18]
      s1_meta_errors_r0_0 <= io_metaArray_fromIMeta_errors_0_0; // @[Reg.scala 17:22]
    end
    if (s1_meta_errors_REG) begin // @[Reg.scala 17:18]
      s1_meta_errors_r0_1 <= io_metaArray_fromIMeta_errors_0_1; // @[Reg.scala 17:22]
    end
    if (s1_meta_errors_REG) begin // @[Reg.scala 17:18]
      s1_meta_errors_r0_2 <= io_metaArray_fromIMeta_errors_0_2; // @[Reg.scala 17:22]
    end
    if (s1_meta_errors_REG) begin // @[Reg.scala 17:18]
      s1_meta_errors_r0_3 <= io_metaArray_fromIMeta_errors_0_3; // @[Reg.scala 17:22]
    end
    if (s1_meta_errors_REG) begin // @[Reg.scala 17:18]
      s1_meta_errors_r0_4 <= io_metaArray_fromIMeta_errors_0_4; // @[Reg.scala 17:22]
    end
    if (s1_meta_errors_REG) begin // @[Reg.scala 17:18]
      s1_meta_errors_r0_5 <= io_metaArray_fromIMeta_errors_0_5; // @[Reg.scala 17:22]
    end
    if (s1_meta_errors_REG) begin // @[Reg.scala 17:18]
      s1_meta_errors_r0_6 <= io_metaArray_fromIMeta_errors_0_6; // @[Reg.scala 17:22]
    end
    if (s1_meta_errors_REG) begin // @[Reg.scala 17:18]
      s1_meta_errors_r0_7 <= io_metaArray_fromIMeta_errors_0_7; // @[Reg.scala 17:22]
    end
    if (s1_meta_errors_REG) begin // @[Reg.scala 17:18]
      s1_meta_errors_r1_0 <= io_metaArray_fromIMeta_errors_1_0; // @[Reg.scala 17:22]
    end
    if (s1_meta_errors_REG) begin // @[Reg.scala 17:18]
      s1_meta_errors_r1_1 <= io_metaArray_fromIMeta_errors_1_1; // @[Reg.scala 17:22]
    end
    if (s1_meta_errors_REG) begin // @[Reg.scala 17:18]
      s1_meta_errors_r1_2 <= io_metaArray_fromIMeta_errors_1_2; // @[Reg.scala 17:22]
    end
    if (s1_meta_errors_REG) begin // @[Reg.scala 17:18]
      s1_meta_errors_r1_3 <= io_metaArray_fromIMeta_errors_1_3; // @[Reg.scala 17:22]
    end
    if (s1_meta_errors_REG) begin // @[Reg.scala 17:18]
      s1_meta_errors_r1_4 <= io_metaArray_fromIMeta_errors_1_4; // @[Reg.scala 17:22]
    end
    if (s1_meta_errors_REG) begin // @[Reg.scala 17:18]
      s1_meta_errors_r1_5 <= io_metaArray_fromIMeta_errors_1_5; // @[Reg.scala 17:22]
    end
    if (s1_meta_errors_REG) begin // @[Reg.scala 17:18]
      s1_meta_errors_r1_6 <= io_metaArray_fromIMeta_errors_1_6; // @[Reg.scala 17:22]
    end
    if (s1_meta_errors_REG) begin // @[Reg.scala 17:18]
      s1_meta_errors_r1_7 <= io_metaArray_fromIMeta_errors_1_7; // @[Reg.scala 17:22]
    end
    s1_data_cacheline_REG <= io_fetch_req_valid & s0_can_go; // @[ICacheMainPipe.scala 215:33]
    if (s1_data_cacheline_REG) begin // @[Reg.scala 17:18]
      s1_data_cacheline_r0_0 <= io_dataArray_fromIData_datas_0_0; // @[Reg.scala 17:22]
    end
    if (s1_data_cacheline_REG) begin // @[Reg.scala 17:18]
      s1_data_cacheline_r0_1 <= io_dataArray_fromIData_datas_0_1; // @[Reg.scala 17:22]
    end
    if (s1_data_cacheline_REG) begin // @[Reg.scala 17:18]
      s1_data_cacheline_r0_2 <= io_dataArray_fromIData_datas_0_2; // @[Reg.scala 17:22]
    end
    if (s1_data_cacheline_REG) begin // @[Reg.scala 17:18]
      s1_data_cacheline_r0_3 <= io_dataArray_fromIData_datas_0_3; // @[Reg.scala 17:22]
    end
    if (s1_data_cacheline_REG) begin // @[Reg.scala 17:18]
      s1_data_cacheline_r0_4 <= io_dataArray_fromIData_datas_0_4; // @[Reg.scala 17:22]
    end
    if (s1_data_cacheline_REG) begin // @[Reg.scala 17:18]
      s1_data_cacheline_r0_5 <= io_dataArray_fromIData_datas_0_5; // @[Reg.scala 17:22]
    end
    if (s1_data_cacheline_REG) begin // @[Reg.scala 17:18]
      s1_data_cacheline_r0_6 <= io_dataArray_fromIData_datas_0_6; // @[Reg.scala 17:22]
    end
    if (s1_data_cacheline_REG) begin // @[Reg.scala 17:18]
      s1_data_cacheline_r0_7 <= io_dataArray_fromIData_datas_0_7; // @[Reg.scala 17:22]
    end
    if (s1_data_cacheline_REG) begin // @[Reg.scala 17:18]
      s1_data_cacheline_r1_0 <= io_dataArray_fromIData_datas_1_0; // @[Reg.scala 17:22]
    end
    if (s1_data_cacheline_REG) begin // @[Reg.scala 17:18]
      s1_data_cacheline_r1_1 <= io_dataArray_fromIData_datas_1_1; // @[Reg.scala 17:22]
    end
    if (s1_data_cacheline_REG) begin // @[Reg.scala 17:18]
      s1_data_cacheline_r1_2 <= io_dataArray_fromIData_datas_1_2; // @[Reg.scala 17:22]
    end
    if (s1_data_cacheline_REG) begin // @[Reg.scala 17:18]
      s1_data_cacheline_r1_3 <= io_dataArray_fromIData_datas_1_3; // @[Reg.scala 17:22]
    end
    if (s1_data_cacheline_REG) begin // @[Reg.scala 17:18]
      s1_data_cacheline_r1_4 <= io_dataArray_fromIData_datas_1_4; // @[Reg.scala 17:22]
    end
    if (s1_data_cacheline_REG) begin // @[Reg.scala 17:18]
      s1_data_cacheline_r1_5 <= io_dataArray_fromIData_datas_1_5; // @[Reg.scala 17:22]
    end
    if (s1_data_cacheline_REG) begin // @[Reg.scala 17:18]
      s1_data_cacheline_r1_6 <= io_dataArray_fromIData_datas_1_6; // @[Reg.scala 17:22]
    end
    if (s1_data_cacheline_REG) begin // @[Reg.scala 17:18]
      s1_data_cacheline_r1_7 <= io_dataArray_fromIData_datas_1_7; // @[Reg.scala 17:22]
    end
    s1_data_errorBits_REG <= io_fetch_req_valid & s0_can_go; // @[ICacheMainPipe.scala 215:33]
    if (s1_data_errorBits_REG) begin // @[Reg.scala 17:18]
      s1_data_errorBits_r0_0 <= io_dataArray_fromIData_codes_0_0; // @[Reg.scala 17:22]
    end
    if (s1_data_errorBits_REG) begin // @[Reg.scala 17:18]
      s1_data_errorBits_r0_1 <= io_dataArray_fromIData_codes_0_1; // @[Reg.scala 17:22]
    end
    if (s1_data_errorBits_REG) begin // @[Reg.scala 17:18]
      s1_data_errorBits_r0_2 <= io_dataArray_fromIData_codes_0_2; // @[Reg.scala 17:22]
    end
    if (s1_data_errorBits_REG) begin // @[Reg.scala 17:18]
      s1_data_errorBits_r0_3 <= io_dataArray_fromIData_codes_0_3; // @[Reg.scala 17:22]
    end
    if (s1_data_errorBits_REG) begin // @[Reg.scala 17:18]
      s1_data_errorBits_r0_4 <= io_dataArray_fromIData_codes_0_4; // @[Reg.scala 17:22]
    end
    if (s1_data_errorBits_REG) begin // @[Reg.scala 17:18]
      s1_data_errorBits_r0_5 <= io_dataArray_fromIData_codes_0_5; // @[Reg.scala 17:22]
    end
    if (s1_data_errorBits_REG) begin // @[Reg.scala 17:18]
      s1_data_errorBits_r0_6 <= io_dataArray_fromIData_codes_0_6; // @[Reg.scala 17:22]
    end
    if (s1_data_errorBits_REG) begin // @[Reg.scala 17:18]
      s1_data_errorBits_r0_7 <= io_dataArray_fromIData_codes_0_7; // @[Reg.scala 17:22]
    end
    if (s1_data_errorBits_REG) begin // @[Reg.scala 17:18]
      s1_data_errorBits_r1_0 <= io_dataArray_fromIData_codes_1_0; // @[Reg.scala 17:22]
    end
    if (s1_data_errorBits_REG) begin // @[Reg.scala 17:18]
      s1_data_errorBits_r1_1 <= io_dataArray_fromIData_codes_1_1; // @[Reg.scala 17:22]
    end
    if (s1_data_errorBits_REG) begin // @[Reg.scala 17:18]
      s1_data_errorBits_r1_2 <= io_dataArray_fromIData_codes_1_2; // @[Reg.scala 17:22]
    end
    if (s1_data_errorBits_REG) begin // @[Reg.scala 17:18]
      s1_data_errorBits_r1_3 <= io_dataArray_fromIData_codes_1_3; // @[Reg.scala 17:22]
    end
    if (s1_data_errorBits_REG) begin // @[Reg.scala 17:18]
      s1_data_errorBits_r1_4 <= io_dataArray_fromIData_codes_1_4; // @[Reg.scala 17:22]
    end
    if (s1_data_errorBits_REG) begin // @[Reg.scala 17:18]
      s1_data_errorBits_r1_5 <= io_dataArray_fromIData_codes_1_5; // @[Reg.scala 17:22]
    end
    if (s1_data_errorBits_REG) begin // @[Reg.scala 17:18]
      s1_data_errorBits_r1_6 <= io_dataArray_fromIData_codes_1_6; // @[Reg.scala 17:22]
    end
    if (s1_data_errorBits_REG) begin // @[Reg.scala 17:18]
      s1_data_errorBits_r1_7 <= io_dataArray_fromIData_codes_1_7; // @[Reg.scala 17:22]
    end
    s1_victim_oh_REG <= io_fetch_req_valid & s0_can_go; // @[ICacheMainPipe.scala 215:33]
    if (s1_victim_oh_REG) begin // @[Reg.scala 17:18]
      s1_victim_oh_r0 <= _s1_victim_oh_T_11; // @[Reg.scala 17:22]
    end
    if (s1_victim_oh_REG) begin // @[Reg.scala 17:18]
      s1_victim_oh_r1 <= _s1_victim_oh_T_23; // @[Reg.scala 17:22]
    end
    if (s1_fire) begin // @[Reg.scala 17:18]
      s2_req_vsetIdx_0 <= s1_req_vsetIdx_0; // @[Reg.scala 17:22]
    end
    if (s1_fire) begin // @[Reg.scala 17:18]
      s2_tag_match_vec_0_7 <= s1_tag_match_vec_0_7; // @[Reg.scala 17:22]
    end
    if (s1_fire) begin // @[Reg.scala 17:18]
      s2_tag_match_vec_0_6 <= s1_tag_match_vec_0_6; // @[Reg.scala 17:22]
    end
    if (s1_fire) begin // @[Reg.scala 17:18]
      s2_tag_match_vec_0_5 <= s1_tag_match_vec_0_5; // @[Reg.scala 17:22]
    end
    if (s1_fire) begin // @[Reg.scala 17:18]
      s2_tag_match_vec_0_4 <= s1_tag_match_vec_0_4; // @[Reg.scala 17:22]
    end
    if (s1_fire) begin // @[Reg.scala 17:18]
      s2_tag_match_vec_0_3 <= s1_tag_match_vec_0_3; // @[Reg.scala 17:22]
    end
    if (s1_fire) begin // @[Reg.scala 17:18]
      s2_tag_match_vec_0_2 <= s1_tag_match_vec_0_2; // @[Reg.scala 17:22]
    end
    if (s1_fire) begin // @[Reg.scala 17:18]
      s2_tag_match_vec_0_1 <= s1_tag_match_vec_0_1; // @[Reg.scala 17:22]
    end
    if (s1_fire) begin // @[Reg.scala 17:18]
      s2_tag_match_vec_0_0 <= s1_tag_match_vec_0_0; // @[Reg.scala 17:22]
    end
    if (s1_fire) begin // @[Reg.scala 17:18]
      if (s1_victim_oh_REG) begin // @[Reg.scala 17:18]
        s2_waymask_0 <= _s1_victim_oh_T_11; // @[Reg.scala 17:22]
      end else begin
        s2_waymask_0 <= s1_victim_oh_r0; // @[Reg.scala 16:16]
      end
    end
    if (s1_fire) begin // @[Reg.scala 17:18]
      s2_req_vsetIdx_1 <= s1_req_vsetIdx_1; // @[Reg.scala 17:22]
    end
    if (s1_fire) begin // @[Reg.scala 17:18]
      s2_tag_match_vec_1_7 <= s1_tag_match_vec_1_7; // @[Reg.scala 17:22]
    end
    if (s1_fire) begin // @[Reg.scala 17:18]
      s2_tag_match_vec_1_6 <= s1_tag_match_vec_1_6; // @[Reg.scala 17:22]
    end
    if (s1_fire) begin // @[Reg.scala 17:18]
      s2_tag_match_vec_1_5 <= s1_tag_match_vec_1_5; // @[Reg.scala 17:22]
    end
    if (s1_fire) begin // @[Reg.scala 17:18]
      s2_tag_match_vec_1_4 <= s1_tag_match_vec_1_4; // @[Reg.scala 17:22]
    end
    if (s1_fire) begin // @[Reg.scala 17:18]
      s2_tag_match_vec_1_3 <= s1_tag_match_vec_1_3; // @[Reg.scala 17:22]
    end
    if (s1_fire) begin // @[Reg.scala 17:18]
      s2_tag_match_vec_1_2 <= s1_tag_match_vec_1_2; // @[Reg.scala 17:22]
    end
    if (s1_fire) begin // @[Reg.scala 17:18]
      s2_tag_match_vec_1_1 <= s1_tag_match_vec_1_1; // @[Reg.scala 17:22]
    end
    if (s1_fire) begin // @[Reg.scala 17:18]
      s2_tag_match_vec_1_0 <= s1_tag_match_vec_1_0; // @[Reg.scala 17:22]
    end
    if (s1_fire) begin // @[Reg.scala 17:18]
      if (s1_victim_oh_REG) begin // @[Reg.scala 17:18]
        s2_waymask_1 <= _s1_victim_oh_T_23; // @[Reg.scala 17:22]
      end else begin
        s2_waymask_1 <= s1_victim_oh_r1; // @[Reg.scala 16:16]
      end
    end
    if (s1_fire) begin // @[Reg.scala 17:18]
      if (tlb_back_0) begin // @[Reg.scala 17:18]
        s2_req_paddr_0 <= io_itlb_0_resp_bits_paddr_0; // @[Reg.scala 17:22]
      end else begin
        s2_req_paddr_0 <= tlbRespPAddr_r; // @[Reg.scala 16:16]
      end
    end
    if (s1_fire) begin // @[Reg.scala 17:18]
      if (tlb_back_1) begin // @[Reg.scala 17:18]
        s2_req_paddr_1 <= io_itlb_1_resp_bits_paddr_0; // @[Reg.scala 17:22]
      end else begin
        s2_req_paddr_1 <= tlbRespPAddr_r1; // @[Reg.scala 16:16]
      end
    end
    if (s1_fire) begin // @[Reg.scala 17:18]
      s2_req_vaddr_0 <= s1_req_vaddr_0; // @[Reg.scala 17:22]
    end
    if (s1_fire) begin // @[Reg.scala 17:18]
      s2_req_vaddr_1 <= s1_req_vaddr_1; // @[Reg.scala 17:22]
    end
    if (s1_fire) begin // @[Reg.scala 17:18]
      if (s1_meta_errors_REG) begin // @[Reg.scala 17:18]
        s2_meta_errors_0_0 <= io_metaArray_fromIMeta_errors_0_0; // @[Reg.scala 17:22]
      end else begin
        s2_meta_errors_0_0 <= s1_meta_errors_r0_0; // @[Reg.scala 16:16]
      end
    end
    if (s1_fire) begin // @[Reg.scala 17:18]
      if (s1_meta_errors_REG) begin // @[Reg.scala 17:18]
        s2_meta_errors_0_1 <= io_metaArray_fromIMeta_errors_0_1; // @[Reg.scala 17:22]
      end else begin
        s2_meta_errors_0_1 <= s1_meta_errors_r0_1; // @[Reg.scala 16:16]
      end
    end
    if (s1_fire) begin // @[Reg.scala 17:18]
      if (s1_meta_errors_REG) begin // @[Reg.scala 17:18]
        s2_meta_errors_0_2 <= io_metaArray_fromIMeta_errors_0_2; // @[Reg.scala 17:22]
      end else begin
        s2_meta_errors_0_2 <= s1_meta_errors_r0_2; // @[Reg.scala 16:16]
      end
    end
    if (s1_fire) begin // @[Reg.scala 17:18]
      if (s1_meta_errors_REG) begin // @[Reg.scala 17:18]
        s2_meta_errors_0_3 <= io_metaArray_fromIMeta_errors_0_3; // @[Reg.scala 17:22]
      end else begin
        s2_meta_errors_0_3 <= s1_meta_errors_r0_3; // @[Reg.scala 16:16]
      end
    end
    if (s1_fire) begin // @[Reg.scala 17:18]
      if (s1_meta_errors_REG) begin // @[Reg.scala 17:18]
        s2_meta_errors_0_4 <= io_metaArray_fromIMeta_errors_0_4; // @[Reg.scala 17:22]
      end else begin
        s2_meta_errors_0_4 <= s1_meta_errors_r0_4; // @[Reg.scala 16:16]
      end
    end
    if (s1_fire) begin // @[Reg.scala 17:18]
      if (s1_meta_errors_REG) begin // @[Reg.scala 17:18]
        s2_meta_errors_0_5 <= io_metaArray_fromIMeta_errors_0_5; // @[Reg.scala 17:22]
      end else begin
        s2_meta_errors_0_5 <= s1_meta_errors_r0_5; // @[Reg.scala 16:16]
      end
    end
    if (s1_fire) begin // @[Reg.scala 17:18]
      if (s1_meta_errors_REG) begin // @[Reg.scala 17:18]
        s2_meta_errors_0_6 <= io_metaArray_fromIMeta_errors_0_6; // @[Reg.scala 17:22]
      end else begin
        s2_meta_errors_0_6 <= s1_meta_errors_r0_6; // @[Reg.scala 16:16]
      end
    end
    if (s1_fire) begin // @[Reg.scala 17:18]
      if (s1_meta_errors_REG) begin // @[Reg.scala 17:18]
        s2_meta_errors_0_7 <= io_metaArray_fromIMeta_errors_0_7; // @[Reg.scala 17:22]
      end else begin
        s2_meta_errors_0_7 <= s1_meta_errors_r0_7; // @[Reg.scala 16:16]
      end
    end
    if (s1_fire) begin // @[Reg.scala 17:18]
      if (s1_meta_errors_REG) begin // @[Reg.scala 17:18]
        s2_meta_errors_1_0 <= io_metaArray_fromIMeta_errors_1_0; // @[Reg.scala 17:22]
      end else begin
        s2_meta_errors_1_0 <= s1_meta_errors_r1_0; // @[Reg.scala 16:16]
      end
    end
    if (s1_fire) begin // @[Reg.scala 17:18]
      if (s1_meta_errors_REG) begin // @[Reg.scala 17:18]
        s2_meta_errors_1_1 <= io_metaArray_fromIMeta_errors_1_1; // @[Reg.scala 17:22]
      end else begin
        s2_meta_errors_1_1 <= s1_meta_errors_r1_1; // @[Reg.scala 16:16]
      end
    end
    if (s1_fire) begin // @[Reg.scala 17:18]
      if (s1_meta_errors_REG) begin // @[Reg.scala 17:18]
        s2_meta_errors_1_2 <= io_metaArray_fromIMeta_errors_1_2; // @[Reg.scala 17:22]
      end else begin
        s2_meta_errors_1_2 <= s1_meta_errors_r1_2; // @[Reg.scala 16:16]
      end
    end
    if (s1_fire) begin // @[Reg.scala 17:18]
      if (s1_meta_errors_REG) begin // @[Reg.scala 17:18]
        s2_meta_errors_1_3 <= io_metaArray_fromIMeta_errors_1_3; // @[Reg.scala 17:22]
      end else begin
        s2_meta_errors_1_3 <= s1_meta_errors_r1_3; // @[Reg.scala 16:16]
      end
    end
    if (s1_fire) begin // @[Reg.scala 17:18]
      if (s1_meta_errors_REG) begin // @[Reg.scala 17:18]
        s2_meta_errors_1_4 <= io_metaArray_fromIMeta_errors_1_4; // @[Reg.scala 17:22]
      end else begin
        s2_meta_errors_1_4 <= s1_meta_errors_r1_4; // @[Reg.scala 16:16]
      end
    end
    if (s1_fire) begin // @[Reg.scala 17:18]
      if (s1_meta_errors_REG) begin // @[Reg.scala 17:18]
        s2_meta_errors_1_5 <= io_metaArray_fromIMeta_errors_1_5; // @[Reg.scala 17:22]
      end else begin
        s2_meta_errors_1_5 <= s1_meta_errors_r1_5; // @[Reg.scala 16:16]
      end
    end
    if (s1_fire) begin // @[Reg.scala 17:18]
      if (s1_meta_errors_REG) begin // @[Reg.scala 17:18]
        s2_meta_errors_1_6 <= io_metaArray_fromIMeta_errors_1_6; // @[Reg.scala 17:22]
      end else begin
        s2_meta_errors_1_6 <= s1_meta_errors_r1_6; // @[Reg.scala 16:16]
      end
    end
    if (s1_fire) begin // @[Reg.scala 17:18]
      if (s1_meta_errors_REG) begin // @[Reg.scala 17:18]
        s2_meta_errors_1_7 <= io_metaArray_fromIMeta_errors_1_7; // @[Reg.scala 17:22]
      end else begin
        s2_meta_errors_1_7 <= s1_meta_errors_r1_7; // @[Reg.scala 16:16]
      end
    end
    if (s1_fire) begin // @[Reg.scala 17:18]
      if (s1_data_errorBits_REG) begin // @[Reg.scala 17:18]
        s2_data_errorBits_0_0 <= io_dataArray_fromIData_codes_0_0; // @[Reg.scala 17:22]
      end else begin
        s2_data_errorBits_0_0 <= s1_data_errorBits_r0_0; // @[Reg.scala 16:16]
      end
    end
    if (s1_fire) begin // @[Reg.scala 17:18]
      if (s1_data_errorBits_REG) begin // @[Reg.scala 17:18]
        s2_data_errorBits_0_1 <= io_dataArray_fromIData_codes_0_1; // @[Reg.scala 17:22]
      end else begin
        s2_data_errorBits_0_1 <= s1_data_errorBits_r0_1; // @[Reg.scala 16:16]
      end
    end
    if (s1_fire) begin // @[Reg.scala 17:18]
      if (s1_data_errorBits_REG) begin // @[Reg.scala 17:18]
        s2_data_errorBits_0_2 <= io_dataArray_fromIData_codes_0_2; // @[Reg.scala 17:22]
      end else begin
        s2_data_errorBits_0_2 <= s1_data_errorBits_r0_2; // @[Reg.scala 16:16]
      end
    end
    if (s1_fire) begin // @[Reg.scala 17:18]
      if (s1_data_errorBits_REG) begin // @[Reg.scala 17:18]
        s2_data_errorBits_0_3 <= io_dataArray_fromIData_codes_0_3; // @[Reg.scala 17:22]
      end else begin
        s2_data_errorBits_0_3 <= s1_data_errorBits_r0_3; // @[Reg.scala 16:16]
      end
    end
    if (s1_fire) begin // @[Reg.scala 17:18]
      if (s1_data_errorBits_REG) begin // @[Reg.scala 17:18]
        s2_data_errorBits_0_4 <= io_dataArray_fromIData_codes_0_4; // @[Reg.scala 17:22]
      end else begin
        s2_data_errorBits_0_4 <= s1_data_errorBits_r0_4; // @[Reg.scala 16:16]
      end
    end
    if (s1_fire) begin // @[Reg.scala 17:18]
      if (s1_data_errorBits_REG) begin // @[Reg.scala 17:18]
        s2_data_errorBits_0_5 <= io_dataArray_fromIData_codes_0_5; // @[Reg.scala 17:22]
      end else begin
        s2_data_errorBits_0_5 <= s1_data_errorBits_r0_5; // @[Reg.scala 16:16]
      end
    end
    if (s1_fire) begin // @[Reg.scala 17:18]
      if (s1_data_errorBits_REG) begin // @[Reg.scala 17:18]
        s2_data_errorBits_0_6 <= io_dataArray_fromIData_codes_0_6; // @[Reg.scala 17:22]
      end else begin
        s2_data_errorBits_0_6 <= s1_data_errorBits_r0_6; // @[Reg.scala 16:16]
      end
    end
    if (s1_fire) begin // @[Reg.scala 17:18]
      if (s1_data_errorBits_REG) begin // @[Reg.scala 17:18]
        s2_data_errorBits_0_7 <= io_dataArray_fromIData_codes_0_7; // @[Reg.scala 17:22]
      end else begin
        s2_data_errorBits_0_7 <= s1_data_errorBits_r0_7; // @[Reg.scala 16:16]
      end
    end
    if (s1_fire) begin // @[Reg.scala 17:18]
      if (s1_data_errorBits_REG) begin // @[Reg.scala 17:18]
        s2_data_errorBits_1_0 <= io_dataArray_fromIData_codes_1_0; // @[Reg.scala 17:22]
      end else begin
        s2_data_errorBits_1_0 <= s1_data_errorBits_r1_0; // @[Reg.scala 16:16]
      end
    end
    if (s1_fire) begin // @[Reg.scala 17:18]
      if (s1_data_errorBits_REG) begin // @[Reg.scala 17:18]
        s2_data_errorBits_1_1 <= io_dataArray_fromIData_codes_1_1; // @[Reg.scala 17:22]
      end else begin
        s2_data_errorBits_1_1 <= s1_data_errorBits_r1_1; // @[Reg.scala 16:16]
      end
    end
    if (s1_fire) begin // @[Reg.scala 17:18]
      if (s1_data_errorBits_REG) begin // @[Reg.scala 17:18]
        s2_data_errorBits_1_2 <= io_dataArray_fromIData_codes_1_2; // @[Reg.scala 17:22]
      end else begin
        s2_data_errorBits_1_2 <= s1_data_errorBits_r1_2; // @[Reg.scala 16:16]
      end
    end
    if (s1_fire) begin // @[Reg.scala 17:18]
      if (s1_data_errorBits_REG) begin // @[Reg.scala 17:18]
        s2_data_errorBits_1_3 <= io_dataArray_fromIData_codes_1_3; // @[Reg.scala 17:22]
      end else begin
        s2_data_errorBits_1_3 <= s1_data_errorBits_r1_3; // @[Reg.scala 16:16]
      end
    end
    if (s1_fire) begin // @[Reg.scala 17:18]
      if (s1_data_errorBits_REG) begin // @[Reg.scala 17:18]
        s2_data_errorBits_1_4 <= io_dataArray_fromIData_codes_1_4; // @[Reg.scala 17:22]
      end else begin
        s2_data_errorBits_1_4 <= s1_data_errorBits_r1_4; // @[Reg.scala 16:16]
      end
    end
    if (s1_fire) begin // @[Reg.scala 17:18]
      if (s1_data_errorBits_REG) begin // @[Reg.scala 17:18]
        s2_data_errorBits_1_5 <= io_dataArray_fromIData_codes_1_5; // @[Reg.scala 17:22]
      end else begin
        s2_data_errorBits_1_5 <= s1_data_errorBits_r1_5; // @[Reg.scala 16:16]
      end
    end
    if (s1_fire) begin // @[Reg.scala 17:18]
      if (s1_data_errorBits_REG) begin // @[Reg.scala 17:18]
        s2_data_errorBits_1_6 <= io_dataArray_fromIData_codes_1_6; // @[Reg.scala 17:22]
      end else begin
        s2_data_errorBits_1_6 <= s1_data_errorBits_r1_6; // @[Reg.scala 16:16]
      end
    end
    if (s1_fire) begin // @[Reg.scala 17:18]
      if (s1_data_errorBits_REG) begin // @[Reg.scala 17:18]
        s2_data_errorBits_1_7 <= io_dataArray_fromIData_codes_1_7; // @[Reg.scala 17:22]
      end else begin
        s2_data_errorBits_1_7 <= s1_data_errorBits_r1_7; // @[Reg.scala 16:16]
      end
    end
    if (s1_fire) begin // @[Reg.scala 17:18]
      if (s1_data_cacheline_REG) begin // @[Reg.scala 17:18]
        s2_data_cacheline_0_0 <= io_dataArray_fromIData_datas_0_0; // @[Reg.scala 17:22]
      end else begin
        s2_data_cacheline_0_0 <= s1_data_cacheline_r0_0; // @[Reg.scala 16:16]
      end
    end
    if (s1_fire) begin // @[Reg.scala 17:18]
      if (s1_data_cacheline_REG) begin // @[Reg.scala 17:18]
        s2_data_cacheline_0_1 <= io_dataArray_fromIData_datas_0_1; // @[Reg.scala 17:22]
      end else begin
        s2_data_cacheline_0_1 <= s1_data_cacheline_r0_1; // @[Reg.scala 16:16]
      end
    end
    if (s1_fire) begin // @[Reg.scala 17:18]
      if (s1_data_cacheline_REG) begin // @[Reg.scala 17:18]
        s2_data_cacheline_0_2 <= io_dataArray_fromIData_datas_0_2; // @[Reg.scala 17:22]
      end else begin
        s2_data_cacheline_0_2 <= s1_data_cacheline_r0_2; // @[Reg.scala 16:16]
      end
    end
    if (s1_fire) begin // @[Reg.scala 17:18]
      if (s1_data_cacheline_REG) begin // @[Reg.scala 17:18]
        s2_data_cacheline_0_3 <= io_dataArray_fromIData_datas_0_3; // @[Reg.scala 17:22]
      end else begin
        s2_data_cacheline_0_3 <= s1_data_cacheline_r0_3; // @[Reg.scala 16:16]
      end
    end
    if (s1_fire) begin // @[Reg.scala 17:18]
      if (s1_data_cacheline_REG) begin // @[Reg.scala 17:18]
        s2_data_cacheline_0_4 <= io_dataArray_fromIData_datas_0_4; // @[Reg.scala 17:22]
      end else begin
        s2_data_cacheline_0_4 <= s1_data_cacheline_r0_4; // @[Reg.scala 16:16]
      end
    end
    if (s1_fire) begin // @[Reg.scala 17:18]
      if (s1_data_cacheline_REG) begin // @[Reg.scala 17:18]
        s2_data_cacheline_0_5 <= io_dataArray_fromIData_datas_0_5; // @[Reg.scala 17:22]
      end else begin
        s2_data_cacheline_0_5 <= s1_data_cacheline_r0_5; // @[Reg.scala 16:16]
      end
    end
    if (s1_fire) begin // @[Reg.scala 17:18]
      if (s1_data_cacheline_REG) begin // @[Reg.scala 17:18]
        s2_data_cacheline_0_6 <= io_dataArray_fromIData_datas_0_6; // @[Reg.scala 17:22]
      end else begin
        s2_data_cacheline_0_6 <= s1_data_cacheline_r0_6; // @[Reg.scala 16:16]
      end
    end
    if (s1_fire) begin // @[Reg.scala 17:18]
      if (s1_data_cacheline_REG) begin // @[Reg.scala 17:18]
        s2_data_cacheline_0_7 <= io_dataArray_fromIData_datas_0_7; // @[Reg.scala 17:22]
      end else begin
        s2_data_cacheline_0_7 <= s1_data_cacheline_r0_7; // @[Reg.scala 16:16]
      end
    end
    if (s1_fire) begin // @[Reg.scala 17:18]
      if (s1_data_cacheline_REG) begin // @[Reg.scala 17:18]
        s2_data_cacheline_1_0 <= io_dataArray_fromIData_datas_1_0; // @[Reg.scala 17:22]
      end else begin
        s2_data_cacheline_1_0 <= s1_data_cacheline_r1_0; // @[Reg.scala 16:16]
      end
    end
    if (s1_fire) begin // @[Reg.scala 17:18]
      if (s1_data_cacheline_REG) begin // @[Reg.scala 17:18]
        s2_data_cacheline_1_1 <= io_dataArray_fromIData_datas_1_1; // @[Reg.scala 17:22]
      end else begin
        s2_data_cacheline_1_1 <= s1_data_cacheline_r1_1; // @[Reg.scala 16:16]
      end
    end
    if (s1_fire) begin // @[Reg.scala 17:18]
      if (s1_data_cacheline_REG) begin // @[Reg.scala 17:18]
        s2_data_cacheline_1_2 <= io_dataArray_fromIData_datas_1_2; // @[Reg.scala 17:22]
      end else begin
        s2_data_cacheline_1_2 <= s1_data_cacheline_r1_2; // @[Reg.scala 16:16]
      end
    end
    if (s1_fire) begin // @[Reg.scala 17:18]
      if (s1_data_cacheline_REG) begin // @[Reg.scala 17:18]
        s2_data_cacheline_1_3 <= io_dataArray_fromIData_datas_1_3; // @[Reg.scala 17:22]
      end else begin
        s2_data_cacheline_1_3 <= s1_data_cacheline_r1_3; // @[Reg.scala 16:16]
      end
    end
    if (s1_fire) begin // @[Reg.scala 17:18]
      if (s1_data_cacheline_REG) begin // @[Reg.scala 17:18]
        s2_data_cacheline_1_4 <= io_dataArray_fromIData_datas_1_4; // @[Reg.scala 17:22]
      end else begin
        s2_data_cacheline_1_4 <= s1_data_cacheline_r1_4; // @[Reg.scala 16:16]
      end
    end
    if (s1_fire) begin // @[Reg.scala 17:18]
      if (s1_data_cacheline_REG) begin // @[Reg.scala 17:18]
        s2_data_cacheline_1_5 <= io_dataArray_fromIData_datas_1_5; // @[Reg.scala 17:22]
      end else begin
        s2_data_cacheline_1_5 <= s1_data_cacheline_r1_5; // @[Reg.scala 16:16]
      end
    end
    if (s1_fire) begin // @[Reg.scala 17:18]
      if (s1_data_cacheline_REG) begin // @[Reg.scala 17:18]
        s2_data_cacheline_1_6 <= io_dataArray_fromIData_datas_1_6; // @[Reg.scala 17:22]
      end else begin
        s2_data_cacheline_1_6 <= s1_data_cacheline_r1_6; // @[Reg.scala 16:16]
      end
    end
    if (s1_fire) begin // @[Reg.scala 17:18]
      if (s1_data_cacheline_REG) begin // @[Reg.scala 17:18]
        s2_data_cacheline_1_7 <= io_dataArray_fromIData_datas_1_7; // @[Reg.scala 17:22]
      end else begin
        s2_data_cacheline_1_7 <= s1_data_cacheline_r1_7; // @[Reg.scala 16:16]
      end
    end
    s2_data_errors_0_0_REG <= s1_valid & tlbRespAllValid & s2_ready; // @[ICacheMainPipe.scala 270:43]
    s2_data_errors_0_0_REG_1 <= s2_data_errors_0_0_REG; // @[ICacheMainPipe.scala 379:40]
    s2_data_errors_0_0_REG_2_0 <= ^data_full_wayBits__0_0; // @[ECC.scala 87:27]
    s2_data_errors_0_0_REG_2_1 <= ^data_full_wayBits__0_1; // @[ECC.scala 87:27]
    s2_data_errors_0_0_REG_2_2 <= ^data_full_wayBits__0_2; // @[ECC.scala 87:27]
    s2_data_errors_0_0_REG_2_3 <= ^data_full_wayBits__0_3; // @[ECC.scala 87:27]
    s2_data_errors_0_0_REG_2_4 <= ^data_full_wayBits__0_4; // @[ECC.scala 87:27]
    s2_data_errors_0_0_REG_2_5 <= ^data_full_wayBits__0_5; // @[ECC.scala 87:27]
    s2_data_errors_0_0_REG_2_6 <= ^data_full_wayBits__0_6; // @[ECC.scala 87:27]
    s2_data_errors_0_0_REG_2_7 <= ^data_full_wayBits__0_7; // @[ECC.scala 87:27]
    s2_data_errors_0_0_REG_2_8 <= ^data_full_wayBits__0_8; // @[ECC.scala 87:27]
    s2_data_errors_0_0_REG_2_9 <= ^data_full_wayBits__0_9; // @[ECC.scala 87:27]
    s2_data_errors_0_0_REG_2_10 <= ^data_full_wayBits__0_10; // @[ECC.scala 87:27]
    s2_data_errors_0_0_REG_2_11 <= ^data_full_wayBits__0_11; // @[ECC.scala 87:27]
    s2_data_errors_0_0_REG_2_12 <= ^data_full_wayBits__0_12; // @[ECC.scala 87:27]
    s2_data_errors_0_0_REG_2_13 <= ^data_full_wayBits__0_13; // @[ECC.scala 87:27]
    s2_data_errors_0_0_REG_2_14 <= ^data_full_wayBits__0_14; // @[ECC.scala 87:27]
    s2_data_errors_0_0_REG_2_15 <= ^data_full_wayBits__0_15; // @[ECC.scala 87:27]
    s2_data_errors_0_0_REG_2_16 <= ^data_full_wayBits__0_16; // @[ECC.scala 87:27]
    s2_data_errors_0_0_REG_2_17 <= ^data_full_wayBits__0_17; // @[ECC.scala 87:27]
    s2_data_errors_0_0_REG_2_18 <= ^data_full_wayBits__0_18; // @[ECC.scala 87:27]
    s2_data_errors_0_0_REG_2_19 <= ^data_full_wayBits__0_19; // @[ECC.scala 87:27]
    s2_data_errors_0_0_REG_2_20 <= ^data_full_wayBits__0_20; // @[ECC.scala 87:27]
    s2_data_errors_0_0_REG_2_21 <= ^data_full_wayBits__0_21; // @[ECC.scala 87:27]
    s2_data_errors_0_0_REG_2_22 <= ^data_full_wayBits__0_22; // @[ECC.scala 87:27]
    s2_data_errors_0_0_REG_2_23 <= ^data_full_wayBits__0_23; // @[ECC.scala 87:27]
    s2_data_errors_0_0_REG_2_24 <= ^data_full_wayBits__0_24; // @[ECC.scala 87:27]
    s2_data_errors_0_0_REG_2_25 <= ^data_full_wayBits__0_25; // @[ECC.scala 87:27]
    s2_data_errors_0_0_REG_2_26 <= ^data_full_wayBits__0_26; // @[ECC.scala 87:27]
    s2_data_errors_0_0_REG_2_27 <= ^data_full_wayBits__0_27; // @[ECC.scala 87:27]
    s2_data_errors_0_0_REG_2_28 <= ^data_full_wayBits__0_28; // @[ECC.scala 87:27]
    s2_data_errors_0_0_REG_2_29 <= ^data_full_wayBits__0_29; // @[ECC.scala 87:27]
    s2_data_errors_0_0_REG_2_30 <= ^data_full_wayBits__0_30; // @[ECC.scala 87:27]
    s2_data_errors_0_0_REG_2_31 <= ^data_full_wayBits__0_31; // @[ECC.scala 87:27]
    s2_data_errors_0_1_REG <= s1_valid & tlbRespAllValid & s2_ready; // @[ICacheMainPipe.scala 270:43]
    s2_data_errors_0_1_REG_1 <= s2_data_errors_0_1_REG; // @[ICacheMainPipe.scala 379:40]
    s2_data_errors_0_1_REG_2_0 <= ^data_full_wayBits__1_0; // @[ECC.scala 87:27]
    s2_data_errors_0_1_REG_2_1 <= ^data_full_wayBits__1_1; // @[ECC.scala 87:27]
    s2_data_errors_0_1_REG_2_2 <= ^data_full_wayBits__1_2; // @[ECC.scala 87:27]
    s2_data_errors_0_1_REG_2_3 <= ^data_full_wayBits__1_3; // @[ECC.scala 87:27]
    s2_data_errors_0_1_REG_2_4 <= ^data_full_wayBits__1_4; // @[ECC.scala 87:27]
    s2_data_errors_0_1_REG_2_5 <= ^data_full_wayBits__1_5; // @[ECC.scala 87:27]
    s2_data_errors_0_1_REG_2_6 <= ^data_full_wayBits__1_6; // @[ECC.scala 87:27]
    s2_data_errors_0_1_REG_2_7 <= ^data_full_wayBits__1_7; // @[ECC.scala 87:27]
    s2_data_errors_0_1_REG_2_8 <= ^data_full_wayBits__1_8; // @[ECC.scala 87:27]
    s2_data_errors_0_1_REG_2_9 <= ^data_full_wayBits__1_9; // @[ECC.scala 87:27]
    s2_data_errors_0_1_REG_2_10 <= ^data_full_wayBits__1_10; // @[ECC.scala 87:27]
    s2_data_errors_0_1_REG_2_11 <= ^data_full_wayBits__1_11; // @[ECC.scala 87:27]
    s2_data_errors_0_1_REG_2_12 <= ^data_full_wayBits__1_12; // @[ECC.scala 87:27]
    s2_data_errors_0_1_REG_2_13 <= ^data_full_wayBits__1_13; // @[ECC.scala 87:27]
    s2_data_errors_0_1_REG_2_14 <= ^data_full_wayBits__1_14; // @[ECC.scala 87:27]
    s2_data_errors_0_1_REG_2_15 <= ^data_full_wayBits__1_15; // @[ECC.scala 87:27]
    s2_data_errors_0_1_REG_2_16 <= ^data_full_wayBits__1_16; // @[ECC.scala 87:27]
    s2_data_errors_0_1_REG_2_17 <= ^data_full_wayBits__1_17; // @[ECC.scala 87:27]
    s2_data_errors_0_1_REG_2_18 <= ^data_full_wayBits__1_18; // @[ECC.scala 87:27]
    s2_data_errors_0_1_REG_2_19 <= ^data_full_wayBits__1_19; // @[ECC.scala 87:27]
    s2_data_errors_0_1_REG_2_20 <= ^data_full_wayBits__1_20; // @[ECC.scala 87:27]
    s2_data_errors_0_1_REG_2_21 <= ^data_full_wayBits__1_21; // @[ECC.scala 87:27]
    s2_data_errors_0_1_REG_2_22 <= ^data_full_wayBits__1_22; // @[ECC.scala 87:27]
    s2_data_errors_0_1_REG_2_23 <= ^data_full_wayBits__1_23; // @[ECC.scala 87:27]
    s2_data_errors_0_1_REG_2_24 <= ^data_full_wayBits__1_24; // @[ECC.scala 87:27]
    s2_data_errors_0_1_REG_2_25 <= ^data_full_wayBits__1_25; // @[ECC.scala 87:27]
    s2_data_errors_0_1_REG_2_26 <= ^data_full_wayBits__1_26; // @[ECC.scala 87:27]
    s2_data_errors_0_1_REG_2_27 <= ^data_full_wayBits__1_27; // @[ECC.scala 87:27]
    s2_data_errors_0_1_REG_2_28 <= ^data_full_wayBits__1_28; // @[ECC.scala 87:27]
    s2_data_errors_0_1_REG_2_29 <= ^data_full_wayBits__1_29; // @[ECC.scala 87:27]
    s2_data_errors_0_1_REG_2_30 <= ^data_full_wayBits__1_30; // @[ECC.scala 87:27]
    s2_data_errors_0_1_REG_2_31 <= ^data_full_wayBits__1_31; // @[ECC.scala 87:27]
    s2_data_errors_0_2_REG <= s1_valid & tlbRespAllValid & s2_ready; // @[ICacheMainPipe.scala 270:43]
    s2_data_errors_0_2_REG_1 <= s2_data_errors_0_2_REG; // @[ICacheMainPipe.scala 379:40]
    s2_data_errors_0_2_REG_2_0 <= ^data_full_wayBits__2_0; // @[ECC.scala 87:27]
    s2_data_errors_0_2_REG_2_1 <= ^data_full_wayBits__2_1; // @[ECC.scala 87:27]
    s2_data_errors_0_2_REG_2_2 <= ^data_full_wayBits__2_2; // @[ECC.scala 87:27]
    s2_data_errors_0_2_REG_2_3 <= ^data_full_wayBits__2_3; // @[ECC.scala 87:27]
    s2_data_errors_0_2_REG_2_4 <= ^data_full_wayBits__2_4; // @[ECC.scala 87:27]
    s2_data_errors_0_2_REG_2_5 <= ^data_full_wayBits__2_5; // @[ECC.scala 87:27]
    s2_data_errors_0_2_REG_2_6 <= ^data_full_wayBits__2_6; // @[ECC.scala 87:27]
    s2_data_errors_0_2_REG_2_7 <= ^data_full_wayBits__2_7; // @[ECC.scala 87:27]
    s2_data_errors_0_2_REG_2_8 <= ^data_full_wayBits__2_8; // @[ECC.scala 87:27]
    s2_data_errors_0_2_REG_2_9 <= ^data_full_wayBits__2_9; // @[ECC.scala 87:27]
    s2_data_errors_0_2_REG_2_10 <= ^data_full_wayBits__2_10; // @[ECC.scala 87:27]
    s2_data_errors_0_2_REG_2_11 <= ^data_full_wayBits__2_11; // @[ECC.scala 87:27]
    s2_data_errors_0_2_REG_2_12 <= ^data_full_wayBits__2_12; // @[ECC.scala 87:27]
    s2_data_errors_0_2_REG_2_13 <= ^data_full_wayBits__2_13; // @[ECC.scala 87:27]
    s2_data_errors_0_2_REG_2_14 <= ^data_full_wayBits__2_14; // @[ECC.scala 87:27]
    s2_data_errors_0_2_REG_2_15 <= ^data_full_wayBits__2_15; // @[ECC.scala 87:27]
    s2_data_errors_0_2_REG_2_16 <= ^data_full_wayBits__2_16; // @[ECC.scala 87:27]
    s2_data_errors_0_2_REG_2_17 <= ^data_full_wayBits__2_17; // @[ECC.scala 87:27]
    s2_data_errors_0_2_REG_2_18 <= ^data_full_wayBits__2_18; // @[ECC.scala 87:27]
    s2_data_errors_0_2_REG_2_19 <= ^data_full_wayBits__2_19; // @[ECC.scala 87:27]
    s2_data_errors_0_2_REG_2_20 <= ^data_full_wayBits__2_20; // @[ECC.scala 87:27]
    s2_data_errors_0_2_REG_2_21 <= ^data_full_wayBits__2_21; // @[ECC.scala 87:27]
    s2_data_errors_0_2_REG_2_22 <= ^data_full_wayBits__2_22; // @[ECC.scala 87:27]
    s2_data_errors_0_2_REG_2_23 <= ^data_full_wayBits__2_23; // @[ECC.scala 87:27]
    s2_data_errors_0_2_REG_2_24 <= ^data_full_wayBits__2_24; // @[ECC.scala 87:27]
    s2_data_errors_0_2_REG_2_25 <= ^data_full_wayBits__2_25; // @[ECC.scala 87:27]
    s2_data_errors_0_2_REG_2_26 <= ^data_full_wayBits__2_26; // @[ECC.scala 87:27]
    s2_data_errors_0_2_REG_2_27 <= ^data_full_wayBits__2_27; // @[ECC.scala 87:27]
    s2_data_errors_0_2_REG_2_28 <= ^data_full_wayBits__2_28; // @[ECC.scala 87:27]
    s2_data_errors_0_2_REG_2_29 <= ^data_full_wayBits__2_29; // @[ECC.scala 87:27]
    s2_data_errors_0_2_REG_2_30 <= ^data_full_wayBits__2_30; // @[ECC.scala 87:27]
    s2_data_errors_0_2_REG_2_31 <= ^data_full_wayBits__2_31; // @[ECC.scala 87:27]
    s2_data_errors_0_3_REG <= s1_valid & tlbRespAllValid & s2_ready; // @[ICacheMainPipe.scala 270:43]
    s2_data_errors_0_3_REG_1 <= s2_data_errors_0_3_REG; // @[ICacheMainPipe.scala 379:40]
    s2_data_errors_0_3_REG_2_0 <= ^data_full_wayBits__3_0; // @[ECC.scala 87:27]
    s2_data_errors_0_3_REG_2_1 <= ^data_full_wayBits__3_1; // @[ECC.scala 87:27]
    s2_data_errors_0_3_REG_2_2 <= ^data_full_wayBits__3_2; // @[ECC.scala 87:27]
    s2_data_errors_0_3_REG_2_3 <= ^data_full_wayBits__3_3; // @[ECC.scala 87:27]
    s2_data_errors_0_3_REG_2_4 <= ^data_full_wayBits__3_4; // @[ECC.scala 87:27]
    s2_data_errors_0_3_REG_2_5 <= ^data_full_wayBits__3_5; // @[ECC.scala 87:27]
    s2_data_errors_0_3_REG_2_6 <= ^data_full_wayBits__3_6; // @[ECC.scala 87:27]
    s2_data_errors_0_3_REG_2_7 <= ^data_full_wayBits__3_7; // @[ECC.scala 87:27]
    s2_data_errors_0_3_REG_2_8 <= ^data_full_wayBits__3_8; // @[ECC.scala 87:27]
    s2_data_errors_0_3_REG_2_9 <= ^data_full_wayBits__3_9; // @[ECC.scala 87:27]
    s2_data_errors_0_3_REG_2_10 <= ^data_full_wayBits__3_10; // @[ECC.scala 87:27]
    s2_data_errors_0_3_REG_2_11 <= ^data_full_wayBits__3_11; // @[ECC.scala 87:27]
    s2_data_errors_0_3_REG_2_12 <= ^data_full_wayBits__3_12; // @[ECC.scala 87:27]
    s2_data_errors_0_3_REG_2_13 <= ^data_full_wayBits__3_13; // @[ECC.scala 87:27]
    s2_data_errors_0_3_REG_2_14 <= ^data_full_wayBits__3_14; // @[ECC.scala 87:27]
    s2_data_errors_0_3_REG_2_15 <= ^data_full_wayBits__3_15; // @[ECC.scala 87:27]
    s2_data_errors_0_3_REG_2_16 <= ^data_full_wayBits__3_16; // @[ECC.scala 87:27]
    s2_data_errors_0_3_REG_2_17 <= ^data_full_wayBits__3_17; // @[ECC.scala 87:27]
    s2_data_errors_0_3_REG_2_18 <= ^data_full_wayBits__3_18; // @[ECC.scala 87:27]
    s2_data_errors_0_3_REG_2_19 <= ^data_full_wayBits__3_19; // @[ECC.scala 87:27]
    s2_data_errors_0_3_REG_2_20 <= ^data_full_wayBits__3_20; // @[ECC.scala 87:27]
    s2_data_errors_0_3_REG_2_21 <= ^data_full_wayBits__3_21; // @[ECC.scala 87:27]
    s2_data_errors_0_3_REG_2_22 <= ^data_full_wayBits__3_22; // @[ECC.scala 87:27]
    s2_data_errors_0_3_REG_2_23 <= ^data_full_wayBits__3_23; // @[ECC.scala 87:27]
    s2_data_errors_0_3_REG_2_24 <= ^data_full_wayBits__3_24; // @[ECC.scala 87:27]
    s2_data_errors_0_3_REG_2_25 <= ^data_full_wayBits__3_25; // @[ECC.scala 87:27]
    s2_data_errors_0_3_REG_2_26 <= ^data_full_wayBits__3_26; // @[ECC.scala 87:27]
    s2_data_errors_0_3_REG_2_27 <= ^data_full_wayBits__3_27; // @[ECC.scala 87:27]
    s2_data_errors_0_3_REG_2_28 <= ^data_full_wayBits__3_28; // @[ECC.scala 87:27]
    s2_data_errors_0_3_REG_2_29 <= ^data_full_wayBits__3_29; // @[ECC.scala 87:27]
    s2_data_errors_0_3_REG_2_30 <= ^data_full_wayBits__3_30; // @[ECC.scala 87:27]
    s2_data_errors_0_3_REG_2_31 <= ^data_full_wayBits__3_31; // @[ECC.scala 87:27]
    s2_data_errors_0_4_REG <= s1_valid & tlbRespAllValid & s2_ready; // @[ICacheMainPipe.scala 270:43]
    s2_data_errors_0_4_REG_1 <= s2_data_errors_0_4_REG; // @[ICacheMainPipe.scala 379:40]
    s2_data_errors_0_4_REG_2_0 <= ^data_full_wayBits__4_0; // @[ECC.scala 87:27]
    s2_data_errors_0_4_REG_2_1 <= ^data_full_wayBits__4_1; // @[ECC.scala 87:27]
    s2_data_errors_0_4_REG_2_2 <= ^data_full_wayBits__4_2; // @[ECC.scala 87:27]
    s2_data_errors_0_4_REG_2_3 <= ^data_full_wayBits__4_3; // @[ECC.scala 87:27]
    s2_data_errors_0_4_REG_2_4 <= ^data_full_wayBits__4_4; // @[ECC.scala 87:27]
    s2_data_errors_0_4_REG_2_5 <= ^data_full_wayBits__4_5; // @[ECC.scala 87:27]
    s2_data_errors_0_4_REG_2_6 <= ^data_full_wayBits__4_6; // @[ECC.scala 87:27]
    s2_data_errors_0_4_REG_2_7 <= ^data_full_wayBits__4_7; // @[ECC.scala 87:27]
    s2_data_errors_0_4_REG_2_8 <= ^data_full_wayBits__4_8; // @[ECC.scala 87:27]
    s2_data_errors_0_4_REG_2_9 <= ^data_full_wayBits__4_9; // @[ECC.scala 87:27]
    s2_data_errors_0_4_REG_2_10 <= ^data_full_wayBits__4_10; // @[ECC.scala 87:27]
    s2_data_errors_0_4_REG_2_11 <= ^data_full_wayBits__4_11; // @[ECC.scala 87:27]
    s2_data_errors_0_4_REG_2_12 <= ^data_full_wayBits__4_12; // @[ECC.scala 87:27]
    s2_data_errors_0_4_REG_2_13 <= ^data_full_wayBits__4_13; // @[ECC.scala 87:27]
    s2_data_errors_0_4_REG_2_14 <= ^data_full_wayBits__4_14; // @[ECC.scala 87:27]
    s2_data_errors_0_4_REG_2_15 <= ^data_full_wayBits__4_15; // @[ECC.scala 87:27]
    s2_data_errors_0_4_REG_2_16 <= ^data_full_wayBits__4_16; // @[ECC.scala 87:27]
    s2_data_errors_0_4_REG_2_17 <= ^data_full_wayBits__4_17; // @[ECC.scala 87:27]
    s2_data_errors_0_4_REG_2_18 <= ^data_full_wayBits__4_18; // @[ECC.scala 87:27]
    s2_data_errors_0_4_REG_2_19 <= ^data_full_wayBits__4_19; // @[ECC.scala 87:27]
    s2_data_errors_0_4_REG_2_20 <= ^data_full_wayBits__4_20; // @[ECC.scala 87:27]
    s2_data_errors_0_4_REG_2_21 <= ^data_full_wayBits__4_21; // @[ECC.scala 87:27]
    s2_data_errors_0_4_REG_2_22 <= ^data_full_wayBits__4_22; // @[ECC.scala 87:27]
    s2_data_errors_0_4_REG_2_23 <= ^data_full_wayBits__4_23; // @[ECC.scala 87:27]
    s2_data_errors_0_4_REG_2_24 <= ^data_full_wayBits__4_24; // @[ECC.scala 87:27]
    s2_data_errors_0_4_REG_2_25 <= ^data_full_wayBits__4_25; // @[ECC.scala 87:27]
    s2_data_errors_0_4_REG_2_26 <= ^data_full_wayBits__4_26; // @[ECC.scala 87:27]
    s2_data_errors_0_4_REG_2_27 <= ^data_full_wayBits__4_27; // @[ECC.scala 87:27]
    s2_data_errors_0_4_REG_2_28 <= ^data_full_wayBits__4_28; // @[ECC.scala 87:27]
    s2_data_errors_0_4_REG_2_29 <= ^data_full_wayBits__4_29; // @[ECC.scala 87:27]
    s2_data_errors_0_4_REG_2_30 <= ^data_full_wayBits__4_30; // @[ECC.scala 87:27]
    s2_data_errors_0_4_REG_2_31 <= ^data_full_wayBits__4_31; // @[ECC.scala 87:27]
    s2_data_errors_0_5_REG <= s1_valid & tlbRespAllValid & s2_ready; // @[ICacheMainPipe.scala 270:43]
    s2_data_errors_0_5_REG_1 <= s2_data_errors_0_5_REG; // @[ICacheMainPipe.scala 379:40]
    s2_data_errors_0_5_REG_2_0 <= ^data_full_wayBits__5_0; // @[ECC.scala 87:27]
    s2_data_errors_0_5_REG_2_1 <= ^data_full_wayBits__5_1; // @[ECC.scala 87:27]
    s2_data_errors_0_5_REG_2_2 <= ^data_full_wayBits__5_2; // @[ECC.scala 87:27]
    s2_data_errors_0_5_REG_2_3 <= ^data_full_wayBits__5_3; // @[ECC.scala 87:27]
    s2_data_errors_0_5_REG_2_4 <= ^data_full_wayBits__5_4; // @[ECC.scala 87:27]
    s2_data_errors_0_5_REG_2_5 <= ^data_full_wayBits__5_5; // @[ECC.scala 87:27]
    s2_data_errors_0_5_REG_2_6 <= ^data_full_wayBits__5_6; // @[ECC.scala 87:27]
    s2_data_errors_0_5_REG_2_7 <= ^data_full_wayBits__5_7; // @[ECC.scala 87:27]
    s2_data_errors_0_5_REG_2_8 <= ^data_full_wayBits__5_8; // @[ECC.scala 87:27]
    s2_data_errors_0_5_REG_2_9 <= ^data_full_wayBits__5_9; // @[ECC.scala 87:27]
    s2_data_errors_0_5_REG_2_10 <= ^data_full_wayBits__5_10; // @[ECC.scala 87:27]
    s2_data_errors_0_5_REG_2_11 <= ^data_full_wayBits__5_11; // @[ECC.scala 87:27]
    s2_data_errors_0_5_REG_2_12 <= ^data_full_wayBits__5_12; // @[ECC.scala 87:27]
    s2_data_errors_0_5_REG_2_13 <= ^data_full_wayBits__5_13; // @[ECC.scala 87:27]
    s2_data_errors_0_5_REG_2_14 <= ^data_full_wayBits__5_14; // @[ECC.scala 87:27]
    s2_data_errors_0_5_REG_2_15 <= ^data_full_wayBits__5_15; // @[ECC.scala 87:27]
    s2_data_errors_0_5_REG_2_16 <= ^data_full_wayBits__5_16; // @[ECC.scala 87:27]
    s2_data_errors_0_5_REG_2_17 <= ^data_full_wayBits__5_17; // @[ECC.scala 87:27]
    s2_data_errors_0_5_REG_2_18 <= ^data_full_wayBits__5_18; // @[ECC.scala 87:27]
    s2_data_errors_0_5_REG_2_19 <= ^data_full_wayBits__5_19; // @[ECC.scala 87:27]
    s2_data_errors_0_5_REG_2_20 <= ^data_full_wayBits__5_20; // @[ECC.scala 87:27]
    s2_data_errors_0_5_REG_2_21 <= ^data_full_wayBits__5_21; // @[ECC.scala 87:27]
    s2_data_errors_0_5_REG_2_22 <= ^data_full_wayBits__5_22; // @[ECC.scala 87:27]
    s2_data_errors_0_5_REG_2_23 <= ^data_full_wayBits__5_23; // @[ECC.scala 87:27]
    s2_data_errors_0_5_REG_2_24 <= ^data_full_wayBits__5_24; // @[ECC.scala 87:27]
    s2_data_errors_0_5_REG_2_25 <= ^data_full_wayBits__5_25; // @[ECC.scala 87:27]
    s2_data_errors_0_5_REG_2_26 <= ^data_full_wayBits__5_26; // @[ECC.scala 87:27]
    s2_data_errors_0_5_REG_2_27 <= ^data_full_wayBits__5_27; // @[ECC.scala 87:27]
    s2_data_errors_0_5_REG_2_28 <= ^data_full_wayBits__5_28; // @[ECC.scala 87:27]
    s2_data_errors_0_5_REG_2_29 <= ^data_full_wayBits__5_29; // @[ECC.scala 87:27]
    s2_data_errors_0_5_REG_2_30 <= ^data_full_wayBits__5_30; // @[ECC.scala 87:27]
    s2_data_errors_0_5_REG_2_31 <= ^data_full_wayBits__5_31; // @[ECC.scala 87:27]
    s2_data_errors_0_6_REG <= s1_valid & tlbRespAllValid & s2_ready; // @[ICacheMainPipe.scala 270:43]
    s2_data_errors_0_6_REG_1 <= s2_data_errors_0_6_REG; // @[ICacheMainPipe.scala 379:40]
    s2_data_errors_0_6_REG_2_0 <= ^data_full_wayBits__6_0; // @[ECC.scala 87:27]
    s2_data_errors_0_6_REG_2_1 <= ^data_full_wayBits__6_1; // @[ECC.scala 87:27]
    s2_data_errors_0_6_REG_2_2 <= ^data_full_wayBits__6_2; // @[ECC.scala 87:27]
    s2_data_errors_0_6_REG_2_3 <= ^data_full_wayBits__6_3; // @[ECC.scala 87:27]
    s2_data_errors_0_6_REG_2_4 <= ^data_full_wayBits__6_4; // @[ECC.scala 87:27]
    s2_data_errors_0_6_REG_2_5 <= ^data_full_wayBits__6_5; // @[ECC.scala 87:27]
    s2_data_errors_0_6_REG_2_6 <= ^data_full_wayBits__6_6; // @[ECC.scala 87:27]
    s2_data_errors_0_6_REG_2_7 <= ^data_full_wayBits__6_7; // @[ECC.scala 87:27]
    s2_data_errors_0_6_REG_2_8 <= ^data_full_wayBits__6_8; // @[ECC.scala 87:27]
    s2_data_errors_0_6_REG_2_9 <= ^data_full_wayBits__6_9; // @[ECC.scala 87:27]
    s2_data_errors_0_6_REG_2_10 <= ^data_full_wayBits__6_10; // @[ECC.scala 87:27]
    s2_data_errors_0_6_REG_2_11 <= ^data_full_wayBits__6_11; // @[ECC.scala 87:27]
    s2_data_errors_0_6_REG_2_12 <= ^data_full_wayBits__6_12; // @[ECC.scala 87:27]
    s2_data_errors_0_6_REG_2_13 <= ^data_full_wayBits__6_13; // @[ECC.scala 87:27]
    s2_data_errors_0_6_REG_2_14 <= ^data_full_wayBits__6_14; // @[ECC.scala 87:27]
    s2_data_errors_0_6_REG_2_15 <= ^data_full_wayBits__6_15; // @[ECC.scala 87:27]
    s2_data_errors_0_6_REG_2_16 <= ^data_full_wayBits__6_16; // @[ECC.scala 87:27]
    s2_data_errors_0_6_REG_2_17 <= ^data_full_wayBits__6_17; // @[ECC.scala 87:27]
    s2_data_errors_0_6_REG_2_18 <= ^data_full_wayBits__6_18; // @[ECC.scala 87:27]
    s2_data_errors_0_6_REG_2_19 <= ^data_full_wayBits__6_19; // @[ECC.scala 87:27]
    s2_data_errors_0_6_REG_2_20 <= ^data_full_wayBits__6_20; // @[ECC.scala 87:27]
    s2_data_errors_0_6_REG_2_21 <= ^data_full_wayBits__6_21; // @[ECC.scala 87:27]
    s2_data_errors_0_6_REG_2_22 <= ^data_full_wayBits__6_22; // @[ECC.scala 87:27]
    s2_data_errors_0_6_REG_2_23 <= ^data_full_wayBits__6_23; // @[ECC.scala 87:27]
    s2_data_errors_0_6_REG_2_24 <= ^data_full_wayBits__6_24; // @[ECC.scala 87:27]
    s2_data_errors_0_6_REG_2_25 <= ^data_full_wayBits__6_25; // @[ECC.scala 87:27]
    s2_data_errors_0_6_REG_2_26 <= ^data_full_wayBits__6_26; // @[ECC.scala 87:27]
    s2_data_errors_0_6_REG_2_27 <= ^data_full_wayBits__6_27; // @[ECC.scala 87:27]
    s2_data_errors_0_6_REG_2_28 <= ^data_full_wayBits__6_28; // @[ECC.scala 87:27]
    s2_data_errors_0_6_REG_2_29 <= ^data_full_wayBits__6_29; // @[ECC.scala 87:27]
    s2_data_errors_0_6_REG_2_30 <= ^data_full_wayBits__6_30; // @[ECC.scala 87:27]
    s2_data_errors_0_6_REG_2_31 <= ^data_full_wayBits__6_31; // @[ECC.scala 87:27]
    s2_data_errors_0_7_REG <= s1_valid & tlbRespAllValid & s2_ready; // @[ICacheMainPipe.scala 270:43]
    s2_data_errors_0_7_REG_1 <= s2_data_errors_0_7_REG; // @[ICacheMainPipe.scala 379:40]
    s2_data_errors_0_7_REG_2_0 <= ^data_full_wayBits__7_0; // @[ECC.scala 87:27]
    s2_data_errors_0_7_REG_2_1 <= ^data_full_wayBits__7_1; // @[ECC.scala 87:27]
    s2_data_errors_0_7_REG_2_2 <= ^data_full_wayBits__7_2; // @[ECC.scala 87:27]
    s2_data_errors_0_7_REG_2_3 <= ^data_full_wayBits__7_3; // @[ECC.scala 87:27]
    s2_data_errors_0_7_REG_2_4 <= ^data_full_wayBits__7_4; // @[ECC.scala 87:27]
    s2_data_errors_0_7_REG_2_5 <= ^data_full_wayBits__7_5; // @[ECC.scala 87:27]
    s2_data_errors_0_7_REG_2_6 <= ^data_full_wayBits__7_6; // @[ECC.scala 87:27]
    s2_data_errors_0_7_REG_2_7 <= ^data_full_wayBits__7_7; // @[ECC.scala 87:27]
    s2_data_errors_0_7_REG_2_8 <= ^data_full_wayBits__7_8; // @[ECC.scala 87:27]
    s2_data_errors_0_7_REG_2_9 <= ^data_full_wayBits__7_9; // @[ECC.scala 87:27]
    s2_data_errors_0_7_REG_2_10 <= ^data_full_wayBits__7_10; // @[ECC.scala 87:27]
    s2_data_errors_0_7_REG_2_11 <= ^data_full_wayBits__7_11; // @[ECC.scala 87:27]
    s2_data_errors_0_7_REG_2_12 <= ^data_full_wayBits__7_12; // @[ECC.scala 87:27]
    s2_data_errors_0_7_REG_2_13 <= ^data_full_wayBits__7_13; // @[ECC.scala 87:27]
    s2_data_errors_0_7_REG_2_14 <= ^data_full_wayBits__7_14; // @[ECC.scala 87:27]
    s2_data_errors_0_7_REG_2_15 <= ^data_full_wayBits__7_15; // @[ECC.scala 87:27]
    s2_data_errors_0_7_REG_2_16 <= ^data_full_wayBits__7_16; // @[ECC.scala 87:27]
    s2_data_errors_0_7_REG_2_17 <= ^data_full_wayBits__7_17; // @[ECC.scala 87:27]
    s2_data_errors_0_7_REG_2_18 <= ^data_full_wayBits__7_18; // @[ECC.scala 87:27]
    s2_data_errors_0_7_REG_2_19 <= ^data_full_wayBits__7_19; // @[ECC.scala 87:27]
    s2_data_errors_0_7_REG_2_20 <= ^data_full_wayBits__7_20; // @[ECC.scala 87:27]
    s2_data_errors_0_7_REG_2_21 <= ^data_full_wayBits__7_21; // @[ECC.scala 87:27]
    s2_data_errors_0_7_REG_2_22 <= ^data_full_wayBits__7_22; // @[ECC.scala 87:27]
    s2_data_errors_0_7_REG_2_23 <= ^data_full_wayBits__7_23; // @[ECC.scala 87:27]
    s2_data_errors_0_7_REG_2_24 <= ^data_full_wayBits__7_24; // @[ECC.scala 87:27]
    s2_data_errors_0_7_REG_2_25 <= ^data_full_wayBits__7_25; // @[ECC.scala 87:27]
    s2_data_errors_0_7_REG_2_26 <= ^data_full_wayBits__7_26; // @[ECC.scala 87:27]
    s2_data_errors_0_7_REG_2_27 <= ^data_full_wayBits__7_27; // @[ECC.scala 87:27]
    s2_data_errors_0_7_REG_2_28 <= ^data_full_wayBits__7_28; // @[ECC.scala 87:27]
    s2_data_errors_0_7_REG_2_29 <= ^data_full_wayBits__7_29; // @[ECC.scala 87:27]
    s2_data_errors_0_7_REG_2_30 <= ^data_full_wayBits__7_30; // @[ECC.scala 87:27]
    s2_data_errors_0_7_REG_2_31 <= ^data_full_wayBits__7_31; // @[ECC.scala 87:27]
    s2_data_errors_1_0_REG <= s1_valid & tlbRespAllValid & s2_ready; // @[ICacheMainPipe.scala 270:43]
    s2_data_errors_1_0_REG_1 <= s2_data_errors_1_0_REG; // @[ICacheMainPipe.scala 383:40]
    s2_data_errors_1_0_REG_2 <= s1_double_line; // @[ICacheMainPipe.scala 383:77]
    s2_data_errors_1_0_REG_3 <= s2_data_errors_1_0_REG_2; // @[ICacheMainPipe.scala 383:69]
    s2_data_errors_1_0_REG_4_0 <= ^data_full_wayBits_1_0_0; // @[ECC.scala 87:27]
    s2_data_errors_1_0_REG_4_1 <= ^data_full_wayBits_1_0_1; // @[ECC.scala 87:27]
    s2_data_errors_1_0_REG_4_2 <= ^data_full_wayBits_1_0_2; // @[ECC.scala 87:27]
    s2_data_errors_1_0_REG_4_3 <= ^data_full_wayBits_1_0_3; // @[ECC.scala 87:27]
    s2_data_errors_1_0_REG_4_4 <= ^data_full_wayBits_1_0_4; // @[ECC.scala 87:27]
    s2_data_errors_1_0_REG_4_5 <= ^data_full_wayBits_1_0_5; // @[ECC.scala 87:27]
    s2_data_errors_1_0_REG_4_6 <= ^data_full_wayBits_1_0_6; // @[ECC.scala 87:27]
    s2_data_errors_1_0_REG_4_7 <= ^data_full_wayBits_1_0_7; // @[ECC.scala 87:27]
    s2_data_errors_1_0_REG_4_8 <= ^data_full_wayBits_1_0_8; // @[ECC.scala 87:27]
    s2_data_errors_1_0_REG_4_9 <= ^data_full_wayBits_1_0_9; // @[ECC.scala 87:27]
    s2_data_errors_1_0_REG_4_10 <= ^data_full_wayBits_1_0_10; // @[ECC.scala 87:27]
    s2_data_errors_1_0_REG_4_11 <= ^data_full_wayBits_1_0_11; // @[ECC.scala 87:27]
    s2_data_errors_1_0_REG_4_12 <= ^data_full_wayBits_1_0_12; // @[ECC.scala 87:27]
    s2_data_errors_1_0_REG_4_13 <= ^data_full_wayBits_1_0_13; // @[ECC.scala 87:27]
    s2_data_errors_1_0_REG_4_14 <= ^data_full_wayBits_1_0_14; // @[ECC.scala 87:27]
    s2_data_errors_1_0_REG_4_15 <= ^data_full_wayBits_1_0_15; // @[ECC.scala 87:27]
    s2_data_errors_1_0_REG_4_16 <= ^data_full_wayBits_1_0_16; // @[ECC.scala 87:27]
    s2_data_errors_1_0_REG_4_17 <= ^data_full_wayBits_1_0_17; // @[ECC.scala 87:27]
    s2_data_errors_1_0_REG_4_18 <= ^data_full_wayBits_1_0_18; // @[ECC.scala 87:27]
    s2_data_errors_1_0_REG_4_19 <= ^data_full_wayBits_1_0_19; // @[ECC.scala 87:27]
    s2_data_errors_1_0_REG_4_20 <= ^data_full_wayBits_1_0_20; // @[ECC.scala 87:27]
    s2_data_errors_1_0_REG_4_21 <= ^data_full_wayBits_1_0_21; // @[ECC.scala 87:27]
    s2_data_errors_1_0_REG_4_22 <= ^data_full_wayBits_1_0_22; // @[ECC.scala 87:27]
    s2_data_errors_1_0_REG_4_23 <= ^data_full_wayBits_1_0_23; // @[ECC.scala 87:27]
    s2_data_errors_1_0_REG_4_24 <= ^data_full_wayBits_1_0_24; // @[ECC.scala 87:27]
    s2_data_errors_1_0_REG_4_25 <= ^data_full_wayBits_1_0_25; // @[ECC.scala 87:27]
    s2_data_errors_1_0_REG_4_26 <= ^data_full_wayBits_1_0_26; // @[ECC.scala 87:27]
    s2_data_errors_1_0_REG_4_27 <= ^data_full_wayBits_1_0_27; // @[ECC.scala 87:27]
    s2_data_errors_1_0_REG_4_28 <= ^data_full_wayBits_1_0_28; // @[ECC.scala 87:27]
    s2_data_errors_1_0_REG_4_29 <= ^data_full_wayBits_1_0_29; // @[ECC.scala 87:27]
    s2_data_errors_1_0_REG_4_30 <= ^data_full_wayBits_1_0_30; // @[ECC.scala 87:27]
    s2_data_errors_1_0_REG_4_31 <= ^data_full_wayBits_1_0_31; // @[ECC.scala 87:27]
    s2_data_errors_1_1_REG <= s1_valid & tlbRespAllValid & s2_ready; // @[ICacheMainPipe.scala 270:43]
    s2_data_errors_1_1_REG_1 <= s2_data_errors_1_1_REG; // @[ICacheMainPipe.scala 383:40]
    s2_data_errors_1_1_REG_2 <= s1_double_line; // @[ICacheMainPipe.scala 383:77]
    s2_data_errors_1_1_REG_3 <= s2_data_errors_1_1_REG_2; // @[ICacheMainPipe.scala 383:69]
    s2_data_errors_1_1_REG_4_0 <= ^data_full_wayBits_1_1_0; // @[ECC.scala 87:27]
    s2_data_errors_1_1_REG_4_1 <= ^data_full_wayBits_1_1_1; // @[ECC.scala 87:27]
    s2_data_errors_1_1_REG_4_2 <= ^data_full_wayBits_1_1_2; // @[ECC.scala 87:27]
    s2_data_errors_1_1_REG_4_3 <= ^data_full_wayBits_1_1_3; // @[ECC.scala 87:27]
    s2_data_errors_1_1_REG_4_4 <= ^data_full_wayBits_1_1_4; // @[ECC.scala 87:27]
    s2_data_errors_1_1_REG_4_5 <= ^data_full_wayBits_1_1_5; // @[ECC.scala 87:27]
    s2_data_errors_1_1_REG_4_6 <= ^data_full_wayBits_1_1_6; // @[ECC.scala 87:27]
    s2_data_errors_1_1_REG_4_7 <= ^data_full_wayBits_1_1_7; // @[ECC.scala 87:27]
    s2_data_errors_1_1_REG_4_8 <= ^data_full_wayBits_1_1_8; // @[ECC.scala 87:27]
    s2_data_errors_1_1_REG_4_9 <= ^data_full_wayBits_1_1_9; // @[ECC.scala 87:27]
    s2_data_errors_1_1_REG_4_10 <= ^data_full_wayBits_1_1_10; // @[ECC.scala 87:27]
    s2_data_errors_1_1_REG_4_11 <= ^data_full_wayBits_1_1_11; // @[ECC.scala 87:27]
    s2_data_errors_1_1_REG_4_12 <= ^data_full_wayBits_1_1_12; // @[ECC.scala 87:27]
    s2_data_errors_1_1_REG_4_13 <= ^data_full_wayBits_1_1_13; // @[ECC.scala 87:27]
    s2_data_errors_1_1_REG_4_14 <= ^data_full_wayBits_1_1_14; // @[ECC.scala 87:27]
    s2_data_errors_1_1_REG_4_15 <= ^data_full_wayBits_1_1_15; // @[ECC.scala 87:27]
    s2_data_errors_1_1_REG_4_16 <= ^data_full_wayBits_1_1_16; // @[ECC.scala 87:27]
    s2_data_errors_1_1_REG_4_17 <= ^data_full_wayBits_1_1_17; // @[ECC.scala 87:27]
    s2_data_errors_1_1_REG_4_18 <= ^data_full_wayBits_1_1_18; // @[ECC.scala 87:27]
    s2_data_errors_1_1_REG_4_19 <= ^data_full_wayBits_1_1_19; // @[ECC.scala 87:27]
    s2_data_errors_1_1_REG_4_20 <= ^data_full_wayBits_1_1_20; // @[ECC.scala 87:27]
    s2_data_errors_1_1_REG_4_21 <= ^data_full_wayBits_1_1_21; // @[ECC.scala 87:27]
    s2_data_errors_1_1_REG_4_22 <= ^data_full_wayBits_1_1_22; // @[ECC.scala 87:27]
    s2_data_errors_1_1_REG_4_23 <= ^data_full_wayBits_1_1_23; // @[ECC.scala 87:27]
    s2_data_errors_1_1_REG_4_24 <= ^data_full_wayBits_1_1_24; // @[ECC.scala 87:27]
    s2_data_errors_1_1_REG_4_25 <= ^data_full_wayBits_1_1_25; // @[ECC.scala 87:27]
    s2_data_errors_1_1_REG_4_26 <= ^data_full_wayBits_1_1_26; // @[ECC.scala 87:27]
    s2_data_errors_1_1_REG_4_27 <= ^data_full_wayBits_1_1_27; // @[ECC.scala 87:27]
    s2_data_errors_1_1_REG_4_28 <= ^data_full_wayBits_1_1_28; // @[ECC.scala 87:27]
    s2_data_errors_1_1_REG_4_29 <= ^data_full_wayBits_1_1_29; // @[ECC.scala 87:27]
    s2_data_errors_1_1_REG_4_30 <= ^data_full_wayBits_1_1_30; // @[ECC.scala 87:27]
    s2_data_errors_1_1_REG_4_31 <= ^data_full_wayBits_1_1_31; // @[ECC.scala 87:27]
    s2_data_errors_1_2_REG <= s1_valid & tlbRespAllValid & s2_ready; // @[ICacheMainPipe.scala 270:43]
    s2_data_errors_1_2_REG_1 <= s2_data_errors_1_2_REG; // @[ICacheMainPipe.scala 383:40]
    s2_data_errors_1_2_REG_2 <= s1_double_line; // @[ICacheMainPipe.scala 383:77]
    s2_data_errors_1_2_REG_3 <= s2_data_errors_1_2_REG_2; // @[ICacheMainPipe.scala 383:69]
    s2_data_errors_1_2_REG_4_0 <= ^data_full_wayBits_1_2_0; // @[ECC.scala 87:27]
    s2_data_errors_1_2_REG_4_1 <= ^data_full_wayBits_1_2_1; // @[ECC.scala 87:27]
    s2_data_errors_1_2_REG_4_2 <= ^data_full_wayBits_1_2_2; // @[ECC.scala 87:27]
    s2_data_errors_1_2_REG_4_3 <= ^data_full_wayBits_1_2_3; // @[ECC.scala 87:27]
    s2_data_errors_1_2_REG_4_4 <= ^data_full_wayBits_1_2_4; // @[ECC.scala 87:27]
    s2_data_errors_1_2_REG_4_5 <= ^data_full_wayBits_1_2_5; // @[ECC.scala 87:27]
    s2_data_errors_1_2_REG_4_6 <= ^data_full_wayBits_1_2_6; // @[ECC.scala 87:27]
    s2_data_errors_1_2_REG_4_7 <= ^data_full_wayBits_1_2_7; // @[ECC.scala 87:27]
    s2_data_errors_1_2_REG_4_8 <= ^data_full_wayBits_1_2_8; // @[ECC.scala 87:27]
    s2_data_errors_1_2_REG_4_9 <= ^data_full_wayBits_1_2_9; // @[ECC.scala 87:27]
    s2_data_errors_1_2_REG_4_10 <= ^data_full_wayBits_1_2_10; // @[ECC.scala 87:27]
    s2_data_errors_1_2_REG_4_11 <= ^data_full_wayBits_1_2_11; // @[ECC.scala 87:27]
    s2_data_errors_1_2_REG_4_12 <= ^data_full_wayBits_1_2_12; // @[ECC.scala 87:27]
    s2_data_errors_1_2_REG_4_13 <= ^data_full_wayBits_1_2_13; // @[ECC.scala 87:27]
    s2_data_errors_1_2_REG_4_14 <= ^data_full_wayBits_1_2_14; // @[ECC.scala 87:27]
    s2_data_errors_1_2_REG_4_15 <= ^data_full_wayBits_1_2_15; // @[ECC.scala 87:27]
    s2_data_errors_1_2_REG_4_16 <= ^data_full_wayBits_1_2_16; // @[ECC.scala 87:27]
    s2_data_errors_1_2_REG_4_17 <= ^data_full_wayBits_1_2_17; // @[ECC.scala 87:27]
    s2_data_errors_1_2_REG_4_18 <= ^data_full_wayBits_1_2_18; // @[ECC.scala 87:27]
    s2_data_errors_1_2_REG_4_19 <= ^data_full_wayBits_1_2_19; // @[ECC.scala 87:27]
    s2_data_errors_1_2_REG_4_20 <= ^data_full_wayBits_1_2_20; // @[ECC.scala 87:27]
    s2_data_errors_1_2_REG_4_21 <= ^data_full_wayBits_1_2_21; // @[ECC.scala 87:27]
    s2_data_errors_1_2_REG_4_22 <= ^data_full_wayBits_1_2_22; // @[ECC.scala 87:27]
    s2_data_errors_1_2_REG_4_23 <= ^data_full_wayBits_1_2_23; // @[ECC.scala 87:27]
    s2_data_errors_1_2_REG_4_24 <= ^data_full_wayBits_1_2_24; // @[ECC.scala 87:27]
    s2_data_errors_1_2_REG_4_25 <= ^data_full_wayBits_1_2_25; // @[ECC.scala 87:27]
    s2_data_errors_1_2_REG_4_26 <= ^data_full_wayBits_1_2_26; // @[ECC.scala 87:27]
    s2_data_errors_1_2_REG_4_27 <= ^data_full_wayBits_1_2_27; // @[ECC.scala 87:27]
    s2_data_errors_1_2_REG_4_28 <= ^data_full_wayBits_1_2_28; // @[ECC.scala 87:27]
    s2_data_errors_1_2_REG_4_29 <= ^data_full_wayBits_1_2_29; // @[ECC.scala 87:27]
    s2_data_errors_1_2_REG_4_30 <= ^data_full_wayBits_1_2_30; // @[ECC.scala 87:27]
    s2_data_errors_1_2_REG_4_31 <= ^data_full_wayBits_1_2_31; // @[ECC.scala 87:27]
    s2_data_errors_1_3_REG <= s1_valid & tlbRespAllValid & s2_ready; // @[ICacheMainPipe.scala 270:43]
    s2_data_errors_1_3_REG_1 <= s2_data_errors_1_3_REG; // @[ICacheMainPipe.scala 383:40]
    s2_data_errors_1_3_REG_2 <= s1_double_line; // @[ICacheMainPipe.scala 383:77]
    s2_data_errors_1_3_REG_3 <= s2_data_errors_1_3_REG_2; // @[ICacheMainPipe.scala 383:69]
    s2_data_errors_1_3_REG_4_0 <= ^data_full_wayBits_1_3_0; // @[ECC.scala 87:27]
    s2_data_errors_1_3_REG_4_1 <= ^data_full_wayBits_1_3_1; // @[ECC.scala 87:27]
    s2_data_errors_1_3_REG_4_2 <= ^data_full_wayBits_1_3_2; // @[ECC.scala 87:27]
    s2_data_errors_1_3_REG_4_3 <= ^data_full_wayBits_1_3_3; // @[ECC.scala 87:27]
    s2_data_errors_1_3_REG_4_4 <= ^data_full_wayBits_1_3_4; // @[ECC.scala 87:27]
    s2_data_errors_1_3_REG_4_5 <= ^data_full_wayBits_1_3_5; // @[ECC.scala 87:27]
    s2_data_errors_1_3_REG_4_6 <= ^data_full_wayBits_1_3_6; // @[ECC.scala 87:27]
    s2_data_errors_1_3_REG_4_7 <= ^data_full_wayBits_1_3_7; // @[ECC.scala 87:27]
    s2_data_errors_1_3_REG_4_8 <= ^data_full_wayBits_1_3_8; // @[ECC.scala 87:27]
    s2_data_errors_1_3_REG_4_9 <= ^data_full_wayBits_1_3_9; // @[ECC.scala 87:27]
    s2_data_errors_1_3_REG_4_10 <= ^data_full_wayBits_1_3_10; // @[ECC.scala 87:27]
    s2_data_errors_1_3_REG_4_11 <= ^data_full_wayBits_1_3_11; // @[ECC.scala 87:27]
    s2_data_errors_1_3_REG_4_12 <= ^data_full_wayBits_1_3_12; // @[ECC.scala 87:27]
    s2_data_errors_1_3_REG_4_13 <= ^data_full_wayBits_1_3_13; // @[ECC.scala 87:27]
    s2_data_errors_1_3_REG_4_14 <= ^data_full_wayBits_1_3_14; // @[ECC.scala 87:27]
    s2_data_errors_1_3_REG_4_15 <= ^data_full_wayBits_1_3_15; // @[ECC.scala 87:27]
    s2_data_errors_1_3_REG_4_16 <= ^data_full_wayBits_1_3_16; // @[ECC.scala 87:27]
    s2_data_errors_1_3_REG_4_17 <= ^data_full_wayBits_1_3_17; // @[ECC.scala 87:27]
    s2_data_errors_1_3_REG_4_18 <= ^data_full_wayBits_1_3_18; // @[ECC.scala 87:27]
    s2_data_errors_1_3_REG_4_19 <= ^data_full_wayBits_1_3_19; // @[ECC.scala 87:27]
    s2_data_errors_1_3_REG_4_20 <= ^data_full_wayBits_1_3_20; // @[ECC.scala 87:27]
    s2_data_errors_1_3_REG_4_21 <= ^data_full_wayBits_1_3_21; // @[ECC.scala 87:27]
    s2_data_errors_1_3_REG_4_22 <= ^data_full_wayBits_1_3_22; // @[ECC.scala 87:27]
    s2_data_errors_1_3_REG_4_23 <= ^data_full_wayBits_1_3_23; // @[ECC.scala 87:27]
    s2_data_errors_1_3_REG_4_24 <= ^data_full_wayBits_1_3_24; // @[ECC.scala 87:27]
    s2_data_errors_1_3_REG_4_25 <= ^data_full_wayBits_1_3_25; // @[ECC.scala 87:27]
    s2_data_errors_1_3_REG_4_26 <= ^data_full_wayBits_1_3_26; // @[ECC.scala 87:27]
    s2_data_errors_1_3_REG_4_27 <= ^data_full_wayBits_1_3_27; // @[ECC.scala 87:27]
    s2_data_errors_1_3_REG_4_28 <= ^data_full_wayBits_1_3_28; // @[ECC.scala 87:27]
    s2_data_errors_1_3_REG_4_29 <= ^data_full_wayBits_1_3_29; // @[ECC.scala 87:27]
    s2_data_errors_1_3_REG_4_30 <= ^data_full_wayBits_1_3_30; // @[ECC.scala 87:27]
    s2_data_errors_1_3_REG_4_31 <= ^data_full_wayBits_1_3_31; // @[ECC.scala 87:27]
    s2_data_errors_1_4_REG <= s1_valid & tlbRespAllValid & s2_ready; // @[ICacheMainPipe.scala 270:43]
    s2_data_errors_1_4_REG_1 <= s2_data_errors_1_4_REG; // @[ICacheMainPipe.scala 383:40]
    s2_data_errors_1_4_REG_2 <= s1_double_line; // @[ICacheMainPipe.scala 383:77]
    s2_data_errors_1_4_REG_3 <= s2_data_errors_1_4_REG_2; // @[ICacheMainPipe.scala 383:69]
    s2_data_errors_1_4_REG_4_0 <= ^data_full_wayBits_1_4_0; // @[ECC.scala 87:27]
    s2_data_errors_1_4_REG_4_1 <= ^data_full_wayBits_1_4_1; // @[ECC.scala 87:27]
    s2_data_errors_1_4_REG_4_2 <= ^data_full_wayBits_1_4_2; // @[ECC.scala 87:27]
    s2_data_errors_1_4_REG_4_3 <= ^data_full_wayBits_1_4_3; // @[ECC.scala 87:27]
    s2_data_errors_1_4_REG_4_4 <= ^data_full_wayBits_1_4_4; // @[ECC.scala 87:27]
    s2_data_errors_1_4_REG_4_5 <= ^data_full_wayBits_1_4_5; // @[ECC.scala 87:27]
    s2_data_errors_1_4_REG_4_6 <= ^data_full_wayBits_1_4_6; // @[ECC.scala 87:27]
    s2_data_errors_1_4_REG_4_7 <= ^data_full_wayBits_1_4_7; // @[ECC.scala 87:27]
    s2_data_errors_1_4_REG_4_8 <= ^data_full_wayBits_1_4_8; // @[ECC.scala 87:27]
    s2_data_errors_1_4_REG_4_9 <= ^data_full_wayBits_1_4_9; // @[ECC.scala 87:27]
    s2_data_errors_1_4_REG_4_10 <= ^data_full_wayBits_1_4_10; // @[ECC.scala 87:27]
    s2_data_errors_1_4_REG_4_11 <= ^data_full_wayBits_1_4_11; // @[ECC.scala 87:27]
    s2_data_errors_1_4_REG_4_12 <= ^data_full_wayBits_1_4_12; // @[ECC.scala 87:27]
    s2_data_errors_1_4_REG_4_13 <= ^data_full_wayBits_1_4_13; // @[ECC.scala 87:27]
    s2_data_errors_1_4_REG_4_14 <= ^data_full_wayBits_1_4_14; // @[ECC.scala 87:27]
    s2_data_errors_1_4_REG_4_15 <= ^data_full_wayBits_1_4_15; // @[ECC.scala 87:27]
    s2_data_errors_1_4_REG_4_16 <= ^data_full_wayBits_1_4_16; // @[ECC.scala 87:27]
    s2_data_errors_1_4_REG_4_17 <= ^data_full_wayBits_1_4_17; // @[ECC.scala 87:27]
    s2_data_errors_1_4_REG_4_18 <= ^data_full_wayBits_1_4_18; // @[ECC.scala 87:27]
    s2_data_errors_1_4_REG_4_19 <= ^data_full_wayBits_1_4_19; // @[ECC.scala 87:27]
    s2_data_errors_1_4_REG_4_20 <= ^data_full_wayBits_1_4_20; // @[ECC.scala 87:27]
    s2_data_errors_1_4_REG_4_21 <= ^data_full_wayBits_1_4_21; // @[ECC.scala 87:27]
    s2_data_errors_1_4_REG_4_22 <= ^data_full_wayBits_1_4_22; // @[ECC.scala 87:27]
    s2_data_errors_1_4_REG_4_23 <= ^data_full_wayBits_1_4_23; // @[ECC.scala 87:27]
    s2_data_errors_1_4_REG_4_24 <= ^data_full_wayBits_1_4_24; // @[ECC.scala 87:27]
    s2_data_errors_1_4_REG_4_25 <= ^data_full_wayBits_1_4_25; // @[ECC.scala 87:27]
    s2_data_errors_1_4_REG_4_26 <= ^data_full_wayBits_1_4_26; // @[ECC.scala 87:27]
    s2_data_errors_1_4_REG_4_27 <= ^data_full_wayBits_1_4_27; // @[ECC.scala 87:27]
    s2_data_errors_1_4_REG_4_28 <= ^data_full_wayBits_1_4_28; // @[ECC.scala 87:27]
    s2_data_errors_1_4_REG_4_29 <= ^data_full_wayBits_1_4_29; // @[ECC.scala 87:27]
    s2_data_errors_1_4_REG_4_30 <= ^data_full_wayBits_1_4_30; // @[ECC.scala 87:27]
    s2_data_errors_1_4_REG_4_31 <= ^data_full_wayBits_1_4_31; // @[ECC.scala 87:27]
    s2_data_errors_1_5_REG <= s1_valid & tlbRespAllValid & s2_ready; // @[ICacheMainPipe.scala 270:43]
    s2_data_errors_1_5_REG_1 <= s2_data_errors_1_5_REG; // @[ICacheMainPipe.scala 383:40]
    s2_data_errors_1_5_REG_2 <= s1_double_line; // @[ICacheMainPipe.scala 383:77]
    s2_data_errors_1_5_REG_3 <= s2_data_errors_1_5_REG_2; // @[ICacheMainPipe.scala 383:69]
    s2_data_errors_1_5_REG_4_0 <= ^data_full_wayBits_1_5_0; // @[ECC.scala 87:27]
    s2_data_errors_1_5_REG_4_1 <= ^data_full_wayBits_1_5_1; // @[ECC.scala 87:27]
    s2_data_errors_1_5_REG_4_2 <= ^data_full_wayBits_1_5_2; // @[ECC.scala 87:27]
    s2_data_errors_1_5_REG_4_3 <= ^data_full_wayBits_1_5_3; // @[ECC.scala 87:27]
    s2_data_errors_1_5_REG_4_4 <= ^data_full_wayBits_1_5_4; // @[ECC.scala 87:27]
    s2_data_errors_1_5_REG_4_5 <= ^data_full_wayBits_1_5_5; // @[ECC.scala 87:27]
    s2_data_errors_1_5_REG_4_6 <= ^data_full_wayBits_1_5_6; // @[ECC.scala 87:27]
    s2_data_errors_1_5_REG_4_7 <= ^data_full_wayBits_1_5_7; // @[ECC.scala 87:27]
    s2_data_errors_1_5_REG_4_8 <= ^data_full_wayBits_1_5_8; // @[ECC.scala 87:27]
    s2_data_errors_1_5_REG_4_9 <= ^data_full_wayBits_1_5_9; // @[ECC.scala 87:27]
    s2_data_errors_1_5_REG_4_10 <= ^data_full_wayBits_1_5_10; // @[ECC.scala 87:27]
    s2_data_errors_1_5_REG_4_11 <= ^data_full_wayBits_1_5_11; // @[ECC.scala 87:27]
    s2_data_errors_1_5_REG_4_12 <= ^data_full_wayBits_1_5_12; // @[ECC.scala 87:27]
    s2_data_errors_1_5_REG_4_13 <= ^data_full_wayBits_1_5_13; // @[ECC.scala 87:27]
    s2_data_errors_1_5_REG_4_14 <= ^data_full_wayBits_1_5_14; // @[ECC.scala 87:27]
    s2_data_errors_1_5_REG_4_15 <= ^data_full_wayBits_1_5_15; // @[ECC.scala 87:27]
    s2_data_errors_1_5_REG_4_16 <= ^data_full_wayBits_1_5_16; // @[ECC.scala 87:27]
    s2_data_errors_1_5_REG_4_17 <= ^data_full_wayBits_1_5_17; // @[ECC.scala 87:27]
    s2_data_errors_1_5_REG_4_18 <= ^data_full_wayBits_1_5_18; // @[ECC.scala 87:27]
    s2_data_errors_1_5_REG_4_19 <= ^data_full_wayBits_1_5_19; // @[ECC.scala 87:27]
    s2_data_errors_1_5_REG_4_20 <= ^data_full_wayBits_1_5_20; // @[ECC.scala 87:27]
    s2_data_errors_1_5_REG_4_21 <= ^data_full_wayBits_1_5_21; // @[ECC.scala 87:27]
    s2_data_errors_1_5_REG_4_22 <= ^data_full_wayBits_1_5_22; // @[ECC.scala 87:27]
    s2_data_errors_1_5_REG_4_23 <= ^data_full_wayBits_1_5_23; // @[ECC.scala 87:27]
    s2_data_errors_1_5_REG_4_24 <= ^data_full_wayBits_1_5_24; // @[ECC.scala 87:27]
    s2_data_errors_1_5_REG_4_25 <= ^data_full_wayBits_1_5_25; // @[ECC.scala 87:27]
    s2_data_errors_1_5_REG_4_26 <= ^data_full_wayBits_1_5_26; // @[ECC.scala 87:27]
    s2_data_errors_1_5_REG_4_27 <= ^data_full_wayBits_1_5_27; // @[ECC.scala 87:27]
    s2_data_errors_1_5_REG_4_28 <= ^data_full_wayBits_1_5_28; // @[ECC.scala 87:27]
    s2_data_errors_1_5_REG_4_29 <= ^data_full_wayBits_1_5_29; // @[ECC.scala 87:27]
    s2_data_errors_1_5_REG_4_30 <= ^data_full_wayBits_1_5_30; // @[ECC.scala 87:27]
    s2_data_errors_1_5_REG_4_31 <= ^data_full_wayBits_1_5_31; // @[ECC.scala 87:27]
    s2_data_errors_1_6_REG <= s1_valid & tlbRespAllValid & s2_ready; // @[ICacheMainPipe.scala 270:43]
    s2_data_errors_1_6_REG_1 <= s2_data_errors_1_6_REG; // @[ICacheMainPipe.scala 383:40]
    s2_data_errors_1_6_REG_2 <= s1_double_line; // @[ICacheMainPipe.scala 383:77]
    s2_data_errors_1_6_REG_3 <= s2_data_errors_1_6_REG_2; // @[ICacheMainPipe.scala 383:69]
    s2_data_errors_1_6_REG_4_0 <= ^data_full_wayBits_1_6_0; // @[ECC.scala 87:27]
    s2_data_errors_1_6_REG_4_1 <= ^data_full_wayBits_1_6_1; // @[ECC.scala 87:27]
    s2_data_errors_1_6_REG_4_2 <= ^data_full_wayBits_1_6_2; // @[ECC.scala 87:27]
    s2_data_errors_1_6_REG_4_3 <= ^data_full_wayBits_1_6_3; // @[ECC.scala 87:27]
    s2_data_errors_1_6_REG_4_4 <= ^data_full_wayBits_1_6_4; // @[ECC.scala 87:27]
    s2_data_errors_1_6_REG_4_5 <= ^data_full_wayBits_1_6_5; // @[ECC.scala 87:27]
    s2_data_errors_1_6_REG_4_6 <= ^data_full_wayBits_1_6_6; // @[ECC.scala 87:27]
    s2_data_errors_1_6_REG_4_7 <= ^data_full_wayBits_1_6_7; // @[ECC.scala 87:27]
    s2_data_errors_1_6_REG_4_8 <= ^data_full_wayBits_1_6_8; // @[ECC.scala 87:27]
    s2_data_errors_1_6_REG_4_9 <= ^data_full_wayBits_1_6_9; // @[ECC.scala 87:27]
    s2_data_errors_1_6_REG_4_10 <= ^data_full_wayBits_1_6_10; // @[ECC.scala 87:27]
    s2_data_errors_1_6_REG_4_11 <= ^data_full_wayBits_1_6_11; // @[ECC.scala 87:27]
    s2_data_errors_1_6_REG_4_12 <= ^data_full_wayBits_1_6_12; // @[ECC.scala 87:27]
    s2_data_errors_1_6_REG_4_13 <= ^data_full_wayBits_1_6_13; // @[ECC.scala 87:27]
    s2_data_errors_1_6_REG_4_14 <= ^data_full_wayBits_1_6_14; // @[ECC.scala 87:27]
    s2_data_errors_1_6_REG_4_15 <= ^data_full_wayBits_1_6_15; // @[ECC.scala 87:27]
    s2_data_errors_1_6_REG_4_16 <= ^data_full_wayBits_1_6_16; // @[ECC.scala 87:27]
    s2_data_errors_1_6_REG_4_17 <= ^data_full_wayBits_1_6_17; // @[ECC.scala 87:27]
    s2_data_errors_1_6_REG_4_18 <= ^data_full_wayBits_1_6_18; // @[ECC.scala 87:27]
    s2_data_errors_1_6_REG_4_19 <= ^data_full_wayBits_1_6_19; // @[ECC.scala 87:27]
    s2_data_errors_1_6_REG_4_20 <= ^data_full_wayBits_1_6_20; // @[ECC.scala 87:27]
    s2_data_errors_1_6_REG_4_21 <= ^data_full_wayBits_1_6_21; // @[ECC.scala 87:27]
    s2_data_errors_1_6_REG_4_22 <= ^data_full_wayBits_1_6_22; // @[ECC.scala 87:27]
    s2_data_errors_1_6_REG_4_23 <= ^data_full_wayBits_1_6_23; // @[ECC.scala 87:27]
    s2_data_errors_1_6_REG_4_24 <= ^data_full_wayBits_1_6_24; // @[ECC.scala 87:27]
    s2_data_errors_1_6_REG_4_25 <= ^data_full_wayBits_1_6_25; // @[ECC.scala 87:27]
    s2_data_errors_1_6_REG_4_26 <= ^data_full_wayBits_1_6_26; // @[ECC.scala 87:27]
    s2_data_errors_1_6_REG_4_27 <= ^data_full_wayBits_1_6_27; // @[ECC.scala 87:27]
    s2_data_errors_1_6_REG_4_28 <= ^data_full_wayBits_1_6_28; // @[ECC.scala 87:27]
    s2_data_errors_1_6_REG_4_29 <= ^data_full_wayBits_1_6_29; // @[ECC.scala 87:27]
    s2_data_errors_1_6_REG_4_30 <= ^data_full_wayBits_1_6_30; // @[ECC.scala 87:27]
    s2_data_errors_1_6_REG_4_31 <= ^data_full_wayBits_1_6_31; // @[ECC.scala 87:27]
    s2_data_errors_1_7_REG <= s1_valid & tlbRespAllValid & s2_ready; // @[ICacheMainPipe.scala 270:43]
    s2_data_errors_1_7_REG_1 <= s2_data_errors_1_7_REG; // @[ICacheMainPipe.scala 383:40]
    s2_data_errors_1_7_REG_2 <= s1_double_line; // @[ICacheMainPipe.scala 383:77]
    s2_data_errors_1_7_REG_3 <= s2_data_errors_1_7_REG_2; // @[ICacheMainPipe.scala 383:69]
    s2_data_errors_1_7_REG_4_0 <= ^data_full_wayBits_1_7_0; // @[ECC.scala 87:27]
    s2_data_errors_1_7_REG_4_1 <= ^data_full_wayBits_1_7_1; // @[ECC.scala 87:27]
    s2_data_errors_1_7_REG_4_2 <= ^data_full_wayBits_1_7_2; // @[ECC.scala 87:27]
    s2_data_errors_1_7_REG_4_3 <= ^data_full_wayBits_1_7_3; // @[ECC.scala 87:27]
    s2_data_errors_1_7_REG_4_4 <= ^data_full_wayBits_1_7_4; // @[ECC.scala 87:27]
    s2_data_errors_1_7_REG_4_5 <= ^data_full_wayBits_1_7_5; // @[ECC.scala 87:27]
    s2_data_errors_1_7_REG_4_6 <= ^data_full_wayBits_1_7_6; // @[ECC.scala 87:27]
    s2_data_errors_1_7_REG_4_7 <= ^data_full_wayBits_1_7_7; // @[ECC.scala 87:27]
    s2_data_errors_1_7_REG_4_8 <= ^data_full_wayBits_1_7_8; // @[ECC.scala 87:27]
    s2_data_errors_1_7_REG_4_9 <= ^data_full_wayBits_1_7_9; // @[ECC.scala 87:27]
    s2_data_errors_1_7_REG_4_10 <= ^data_full_wayBits_1_7_10; // @[ECC.scala 87:27]
    s2_data_errors_1_7_REG_4_11 <= ^data_full_wayBits_1_7_11; // @[ECC.scala 87:27]
    s2_data_errors_1_7_REG_4_12 <= ^data_full_wayBits_1_7_12; // @[ECC.scala 87:27]
    s2_data_errors_1_7_REG_4_13 <= ^data_full_wayBits_1_7_13; // @[ECC.scala 87:27]
    s2_data_errors_1_7_REG_4_14 <= ^data_full_wayBits_1_7_14; // @[ECC.scala 87:27]
    s2_data_errors_1_7_REG_4_15 <= ^data_full_wayBits_1_7_15; // @[ECC.scala 87:27]
    s2_data_errors_1_7_REG_4_16 <= ^data_full_wayBits_1_7_16; // @[ECC.scala 87:27]
    s2_data_errors_1_7_REG_4_17 <= ^data_full_wayBits_1_7_17; // @[ECC.scala 87:27]
    s2_data_errors_1_7_REG_4_18 <= ^data_full_wayBits_1_7_18; // @[ECC.scala 87:27]
    s2_data_errors_1_7_REG_4_19 <= ^data_full_wayBits_1_7_19; // @[ECC.scala 87:27]
    s2_data_errors_1_7_REG_4_20 <= ^data_full_wayBits_1_7_20; // @[ECC.scala 87:27]
    s2_data_errors_1_7_REG_4_21 <= ^data_full_wayBits_1_7_21; // @[ECC.scala 87:27]
    s2_data_errors_1_7_REG_4_22 <= ^data_full_wayBits_1_7_22; // @[ECC.scala 87:27]
    s2_data_errors_1_7_REG_4_23 <= ^data_full_wayBits_1_7_23; // @[ECC.scala 87:27]
    s2_data_errors_1_7_REG_4_24 <= ^data_full_wayBits_1_7_24; // @[ECC.scala 87:27]
    s2_data_errors_1_7_REG_4_25 <= ^data_full_wayBits_1_7_25; // @[ECC.scala 87:27]
    s2_data_errors_1_7_REG_4_26 <= ^data_full_wayBits_1_7_26; // @[ECC.scala 87:27]
    s2_data_errors_1_7_REG_4_27 <= ^data_full_wayBits_1_7_27; // @[ECC.scala 87:27]
    s2_data_errors_1_7_REG_4_28 <= ^data_full_wayBits_1_7_28; // @[ECC.scala 87:27]
    s2_data_errors_1_7_REG_4_29 <= ^data_full_wayBits_1_7_29; // @[ECC.scala 87:27]
    s2_data_errors_1_7_REG_4_30 <= ^data_full_wayBits_1_7_30; // @[ECC.scala 87:27]
    s2_data_errors_1_7_REG_4_31 <= ^data_full_wayBits_1_7_31; // @[ECC.scala 87:27]
    s2_parity_error_REG <= (s2_meta_errors_0_0 | s2_meta_errors_0_1 | s2_meta_errors_0_2 | s2_meta_errors_0_3 |
      s2_meta_errors_0_4 | s2_meta_errors_0_5 | s2_meta_errors_0_6 | s2_meta_errors_0_7) & io_csr_parity_enable; // @[ICacheMainPipe.scala 388:100]
    s2_parity_error_REG_1 <= (s2_meta_errors_1_0 | s2_meta_errors_1_1 | s2_meta_errors_1_2 | s2_meta_errors_1_3 |
      s2_meta_errors_1_4 | s2_meta_errors_1_5 | s2_meta_errors_1_6 | s2_meta_errors_1_7) & io_csr_parity_enable; // @[ICacheMainPipe.scala 388:100]
    io_errors_0_valid_REG <= s1_valid & tlbRespAllValid & s2_ready; // @[ICacheMainPipe.scala 270:43]
    io_errors_0_valid_REG_1 <= io_errors_0_valid_REG; // @[ICacheMainPipe.scala 393:75]
    io_errors_0_valid_REG_2 <= s2_parity_error_0 & io_errors_0_valid_REG_1; // @[ICacheMainPipe.scala 393:65]
    io_errors_0_report_to_beu_REG <= s1_valid & tlbRespAllValid & s2_ready; // @[ICacheMainPipe.scala 270:43]
    io_errors_0_report_to_beu_REG_1 <= io_errors_0_report_to_beu_REG; // @[ICacheMainPipe.scala 394:75]
    io_errors_0_report_to_beu_REG_2 <= s2_parity_error_0 & io_errors_0_report_to_beu_REG_1; // @[ICacheMainPipe.scala 394:65]
    io_errors_0_paddr_REG <= s2_req_paddr_0; // @[ICacheMainPipe.scala 395:53]
    io_errors_0_paddr_REG_1 <= io_errors_0_paddr_REG; // @[ICacheMainPipe.scala 395:45]
    io_errors_0_source_tag_REG <= (s2_meta_errors_0_0 | s2_meta_errors_0_1 | s2_meta_errors_0_2 | s2_meta_errors_0_3 |
      s2_meta_errors_0_4 | s2_meta_errors_0_5 | s2_meta_errors_0_6 | s2_meta_errors_0_7) & io_csr_parity_enable; // @[ICacheMainPipe.scala 388:100]
    io_errors_0_source_tag_REG_1 <= io_errors_0_source_tag_REG; // @[ICacheMainPipe.scala 397:45]
    io_errors_0_source_data_REG <= (s2_data_errors_0_0 | s2_data_errors_0_1 | s2_data_errors_0_2 | s2_data_errors_0_3 |
      s2_data_errors_0_4 | s2_data_errors_0_5 | s2_data_errors_0_6 | s2_data_errors_0_7) & io_csr_parity_enable; // @[ICacheMainPipe.scala 389:100]
    io_errors_1_valid_REG <= s1_valid & tlbRespAllValid & s2_ready; // @[ICacheMainPipe.scala 270:43]
    io_errors_1_valid_REG_1 <= io_errors_1_valid_REG; // @[ICacheMainPipe.scala 393:75]
    io_errors_1_valid_REG_2 <= s2_parity_error_1 & io_errors_1_valid_REG_1; // @[ICacheMainPipe.scala 393:65]
    io_errors_1_report_to_beu_REG <= s1_valid & tlbRespAllValid & s2_ready; // @[ICacheMainPipe.scala 270:43]
    io_errors_1_report_to_beu_REG_1 <= io_errors_1_report_to_beu_REG; // @[ICacheMainPipe.scala 394:75]
    io_errors_1_report_to_beu_REG_2 <= s2_parity_error_1 & io_errors_1_report_to_beu_REG_1; // @[ICacheMainPipe.scala 394:65]
    io_errors_1_paddr_REG <= s2_req_paddr_1; // @[ICacheMainPipe.scala 395:53]
    io_errors_1_paddr_REG_1 <= io_errors_1_paddr_REG; // @[ICacheMainPipe.scala 395:45]
    io_errors_1_source_tag_REG <= (s2_meta_errors_1_0 | s2_meta_errors_1_1 | s2_meta_errors_1_2 | s2_meta_errors_1_3 |
      s2_meta_errors_1_4 | s2_meta_errors_1_5 | s2_meta_errors_1_6 | s2_meta_errors_1_7) & io_csr_parity_enable; // @[ICacheMainPipe.scala 388:100]
    io_errors_1_source_tag_REG_1 <= io_errors_1_source_tag_REG; // @[ICacheMainPipe.scala 397:45]
    io_errors_1_source_data_REG <= (s2_data_errors_1_0 | s2_data_errors_1_1 | s2_data_errors_1_2 | s2_data_errors_1_3 |
      s2_data_errors_1_4 | s2_data_errors_1_5 | s2_data_errors_1_6 | s2_data_errors_1_7) & io_csr_parity_enable; // @[ICacheMainPipe.scala 389:100]
    s2_except_pmp_af_REG <= s1_valid & tlbRespAllValid & s2_ready; // @[ICacheMainPipe.scala 270:43]
    if (s2_except_pmp_af_REG) begin // @[Reg.scala 17:18]
      s2_except_pmp_af_r0 <= pmpExcpAF_0; // @[Reg.scala 17:22]
    end
    if (s2_except_pmp_af_REG) begin // @[Reg.scala 17:18]
      s2_except_pmp_af_r1 <= pmpExcpAF_1; // @[Reg.scala 17:22]
    end
    s2_mmio_REG <= s1_valid & tlbRespAllValid & s2_ready; // @[ICacheMainPipe.scala 270:43]
    if (s2_mmio_REG) begin // @[Reg.scala 17:18]
      s2_mmio_r <= _s2_mmio_T_5; // @[Reg.scala 17:22]
    end
    only_0_miss_REG <= s1_valid & tlbRespAllValid & s2_ready; // @[ICacheMainPipe.scala 270:43]
    only_0_hit_REG <= s1_valid & tlbRespAllValid & s2_ready; // @[ICacheMainPipe.scala 270:43]
    hit_0_hit_1_REG <= s1_valid & tlbRespAllValid & s2_ready; // @[ICacheMainPipe.scala 270:43]
    hit_0_miss_1_REG <= s1_valid & tlbRespAllValid & s2_ready; // @[ICacheMainPipe.scala 270:43]
    miss_0_hit_1_REG <= s1_valid & tlbRespAllValid & s2_ready; // @[ICacheMainPipe.scala 270:43]
    miss_0_miss_1_REG <= s1_valid & tlbRespAllValid & s2_ready; // @[ICacheMainPipe.scala 270:43]
    miss_0_except_1_REG <= s1_valid & tlbRespAllValid & s2_ready; // @[ICacheMainPipe.scala 270:43]
    if (_reservedRefillData_0_T) begin // @[Reg.scala 17:18]
      reservedRefillData_0_r <= missSlot_0_m_data; // @[Reg.scala 17:22]
    end
    if (_reservedRefillData_1_T) begin // @[Reg.scala 17:18]
      reservedRefillData_1_r <= missSlot_1_m_data; // @[Reg.scala 17:22]
    end
    REG_8 <= _s2_ready_T_2 & missSlot_0_m_corrupt; // @[ICacheMainPipe.scala 710:26]
    io_errors_0_paddr_REG_2 <= s2_req_paddr_0; // @[ICacheMainPipe.scala 713:47]
    REG_9 <= _s2_ready_T_2 & missSlot_1_m_corrupt; // @[ICacheMainPipe.scala 710:26]
    io_errors_1_paddr_REG_2 <= s2_req_paddr_1; // @[ICacheMainPipe.scala 713:47]
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ICacheMainPipe.scala 656:41]
      missSwitchBit <= 1'h0; // @[ICacheMainPipe.scala 657:19]
    end else begin
      missSwitchBit <= io_mshr_0_toMSHR_valid | io_mshr_1_toMSHR_valid | _GEN_426;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ICache.scala 100:42]
      s2_valid <= 1'h0; // @[ICache.scala 100:50]
    end else begin
      s2_valid <= s1_fire | _GEN_235;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ICacheMainPipe.scala 480:35]
      miss_0_s2_0_latch_bit <= 1'h0; // @[ICacheMainPipe.scala 480:41]
    end else begin
      miss_0_s2_0_latch_bit <= miss_0_s2_0 & ~_s2_ready_T_2 | _GEN_361;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ICacheMainPipe.scala 645:66]
      missStateQueue_0 <= 3'h0; // @[ICacheMainPipe.scala 646:29]
    end else if (missStateQueue_0 == 3'h5 & _T_544) begin // @[ICacheMainPipe.scala 649:53]
      missStateQueue_0 <= 3'h1; // @[ICacheMainPipe.scala 650:29]
    end else if (_T_564) begin // @[ICacheMainPipe.scala 634:48]
      missStateQueue_0 <= 3'h0; // @[ICacheMainPipe.scala 636:72 637:31]
    end else if (_miss_0_s2_0_T_6) begin // @[ICacheMainPipe.scala 629:54]
      if (slot_0_solve & _s2_ready_T_2 | ~slot_0_solve & _s2_ready_T_2) begin // @[ICacheMainPipe.scala 630:29]
        missStateQueue_0 <= 3'h0;
      end else begin
        missStateQueue_0 <= _GEN_405;
      end
    end else if (_s2_ready_T_2 & missStateQueue_0 == 3'h2) begin
      missStateQueue_0 <= 3'h4;
    end else begin
      missStateQueue_0 <= _GEN_401;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ICacheMainPipe.scala 480:35]
      miss_1_s2_0_latch_bit <= 1'h0; // @[ICacheMainPipe.scala 480:41]
    end else begin
      miss_1_s2_0_latch_bit <= miss_1_s2_0 & ~_s2_ready_T_2 | _GEN_367;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ICacheMainPipe.scala 645:66]
      missStateQueue_1 <= 3'h0; // @[ICacheMainPipe.scala 646:29]
    end else if (missStateQueue_1 == 3'h5 & _T_568) begin // @[ICacheMainPipe.scala 649:53]
      missStateQueue_1 <= 3'h1; // @[ICacheMainPipe.scala 650:29]
    end else if (_T_588) begin // @[ICacheMainPipe.scala 634:48]
      missStateQueue_1 <= 3'h0; // @[ICacheMainPipe.scala 636:72 637:31]
    end else if (_miss_1_s2_0_T_6) begin // @[ICacheMainPipe.scala 629:54]
      if (slot_1_solve & _s2_ready_T_2 | ~slot_1_solve & _s2_ready_T_2) begin // @[ICacheMainPipe.scala 630:29]
        missStateQueue_1 <= 3'h0;
      end else begin
        missStateQueue_1 <= _GEN_419;
      end
    end else if (_s2_ready_T_2 & missStateQueue_1 == 3'h2) begin
      missStateQueue_1 <= 3'h4;
    end else begin
      missStateQueue_1 <= _GEN_415;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ICacheMainPipe.scala 480:35]
      miss_0_s2_1_latch_bit <= 1'h0; // @[ICacheMainPipe.scala 480:41]
    end else begin
      miss_0_s2_1_latch_bit <= miss_0_s2_1 & ~_s2_ready_T_2 | _GEN_364;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ICacheMainPipe.scala 480:35]
      miss_1_s2_1_latch_bit <= 1'h0; // @[ICacheMainPipe.scala 480:41]
    end else begin
      miss_1_s2_1_latch_bit <= miss_1_s2_1 & ~_s2_ready_T_2 | _GEN_370;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ICacheMainPipe.scala 540:21]
      wait_state <= 4'h0; // @[ICacheMainPipe.scala 542:56 546:20 547:40 548:20 549:60 550:20]
    end else if (4'h0 == wait_state) begin // @[ICacheMainPipe.scala 540:21]
      if (only_pmp_af_0 | only_pmp_af_1 | s2_mmio) begin // @[ICacheMainPipe.scala 559:18]
        wait_state <= 4'h7;
      end else if (miss_0_except_1_latch) begin
        wait_state <= _wait_state_T;
      end else if (only_0_miss_latch | miss_0_hit_1_latch) begin
        wait_state <= _wait_state_T;
      end else begin
        wait_state <= _GEN_376;
      end
    end else if (4'h1 == wait_state) begin // @[ICacheMainPipe.scala 540:21]
      wait_state <= 4'h2; // @[ICacheMainPipe.scala 563:99 564:20]
    end else if (4'h2 == wait_state) begin // @[ICacheMainPipe.scala 540:21]
      if (miss_0_except_1_latch | only_0_miss_latch | hit_0_miss_1_latch | miss_0_hit_1_latch) begin
        wait_state <= 4'h6;
      end else begin
        wait_state <= _GEN_380;
      end
    end else if (4'h6 == wait_state) begin
      wait_state <= _GEN_383;
    end else begin
      wait_state <= _GEN_393;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ICacheMainPipe.scala 480:35]
      hit_0_except_1_latch_bit <= 1'h0; // @[ICacheMainPipe.scala 480:41]
    end else begin
      hit_0_except_1_latch_bit <= hit_0_except_1 & ~_s2_ready_T_2 | _GEN_352;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ICacheMainPipe.scala 480:35]
      except_0_latch_bit <= 1'h0; // @[ICacheMainPipe.scala 480:41]
    end else begin
      except_0_latch_bit <= except_0 & ~_s2_ready_T_2 | _GEN_349;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Hold.scala 42:19]
      tlb_need_back_valid <= 1'h0; // @[Hold.scala 42:27]
    end else begin
      tlb_need_back_valid <= _tlb_need_back_T_1 | _GEN_9;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ICacheMainPipe.scala 251:57]
      tlb_already_recv_0 <= 1'h0; // @[ICacheMainPipe.scala 252:27]
    end else begin
      tlb_already_recv_0 <= tlb_back_0 & tlb_ready_recv_0 & ~s1_fire | _GEN_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ICacheMainPipe.scala 215:33]
      tlb_ready_recv_REG <= 1'h0;
    end else begin
      tlb_ready_recv_REG <= io_fetch_req_valid & s0_can_go;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ICache.scala 100:42]
      s1_valid <= 1'h0; // @[ICache.scala 100:50]
    end else begin
      s1_valid <= s0_fetch_fire | _GEN_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Hold.scala 42:19]
      tlb_need_back_valid_1 <= 1'h0; // @[Hold.scala 42:27]
    end else begin
      tlb_need_back_valid_1 <= _tlb_need_back_T_3 | _GEN_12;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ICacheMainPipe.scala 251:57]
      tlb_already_recv_1 <= 1'h0; // @[ICacheMainPipe.scala 252:27]
    end else begin
      tlb_already_recv_1 <= tlb_back_1 & tlb_ready_recv_1 & ~s1_fire | _GEN_17;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ICacheMainPipe.scala 215:33]
      tlb_ready_recv_REG_1 <= 1'h0;
    end else begin
      tlb_ready_recv_REG_1 <= io_fetch_req_valid & s0_can_go;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec__0 <= 7'h0; // @[Replacement.scala 22:{56,56}]
    end else if (_T_79) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_1_valid) begin
        state_vec__0 <= _state_vec_0_T_46;
      end else if (set_touch_ways_0_valid) begin
        state_vec__0 <= _state_vec_0_T_22;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec__1 <= 7'h0; // @[Replacement.scala 22:{56,56}]
    end else if (_T_80) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_1_1_valid) begin
        state_vec__1 <= _state_vec_1_T_46;
      end else if (set_touch_ways_0_1_valid) begin
        state_vec__1 <= _state_vec_1_T_22;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec__2 <= 7'h0; // @[Replacement.scala 22:{56,56}]
    end else if (_T_81) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_1_2_valid) begin
        state_vec__2 <= _state_vec_2_T_46;
      end else if (set_touch_ways_0_2_valid) begin
        state_vec__2 <= _state_vec_2_T_22;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec__3 <= 7'h0; // @[Replacement.scala 22:{56,56}]
    end else if (_T_82) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_1_3_valid) begin
        state_vec__3 <= _state_vec_3_T_46;
      end else if (set_touch_ways_0_3_valid) begin
        state_vec__3 <= _state_vec_3_T_22;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec__4 <= 7'h0; // @[Replacement.scala 22:{56,56}]
    end else if (_T_83) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_1_4_valid) begin
        state_vec__4 <= _state_vec_4_T_46;
      end else if (set_touch_ways_0_4_valid) begin
        state_vec__4 <= _state_vec_4_T_22;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec__5 <= 7'h0; // @[Replacement.scala 22:{56,56}]
    end else if (_T_84) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_1_5_valid) begin
        state_vec__5 <= _state_vec_5_T_46;
      end else if (set_touch_ways_0_5_valid) begin
        state_vec__5 <= _state_vec_5_T_22;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec__6 <= 7'h0; // @[Replacement.scala 22:{56,56}]
    end else if (_T_85) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_1_6_valid) begin
        state_vec__6 <= _state_vec_6_T_46;
      end else if (set_touch_ways_0_6_valid) begin
        state_vec__6 <= _state_vec_6_T_22;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec__7 <= 7'h0; // @[Replacement.scala 22:{56,56}]
    end else if (_T_86) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_1_7_valid) begin
        state_vec__7 <= _state_vec_7_T_46;
      end else if (set_touch_ways_0_7_valid) begin
        state_vec__7 <= _state_vec_7_T_22;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec__8 <= 7'h0; // @[Replacement.scala 22:{56,56}]
    end else if (_T_87) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_1_8_valid) begin
        state_vec__8 <= _state_vec_8_T_46;
      end else if (set_touch_ways_0_8_valid) begin
        state_vec__8 <= _state_vec_8_T_22;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec__9 <= 7'h0; // @[Replacement.scala 22:{56,56}]
    end else if (_T_88) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_1_9_valid) begin
        state_vec__9 <= _state_vec_9_T_46;
      end else if (set_touch_ways_0_9_valid) begin
        state_vec__9 <= _state_vec_9_T_22;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec__10 <= 7'h0; // @[Replacement.scala 22:{56,56}]
    end else if (_T_89) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_1_10_valid) begin
        state_vec__10 <= _state_vec_10_T_46;
      end else if (set_touch_ways_0_10_valid) begin
        state_vec__10 <= _state_vec_10_T_22;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec__11 <= 7'h0; // @[Replacement.scala 22:{56,56}]
    end else if (_T_90) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_1_11_valid) begin
        state_vec__11 <= _state_vec_11_T_46;
      end else if (set_touch_ways_0_11_valid) begin
        state_vec__11 <= _state_vec_11_T_22;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec__12 <= 7'h0; // @[Replacement.scala 22:{56,56}]
    end else if (_T_91) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_1_12_valid) begin
        state_vec__12 <= _state_vec_12_T_46;
      end else if (set_touch_ways_0_12_valid) begin
        state_vec__12 <= _state_vec_12_T_22;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec__13 <= 7'h0; // @[Replacement.scala 22:{56,56}]
    end else if (_T_92) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_1_13_valid) begin
        state_vec__13 <= _state_vec_13_T_46;
      end else if (set_touch_ways_0_13_valid) begin
        state_vec__13 <= _state_vec_13_T_22;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec__14 <= 7'h0; // @[Replacement.scala 22:{56,56}]
    end else if (_T_93) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_1_14_valid) begin
        state_vec__14 <= _state_vec_14_T_46;
      end else if (set_touch_ways_0_14_valid) begin
        state_vec__14 <= _state_vec_14_T_22;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec__15 <= 7'h0; // @[Replacement.scala 22:{56,56}]
    end else if (_T_94) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_1_15_valid) begin
        state_vec__15 <= _state_vec_15_T_46;
      end else if (set_touch_ways_0_15_valid) begin
        state_vec__15 <= _state_vec_15_T_22;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec__16 <= 7'h0; // @[Replacement.scala 22:{56,56}]
    end else if (_T_95) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_1_16_valid) begin
        state_vec__16 <= _state_vec_16_T_46;
      end else if (set_touch_ways_0_16_valid) begin
        state_vec__16 <= _state_vec_16_T_22;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec__17 <= 7'h0; // @[Replacement.scala 22:{56,56}]
    end else if (_T_96) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_1_17_valid) begin
        state_vec__17 <= _state_vec_17_T_46;
      end else if (set_touch_ways_0_17_valid) begin
        state_vec__17 <= _state_vec_17_T_22;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec__18 <= 7'h0; // @[Replacement.scala 22:{56,56}]
    end else if (_T_97) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_1_18_valid) begin
        state_vec__18 <= _state_vec_18_T_46;
      end else if (set_touch_ways_0_18_valid) begin
        state_vec__18 <= _state_vec_18_T_22;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec__19 <= 7'h0; // @[Replacement.scala 22:{56,56}]
    end else if (_T_98) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_1_19_valid) begin
        state_vec__19 <= _state_vec_19_T_46;
      end else if (set_touch_ways_0_19_valid) begin
        state_vec__19 <= _state_vec_19_T_22;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec__20 <= 7'h0; // @[Replacement.scala 22:{56,56}]
    end else if (_T_99) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_1_20_valid) begin
        state_vec__20 <= _state_vec_20_T_46;
      end else if (set_touch_ways_0_20_valid) begin
        state_vec__20 <= _state_vec_20_T_22;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec__21 <= 7'h0; // @[Replacement.scala 22:{56,56}]
    end else if (_T_100) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_1_21_valid) begin
        state_vec__21 <= _state_vec_21_T_46;
      end else if (set_touch_ways_0_21_valid) begin
        state_vec__21 <= _state_vec_21_T_22;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec__22 <= 7'h0; // @[Replacement.scala 22:{56,56}]
    end else if (_T_101) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_1_22_valid) begin
        state_vec__22 <= _state_vec_22_T_46;
      end else if (set_touch_ways_0_22_valid) begin
        state_vec__22 <= _state_vec_22_T_22;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec__23 <= 7'h0; // @[Replacement.scala 22:{56,56}]
    end else if (_T_102) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_1_23_valid) begin
        state_vec__23 <= _state_vec_23_T_46;
      end else if (set_touch_ways_0_23_valid) begin
        state_vec__23 <= _state_vec_23_T_22;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec__24 <= 7'h0; // @[Replacement.scala 22:{56,56}]
    end else if (_T_103) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_1_24_valid) begin
        state_vec__24 <= _state_vec_24_T_46;
      end else if (set_touch_ways_0_24_valid) begin
        state_vec__24 <= _state_vec_24_T_22;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec__25 <= 7'h0; // @[Replacement.scala 22:{56,56}]
    end else if (_T_104) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_1_25_valid) begin
        state_vec__25 <= _state_vec_25_T_46;
      end else if (set_touch_ways_0_25_valid) begin
        state_vec__25 <= _state_vec_25_T_22;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec__26 <= 7'h0; // @[Replacement.scala 22:{56,56}]
    end else if (_T_105) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_1_26_valid) begin
        state_vec__26 <= _state_vec_26_T_46;
      end else if (set_touch_ways_0_26_valid) begin
        state_vec__26 <= _state_vec_26_T_22;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec__27 <= 7'h0; // @[Replacement.scala 22:{56,56}]
    end else if (_T_106) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_1_27_valid) begin
        state_vec__27 <= _state_vec_27_T_46;
      end else if (set_touch_ways_0_27_valid) begin
        state_vec__27 <= _state_vec_27_T_22;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec__28 <= 7'h0; // @[Replacement.scala 22:{56,56}]
    end else if (_T_107) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_1_28_valid) begin
        state_vec__28 <= _state_vec_28_T_46;
      end else if (set_touch_ways_0_28_valid) begin
        state_vec__28 <= _state_vec_28_T_22;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec__29 <= 7'h0; // @[Replacement.scala 22:{56,56}]
    end else if (_T_108) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_1_29_valid) begin
        state_vec__29 <= _state_vec_29_T_46;
      end else if (set_touch_ways_0_29_valid) begin
        state_vec__29 <= _state_vec_29_T_22;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec__30 <= 7'h0; // @[Replacement.scala 22:{56,56}]
    end else if (_T_109) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_1_30_valid) begin
        state_vec__30 <= _state_vec_30_T_46;
      end else if (set_touch_ways_0_30_valid) begin
        state_vec__30 <= _state_vec_30_T_22;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec__31 <= 7'h0; // @[Replacement.scala 22:{56,56}]
    end else if (_T_110) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_1_31_valid) begin
        state_vec__31 <= _state_vec_31_T_46;
      end else if (set_touch_ways_0_31_valid) begin
        state_vec__31 <= _state_vec_31_T_22;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_1_0 <= 7'h0; // @[Replacement.scala 22:{56,56}]
    end else if (_T_111) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_1_32_valid) begin
        state_vec_1_0 <= _state_vec_0_T_94;
      end else if (set_touch_ways_0_32_valid) begin
        state_vec_1_0 <= _state_vec_0_T_70;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_1_1 <= 7'h0; // @[Replacement.scala 22:{56,56}]
    end else if (_T_112) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_1_33_valid) begin
        state_vec_1_1 <= _state_vec_1_T_94;
      end else if (set_touch_ways_0_33_valid) begin
        state_vec_1_1 <= _state_vec_1_T_70;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_1_2 <= 7'h0; // @[Replacement.scala 22:{56,56}]
    end else if (_T_113) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_1_34_valid) begin
        state_vec_1_2 <= _state_vec_2_T_94;
      end else if (set_touch_ways_0_34_valid) begin
        state_vec_1_2 <= _state_vec_2_T_70;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_1_3 <= 7'h0; // @[Replacement.scala 22:{56,56}]
    end else if (_T_114) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_1_35_valid) begin
        state_vec_1_3 <= _state_vec_3_T_94;
      end else if (set_touch_ways_0_35_valid) begin
        state_vec_1_3 <= _state_vec_3_T_70;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_1_4 <= 7'h0; // @[Replacement.scala 22:{56,56}]
    end else if (_T_115) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_1_36_valid) begin
        state_vec_1_4 <= _state_vec_4_T_94;
      end else if (set_touch_ways_0_36_valid) begin
        state_vec_1_4 <= _state_vec_4_T_70;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_1_5 <= 7'h0; // @[Replacement.scala 22:{56,56}]
    end else if (_T_116) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_1_37_valid) begin
        state_vec_1_5 <= _state_vec_5_T_94;
      end else if (set_touch_ways_0_37_valid) begin
        state_vec_1_5 <= _state_vec_5_T_70;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_1_6 <= 7'h0; // @[Replacement.scala 22:{56,56}]
    end else if (_T_117) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_1_38_valid) begin
        state_vec_1_6 <= _state_vec_6_T_94;
      end else if (set_touch_ways_0_38_valid) begin
        state_vec_1_6 <= _state_vec_6_T_70;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_1_7 <= 7'h0; // @[Replacement.scala 22:{56,56}]
    end else if (_T_118) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_1_39_valid) begin
        state_vec_1_7 <= _state_vec_7_T_94;
      end else if (set_touch_ways_0_39_valid) begin
        state_vec_1_7 <= _state_vec_7_T_70;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_1_8 <= 7'h0; // @[Replacement.scala 22:{56,56}]
    end else if (_T_119) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_1_40_valid) begin
        state_vec_1_8 <= _state_vec_8_T_94;
      end else if (set_touch_ways_0_40_valid) begin
        state_vec_1_8 <= _state_vec_8_T_70;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_1_9 <= 7'h0; // @[Replacement.scala 22:{56,56}]
    end else if (_T_120) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_1_41_valid) begin
        state_vec_1_9 <= _state_vec_9_T_94;
      end else if (set_touch_ways_0_41_valid) begin
        state_vec_1_9 <= _state_vec_9_T_70;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_1_10 <= 7'h0; // @[Replacement.scala 22:{56,56}]
    end else if (_T_121) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_1_42_valid) begin
        state_vec_1_10 <= _state_vec_10_T_94;
      end else if (set_touch_ways_0_42_valid) begin
        state_vec_1_10 <= _state_vec_10_T_70;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_1_11 <= 7'h0; // @[Replacement.scala 22:{56,56}]
    end else if (_T_122) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_1_43_valid) begin
        state_vec_1_11 <= _state_vec_11_T_94;
      end else if (set_touch_ways_0_43_valid) begin
        state_vec_1_11 <= _state_vec_11_T_70;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_1_12 <= 7'h0; // @[Replacement.scala 22:{56,56}]
    end else if (_T_123) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_1_44_valid) begin
        state_vec_1_12 <= _state_vec_12_T_94;
      end else if (set_touch_ways_0_44_valid) begin
        state_vec_1_12 <= _state_vec_12_T_70;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_1_13 <= 7'h0; // @[Replacement.scala 22:{56,56}]
    end else if (_T_124) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_1_45_valid) begin
        state_vec_1_13 <= _state_vec_13_T_94;
      end else if (set_touch_ways_0_45_valid) begin
        state_vec_1_13 <= _state_vec_13_T_70;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_1_14 <= 7'h0; // @[Replacement.scala 22:{56,56}]
    end else if (_T_125) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_1_46_valid) begin
        state_vec_1_14 <= _state_vec_14_T_94;
      end else if (set_touch_ways_0_46_valid) begin
        state_vec_1_14 <= _state_vec_14_T_70;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_1_15 <= 7'h0; // @[Replacement.scala 22:{56,56}]
    end else if (_T_126) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_1_47_valid) begin
        state_vec_1_15 <= _state_vec_15_T_94;
      end else if (set_touch_ways_0_47_valid) begin
        state_vec_1_15 <= _state_vec_15_T_70;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_1_16 <= 7'h0; // @[Replacement.scala 22:{56,56}]
    end else if (_T_127) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_1_48_valid) begin
        state_vec_1_16 <= _state_vec_16_T_94;
      end else if (set_touch_ways_0_48_valid) begin
        state_vec_1_16 <= _state_vec_16_T_70;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_1_17 <= 7'h0; // @[Replacement.scala 22:{56,56}]
    end else if (_T_128) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_1_49_valid) begin
        state_vec_1_17 <= _state_vec_17_T_94;
      end else if (set_touch_ways_0_49_valid) begin
        state_vec_1_17 <= _state_vec_17_T_70;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_1_18 <= 7'h0; // @[Replacement.scala 22:{56,56}]
    end else if (_T_129) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_1_50_valid) begin
        state_vec_1_18 <= _state_vec_18_T_94;
      end else if (set_touch_ways_0_50_valid) begin
        state_vec_1_18 <= _state_vec_18_T_70;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_1_19 <= 7'h0; // @[Replacement.scala 22:{56,56}]
    end else if (_T_130) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_1_51_valid) begin
        state_vec_1_19 <= _state_vec_19_T_94;
      end else if (set_touch_ways_0_51_valid) begin
        state_vec_1_19 <= _state_vec_19_T_70;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_1_20 <= 7'h0; // @[Replacement.scala 22:{56,56}]
    end else if (_T_131) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_1_52_valid) begin
        state_vec_1_20 <= _state_vec_20_T_94;
      end else if (set_touch_ways_0_52_valid) begin
        state_vec_1_20 <= _state_vec_20_T_70;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_1_21 <= 7'h0; // @[Replacement.scala 22:{56,56}]
    end else if (_T_132) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_1_53_valid) begin
        state_vec_1_21 <= _state_vec_21_T_94;
      end else if (set_touch_ways_0_53_valid) begin
        state_vec_1_21 <= _state_vec_21_T_70;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_1_22 <= 7'h0; // @[Replacement.scala 22:{56,56}]
    end else if (_T_133) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_1_54_valid) begin
        state_vec_1_22 <= _state_vec_22_T_94;
      end else if (set_touch_ways_0_54_valid) begin
        state_vec_1_22 <= _state_vec_22_T_70;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_1_23 <= 7'h0; // @[Replacement.scala 22:{56,56}]
    end else if (_T_134) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_1_55_valid) begin
        state_vec_1_23 <= _state_vec_23_T_94;
      end else if (set_touch_ways_0_55_valid) begin
        state_vec_1_23 <= _state_vec_23_T_70;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_1_24 <= 7'h0; // @[Replacement.scala 22:{56,56}]
    end else if (_T_135) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_1_56_valid) begin
        state_vec_1_24 <= _state_vec_24_T_94;
      end else if (set_touch_ways_0_56_valid) begin
        state_vec_1_24 <= _state_vec_24_T_70;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_1_25 <= 7'h0; // @[Replacement.scala 22:{56,56}]
    end else if (_T_136) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_1_57_valid) begin
        state_vec_1_25 <= _state_vec_25_T_94;
      end else if (set_touch_ways_0_57_valid) begin
        state_vec_1_25 <= _state_vec_25_T_70;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_1_26 <= 7'h0; // @[Replacement.scala 22:{56,56}]
    end else if (_T_137) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_1_58_valid) begin
        state_vec_1_26 <= _state_vec_26_T_94;
      end else if (set_touch_ways_0_58_valid) begin
        state_vec_1_26 <= _state_vec_26_T_70;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_1_27 <= 7'h0; // @[Replacement.scala 22:{56,56}]
    end else if (_T_138) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_1_59_valid) begin
        state_vec_1_27 <= _state_vec_27_T_94;
      end else if (set_touch_ways_0_59_valid) begin
        state_vec_1_27 <= _state_vec_27_T_70;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_1_28 <= 7'h0; // @[Replacement.scala 22:{56,56}]
    end else if (_T_139) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_1_60_valid) begin
        state_vec_1_28 <= _state_vec_28_T_94;
      end else if (set_touch_ways_0_60_valid) begin
        state_vec_1_28 <= _state_vec_28_T_70;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_1_29 <= 7'h0; // @[Replacement.scala 22:{56,56}]
    end else if (_T_140) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_1_61_valid) begin
        state_vec_1_29 <= _state_vec_29_T_94;
      end else if (set_touch_ways_0_61_valid) begin
        state_vec_1_29 <= _state_vec_29_T_70;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_1_30 <= 7'h0; // @[Replacement.scala 22:{56,56}]
    end else if (_T_141) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_1_62_valid) begin
        state_vec_1_30 <= _state_vec_30_T_94;
      end else if (set_touch_ways_0_62_valid) begin
        state_vec_1_30 <= _state_vec_30_T_70;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_1_31 <= 7'h0; // @[Replacement.scala 22:{56,56}]
    end else if (_T_142) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_1_63_valid) begin
        state_vec_1_31 <= _state_vec_31_T_94;
      end else if (set_touch_ways_0_63_valid) begin
        state_vec_1_31 <= _state_vec_31_T_70;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Hold.scala 42:19]
      s2_tlb_need_back_valid <= 1'h0; // @[Hold.scala 42:27]
    end else begin
      s2_tlb_need_back_valid <= _s2_tlb_need_back_T | _GEN_321;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Hold.scala 42:19]
      s2_tlb_need_back_valid_1 <= 1'h0; // @[Hold.scala 42:27]
    end else begin
      s2_tlb_need_back_valid_1 <= _s2_tlb_need_back_T_1 | _GEN_324;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ICacheMainPipe.scala 645:66]
      missSlot_0_m_vSetIdx <= 6'h0; // @[ICacheMainPipe.scala 647:29]
    end else if (missStateQueue_0 == 3'h5 & _T_544) begin // @[ICacheMainPipe.scala 616:62]
      missSlot_0_m_vSetIdx <= s2_req_vsetIdx_0; // @[ICacheMainPipe.scala 618:29]
    end else if (_T_544 & _s2_miss_available_T) begin // @[ICacheMainPipe.scala 447:40]
      missSlot_0_m_vSetIdx <= s2_req_vsetIdx_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ICacheMainPipe.scala 645:66]
      missSlot_0_m_pTag <= 24'h0; // @[ICacheMainPipe.scala 648:29]
    end else if (missStateQueue_0 == 3'h5 & _T_544) begin // @[ICacheMainPipe.scala 616:62]
      missSlot_0_m_pTag <= s2_req_paddr_0[35:12]; // @[ICacheMainPipe.scala 619:29]
    end else if (_T_544 & _s2_miss_available_T) begin // @[ICacheMainPipe.scala 447:40]
      missSlot_0_m_pTag <= s2_req_paddr_0[35:12];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ICacheMainPipe.scala 622:63]
      missSlot_0_m_data <= 512'h0; // @[ICacheMainPipe.scala 624:33]
    end else if (io_mshr_0_fromMSHR_valid & missStateQueue_0 == 3'h1) begin // @[ICacheMainPipe.scala 447:40]
      missSlot_0_m_data <= io_mshr_0_fromMSHR_bits_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ICacheMainPipe.scala 622:63]
      missSlot_0_m_corrupt <= 1'h0; // @[ICacheMainPipe.scala 625:33]
    end else if (io_mshr_0_fromMSHR_valid & missStateQueue_0 == 3'h1) begin // @[ICacheMainPipe.scala 447:40]
      missSlot_0_m_corrupt <= io_mshr_0_fromMSHR_bits_corrupt;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ICacheMainPipe.scala 645:66]
      missSlot_1_m_vSetIdx <= 6'h0; // @[ICacheMainPipe.scala 647:29]
    end else if (missStateQueue_1 == 3'h5 & _T_568) begin // @[ICacheMainPipe.scala 616:62]
      missSlot_1_m_vSetIdx <= s2_req_vsetIdx_1; // @[ICacheMainPipe.scala 618:29]
    end else if (_T_568 & _s2_miss_available_T_3) begin // @[ICacheMainPipe.scala 447:40]
      missSlot_1_m_vSetIdx <= s2_req_vsetIdx_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ICacheMainPipe.scala 645:66]
      missSlot_1_m_pTag <= 24'h0; // @[ICacheMainPipe.scala 648:29]
    end else if (missStateQueue_1 == 3'h5 & _T_568) begin // @[ICacheMainPipe.scala 616:62]
      missSlot_1_m_pTag <= s2_req_paddr_1[35:12]; // @[ICacheMainPipe.scala 619:29]
    end else if (_T_568 & _s2_miss_available_T_3) begin // @[ICacheMainPipe.scala 447:40]
      missSlot_1_m_pTag <= s2_req_paddr_1[35:12];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ICacheMainPipe.scala 622:63]
      missSlot_1_m_data <= 512'h0; // @[ICacheMainPipe.scala 624:33]
    end else if (io_mshr_1_fromMSHR_valid & missStateQueue_1 == 3'h1) begin // @[ICacheMainPipe.scala 447:40]
      missSlot_1_m_data <= io_mshr_1_fromMSHR_bits_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ICacheMainPipe.scala 622:63]
      missSlot_1_m_corrupt <= 1'h0; // @[ICacheMainPipe.scala 625:33]
    end else if (io_mshr_1_fromMSHR_valid & missStateQueue_1 == 3'h1) begin // @[ICacheMainPipe.scala 447:40]
      missSlot_1_m_corrupt <= io_mshr_1_fromMSHR_bits_corrupt;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ICacheMainPipe.scala 480:35]
      miss_0_hit_1_latch_bit <= 1'h0; // @[ICacheMainPipe.scala 480:41]
    end else begin
      miss_0_hit_1_latch_bit <= miss_0_hit_1 & ~_s2_ready_T_2 | _GEN_334;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ICacheMainPipe.scala 480:35]
      miss_0_miss_1_latch_bit <= 1'h0; // @[ICacheMainPipe.scala 480:41]
    end else begin
      miss_0_miss_1_latch_bit <= miss_0_miss_1 & ~_s2_ready_T_2 | _GEN_337;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ICacheMainPipe.scala 480:35]
      only_0_miss_latch_bit <= 1'h0; // @[ICacheMainPipe.scala 480:41]
    end else begin
      only_0_miss_latch_bit <= only_0_miss & ~_s2_ready_T_2 | _GEN_340;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ICacheMainPipe.scala 480:35]
      hit_0_miss_1_latch_bit <= 1'h0; // @[ICacheMainPipe.scala 480:41]
    end else begin
      hit_0_miss_1_latch_bit <= hit_0_miss_1 & ~_s2_ready_T_2 | _GEN_343;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ICacheMainPipe.scala 480:35]
      miss_0_except_1_latch_bit <= 1'h0; // @[ICacheMainPipe.scala 480:41]
    end else begin
      miss_0_except_1_latch_bit <= miss_0_except_1 & ~_s2_ready_T_2 | _GEN_346;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ICacheMainPipe.scala 480:35]
      only_0_hit_latch_bit <= 1'h0; // @[ICacheMainPipe.scala 480:41]
    end else begin
      only_0_hit_latch_bit <= only_0_hit & ~_s2_ready_T_2 | _GEN_355;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ICacheMainPipe.scala 480:35]
      hit_0_hit_1_latch_bit <= 1'h0; // @[ICacheMainPipe.scala 480:41]
    end else begin
      hit_0_hit_1_latch_bit <= hit_0_hit_1 & ~_s2_ready_T_2 | _GEN_358;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  missSwitchBit = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  s2_valid = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  s2_port_hit_0 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  miss_0_s2_0_latch_bit = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  miss_0_s2_0_REG = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  miss_0_s2_0_REG_1 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  miss_0_s2_0_REG_2 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  missStateQueue_0 = _RAND_7[2:0];
  _RAND_8 = {1{`RANDOM}};
  miss_1_s2_0_latch_bit = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  miss_1_s2_0_REG = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  miss_1_s2_0_REG_1 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  miss_1_s2_0_REG_2 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  missStateQueue_1 = _RAND_12[2:0];
  _RAND_13 = {1{`RANDOM}};
  s2_port_hit_1 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  miss_0_s2_1_latch_bit = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  miss_0_s2_1_REG = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  miss_0_s2_1_REG_1 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  miss_0_s2_1_REG_2 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  miss_1_s2_1_latch_bit = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  miss_1_s2_1_REG = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  miss_1_s2_1_REG_1 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  miss_1_s2_1_REG_2 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  s2_double_line = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  wait_state = _RAND_23[3:0];
  _RAND_24 = {1{`RANDOM}};
  hit_0_except_1_latch_bit = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  hit_0_except_1_REG = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  s2_except_pf_0 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  s2_except_tlb_af_0 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  s2_except_pf_1 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  s2_except_tlb_af_1 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  except_0_latch_bit = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  except_0_REG = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  tlb_need_back_valid = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  tlb_already_recv_0 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  tlb_ready_recv_REG = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  s1_valid = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  tlb_need_back_valid_1 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  tlb_already_recv_1 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  tlb_ready_recv_REG_1 = _RAND_38[0:0];
  _RAND_39 = {2{`RANDOM}};
  s1_req_vaddr_0 = _RAND_39[38:0];
  _RAND_40 = {2{`RANDOM}};
  s1_req_vaddr_1 = _RAND_40[38:0];
  _RAND_41 = {1{`RANDOM}};
  s1_req_vsetIdx_0 = _RAND_41[5:0];
  _RAND_42 = {1{`RANDOM}};
  s1_req_vsetIdx_1 = _RAND_42[5:0];
  _RAND_43 = {1{`RANDOM}};
  s1_double_line = _RAND_43[0:0];
  _RAND_44 = {2{`RANDOM}};
  tlbRespPAddr_r = _RAND_44[35:0];
  _RAND_45 = {2{`RANDOM}};
  tlbRespPAddr_r1 = _RAND_45[35:0];
  _RAND_46 = {1{`RANDOM}};
  tlbExcpPF_r = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  tlbExcpPF_r1 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  tlbExcpAF_r = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  tlbExcpAF_r1 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  s1_meta_ptags_REG = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  s1_meta_ptags_r0_0 = _RAND_51[23:0];
  _RAND_52 = {1{`RANDOM}};
  s1_meta_ptags_r0_1 = _RAND_52[23:0];
  _RAND_53 = {1{`RANDOM}};
  s1_meta_ptags_r0_2 = _RAND_53[23:0];
  _RAND_54 = {1{`RANDOM}};
  s1_meta_ptags_r0_3 = _RAND_54[23:0];
  _RAND_55 = {1{`RANDOM}};
  s1_meta_ptags_r0_4 = _RAND_55[23:0];
  _RAND_56 = {1{`RANDOM}};
  s1_meta_ptags_r0_5 = _RAND_56[23:0];
  _RAND_57 = {1{`RANDOM}};
  s1_meta_ptags_r0_6 = _RAND_57[23:0];
  _RAND_58 = {1{`RANDOM}};
  s1_meta_ptags_r0_7 = _RAND_58[23:0];
  _RAND_59 = {1{`RANDOM}};
  s1_meta_ptags_r1_0 = _RAND_59[23:0];
  _RAND_60 = {1{`RANDOM}};
  s1_meta_ptags_r1_1 = _RAND_60[23:0];
  _RAND_61 = {1{`RANDOM}};
  s1_meta_ptags_r1_2 = _RAND_61[23:0];
  _RAND_62 = {1{`RANDOM}};
  s1_meta_ptags_r1_3 = _RAND_62[23:0];
  _RAND_63 = {1{`RANDOM}};
  s1_meta_ptags_r1_4 = _RAND_63[23:0];
  _RAND_64 = {1{`RANDOM}};
  s1_meta_ptags_r1_5 = _RAND_64[23:0];
  _RAND_65 = {1{`RANDOM}};
  s1_meta_ptags_r1_6 = _RAND_65[23:0];
  _RAND_66 = {1{`RANDOM}};
  s1_meta_ptags_r1_7 = _RAND_66[23:0];
  _RAND_67 = {1{`RANDOM}};
  s1_meta_cohs_REG = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  s1_meta_cohs_r0_0_state = _RAND_68[1:0];
  _RAND_69 = {1{`RANDOM}};
  s1_meta_cohs_r0_1_state = _RAND_69[1:0];
  _RAND_70 = {1{`RANDOM}};
  s1_meta_cohs_r0_2_state = _RAND_70[1:0];
  _RAND_71 = {1{`RANDOM}};
  s1_meta_cohs_r0_3_state = _RAND_71[1:0];
  _RAND_72 = {1{`RANDOM}};
  s1_meta_cohs_r0_4_state = _RAND_72[1:0];
  _RAND_73 = {1{`RANDOM}};
  s1_meta_cohs_r0_5_state = _RAND_73[1:0];
  _RAND_74 = {1{`RANDOM}};
  s1_meta_cohs_r0_6_state = _RAND_74[1:0];
  _RAND_75 = {1{`RANDOM}};
  s1_meta_cohs_r0_7_state = _RAND_75[1:0];
  _RAND_76 = {1{`RANDOM}};
  s1_meta_cohs_r1_0_state = _RAND_76[1:0];
  _RAND_77 = {1{`RANDOM}};
  s1_meta_cohs_r1_1_state = _RAND_77[1:0];
  _RAND_78 = {1{`RANDOM}};
  s1_meta_cohs_r1_2_state = _RAND_78[1:0];
  _RAND_79 = {1{`RANDOM}};
  s1_meta_cohs_r1_3_state = _RAND_79[1:0];
  _RAND_80 = {1{`RANDOM}};
  s1_meta_cohs_r1_4_state = _RAND_80[1:0];
  _RAND_81 = {1{`RANDOM}};
  s1_meta_cohs_r1_5_state = _RAND_81[1:0];
  _RAND_82 = {1{`RANDOM}};
  s1_meta_cohs_r1_6_state = _RAND_82[1:0];
  _RAND_83 = {1{`RANDOM}};
  s1_meta_cohs_r1_7_state = _RAND_83[1:0];
  _RAND_84 = {1{`RANDOM}};
  s1_meta_errors_REG = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  s1_meta_errors_r0_0 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  s1_meta_errors_r0_1 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  s1_meta_errors_r0_2 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  s1_meta_errors_r0_3 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  s1_meta_errors_r0_4 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  s1_meta_errors_r0_5 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  s1_meta_errors_r0_6 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  s1_meta_errors_r0_7 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  s1_meta_errors_r1_0 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  s1_meta_errors_r1_1 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  s1_meta_errors_r1_2 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  s1_meta_errors_r1_3 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  s1_meta_errors_r1_4 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  s1_meta_errors_r1_5 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  s1_meta_errors_r1_6 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  s1_meta_errors_r1_7 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  s1_data_cacheline_REG = _RAND_101[0:0];
  _RAND_102 = {16{`RANDOM}};
  s1_data_cacheline_r0_0 = _RAND_102[511:0];
  _RAND_103 = {16{`RANDOM}};
  s1_data_cacheline_r0_1 = _RAND_103[511:0];
  _RAND_104 = {16{`RANDOM}};
  s1_data_cacheline_r0_2 = _RAND_104[511:0];
  _RAND_105 = {16{`RANDOM}};
  s1_data_cacheline_r0_3 = _RAND_105[511:0];
  _RAND_106 = {16{`RANDOM}};
  s1_data_cacheline_r0_4 = _RAND_106[511:0];
  _RAND_107 = {16{`RANDOM}};
  s1_data_cacheline_r0_5 = _RAND_107[511:0];
  _RAND_108 = {16{`RANDOM}};
  s1_data_cacheline_r0_6 = _RAND_108[511:0];
  _RAND_109 = {16{`RANDOM}};
  s1_data_cacheline_r0_7 = _RAND_109[511:0];
  _RAND_110 = {16{`RANDOM}};
  s1_data_cacheline_r1_0 = _RAND_110[511:0];
  _RAND_111 = {16{`RANDOM}};
  s1_data_cacheline_r1_1 = _RAND_111[511:0];
  _RAND_112 = {16{`RANDOM}};
  s1_data_cacheline_r1_2 = _RAND_112[511:0];
  _RAND_113 = {16{`RANDOM}};
  s1_data_cacheline_r1_3 = _RAND_113[511:0];
  _RAND_114 = {16{`RANDOM}};
  s1_data_cacheline_r1_4 = _RAND_114[511:0];
  _RAND_115 = {16{`RANDOM}};
  s1_data_cacheline_r1_5 = _RAND_115[511:0];
  _RAND_116 = {16{`RANDOM}};
  s1_data_cacheline_r1_6 = _RAND_116[511:0];
  _RAND_117 = {16{`RANDOM}};
  s1_data_cacheline_r1_7 = _RAND_117[511:0];
  _RAND_118 = {1{`RANDOM}};
  s1_data_errorBits_REG = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  s1_data_errorBits_r0_0 = _RAND_119[31:0];
  _RAND_120 = {1{`RANDOM}};
  s1_data_errorBits_r0_1 = _RAND_120[31:0];
  _RAND_121 = {1{`RANDOM}};
  s1_data_errorBits_r0_2 = _RAND_121[31:0];
  _RAND_122 = {1{`RANDOM}};
  s1_data_errorBits_r0_3 = _RAND_122[31:0];
  _RAND_123 = {1{`RANDOM}};
  s1_data_errorBits_r0_4 = _RAND_123[31:0];
  _RAND_124 = {1{`RANDOM}};
  s1_data_errorBits_r0_5 = _RAND_124[31:0];
  _RAND_125 = {1{`RANDOM}};
  s1_data_errorBits_r0_6 = _RAND_125[31:0];
  _RAND_126 = {1{`RANDOM}};
  s1_data_errorBits_r0_7 = _RAND_126[31:0];
  _RAND_127 = {1{`RANDOM}};
  s1_data_errorBits_r1_0 = _RAND_127[31:0];
  _RAND_128 = {1{`RANDOM}};
  s1_data_errorBits_r1_1 = _RAND_128[31:0];
  _RAND_129 = {1{`RANDOM}};
  s1_data_errorBits_r1_2 = _RAND_129[31:0];
  _RAND_130 = {1{`RANDOM}};
  s1_data_errorBits_r1_3 = _RAND_130[31:0];
  _RAND_131 = {1{`RANDOM}};
  s1_data_errorBits_r1_4 = _RAND_131[31:0];
  _RAND_132 = {1{`RANDOM}};
  s1_data_errorBits_r1_5 = _RAND_132[31:0];
  _RAND_133 = {1{`RANDOM}};
  s1_data_errorBits_r1_6 = _RAND_133[31:0];
  _RAND_134 = {1{`RANDOM}};
  s1_data_errorBits_r1_7 = _RAND_134[31:0];
  _RAND_135 = {1{`RANDOM}};
  state_vec__0 = _RAND_135[6:0];
  _RAND_136 = {1{`RANDOM}};
  state_vec__1 = _RAND_136[6:0];
  _RAND_137 = {1{`RANDOM}};
  state_vec__2 = _RAND_137[6:0];
  _RAND_138 = {1{`RANDOM}};
  state_vec__3 = _RAND_138[6:0];
  _RAND_139 = {1{`RANDOM}};
  state_vec__4 = _RAND_139[6:0];
  _RAND_140 = {1{`RANDOM}};
  state_vec__5 = _RAND_140[6:0];
  _RAND_141 = {1{`RANDOM}};
  state_vec__6 = _RAND_141[6:0];
  _RAND_142 = {1{`RANDOM}};
  state_vec__7 = _RAND_142[6:0];
  _RAND_143 = {1{`RANDOM}};
  state_vec__8 = _RAND_143[6:0];
  _RAND_144 = {1{`RANDOM}};
  state_vec__9 = _RAND_144[6:0];
  _RAND_145 = {1{`RANDOM}};
  state_vec__10 = _RAND_145[6:0];
  _RAND_146 = {1{`RANDOM}};
  state_vec__11 = _RAND_146[6:0];
  _RAND_147 = {1{`RANDOM}};
  state_vec__12 = _RAND_147[6:0];
  _RAND_148 = {1{`RANDOM}};
  state_vec__13 = _RAND_148[6:0];
  _RAND_149 = {1{`RANDOM}};
  state_vec__14 = _RAND_149[6:0];
  _RAND_150 = {1{`RANDOM}};
  state_vec__15 = _RAND_150[6:0];
  _RAND_151 = {1{`RANDOM}};
  state_vec__16 = _RAND_151[6:0];
  _RAND_152 = {1{`RANDOM}};
  state_vec__17 = _RAND_152[6:0];
  _RAND_153 = {1{`RANDOM}};
  state_vec__18 = _RAND_153[6:0];
  _RAND_154 = {1{`RANDOM}};
  state_vec__19 = _RAND_154[6:0];
  _RAND_155 = {1{`RANDOM}};
  state_vec__20 = _RAND_155[6:0];
  _RAND_156 = {1{`RANDOM}};
  state_vec__21 = _RAND_156[6:0];
  _RAND_157 = {1{`RANDOM}};
  state_vec__22 = _RAND_157[6:0];
  _RAND_158 = {1{`RANDOM}};
  state_vec__23 = _RAND_158[6:0];
  _RAND_159 = {1{`RANDOM}};
  state_vec__24 = _RAND_159[6:0];
  _RAND_160 = {1{`RANDOM}};
  state_vec__25 = _RAND_160[6:0];
  _RAND_161 = {1{`RANDOM}};
  state_vec__26 = _RAND_161[6:0];
  _RAND_162 = {1{`RANDOM}};
  state_vec__27 = _RAND_162[6:0];
  _RAND_163 = {1{`RANDOM}};
  state_vec__28 = _RAND_163[6:0];
  _RAND_164 = {1{`RANDOM}};
  state_vec__29 = _RAND_164[6:0];
  _RAND_165 = {1{`RANDOM}};
  state_vec__30 = _RAND_165[6:0];
  _RAND_166 = {1{`RANDOM}};
  state_vec__31 = _RAND_166[6:0];
  _RAND_167 = {1{`RANDOM}};
  state_vec_1_0 = _RAND_167[6:0];
  _RAND_168 = {1{`RANDOM}};
  state_vec_1_1 = _RAND_168[6:0];
  _RAND_169 = {1{`RANDOM}};
  state_vec_1_2 = _RAND_169[6:0];
  _RAND_170 = {1{`RANDOM}};
  state_vec_1_3 = _RAND_170[6:0];
  _RAND_171 = {1{`RANDOM}};
  state_vec_1_4 = _RAND_171[6:0];
  _RAND_172 = {1{`RANDOM}};
  state_vec_1_5 = _RAND_172[6:0];
  _RAND_173 = {1{`RANDOM}};
  state_vec_1_6 = _RAND_173[6:0];
  _RAND_174 = {1{`RANDOM}};
  state_vec_1_7 = _RAND_174[6:0];
  _RAND_175 = {1{`RANDOM}};
  state_vec_1_8 = _RAND_175[6:0];
  _RAND_176 = {1{`RANDOM}};
  state_vec_1_9 = _RAND_176[6:0];
  _RAND_177 = {1{`RANDOM}};
  state_vec_1_10 = _RAND_177[6:0];
  _RAND_178 = {1{`RANDOM}};
  state_vec_1_11 = _RAND_178[6:0];
  _RAND_179 = {1{`RANDOM}};
  state_vec_1_12 = _RAND_179[6:0];
  _RAND_180 = {1{`RANDOM}};
  state_vec_1_13 = _RAND_180[6:0];
  _RAND_181 = {1{`RANDOM}};
  state_vec_1_14 = _RAND_181[6:0];
  _RAND_182 = {1{`RANDOM}};
  state_vec_1_15 = _RAND_182[6:0];
  _RAND_183 = {1{`RANDOM}};
  state_vec_1_16 = _RAND_183[6:0];
  _RAND_184 = {1{`RANDOM}};
  state_vec_1_17 = _RAND_184[6:0];
  _RAND_185 = {1{`RANDOM}};
  state_vec_1_18 = _RAND_185[6:0];
  _RAND_186 = {1{`RANDOM}};
  state_vec_1_19 = _RAND_186[6:0];
  _RAND_187 = {1{`RANDOM}};
  state_vec_1_20 = _RAND_187[6:0];
  _RAND_188 = {1{`RANDOM}};
  state_vec_1_21 = _RAND_188[6:0];
  _RAND_189 = {1{`RANDOM}};
  state_vec_1_22 = _RAND_189[6:0];
  _RAND_190 = {1{`RANDOM}};
  state_vec_1_23 = _RAND_190[6:0];
  _RAND_191 = {1{`RANDOM}};
  state_vec_1_24 = _RAND_191[6:0];
  _RAND_192 = {1{`RANDOM}};
  state_vec_1_25 = _RAND_192[6:0];
  _RAND_193 = {1{`RANDOM}};
  state_vec_1_26 = _RAND_193[6:0];
  _RAND_194 = {1{`RANDOM}};
  state_vec_1_27 = _RAND_194[6:0];
  _RAND_195 = {1{`RANDOM}};
  state_vec_1_28 = _RAND_195[6:0];
  _RAND_196 = {1{`RANDOM}};
  state_vec_1_29 = _RAND_196[6:0];
  _RAND_197 = {1{`RANDOM}};
  state_vec_1_30 = _RAND_197[6:0];
  _RAND_198 = {1{`RANDOM}};
  state_vec_1_31 = _RAND_198[6:0];
  _RAND_199 = {1{`RANDOM}};
  s1_victim_oh_REG = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  s1_victim_oh_r0 = _RAND_200[7:0];
  _RAND_201 = {1{`RANDOM}};
  s1_victim_oh_r1 = _RAND_201[7:0];
  _RAND_202 = {1{`RANDOM}};
  s2_req_vsetIdx_0 = _RAND_202[5:0];
  _RAND_203 = {1{`RANDOM}};
  s2_tag_match_vec_0_7 = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  s2_tag_match_vec_0_6 = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  s2_tag_match_vec_0_5 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  s2_tag_match_vec_0_4 = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  s2_tag_match_vec_0_3 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  s2_tag_match_vec_0_2 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  s2_tag_match_vec_0_1 = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  s2_tag_match_vec_0_0 = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  s2_waymask_0 = _RAND_211[7:0];
  _RAND_212 = {1{`RANDOM}};
  s2_req_vsetIdx_1 = _RAND_212[5:0];
  _RAND_213 = {1{`RANDOM}};
  s2_tag_match_vec_1_7 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  s2_tag_match_vec_1_6 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  s2_tag_match_vec_1_5 = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  s2_tag_match_vec_1_4 = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  s2_tag_match_vec_1_3 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  s2_tag_match_vec_1_2 = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  s2_tag_match_vec_1_1 = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  s2_tag_match_vec_1_0 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  s2_waymask_1 = _RAND_221[7:0];
  _RAND_222 = {2{`RANDOM}};
  s2_req_paddr_0 = _RAND_222[35:0];
  _RAND_223 = {2{`RANDOM}};
  s2_req_paddr_1 = _RAND_223[35:0];
  _RAND_224 = {2{`RANDOM}};
  s2_req_vaddr_0 = _RAND_224[38:0];
  _RAND_225 = {2{`RANDOM}};
  s2_req_vaddr_1 = _RAND_225[38:0];
  _RAND_226 = {1{`RANDOM}};
  s2_meta_errors_0_0 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  s2_meta_errors_0_1 = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  s2_meta_errors_0_2 = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  s2_meta_errors_0_3 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  s2_meta_errors_0_4 = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  s2_meta_errors_0_5 = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  s2_meta_errors_0_6 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  s2_meta_errors_0_7 = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  s2_meta_errors_1_0 = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  s2_meta_errors_1_1 = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  s2_meta_errors_1_2 = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  s2_meta_errors_1_3 = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  s2_meta_errors_1_4 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  s2_meta_errors_1_5 = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  s2_meta_errors_1_6 = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  s2_meta_errors_1_7 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  s2_data_errorBits_0_0 = _RAND_242[31:0];
  _RAND_243 = {1{`RANDOM}};
  s2_data_errorBits_0_1 = _RAND_243[31:0];
  _RAND_244 = {1{`RANDOM}};
  s2_data_errorBits_0_2 = _RAND_244[31:0];
  _RAND_245 = {1{`RANDOM}};
  s2_data_errorBits_0_3 = _RAND_245[31:0];
  _RAND_246 = {1{`RANDOM}};
  s2_data_errorBits_0_4 = _RAND_246[31:0];
  _RAND_247 = {1{`RANDOM}};
  s2_data_errorBits_0_5 = _RAND_247[31:0];
  _RAND_248 = {1{`RANDOM}};
  s2_data_errorBits_0_6 = _RAND_248[31:0];
  _RAND_249 = {1{`RANDOM}};
  s2_data_errorBits_0_7 = _RAND_249[31:0];
  _RAND_250 = {1{`RANDOM}};
  s2_data_errorBits_1_0 = _RAND_250[31:0];
  _RAND_251 = {1{`RANDOM}};
  s2_data_errorBits_1_1 = _RAND_251[31:0];
  _RAND_252 = {1{`RANDOM}};
  s2_data_errorBits_1_2 = _RAND_252[31:0];
  _RAND_253 = {1{`RANDOM}};
  s2_data_errorBits_1_3 = _RAND_253[31:0];
  _RAND_254 = {1{`RANDOM}};
  s2_data_errorBits_1_4 = _RAND_254[31:0];
  _RAND_255 = {1{`RANDOM}};
  s2_data_errorBits_1_5 = _RAND_255[31:0];
  _RAND_256 = {1{`RANDOM}};
  s2_data_errorBits_1_6 = _RAND_256[31:0];
  _RAND_257 = {1{`RANDOM}};
  s2_data_errorBits_1_7 = _RAND_257[31:0];
  _RAND_258 = {16{`RANDOM}};
  s2_data_cacheline_0_0 = _RAND_258[511:0];
  _RAND_259 = {16{`RANDOM}};
  s2_data_cacheline_0_1 = _RAND_259[511:0];
  _RAND_260 = {16{`RANDOM}};
  s2_data_cacheline_0_2 = _RAND_260[511:0];
  _RAND_261 = {16{`RANDOM}};
  s2_data_cacheline_0_3 = _RAND_261[511:0];
  _RAND_262 = {16{`RANDOM}};
  s2_data_cacheline_0_4 = _RAND_262[511:0];
  _RAND_263 = {16{`RANDOM}};
  s2_data_cacheline_0_5 = _RAND_263[511:0];
  _RAND_264 = {16{`RANDOM}};
  s2_data_cacheline_0_6 = _RAND_264[511:0];
  _RAND_265 = {16{`RANDOM}};
  s2_data_cacheline_0_7 = _RAND_265[511:0];
  _RAND_266 = {16{`RANDOM}};
  s2_data_cacheline_1_0 = _RAND_266[511:0];
  _RAND_267 = {16{`RANDOM}};
  s2_data_cacheline_1_1 = _RAND_267[511:0];
  _RAND_268 = {16{`RANDOM}};
  s2_data_cacheline_1_2 = _RAND_268[511:0];
  _RAND_269 = {16{`RANDOM}};
  s2_data_cacheline_1_3 = _RAND_269[511:0];
  _RAND_270 = {16{`RANDOM}};
  s2_data_cacheline_1_4 = _RAND_270[511:0];
  _RAND_271 = {16{`RANDOM}};
  s2_data_cacheline_1_5 = _RAND_271[511:0];
  _RAND_272 = {16{`RANDOM}};
  s2_data_cacheline_1_6 = _RAND_272[511:0];
  _RAND_273 = {16{`RANDOM}};
  s2_data_cacheline_1_7 = _RAND_273[511:0];
  _RAND_274 = {1{`RANDOM}};
  s2_data_errors_0_0_REG = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  s2_data_errors_0_0_REG_1 = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  s2_data_errors_0_0_REG_2_0 = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  s2_data_errors_0_0_REG_2_1 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  s2_data_errors_0_0_REG_2_2 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  s2_data_errors_0_0_REG_2_3 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  s2_data_errors_0_0_REG_2_4 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  s2_data_errors_0_0_REG_2_5 = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  s2_data_errors_0_0_REG_2_6 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  s2_data_errors_0_0_REG_2_7 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  s2_data_errors_0_0_REG_2_8 = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  s2_data_errors_0_0_REG_2_9 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  s2_data_errors_0_0_REG_2_10 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  s2_data_errors_0_0_REG_2_11 = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  s2_data_errors_0_0_REG_2_12 = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  s2_data_errors_0_0_REG_2_13 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  s2_data_errors_0_0_REG_2_14 = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  s2_data_errors_0_0_REG_2_15 = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  s2_data_errors_0_0_REG_2_16 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  s2_data_errors_0_0_REG_2_17 = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  s2_data_errors_0_0_REG_2_18 = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  s2_data_errors_0_0_REG_2_19 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  s2_data_errors_0_0_REG_2_20 = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  s2_data_errors_0_0_REG_2_21 = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  s2_data_errors_0_0_REG_2_22 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  s2_data_errors_0_0_REG_2_23 = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  s2_data_errors_0_0_REG_2_24 = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  s2_data_errors_0_0_REG_2_25 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  s2_data_errors_0_0_REG_2_26 = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  s2_data_errors_0_0_REG_2_27 = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  s2_data_errors_0_0_REG_2_28 = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  s2_data_errors_0_0_REG_2_29 = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  s2_data_errors_0_0_REG_2_30 = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  s2_data_errors_0_0_REG_2_31 = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  s2_data_errors_0_1_REG = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  s2_data_errors_0_1_REG_1 = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  s2_data_errors_0_1_REG_2_0 = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  s2_data_errors_0_1_REG_2_1 = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  s2_data_errors_0_1_REG_2_2 = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  s2_data_errors_0_1_REG_2_3 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  s2_data_errors_0_1_REG_2_4 = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  s2_data_errors_0_1_REG_2_5 = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  s2_data_errors_0_1_REG_2_6 = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  s2_data_errors_0_1_REG_2_7 = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  s2_data_errors_0_1_REG_2_8 = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  s2_data_errors_0_1_REG_2_9 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  s2_data_errors_0_1_REG_2_10 = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  s2_data_errors_0_1_REG_2_11 = _RAND_321[0:0];
  _RAND_322 = {1{`RANDOM}};
  s2_data_errors_0_1_REG_2_12 = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  s2_data_errors_0_1_REG_2_13 = _RAND_323[0:0];
  _RAND_324 = {1{`RANDOM}};
  s2_data_errors_0_1_REG_2_14 = _RAND_324[0:0];
  _RAND_325 = {1{`RANDOM}};
  s2_data_errors_0_1_REG_2_15 = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  s2_data_errors_0_1_REG_2_16 = _RAND_326[0:0];
  _RAND_327 = {1{`RANDOM}};
  s2_data_errors_0_1_REG_2_17 = _RAND_327[0:0];
  _RAND_328 = {1{`RANDOM}};
  s2_data_errors_0_1_REG_2_18 = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  s2_data_errors_0_1_REG_2_19 = _RAND_329[0:0];
  _RAND_330 = {1{`RANDOM}};
  s2_data_errors_0_1_REG_2_20 = _RAND_330[0:0];
  _RAND_331 = {1{`RANDOM}};
  s2_data_errors_0_1_REG_2_21 = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  s2_data_errors_0_1_REG_2_22 = _RAND_332[0:0];
  _RAND_333 = {1{`RANDOM}};
  s2_data_errors_0_1_REG_2_23 = _RAND_333[0:0];
  _RAND_334 = {1{`RANDOM}};
  s2_data_errors_0_1_REG_2_24 = _RAND_334[0:0];
  _RAND_335 = {1{`RANDOM}};
  s2_data_errors_0_1_REG_2_25 = _RAND_335[0:0];
  _RAND_336 = {1{`RANDOM}};
  s2_data_errors_0_1_REG_2_26 = _RAND_336[0:0];
  _RAND_337 = {1{`RANDOM}};
  s2_data_errors_0_1_REG_2_27 = _RAND_337[0:0];
  _RAND_338 = {1{`RANDOM}};
  s2_data_errors_0_1_REG_2_28 = _RAND_338[0:0];
  _RAND_339 = {1{`RANDOM}};
  s2_data_errors_0_1_REG_2_29 = _RAND_339[0:0];
  _RAND_340 = {1{`RANDOM}};
  s2_data_errors_0_1_REG_2_30 = _RAND_340[0:0];
  _RAND_341 = {1{`RANDOM}};
  s2_data_errors_0_1_REG_2_31 = _RAND_341[0:0];
  _RAND_342 = {1{`RANDOM}};
  s2_data_errors_0_2_REG = _RAND_342[0:0];
  _RAND_343 = {1{`RANDOM}};
  s2_data_errors_0_2_REG_1 = _RAND_343[0:0];
  _RAND_344 = {1{`RANDOM}};
  s2_data_errors_0_2_REG_2_0 = _RAND_344[0:0];
  _RAND_345 = {1{`RANDOM}};
  s2_data_errors_0_2_REG_2_1 = _RAND_345[0:0];
  _RAND_346 = {1{`RANDOM}};
  s2_data_errors_0_2_REG_2_2 = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  s2_data_errors_0_2_REG_2_3 = _RAND_347[0:0];
  _RAND_348 = {1{`RANDOM}};
  s2_data_errors_0_2_REG_2_4 = _RAND_348[0:0];
  _RAND_349 = {1{`RANDOM}};
  s2_data_errors_0_2_REG_2_5 = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  s2_data_errors_0_2_REG_2_6 = _RAND_350[0:0];
  _RAND_351 = {1{`RANDOM}};
  s2_data_errors_0_2_REG_2_7 = _RAND_351[0:0];
  _RAND_352 = {1{`RANDOM}};
  s2_data_errors_0_2_REG_2_8 = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  s2_data_errors_0_2_REG_2_9 = _RAND_353[0:0];
  _RAND_354 = {1{`RANDOM}};
  s2_data_errors_0_2_REG_2_10 = _RAND_354[0:0];
  _RAND_355 = {1{`RANDOM}};
  s2_data_errors_0_2_REG_2_11 = _RAND_355[0:0];
  _RAND_356 = {1{`RANDOM}};
  s2_data_errors_0_2_REG_2_12 = _RAND_356[0:0];
  _RAND_357 = {1{`RANDOM}};
  s2_data_errors_0_2_REG_2_13 = _RAND_357[0:0];
  _RAND_358 = {1{`RANDOM}};
  s2_data_errors_0_2_REG_2_14 = _RAND_358[0:0];
  _RAND_359 = {1{`RANDOM}};
  s2_data_errors_0_2_REG_2_15 = _RAND_359[0:0];
  _RAND_360 = {1{`RANDOM}};
  s2_data_errors_0_2_REG_2_16 = _RAND_360[0:0];
  _RAND_361 = {1{`RANDOM}};
  s2_data_errors_0_2_REG_2_17 = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  s2_data_errors_0_2_REG_2_18 = _RAND_362[0:0];
  _RAND_363 = {1{`RANDOM}};
  s2_data_errors_0_2_REG_2_19 = _RAND_363[0:0];
  _RAND_364 = {1{`RANDOM}};
  s2_data_errors_0_2_REG_2_20 = _RAND_364[0:0];
  _RAND_365 = {1{`RANDOM}};
  s2_data_errors_0_2_REG_2_21 = _RAND_365[0:0];
  _RAND_366 = {1{`RANDOM}};
  s2_data_errors_0_2_REG_2_22 = _RAND_366[0:0];
  _RAND_367 = {1{`RANDOM}};
  s2_data_errors_0_2_REG_2_23 = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  s2_data_errors_0_2_REG_2_24 = _RAND_368[0:0];
  _RAND_369 = {1{`RANDOM}};
  s2_data_errors_0_2_REG_2_25 = _RAND_369[0:0];
  _RAND_370 = {1{`RANDOM}};
  s2_data_errors_0_2_REG_2_26 = _RAND_370[0:0];
  _RAND_371 = {1{`RANDOM}};
  s2_data_errors_0_2_REG_2_27 = _RAND_371[0:0];
  _RAND_372 = {1{`RANDOM}};
  s2_data_errors_0_2_REG_2_28 = _RAND_372[0:0];
  _RAND_373 = {1{`RANDOM}};
  s2_data_errors_0_2_REG_2_29 = _RAND_373[0:0];
  _RAND_374 = {1{`RANDOM}};
  s2_data_errors_0_2_REG_2_30 = _RAND_374[0:0];
  _RAND_375 = {1{`RANDOM}};
  s2_data_errors_0_2_REG_2_31 = _RAND_375[0:0];
  _RAND_376 = {1{`RANDOM}};
  s2_data_errors_0_3_REG = _RAND_376[0:0];
  _RAND_377 = {1{`RANDOM}};
  s2_data_errors_0_3_REG_1 = _RAND_377[0:0];
  _RAND_378 = {1{`RANDOM}};
  s2_data_errors_0_3_REG_2_0 = _RAND_378[0:0];
  _RAND_379 = {1{`RANDOM}};
  s2_data_errors_0_3_REG_2_1 = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  s2_data_errors_0_3_REG_2_2 = _RAND_380[0:0];
  _RAND_381 = {1{`RANDOM}};
  s2_data_errors_0_3_REG_2_3 = _RAND_381[0:0];
  _RAND_382 = {1{`RANDOM}};
  s2_data_errors_0_3_REG_2_4 = _RAND_382[0:0];
  _RAND_383 = {1{`RANDOM}};
  s2_data_errors_0_3_REG_2_5 = _RAND_383[0:0];
  _RAND_384 = {1{`RANDOM}};
  s2_data_errors_0_3_REG_2_6 = _RAND_384[0:0];
  _RAND_385 = {1{`RANDOM}};
  s2_data_errors_0_3_REG_2_7 = _RAND_385[0:0];
  _RAND_386 = {1{`RANDOM}};
  s2_data_errors_0_3_REG_2_8 = _RAND_386[0:0];
  _RAND_387 = {1{`RANDOM}};
  s2_data_errors_0_3_REG_2_9 = _RAND_387[0:0];
  _RAND_388 = {1{`RANDOM}};
  s2_data_errors_0_3_REG_2_10 = _RAND_388[0:0];
  _RAND_389 = {1{`RANDOM}};
  s2_data_errors_0_3_REG_2_11 = _RAND_389[0:0];
  _RAND_390 = {1{`RANDOM}};
  s2_data_errors_0_3_REG_2_12 = _RAND_390[0:0];
  _RAND_391 = {1{`RANDOM}};
  s2_data_errors_0_3_REG_2_13 = _RAND_391[0:0];
  _RAND_392 = {1{`RANDOM}};
  s2_data_errors_0_3_REG_2_14 = _RAND_392[0:0];
  _RAND_393 = {1{`RANDOM}};
  s2_data_errors_0_3_REG_2_15 = _RAND_393[0:0];
  _RAND_394 = {1{`RANDOM}};
  s2_data_errors_0_3_REG_2_16 = _RAND_394[0:0];
  _RAND_395 = {1{`RANDOM}};
  s2_data_errors_0_3_REG_2_17 = _RAND_395[0:0];
  _RAND_396 = {1{`RANDOM}};
  s2_data_errors_0_3_REG_2_18 = _RAND_396[0:0];
  _RAND_397 = {1{`RANDOM}};
  s2_data_errors_0_3_REG_2_19 = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  s2_data_errors_0_3_REG_2_20 = _RAND_398[0:0];
  _RAND_399 = {1{`RANDOM}};
  s2_data_errors_0_3_REG_2_21 = _RAND_399[0:0];
  _RAND_400 = {1{`RANDOM}};
  s2_data_errors_0_3_REG_2_22 = _RAND_400[0:0];
  _RAND_401 = {1{`RANDOM}};
  s2_data_errors_0_3_REG_2_23 = _RAND_401[0:0];
  _RAND_402 = {1{`RANDOM}};
  s2_data_errors_0_3_REG_2_24 = _RAND_402[0:0];
  _RAND_403 = {1{`RANDOM}};
  s2_data_errors_0_3_REG_2_25 = _RAND_403[0:0];
  _RAND_404 = {1{`RANDOM}};
  s2_data_errors_0_3_REG_2_26 = _RAND_404[0:0];
  _RAND_405 = {1{`RANDOM}};
  s2_data_errors_0_3_REG_2_27 = _RAND_405[0:0];
  _RAND_406 = {1{`RANDOM}};
  s2_data_errors_0_3_REG_2_28 = _RAND_406[0:0];
  _RAND_407 = {1{`RANDOM}};
  s2_data_errors_0_3_REG_2_29 = _RAND_407[0:0];
  _RAND_408 = {1{`RANDOM}};
  s2_data_errors_0_3_REG_2_30 = _RAND_408[0:0];
  _RAND_409 = {1{`RANDOM}};
  s2_data_errors_0_3_REG_2_31 = _RAND_409[0:0];
  _RAND_410 = {1{`RANDOM}};
  s2_data_errors_0_4_REG = _RAND_410[0:0];
  _RAND_411 = {1{`RANDOM}};
  s2_data_errors_0_4_REG_1 = _RAND_411[0:0];
  _RAND_412 = {1{`RANDOM}};
  s2_data_errors_0_4_REG_2_0 = _RAND_412[0:0];
  _RAND_413 = {1{`RANDOM}};
  s2_data_errors_0_4_REG_2_1 = _RAND_413[0:0];
  _RAND_414 = {1{`RANDOM}};
  s2_data_errors_0_4_REG_2_2 = _RAND_414[0:0];
  _RAND_415 = {1{`RANDOM}};
  s2_data_errors_0_4_REG_2_3 = _RAND_415[0:0];
  _RAND_416 = {1{`RANDOM}};
  s2_data_errors_0_4_REG_2_4 = _RAND_416[0:0];
  _RAND_417 = {1{`RANDOM}};
  s2_data_errors_0_4_REG_2_5 = _RAND_417[0:0];
  _RAND_418 = {1{`RANDOM}};
  s2_data_errors_0_4_REG_2_6 = _RAND_418[0:0];
  _RAND_419 = {1{`RANDOM}};
  s2_data_errors_0_4_REG_2_7 = _RAND_419[0:0];
  _RAND_420 = {1{`RANDOM}};
  s2_data_errors_0_4_REG_2_8 = _RAND_420[0:0];
  _RAND_421 = {1{`RANDOM}};
  s2_data_errors_0_4_REG_2_9 = _RAND_421[0:0];
  _RAND_422 = {1{`RANDOM}};
  s2_data_errors_0_4_REG_2_10 = _RAND_422[0:0];
  _RAND_423 = {1{`RANDOM}};
  s2_data_errors_0_4_REG_2_11 = _RAND_423[0:0];
  _RAND_424 = {1{`RANDOM}};
  s2_data_errors_0_4_REG_2_12 = _RAND_424[0:0];
  _RAND_425 = {1{`RANDOM}};
  s2_data_errors_0_4_REG_2_13 = _RAND_425[0:0];
  _RAND_426 = {1{`RANDOM}};
  s2_data_errors_0_4_REG_2_14 = _RAND_426[0:0];
  _RAND_427 = {1{`RANDOM}};
  s2_data_errors_0_4_REG_2_15 = _RAND_427[0:0];
  _RAND_428 = {1{`RANDOM}};
  s2_data_errors_0_4_REG_2_16 = _RAND_428[0:0];
  _RAND_429 = {1{`RANDOM}};
  s2_data_errors_0_4_REG_2_17 = _RAND_429[0:0];
  _RAND_430 = {1{`RANDOM}};
  s2_data_errors_0_4_REG_2_18 = _RAND_430[0:0];
  _RAND_431 = {1{`RANDOM}};
  s2_data_errors_0_4_REG_2_19 = _RAND_431[0:0];
  _RAND_432 = {1{`RANDOM}};
  s2_data_errors_0_4_REG_2_20 = _RAND_432[0:0];
  _RAND_433 = {1{`RANDOM}};
  s2_data_errors_0_4_REG_2_21 = _RAND_433[0:0];
  _RAND_434 = {1{`RANDOM}};
  s2_data_errors_0_4_REG_2_22 = _RAND_434[0:0];
  _RAND_435 = {1{`RANDOM}};
  s2_data_errors_0_4_REG_2_23 = _RAND_435[0:0];
  _RAND_436 = {1{`RANDOM}};
  s2_data_errors_0_4_REG_2_24 = _RAND_436[0:0];
  _RAND_437 = {1{`RANDOM}};
  s2_data_errors_0_4_REG_2_25 = _RAND_437[0:0];
  _RAND_438 = {1{`RANDOM}};
  s2_data_errors_0_4_REG_2_26 = _RAND_438[0:0];
  _RAND_439 = {1{`RANDOM}};
  s2_data_errors_0_4_REG_2_27 = _RAND_439[0:0];
  _RAND_440 = {1{`RANDOM}};
  s2_data_errors_0_4_REG_2_28 = _RAND_440[0:0];
  _RAND_441 = {1{`RANDOM}};
  s2_data_errors_0_4_REG_2_29 = _RAND_441[0:0];
  _RAND_442 = {1{`RANDOM}};
  s2_data_errors_0_4_REG_2_30 = _RAND_442[0:0];
  _RAND_443 = {1{`RANDOM}};
  s2_data_errors_0_4_REG_2_31 = _RAND_443[0:0];
  _RAND_444 = {1{`RANDOM}};
  s2_data_errors_0_5_REG = _RAND_444[0:0];
  _RAND_445 = {1{`RANDOM}};
  s2_data_errors_0_5_REG_1 = _RAND_445[0:0];
  _RAND_446 = {1{`RANDOM}};
  s2_data_errors_0_5_REG_2_0 = _RAND_446[0:0];
  _RAND_447 = {1{`RANDOM}};
  s2_data_errors_0_5_REG_2_1 = _RAND_447[0:0];
  _RAND_448 = {1{`RANDOM}};
  s2_data_errors_0_5_REG_2_2 = _RAND_448[0:0];
  _RAND_449 = {1{`RANDOM}};
  s2_data_errors_0_5_REG_2_3 = _RAND_449[0:0];
  _RAND_450 = {1{`RANDOM}};
  s2_data_errors_0_5_REG_2_4 = _RAND_450[0:0];
  _RAND_451 = {1{`RANDOM}};
  s2_data_errors_0_5_REG_2_5 = _RAND_451[0:0];
  _RAND_452 = {1{`RANDOM}};
  s2_data_errors_0_5_REG_2_6 = _RAND_452[0:0];
  _RAND_453 = {1{`RANDOM}};
  s2_data_errors_0_5_REG_2_7 = _RAND_453[0:0];
  _RAND_454 = {1{`RANDOM}};
  s2_data_errors_0_5_REG_2_8 = _RAND_454[0:0];
  _RAND_455 = {1{`RANDOM}};
  s2_data_errors_0_5_REG_2_9 = _RAND_455[0:0];
  _RAND_456 = {1{`RANDOM}};
  s2_data_errors_0_5_REG_2_10 = _RAND_456[0:0];
  _RAND_457 = {1{`RANDOM}};
  s2_data_errors_0_5_REG_2_11 = _RAND_457[0:0];
  _RAND_458 = {1{`RANDOM}};
  s2_data_errors_0_5_REG_2_12 = _RAND_458[0:0];
  _RAND_459 = {1{`RANDOM}};
  s2_data_errors_0_5_REG_2_13 = _RAND_459[0:0];
  _RAND_460 = {1{`RANDOM}};
  s2_data_errors_0_5_REG_2_14 = _RAND_460[0:0];
  _RAND_461 = {1{`RANDOM}};
  s2_data_errors_0_5_REG_2_15 = _RAND_461[0:0];
  _RAND_462 = {1{`RANDOM}};
  s2_data_errors_0_5_REG_2_16 = _RAND_462[0:0];
  _RAND_463 = {1{`RANDOM}};
  s2_data_errors_0_5_REG_2_17 = _RAND_463[0:0];
  _RAND_464 = {1{`RANDOM}};
  s2_data_errors_0_5_REG_2_18 = _RAND_464[0:0];
  _RAND_465 = {1{`RANDOM}};
  s2_data_errors_0_5_REG_2_19 = _RAND_465[0:0];
  _RAND_466 = {1{`RANDOM}};
  s2_data_errors_0_5_REG_2_20 = _RAND_466[0:0];
  _RAND_467 = {1{`RANDOM}};
  s2_data_errors_0_5_REG_2_21 = _RAND_467[0:0];
  _RAND_468 = {1{`RANDOM}};
  s2_data_errors_0_5_REG_2_22 = _RAND_468[0:0];
  _RAND_469 = {1{`RANDOM}};
  s2_data_errors_0_5_REG_2_23 = _RAND_469[0:0];
  _RAND_470 = {1{`RANDOM}};
  s2_data_errors_0_5_REG_2_24 = _RAND_470[0:0];
  _RAND_471 = {1{`RANDOM}};
  s2_data_errors_0_5_REG_2_25 = _RAND_471[0:0];
  _RAND_472 = {1{`RANDOM}};
  s2_data_errors_0_5_REG_2_26 = _RAND_472[0:0];
  _RAND_473 = {1{`RANDOM}};
  s2_data_errors_0_5_REG_2_27 = _RAND_473[0:0];
  _RAND_474 = {1{`RANDOM}};
  s2_data_errors_0_5_REG_2_28 = _RAND_474[0:0];
  _RAND_475 = {1{`RANDOM}};
  s2_data_errors_0_5_REG_2_29 = _RAND_475[0:0];
  _RAND_476 = {1{`RANDOM}};
  s2_data_errors_0_5_REG_2_30 = _RAND_476[0:0];
  _RAND_477 = {1{`RANDOM}};
  s2_data_errors_0_5_REG_2_31 = _RAND_477[0:0];
  _RAND_478 = {1{`RANDOM}};
  s2_data_errors_0_6_REG = _RAND_478[0:0];
  _RAND_479 = {1{`RANDOM}};
  s2_data_errors_0_6_REG_1 = _RAND_479[0:0];
  _RAND_480 = {1{`RANDOM}};
  s2_data_errors_0_6_REG_2_0 = _RAND_480[0:0];
  _RAND_481 = {1{`RANDOM}};
  s2_data_errors_0_6_REG_2_1 = _RAND_481[0:0];
  _RAND_482 = {1{`RANDOM}};
  s2_data_errors_0_6_REG_2_2 = _RAND_482[0:0];
  _RAND_483 = {1{`RANDOM}};
  s2_data_errors_0_6_REG_2_3 = _RAND_483[0:0];
  _RAND_484 = {1{`RANDOM}};
  s2_data_errors_0_6_REG_2_4 = _RAND_484[0:0];
  _RAND_485 = {1{`RANDOM}};
  s2_data_errors_0_6_REG_2_5 = _RAND_485[0:0];
  _RAND_486 = {1{`RANDOM}};
  s2_data_errors_0_6_REG_2_6 = _RAND_486[0:0];
  _RAND_487 = {1{`RANDOM}};
  s2_data_errors_0_6_REG_2_7 = _RAND_487[0:0];
  _RAND_488 = {1{`RANDOM}};
  s2_data_errors_0_6_REG_2_8 = _RAND_488[0:0];
  _RAND_489 = {1{`RANDOM}};
  s2_data_errors_0_6_REG_2_9 = _RAND_489[0:0];
  _RAND_490 = {1{`RANDOM}};
  s2_data_errors_0_6_REG_2_10 = _RAND_490[0:0];
  _RAND_491 = {1{`RANDOM}};
  s2_data_errors_0_6_REG_2_11 = _RAND_491[0:0];
  _RAND_492 = {1{`RANDOM}};
  s2_data_errors_0_6_REG_2_12 = _RAND_492[0:0];
  _RAND_493 = {1{`RANDOM}};
  s2_data_errors_0_6_REG_2_13 = _RAND_493[0:0];
  _RAND_494 = {1{`RANDOM}};
  s2_data_errors_0_6_REG_2_14 = _RAND_494[0:0];
  _RAND_495 = {1{`RANDOM}};
  s2_data_errors_0_6_REG_2_15 = _RAND_495[0:0];
  _RAND_496 = {1{`RANDOM}};
  s2_data_errors_0_6_REG_2_16 = _RAND_496[0:0];
  _RAND_497 = {1{`RANDOM}};
  s2_data_errors_0_6_REG_2_17 = _RAND_497[0:0];
  _RAND_498 = {1{`RANDOM}};
  s2_data_errors_0_6_REG_2_18 = _RAND_498[0:0];
  _RAND_499 = {1{`RANDOM}};
  s2_data_errors_0_6_REG_2_19 = _RAND_499[0:0];
  _RAND_500 = {1{`RANDOM}};
  s2_data_errors_0_6_REG_2_20 = _RAND_500[0:0];
  _RAND_501 = {1{`RANDOM}};
  s2_data_errors_0_6_REG_2_21 = _RAND_501[0:0];
  _RAND_502 = {1{`RANDOM}};
  s2_data_errors_0_6_REG_2_22 = _RAND_502[0:0];
  _RAND_503 = {1{`RANDOM}};
  s2_data_errors_0_6_REG_2_23 = _RAND_503[0:0];
  _RAND_504 = {1{`RANDOM}};
  s2_data_errors_0_6_REG_2_24 = _RAND_504[0:0];
  _RAND_505 = {1{`RANDOM}};
  s2_data_errors_0_6_REG_2_25 = _RAND_505[0:0];
  _RAND_506 = {1{`RANDOM}};
  s2_data_errors_0_6_REG_2_26 = _RAND_506[0:0];
  _RAND_507 = {1{`RANDOM}};
  s2_data_errors_0_6_REG_2_27 = _RAND_507[0:0];
  _RAND_508 = {1{`RANDOM}};
  s2_data_errors_0_6_REG_2_28 = _RAND_508[0:0];
  _RAND_509 = {1{`RANDOM}};
  s2_data_errors_0_6_REG_2_29 = _RAND_509[0:0];
  _RAND_510 = {1{`RANDOM}};
  s2_data_errors_0_6_REG_2_30 = _RAND_510[0:0];
  _RAND_511 = {1{`RANDOM}};
  s2_data_errors_0_6_REG_2_31 = _RAND_511[0:0];
  _RAND_512 = {1{`RANDOM}};
  s2_data_errors_0_7_REG = _RAND_512[0:0];
  _RAND_513 = {1{`RANDOM}};
  s2_data_errors_0_7_REG_1 = _RAND_513[0:0];
  _RAND_514 = {1{`RANDOM}};
  s2_data_errors_0_7_REG_2_0 = _RAND_514[0:0];
  _RAND_515 = {1{`RANDOM}};
  s2_data_errors_0_7_REG_2_1 = _RAND_515[0:0];
  _RAND_516 = {1{`RANDOM}};
  s2_data_errors_0_7_REG_2_2 = _RAND_516[0:0];
  _RAND_517 = {1{`RANDOM}};
  s2_data_errors_0_7_REG_2_3 = _RAND_517[0:0];
  _RAND_518 = {1{`RANDOM}};
  s2_data_errors_0_7_REG_2_4 = _RAND_518[0:0];
  _RAND_519 = {1{`RANDOM}};
  s2_data_errors_0_7_REG_2_5 = _RAND_519[0:0];
  _RAND_520 = {1{`RANDOM}};
  s2_data_errors_0_7_REG_2_6 = _RAND_520[0:0];
  _RAND_521 = {1{`RANDOM}};
  s2_data_errors_0_7_REG_2_7 = _RAND_521[0:0];
  _RAND_522 = {1{`RANDOM}};
  s2_data_errors_0_7_REG_2_8 = _RAND_522[0:0];
  _RAND_523 = {1{`RANDOM}};
  s2_data_errors_0_7_REG_2_9 = _RAND_523[0:0];
  _RAND_524 = {1{`RANDOM}};
  s2_data_errors_0_7_REG_2_10 = _RAND_524[0:0];
  _RAND_525 = {1{`RANDOM}};
  s2_data_errors_0_7_REG_2_11 = _RAND_525[0:0];
  _RAND_526 = {1{`RANDOM}};
  s2_data_errors_0_7_REG_2_12 = _RAND_526[0:0];
  _RAND_527 = {1{`RANDOM}};
  s2_data_errors_0_7_REG_2_13 = _RAND_527[0:0];
  _RAND_528 = {1{`RANDOM}};
  s2_data_errors_0_7_REG_2_14 = _RAND_528[0:0];
  _RAND_529 = {1{`RANDOM}};
  s2_data_errors_0_7_REG_2_15 = _RAND_529[0:0];
  _RAND_530 = {1{`RANDOM}};
  s2_data_errors_0_7_REG_2_16 = _RAND_530[0:0];
  _RAND_531 = {1{`RANDOM}};
  s2_data_errors_0_7_REG_2_17 = _RAND_531[0:0];
  _RAND_532 = {1{`RANDOM}};
  s2_data_errors_0_7_REG_2_18 = _RAND_532[0:0];
  _RAND_533 = {1{`RANDOM}};
  s2_data_errors_0_7_REG_2_19 = _RAND_533[0:0];
  _RAND_534 = {1{`RANDOM}};
  s2_data_errors_0_7_REG_2_20 = _RAND_534[0:0];
  _RAND_535 = {1{`RANDOM}};
  s2_data_errors_0_7_REG_2_21 = _RAND_535[0:0];
  _RAND_536 = {1{`RANDOM}};
  s2_data_errors_0_7_REG_2_22 = _RAND_536[0:0];
  _RAND_537 = {1{`RANDOM}};
  s2_data_errors_0_7_REG_2_23 = _RAND_537[0:0];
  _RAND_538 = {1{`RANDOM}};
  s2_data_errors_0_7_REG_2_24 = _RAND_538[0:0];
  _RAND_539 = {1{`RANDOM}};
  s2_data_errors_0_7_REG_2_25 = _RAND_539[0:0];
  _RAND_540 = {1{`RANDOM}};
  s2_data_errors_0_7_REG_2_26 = _RAND_540[0:0];
  _RAND_541 = {1{`RANDOM}};
  s2_data_errors_0_7_REG_2_27 = _RAND_541[0:0];
  _RAND_542 = {1{`RANDOM}};
  s2_data_errors_0_7_REG_2_28 = _RAND_542[0:0];
  _RAND_543 = {1{`RANDOM}};
  s2_data_errors_0_7_REG_2_29 = _RAND_543[0:0];
  _RAND_544 = {1{`RANDOM}};
  s2_data_errors_0_7_REG_2_30 = _RAND_544[0:0];
  _RAND_545 = {1{`RANDOM}};
  s2_data_errors_0_7_REG_2_31 = _RAND_545[0:0];
  _RAND_546 = {1{`RANDOM}};
  s2_data_errors_1_0_REG = _RAND_546[0:0];
  _RAND_547 = {1{`RANDOM}};
  s2_data_errors_1_0_REG_1 = _RAND_547[0:0];
  _RAND_548 = {1{`RANDOM}};
  s2_data_errors_1_0_REG_2 = _RAND_548[0:0];
  _RAND_549 = {1{`RANDOM}};
  s2_data_errors_1_0_REG_3 = _RAND_549[0:0];
  _RAND_550 = {1{`RANDOM}};
  s2_data_errors_1_0_REG_4_0 = _RAND_550[0:0];
  _RAND_551 = {1{`RANDOM}};
  s2_data_errors_1_0_REG_4_1 = _RAND_551[0:0];
  _RAND_552 = {1{`RANDOM}};
  s2_data_errors_1_0_REG_4_2 = _RAND_552[0:0];
  _RAND_553 = {1{`RANDOM}};
  s2_data_errors_1_0_REG_4_3 = _RAND_553[0:0];
  _RAND_554 = {1{`RANDOM}};
  s2_data_errors_1_0_REG_4_4 = _RAND_554[0:0];
  _RAND_555 = {1{`RANDOM}};
  s2_data_errors_1_0_REG_4_5 = _RAND_555[0:0];
  _RAND_556 = {1{`RANDOM}};
  s2_data_errors_1_0_REG_4_6 = _RAND_556[0:0];
  _RAND_557 = {1{`RANDOM}};
  s2_data_errors_1_0_REG_4_7 = _RAND_557[0:0];
  _RAND_558 = {1{`RANDOM}};
  s2_data_errors_1_0_REG_4_8 = _RAND_558[0:0];
  _RAND_559 = {1{`RANDOM}};
  s2_data_errors_1_0_REG_4_9 = _RAND_559[0:0];
  _RAND_560 = {1{`RANDOM}};
  s2_data_errors_1_0_REG_4_10 = _RAND_560[0:0];
  _RAND_561 = {1{`RANDOM}};
  s2_data_errors_1_0_REG_4_11 = _RAND_561[0:0];
  _RAND_562 = {1{`RANDOM}};
  s2_data_errors_1_0_REG_4_12 = _RAND_562[0:0];
  _RAND_563 = {1{`RANDOM}};
  s2_data_errors_1_0_REG_4_13 = _RAND_563[0:0];
  _RAND_564 = {1{`RANDOM}};
  s2_data_errors_1_0_REG_4_14 = _RAND_564[0:0];
  _RAND_565 = {1{`RANDOM}};
  s2_data_errors_1_0_REG_4_15 = _RAND_565[0:0];
  _RAND_566 = {1{`RANDOM}};
  s2_data_errors_1_0_REG_4_16 = _RAND_566[0:0];
  _RAND_567 = {1{`RANDOM}};
  s2_data_errors_1_0_REG_4_17 = _RAND_567[0:0];
  _RAND_568 = {1{`RANDOM}};
  s2_data_errors_1_0_REG_4_18 = _RAND_568[0:0];
  _RAND_569 = {1{`RANDOM}};
  s2_data_errors_1_0_REG_4_19 = _RAND_569[0:0];
  _RAND_570 = {1{`RANDOM}};
  s2_data_errors_1_0_REG_4_20 = _RAND_570[0:0];
  _RAND_571 = {1{`RANDOM}};
  s2_data_errors_1_0_REG_4_21 = _RAND_571[0:0];
  _RAND_572 = {1{`RANDOM}};
  s2_data_errors_1_0_REG_4_22 = _RAND_572[0:0];
  _RAND_573 = {1{`RANDOM}};
  s2_data_errors_1_0_REG_4_23 = _RAND_573[0:0];
  _RAND_574 = {1{`RANDOM}};
  s2_data_errors_1_0_REG_4_24 = _RAND_574[0:0];
  _RAND_575 = {1{`RANDOM}};
  s2_data_errors_1_0_REG_4_25 = _RAND_575[0:0];
  _RAND_576 = {1{`RANDOM}};
  s2_data_errors_1_0_REG_4_26 = _RAND_576[0:0];
  _RAND_577 = {1{`RANDOM}};
  s2_data_errors_1_0_REG_4_27 = _RAND_577[0:0];
  _RAND_578 = {1{`RANDOM}};
  s2_data_errors_1_0_REG_4_28 = _RAND_578[0:0];
  _RAND_579 = {1{`RANDOM}};
  s2_data_errors_1_0_REG_4_29 = _RAND_579[0:0];
  _RAND_580 = {1{`RANDOM}};
  s2_data_errors_1_0_REG_4_30 = _RAND_580[0:0];
  _RAND_581 = {1{`RANDOM}};
  s2_data_errors_1_0_REG_4_31 = _RAND_581[0:0];
  _RAND_582 = {1{`RANDOM}};
  s2_data_errors_1_1_REG = _RAND_582[0:0];
  _RAND_583 = {1{`RANDOM}};
  s2_data_errors_1_1_REG_1 = _RAND_583[0:0];
  _RAND_584 = {1{`RANDOM}};
  s2_data_errors_1_1_REG_2 = _RAND_584[0:0];
  _RAND_585 = {1{`RANDOM}};
  s2_data_errors_1_1_REG_3 = _RAND_585[0:0];
  _RAND_586 = {1{`RANDOM}};
  s2_data_errors_1_1_REG_4_0 = _RAND_586[0:0];
  _RAND_587 = {1{`RANDOM}};
  s2_data_errors_1_1_REG_4_1 = _RAND_587[0:0];
  _RAND_588 = {1{`RANDOM}};
  s2_data_errors_1_1_REG_4_2 = _RAND_588[0:0];
  _RAND_589 = {1{`RANDOM}};
  s2_data_errors_1_1_REG_4_3 = _RAND_589[0:0];
  _RAND_590 = {1{`RANDOM}};
  s2_data_errors_1_1_REG_4_4 = _RAND_590[0:0];
  _RAND_591 = {1{`RANDOM}};
  s2_data_errors_1_1_REG_4_5 = _RAND_591[0:0];
  _RAND_592 = {1{`RANDOM}};
  s2_data_errors_1_1_REG_4_6 = _RAND_592[0:0];
  _RAND_593 = {1{`RANDOM}};
  s2_data_errors_1_1_REG_4_7 = _RAND_593[0:0];
  _RAND_594 = {1{`RANDOM}};
  s2_data_errors_1_1_REG_4_8 = _RAND_594[0:0];
  _RAND_595 = {1{`RANDOM}};
  s2_data_errors_1_1_REG_4_9 = _RAND_595[0:0];
  _RAND_596 = {1{`RANDOM}};
  s2_data_errors_1_1_REG_4_10 = _RAND_596[0:0];
  _RAND_597 = {1{`RANDOM}};
  s2_data_errors_1_1_REG_4_11 = _RAND_597[0:0];
  _RAND_598 = {1{`RANDOM}};
  s2_data_errors_1_1_REG_4_12 = _RAND_598[0:0];
  _RAND_599 = {1{`RANDOM}};
  s2_data_errors_1_1_REG_4_13 = _RAND_599[0:0];
  _RAND_600 = {1{`RANDOM}};
  s2_data_errors_1_1_REG_4_14 = _RAND_600[0:0];
  _RAND_601 = {1{`RANDOM}};
  s2_data_errors_1_1_REG_4_15 = _RAND_601[0:0];
  _RAND_602 = {1{`RANDOM}};
  s2_data_errors_1_1_REG_4_16 = _RAND_602[0:0];
  _RAND_603 = {1{`RANDOM}};
  s2_data_errors_1_1_REG_4_17 = _RAND_603[0:0];
  _RAND_604 = {1{`RANDOM}};
  s2_data_errors_1_1_REG_4_18 = _RAND_604[0:0];
  _RAND_605 = {1{`RANDOM}};
  s2_data_errors_1_1_REG_4_19 = _RAND_605[0:0];
  _RAND_606 = {1{`RANDOM}};
  s2_data_errors_1_1_REG_4_20 = _RAND_606[0:0];
  _RAND_607 = {1{`RANDOM}};
  s2_data_errors_1_1_REG_4_21 = _RAND_607[0:0];
  _RAND_608 = {1{`RANDOM}};
  s2_data_errors_1_1_REG_4_22 = _RAND_608[0:0];
  _RAND_609 = {1{`RANDOM}};
  s2_data_errors_1_1_REG_4_23 = _RAND_609[0:0];
  _RAND_610 = {1{`RANDOM}};
  s2_data_errors_1_1_REG_4_24 = _RAND_610[0:0];
  _RAND_611 = {1{`RANDOM}};
  s2_data_errors_1_1_REG_4_25 = _RAND_611[0:0];
  _RAND_612 = {1{`RANDOM}};
  s2_data_errors_1_1_REG_4_26 = _RAND_612[0:0];
  _RAND_613 = {1{`RANDOM}};
  s2_data_errors_1_1_REG_4_27 = _RAND_613[0:0];
  _RAND_614 = {1{`RANDOM}};
  s2_data_errors_1_1_REG_4_28 = _RAND_614[0:0];
  _RAND_615 = {1{`RANDOM}};
  s2_data_errors_1_1_REG_4_29 = _RAND_615[0:0];
  _RAND_616 = {1{`RANDOM}};
  s2_data_errors_1_1_REG_4_30 = _RAND_616[0:0];
  _RAND_617 = {1{`RANDOM}};
  s2_data_errors_1_1_REG_4_31 = _RAND_617[0:0];
  _RAND_618 = {1{`RANDOM}};
  s2_data_errors_1_2_REG = _RAND_618[0:0];
  _RAND_619 = {1{`RANDOM}};
  s2_data_errors_1_2_REG_1 = _RAND_619[0:0];
  _RAND_620 = {1{`RANDOM}};
  s2_data_errors_1_2_REG_2 = _RAND_620[0:0];
  _RAND_621 = {1{`RANDOM}};
  s2_data_errors_1_2_REG_3 = _RAND_621[0:0];
  _RAND_622 = {1{`RANDOM}};
  s2_data_errors_1_2_REG_4_0 = _RAND_622[0:0];
  _RAND_623 = {1{`RANDOM}};
  s2_data_errors_1_2_REG_4_1 = _RAND_623[0:0];
  _RAND_624 = {1{`RANDOM}};
  s2_data_errors_1_2_REG_4_2 = _RAND_624[0:0];
  _RAND_625 = {1{`RANDOM}};
  s2_data_errors_1_2_REG_4_3 = _RAND_625[0:0];
  _RAND_626 = {1{`RANDOM}};
  s2_data_errors_1_2_REG_4_4 = _RAND_626[0:0];
  _RAND_627 = {1{`RANDOM}};
  s2_data_errors_1_2_REG_4_5 = _RAND_627[0:0];
  _RAND_628 = {1{`RANDOM}};
  s2_data_errors_1_2_REG_4_6 = _RAND_628[0:0];
  _RAND_629 = {1{`RANDOM}};
  s2_data_errors_1_2_REG_4_7 = _RAND_629[0:0];
  _RAND_630 = {1{`RANDOM}};
  s2_data_errors_1_2_REG_4_8 = _RAND_630[0:0];
  _RAND_631 = {1{`RANDOM}};
  s2_data_errors_1_2_REG_4_9 = _RAND_631[0:0];
  _RAND_632 = {1{`RANDOM}};
  s2_data_errors_1_2_REG_4_10 = _RAND_632[0:0];
  _RAND_633 = {1{`RANDOM}};
  s2_data_errors_1_2_REG_4_11 = _RAND_633[0:0];
  _RAND_634 = {1{`RANDOM}};
  s2_data_errors_1_2_REG_4_12 = _RAND_634[0:0];
  _RAND_635 = {1{`RANDOM}};
  s2_data_errors_1_2_REG_4_13 = _RAND_635[0:0];
  _RAND_636 = {1{`RANDOM}};
  s2_data_errors_1_2_REG_4_14 = _RAND_636[0:0];
  _RAND_637 = {1{`RANDOM}};
  s2_data_errors_1_2_REG_4_15 = _RAND_637[0:0];
  _RAND_638 = {1{`RANDOM}};
  s2_data_errors_1_2_REG_4_16 = _RAND_638[0:0];
  _RAND_639 = {1{`RANDOM}};
  s2_data_errors_1_2_REG_4_17 = _RAND_639[0:0];
  _RAND_640 = {1{`RANDOM}};
  s2_data_errors_1_2_REG_4_18 = _RAND_640[0:0];
  _RAND_641 = {1{`RANDOM}};
  s2_data_errors_1_2_REG_4_19 = _RAND_641[0:0];
  _RAND_642 = {1{`RANDOM}};
  s2_data_errors_1_2_REG_4_20 = _RAND_642[0:0];
  _RAND_643 = {1{`RANDOM}};
  s2_data_errors_1_2_REG_4_21 = _RAND_643[0:0];
  _RAND_644 = {1{`RANDOM}};
  s2_data_errors_1_2_REG_4_22 = _RAND_644[0:0];
  _RAND_645 = {1{`RANDOM}};
  s2_data_errors_1_2_REG_4_23 = _RAND_645[0:0];
  _RAND_646 = {1{`RANDOM}};
  s2_data_errors_1_2_REG_4_24 = _RAND_646[0:0];
  _RAND_647 = {1{`RANDOM}};
  s2_data_errors_1_2_REG_4_25 = _RAND_647[0:0];
  _RAND_648 = {1{`RANDOM}};
  s2_data_errors_1_2_REG_4_26 = _RAND_648[0:0];
  _RAND_649 = {1{`RANDOM}};
  s2_data_errors_1_2_REG_4_27 = _RAND_649[0:0];
  _RAND_650 = {1{`RANDOM}};
  s2_data_errors_1_2_REG_4_28 = _RAND_650[0:0];
  _RAND_651 = {1{`RANDOM}};
  s2_data_errors_1_2_REG_4_29 = _RAND_651[0:0];
  _RAND_652 = {1{`RANDOM}};
  s2_data_errors_1_2_REG_4_30 = _RAND_652[0:0];
  _RAND_653 = {1{`RANDOM}};
  s2_data_errors_1_2_REG_4_31 = _RAND_653[0:0];
  _RAND_654 = {1{`RANDOM}};
  s2_data_errors_1_3_REG = _RAND_654[0:0];
  _RAND_655 = {1{`RANDOM}};
  s2_data_errors_1_3_REG_1 = _RAND_655[0:0];
  _RAND_656 = {1{`RANDOM}};
  s2_data_errors_1_3_REG_2 = _RAND_656[0:0];
  _RAND_657 = {1{`RANDOM}};
  s2_data_errors_1_3_REG_3 = _RAND_657[0:0];
  _RAND_658 = {1{`RANDOM}};
  s2_data_errors_1_3_REG_4_0 = _RAND_658[0:0];
  _RAND_659 = {1{`RANDOM}};
  s2_data_errors_1_3_REG_4_1 = _RAND_659[0:0];
  _RAND_660 = {1{`RANDOM}};
  s2_data_errors_1_3_REG_4_2 = _RAND_660[0:0];
  _RAND_661 = {1{`RANDOM}};
  s2_data_errors_1_3_REG_4_3 = _RAND_661[0:0];
  _RAND_662 = {1{`RANDOM}};
  s2_data_errors_1_3_REG_4_4 = _RAND_662[0:0];
  _RAND_663 = {1{`RANDOM}};
  s2_data_errors_1_3_REG_4_5 = _RAND_663[0:0];
  _RAND_664 = {1{`RANDOM}};
  s2_data_errors_1_3_REG_4_6 = _RAND_664[0:0];
  _RAND_665 = {1{`RANDOM}};
  s2_data_errors_1_3_REG_4_7 = _RAND_665[0:0];
  _RAND_666 = {1{`RANDOM}};
  s2_data_errors_1_3_REG_4_8 = _RAND_666[0:0];
  _RAND_667 = {1{`RANDOM}};
  s2_data_errors_1_3_REG_4_9 = _RAND_667[0:0];
  _RAND_668 = {1{`RANDOM}};
  s2_data_errors_1_3_REG_4_10 = _RAND_668[0:0];
  _RAND_669 = {1{`RANDOM}};
  s2_data_errors_1_3_REG_4_11 = _RAND_669[0:0];
  _RAND_670 = {1{`RANDOM}};
  s2_data_errors_1_3_REG_4_12 = _RAND_670[0:0];
  _RAND_671 = {1{`RANDOM}};
  s2_data_errors_1_3_REG_4_13 = _RAND_671[0:0];
  _RAND_672 = {1{`RANDOM}};
  s2_data_errors_1_3_REG_4_14 = _RAND_672[0:0];
  _RAND_673 = {1{`RANDOM}};
  s2_data_errors_1_3_REG_4_15 = _RAND_673[0:0];
  _RAND_674 = {1{`RANDOM}};
  s2_data_errors_1_3_REG_4_16 = _RAND_674[0:0];
  _RAND_675 = {1{`RANDOM}};
  s2_data_errors_1_3_REG_4_17 = _RAND_675[0:0];
  _RAND_676 = {1{`RANDOM}};
  s2_data_errors_1_3_REG_4_18 = _RAND_676[0:0];
  _RAND_677 = {1{`RANDOM}};
  s2_data_errors_1_3_REG_4_19 = _RAND_677[0:0];
  _RAND_678 = {1{`RANDOM}};
  s2_data_errors_1_3_REG_4_20 = _RAND_678[0:0];
  _RAND_679 = {1{`RANDOM}};
  s2_data_errors_1_3_REG_4_21 = _RAND_679[0:0];
  _RAND_680 = {1{`RANDOM}};
  s2_data_errors_1_3_REG_4_22 = _RAND_680[0:0];
  _RAND_681 = {1{`RANDOM}};
  s2_data_errors_1_3_REG_4_23 = _RAND_681[0:0];
  _RAND_682 = {1{`RANDOM}};
  s2_data_errors_1_3_REG_4_24 = _RAND_682[0:0];
  _RAND_683 = {1{`RANDOM}};
  s2_data_errors_1_3_REG_4_25 = _RAND_683[0:0];
  _RAND_684 = {1{`RANDOM}};
  s2_data_errors_1_3_REG_4_26 = _RAND_684[0:0];
  _RAND_685 = {1{`RANDOM}};
  s2_data_errors_1_3_REG_4_27 = _RAND_685[0:0];
  _RAND_686 = {1{`RANDOM}};
  s2_data_errors_1_3_REG_4_28 = _RAND_686[0:0];
  _RAND_687 = {1{`RANDOM}};
  s2_data_errors_1_3_REG_4_29 = _RAND_687[0:0];
  _RAND_688 = {1{`RANDOM}};
  s2_data_errors_1_3_REG_4_30 = _RAND_688[0:0];
  _RAND_689 = {1{`RANDOM}};
  s2_data_errors_1_3_REG_4_31 = _RAND_689[0:0];
  _RAND_690 = {1{`RANDOM}};
  s2_data_errors_1_4_REG = _RAND_690[0:0];
  _RAND_691 = {1{`RANDOM}};
  s2_data_errors_1_4_REG_1 = _RAND_691[0:0];
  _RAND_692 = {1{`RANDOM}};
  s2_data_errors_1_4_REG_2 = _RAND_692[0:0];
  _RAND_693 = {1{`RANDOM}};
  s2_data_errors_1_4_REG_3 = _RAND_693[0:0];
  _RAND_694 = {1{`RANDOM}};
  s2_data_errors_1_4_REG_4_0 = _RAND_694[0:0];
  _RAND_695 = {1{`RANDOM}};
  s2_data_errors_1_4_REG_4_1 = _RAND_695[0:0];
  _RAND_696 = {1{`RANDOM}};
  s2_data_errors_1_4_REG_4_2 = _RAND_696[0:0];
  _RAND_697 = {1{`RANDOM}};
  s2_data_errors_1_4_REG_4_3 = _RAND_697[0:0];
  _RAND_698 = {1{`RANDOM}};
  s2_data_errors_1_4_REG_4_4 = _RAND_698[0:0];
  _RAND_699 = {1{`RANDOM}};
  s2_data_errors_1_4_REG_4_5 = _RAND_699[0:0];
  _RAND_700 = {1{`RANDOM}};
  s2_data_errors_1_4_REG_4_6 = _RAND_700[0:0];
  _RAND_701 = {1{`RANDOM}};
  s2_data_errors_1_4_REG_4_7 = _RAND_701[0:0];
  _RAND_702 = {1{`RANDOM}};
  s2_data_errors_1_4_REG_4_8 = _RAND_702[0:0];
  _RAND_703 = {1{`RANDOM}};
  s2_data_errors_1_4_REG_4_9 = _RAND_703[0:0];
  _RAND_704 = {1{`RANDOM}};
  s2_data_errors_1_4_REG_4_10 = _RAND_704[0:0];
  _RAND_705 = {1{`RANDOM}};
  s2_data_errors_1_4_REG_4_11 = _RAND_705[0:0];
  _RAND_706 = {1{`RANDOM}};
  s2_data_errors_1_4_REG_4_12 = _RAND_706[0:0];
  _RAND_707 = {1{`RANDOM}};
  s2_data_errors_1_4_REG_4_13 = _RAND_707[0:0];
  _RAND_708 = {1{`RANDOM}};
  s2_data_errors_1_4_REG_4_14 = _RAND_708[0:0];
  _RAND_709 = {1{`RANDOM}};
  s2_data_errors_1_4_REG_4_15 = _RAND_709[0:0];
  _RAND_710 = {1{`RANDOM}};
  s2_data_errors_1_4_REG_4_16 = _RAND_710[0:0];
  _RAND_711 = {1{`RANDOM}};
  s2_data_errors_1_4_REG_4_17 = _RAND_711[0:0];
  _RAND_712 = {1{`RANDOM}};
  s2_data_errors_1_4_REG_4_18 = _RAND_712[0:0];
  _RAND_713 = {1{`RANDOM}};
  s2_data_errors_1_4_REG_4_19 = _RAND_713[0:0];
  _RAND_714 = {1{`RANDOM}};
  s2_data_errors_1_4_REG_4_20 = _RAND_714[0:0];
  _RAND_715 = {1{`RANDOM}};
  s2_data_errors_1_4_REG_4_21 = _RAND_715[0:0];
  _RAND_716 = {1{`RANDOM}};
  s2_data_errors_1_4_REG_4_22 = _RAND_716[0:0];
  _RAND_717 = {1{`RANDOM}};
  s2_data_errors_1_4_REG_4_23 = _RAND_717[0:0];
  _RAND_718 = {1{`RANDOM}};
  s2_data_errors_1_4_REG_4_24 = _RAND_718[0:0];
  _RAND_719 = {1{`RANDOM}};
  s2_data_errors_1_4_REG_4_25 = _RAND_719[0:0];
  _RAND_720 = {1{`RANDOM}};
  s2_data_errors_1_4_REG_4_26 = _RAND_720[0:0];
  _RAND_721 = {1{`RANDOM}};
  s2_data_errors_1_4_REG_4_27 = _RAND_721[0:0];
  _RAND_722 = {1{`RANDOM}};
  s2_data_errors_1_4_REG_4_28 = _RAND_722[0:0];
  _RAND_723 = {1{`RANDOM}};
  s2_data_errors_1_4_REG_4_29 = _RAND_723[0:0];
  _RAND_724 = {1{`RANDOM}};
  s2_data_errors_1_4_REG_4_30 = _RAND_724[0:0];
  _RAND_725 = {1{`RANDOM}};
  s2_data_errors_1_4_REG_4_31 = _RAND_725[0:0];
  _RAND_726 = {1{`RANDOM}};
  s2_data_errors_1_5_REG = _RAND_726[0:0];
  _RAND_727 = {1{`RANDOM}};
  s2_data_errors_1_5_REG_1 = _RAND_727[0:0];
  _RAND_728 = {1{`RANDOM}};
  s2_data_errors_1_5_REG_2 = _RAND_728[0:0];
  _RAND_729 = {1{`RANDOM}};
  s2_data_errors_1_5_REG_3 = _RAND_729[0:0];
  _RAND_730 = {1{`RANDOM}};
  s2_data_errors_1_5_REG_4_0 = _RAND_730[0:0];
  _RAND_731 = {1{`RANDOM}};
  s2_data_errors_1_5_REG_4_1 = _RAND_731[0:0];
  _RAND_732 = {1{`RANDOM}};
  s2_data_errors_1_5_REG_4_2 = _RAND_732[0:0];
  _RAND_733 = {1{`RANDOM}};
  s2_data_errors_1_5_REG_4_3 = _RAND_733[0:0];
  _RAND_734 = {1{`RANDOM}};
  s2_data_errors_1_5_REG_4_4 = _RAND_734[0:0];
  _RAND_735 = {1{`RANDOM}};
  s2_data_errors_1_5_REG_4_5 = _RAND_735[0:0];
  _RAND_736 = {1{`RANDOM}};
  s2_data_errors_1_5_REG_4_6 = _RAND_736[0:0];
  _RAND_737 = {1{`RANDOM}};
  s2_data_errors_1_5_REG_4_7 = _RAND_737[0:0];
  _RAND_738 = {1{`RANDOM}};
  s2_data_errors_1_5_REG_4_8 = _RAND_738[0:0];
  _RAND_739 = {1{`RANDOM}};
  s2_data_errors_1_5_REG_4_9 = _RAND_739[0:0];
  _RAND_740 = {1{`RANDOM}};
  s2_data_errors_1_5_REG_4_10 = _RAND_740[0:0];
  _RAND_741 = {1{`RANDOM}};
  s2_data_errors_1_5_REG_4_11 = _RAND_741[0:0];
  _RAND_742 = {1{`RANDOM}};
  s2_data_errors_1_5_REG_4_12 = _RAND_742[0:0];
  _RAND_743 = {1{`RANDOM}};
  s2_data_errors_1_5_REG_4_13 = _RAND_743[0:0];
  _RAND_744 = {1{`RANDOM}};
  s2_data_errors_1_5_REG_4_14 = _RAND_744[0:0];
  _RAND_745 = {1{`RANDOM}};
  s2_data_errors_1_5_REG_4_15 = _RAND_745[0:0];
  _RAND_746 = {1{`RANDOM}};
  s2_data_errors_1_5_REG_4_16 = _RAND_746[0:0];
  _RAND_747 = {1{`RANDOM}};
  s2_data_errors_1_5_REG_4_17 = _RAND_747[0:0];
  _RAND_748 = {1{`RANDOM}};
  s2_data_errors_1_5_REG_4_18 = _RAND_748[0:0];
  _RAND_749 = {1{`RANDOM}};
  s2_data_errors_1_5_REG_4_19 = _RAND_749[0:0];
  _RAND_750 = {1{`RANDOM}};
  s2_data_errors_1_5_REG_4_20 = _RAND_750[0:0];
  _RAND_751 = {1{`RANDOM}};
  s2_data_errors_1_5_REG_4_21 = _RAND_751[0:0];
  _RAND_752 = {1{`RANDOM}};
  s2_data_errors_1_5_REG_4_22 = _RAND_752[0:0];
  _RAND_753 = {1{`RANDOM}};
  s2_data_errors_1_5_REG_4_23 = _RAND_753[0:0];
  _RAND_754 = {1{`RANDOM}};
  s2_data_errors_1_5_REG_4_24 = _RAND_754[0:0];
  _RAND_755 = {1{`RANDOM}};
  s2_data_errors_1_5_REG_4_25 = _RAND_755[0:0];
  _RAND_756 = {1{`RANDOM}};
  s2_data_errors_1_5_REG_4_26 = _RAND_756[0:0];
  _RAND_757 = {1{`RANDOM}};
  s2_data_errors_1_5_REG_4_27 = _RAND_757[0:0];
  _RAND_758 = {1{`RANDOM}};
  s2_data_errors_1_5_REG_4_28 = _RAND_758[0:0];
  _RAND_759 = {1{`RANDOM}};
  s2_data_errors_1_5_REG_4_29 = _RAND_759[0:0];
  _RAND_760 = {1{`RANDOM}};
  s2_data_errors_1_5_REG_4_30 = _RAND_760[0:0];
  _RAND_761 = {1{`RANDOM}};
  s2_data_errors_1_5_REG_4_31 = _RAND_761[0:0];
  _RAND_762 = {1{`RANDOM}};
  s2_data_errors_1_6_REG = _RAND_762[0:0];
  _RAND_763 = {1{`RANDOM}};
  s2_data_errors_1_6_REG_1 = _RAND_763[0:0];
  _RAND_764 = {1{`RANDOM}};
  s2_data_errors_1_6_REG_2 = _RAND_764[0:0];
  _RAND_765 = {1{`RANDOM}};
  s2_data_errors_1_6_REG_3 = _RAND_765[0:0];
  _RAND_766 = {1{`RANDOM}};
  s2_data_errors_1_6_REG_4_0 = _RAND_766[0:0];
  _RAND_767 = {1{`RANDOM}};
  s2_data_errors_1_6_REG_4_1 = _RAND_767[0:0];
  _RAND_768 = {1{`RANDOM}};
  s2_data_errors_1_6_REG_4_2 = _RAND_768[0:0];
  _RAND_769 = {1{`RANDOM}};
  s2_data_errors_1_6_REG_4_3 = _RAND_769[0:0];
  _RAND_770 = {1{`RANDOM}};
  s2_data_errors_1_6_REG_4_4 = _RAND_770[0:0];
  _RAND_771 = {1{`RANDOM}};
  s2_data_errors_1_6_REG_4_5 = _RAND_771[0:0];
  _RAND_772 = {1{`RANDOM}};
  s2_data_errors_1_6_REG_4_6 = _RAND_772[0:0];
  _RAND_773 = {1{`RANDOM}};
  s2_data_errors_1_6_REG_4_7 = _RAND_773[0:0];
  _RAND_774 = {1{`RANDOM}};
  s2_data_errors_1_6_REG_4_8 = _RAND_774[0:0];
  _RAND_775 = {1{`RANDOM}};
  s2_data_errors_1_6_REG_4_9 = _RAND_775[0:0];
  _RAND_776 = {1{`RANDOM}};
  s2_data_errors_1_6_REG_4_10 = _RAND_776[0:0];
  _RAND_777 = {1{`RANDOM}};
  s2_data_errors_1_6_REG_4_11 = _RAND_777[0:0];
  _RAND_778 = {1{`RANDOM}};
  s2_data_errors_1_6_REG_4_12 = _RAND_778[0:0];
  _RAND_779 = {1{`RANDOM}};
  s2_data_errors_1_6_REG_4_13 = _RAND_779[0:0];
  _RAND_780 = {1{`RANDOM}};
  s2_data_errors_1_6_REG_4_14 = _RAND_780[0:0];
  _RAND_781 = {1{`RANDOM}};
  s2_data_errors_1_6_REG_4_15 = _RAND_781[0:0];
  _RAND_782 = {1{`RANDOM}};
  s2_data_errors_1_6_REG_4_16 = _RAND_782[0:0];
  _RAND_783 = {1{`RANDOM}};
  s2_data_errors_1_6_REG_4_17 = _RAND_783[0:0];
  _RAND_784 = {1{`RANDOM}};
  s2_data_errors_1_6_REG_4_18 = _RAND_784[0:0];
  _RAND_785 = {1{`RANDOM}};
  s2_data_errors_1_6_REG_4_19 = _RAND_785[0:0];
  _RAND_786 = {1{`RANDOM}};
  s2_data_errors_1_6_REG_4_20 = _RAND_786[0:0];
  _RAND_787 = {1{`RANDOM}};
  s2_data_errors_1_6_REG_4_21 = _RAND_787[0:0];
  _RAND_788 = {1{`RANDOM}};
  s2_data_errors_1_6_REG_4_22 = _RAND_788[0:0];
  _RAND_789 = {1{`RANDOM}};
  s2_data_errors_1_6_REG_4_23 = _RAND_789[0:0];
  _RAND_790 = {1{`RANDOM}};
  s2_data_errors_1_6_REG_4_24 = _RAND_790[0:0];
  _RAND_791 = {1{`RANDOM}};
  s2_data_errors_1_6_REG_4_25 = _RAND_791[0:0];
  _RAND_792 = {1{`RANDOM}};
  s2_data_errors_1_6_REG_4_26 = _RAND_792[0:0];
  _RAND_793 = {1{`RANDOM}};
  s2_data_errors_1_6_REG_4_27 = _RAND_793[0:0];
  _RAND_794 = {1{`RANDOM}};
  s2_data_errors_1_6_REG_4_28 = _RAND_794[0:0];
  _RAND_795 = {1{`RANDOM}};
  s2_data_errors_1_6_REG_4_29 = _RAND_795[0:0];
  _RAND_796 = {1{`RANDOM}};
  s2_data_errors_1_6_REG_4_30 = _RAND_796[0:0];
  _RAND_797 = {1{`RANDOM}};
  s2_data_errors_1_6_REG_4_31 = _RAND_797[0:0];
  _RAND_798 = {1{`RANDOM}};
  s2_data_errors_1_7_REG = _RAND_798[0:0];
  _RAND_799 = {1{`RANDOM}};
  s2_data_errors_1_7_REG_1 = _RAND_799[0:0];
  _RAND_800 = {1{`RANDOM}};
  s2_data_errors_1_7_REG_2 = _RAND_800[0:0];
  _RAND_801 = {1{`RANDOM}};
  s2_data_errors_1_7_REG_3 = _RAND_801[0:0];
  _RAND_802 = {1{`RANDOM}};
  s2_data_errors_1_7_REG_4_0 = _RAND_802[0:0];
  _RAND_803 = {1{`RANDOM}};
  s2_data_errors_1_7_REG_4_1 = _RAND_803[0:0];
  _RAND_804 = {1{`RANDOM}};
  s2_data_errors_1_7_REG_4_2 = _RAND_804[0:0];
  _RAND_805 = {1{`RANDOM}};
  s2_data_errors_1_7_REG_4_3 = _RAND_805[0:0];
  _RAND_806 = {1{`RANDOM}};
  s2_data_errors_1_7_REG_4_4 = _RAND_806[0:0];
  _RAND_807 = {1{`RANDOM}};
  s2_data_errors_1_7_REG_4_5 = _RAND_807[0:0];
  _RAND_808 = {1{`RANDOM}};
  s2_data_errors_1_7_REG_4_6 = _RAND_808[0:0];
  _RAND_809 = {1{`RANDOM}};
  s2_data_errors_1_7_REG_4_7 = _RAND_809[0:0];
  _RAND_810 = {1{`RANDOM}};
  s2_data_errors_1_7_REG_4_8 = _RAND_810[0:0];
  _RAND_811 = {1{`RANDOM}};
  s2_data_errors_1_7_REG_4_9 = _RAND_811[0:0];
  _RAND_812 = {1{`RANDOM}};
  s2_data_errors_1_7_REG_4_10 = _RAND_812[0:0];
  _RAND_813 = {1{`RANDOM}};
  s2_data_errors_1_7_REG_4_11 = _RAND_813[0:0];
  _RAND_814 = {1{`RANDOM}};
  s2_data_errors_1_7_REG_4_12 = _RAND_814[0:0];
  _RAND_815 = {1{`RANDOM}};
  s2_data_errors_1_7_REG_4_13 = _RAND_815[0:0];
  _RAND_816 = {1{`RANDOM}};
  s2_data_errors_1_7_REG_4_14 = _RAND_816[0:0];
  _RAND_817 = {1{`RANDOM}};
  s2_data_errors_1_7_REG_4_15 = _RAND_817[0:0];
  _RAND_818 = {1{`RANDOM}};
  s2_data_errors_1_7_REG_4_16 = _RAND_818[0:0];
  _RAND_819 = {1{`RANDOM}};
  s2_data_errors_1_7_REG_4_17 = _RAND_819[0:0];
  _RAND_820 = {1{`RANDOM}};
  s2_data_errors_1_7_REG_4_18 = _RAND_820[0:0];
  _RAND_821 = {1{`RANDOM}};
  s2_data_errors_1_7_REG_4_19 = _RAND_821[0:0];
  _RAND_822 = {1{`RANDOM}};
  s2_data_errors_1_7_REG_4_20 = _RAND_822[0:0];
  _RAND_823 = {1{`RANDOM}};
  s2_data_errors_1_7_REG_4_21 = _RAND_823[0:0];
  _RAND_824 = {1{`RANDOM}};
  s2_data_errors_1_7_REG_4_22 = _RAND_824[0:0];
  _RAND_825 = {1{`RANDOM}};
  s2_data_errors_1_7_REG_4_23 = _RAND_825[0:0];
  _RAND_826 = {1{`RANDOM}};
  s2_data_errors_1_7_REG_4_24 = _RAND_826[0:0];
  _RAND_827 = {1{`RANDOM}};
  s2_data_errors_1_7_REG_4_25 = _RAND_827[0:0];
  _RAND_828 = {1{`RANDOM}};
  s2_data_errors_1_7_REG_4_26 = _RAND_828[0:0];
  _RAND_829 = {1{`RANDOM}};
  s2_data_errors_1_7_REG_4_27 = _RAND_829[0:0];
  _RAND_830 = {1{`RANDOM}};
  s2_data_errors_1_7_REG_4_28 = _RAND_830[0:0];
  _RAND_831 = {1{`RANDOM}};
  s2_data_errors_1_7_REG_4_29 = _RAND_831[0:0];
  _RAND_832 = {1{`RANDOM}};
  s2_data_errors_1_7_REG_4_30 = _RAND_832[0:0];
  _RAND_833 = {1{`RANDOM}};
  s2_data_errors_1_7_REG_4_31 = _RAND_833[0:0];
  _RAND_834 = {1{`RANDOM}};
  s2_parity_error_REG = _RAND_834[0:0];
  _RAND_835 = {1{`RANDOM}};
  s2_parity_error_REG_1 = _RAND_835[0:0];
  _RAND_836 = {1{`RANDOM}};
  io_errors_0_valid_REG = _RAND_836[0:0];
  _RAND_837 = {1{`RANDOM}};
  io_errors_0_valid_REG_1 = _RAND_837[0:0];
  _RAND_838 = {1{`RANDOM}};
  io_errors_0_valid_REG_2 = _RAND_838[0:0];
  _RAND_839 = {1{`RANDOM}};
  io_errors_0_report_to_beu_REG = _RAND_839[0:0];
  _RAND_840 = {1{`RANDOM}};
  io_errors_0_report_to_beu_REG_1 = _RAND_840[0:0];
  _RAND_841 = {1{`RANDOM}};
  io_errors_0_report_to_beu_REG_2 = _RAND_841[0:0];
  _RAND_842 = {2{`RANDOM}};
  io_errors_0_paddr_REG = _RAND_842[35:0];
  _RAND_843 = {2{`RANDOM}};
  io_errors_0_paddr_REG_1 = _RAND_843[35:0];
  _RAND_844 = {1{`RANDOM}};
  io_errors_0_source_tag_REG = _RAND_844[0:0];
  _RAND_845 = {1{`RANDOM}};
  io_errors_0_source_tag_REG_1 = _RAND_845[0:0];
  _RAND_846 = {1{`RANDOM}};
  io_errors_0_source_data_REG = _RAND_846[0:0];
  _RAND_847 = {1{`RANDOM}};
  io_errors_1_valid_REG = _RAND_847[0:0];
  _RAND_848 = {1{`RANDOM}};
  io_errors_1_valid_REG_1 = _RAND_848[0:0];
  _RAND_849 = {1{`RANDOM}};
  io_errors_1_valid_REG_2 = _RAND_849[0:0];
  _RAND_850 = {1{`RANDOM}};
  io_errors_1_report_to_beu_REG = _RAND_850[0:0];
  _RAND_851 = {1{`RANDOM}};
  io_errors_1_report_to_beu_REG_1 = _RAND_851[0:0];
  _RAND_852 = {1{`RANDOM}};
  io_errors_1_report_to_beu_REG_2 = _RAND_852[0:0];
  _RAND_853 = {2{`RANDOM}};
  io_errors_1_paddr_REG = _RAND_853[35:0];
  _RAND_854 = {2{`RANDOM}};
  io_errors_1_paddr_REG_1 = _RAND_854[35:0];
  _RAND_855 = {1{`RANDOM}};
  io_errors_1_source_tag_REG = _RAND_855[0:0];
  _RAND_856 = {1{`RANDOM}};
  io_errors_1_source_tag_REG_1 = _RAND_856[0:0];
  _RAND_857 = {1{`RANDOM}};
  io_errors_1_source_data_REG = _RAND_857[0:0];
  _RAND_858 = {1{`RANDOM}};
  s2_tlb_need_back_valid = _RAND_858[0:0];
  _RAND_859 = {1{`RANDOM}};
  s2_tlb_need_back_valid_1 = _RAND_859[0:0];
  _RAND_860 = {1{`RANDOM}};
  s2_except_pmp_af_REG = _RAND_860[0:0];
  _RAND_861 = {1{`RANDOM}};
  s2_except_pmp_af_r0 = _RAND_861[0:0];
  _RAND_862 = {1{`RANDOM}};
  s2_except_pmp_af_r1 = _RAND_862[0:0];
  _RAND_863 = {1{`RANDOM}};
  s2_mmio_REG = _RAND_863[0:0];
  _RAND_864 = {1{`RANDOM}};
  s2_mmio_r = _RAND_864[0:0];
  _RAND_865 = {1{`RANDOM}};
  missSlot_0_m_vSetIdx = _RAND_865[5:0];
  _RAND_866 = {1{`RANDOM}};
  missSlot_0_m_pTag = _RAND_866[23:0];
  _RAND_867 = {16{`RANDOM}};
  missSlot_0_m_data = _RAND_867[511:0];
  _RAND_868 = {1{`RANDOM}};
  missSlot_0_m_corrupt = _RAND_868[0:0];
  _RAND_869 = {1{`RANDOM}};
  missSlot_1_m_vSetIdx = _RAND_869[5:0];
  _RAND_870 = {1{`RANDOM}};
  missSlot_1_m_pTag = _RAND_870[23:0];
  _RAND_871 = {16{`RANDOM}};
  missSlot_1_m_data = _RAND_871[511:0];
  _RAND_872 = {1{`RANDOM}};
  missSlot_1_m_corrupt = _RAND_872[0:0];
  _RAND_873 = {1{`RANDOM}};
  only_0_miss_REG = _RAND_873[0:0];
  _RAND_874 = {1{`RANDOM}};
  only_0_hit_REG = _RAND_874[0:0];
  _RAND_875 = {1{`RANDOM}};
  hit_0_hit_1_REG = _RAND_875[0:0];
  _RAND_876 = {1{`RANDOM}};
  hit_0_miss_1_REG = _RAND_876[0:0];
  _RAND_877 = {1{`RANDOM}};
  miss_0_hit_1_REG = _RAND_877[0:0];
  _RAND_878 = {1{`RANDOM}};
  miss_0_miss_1_REG = _RAND_878[0:0];
  _RAND_879 = {1{`RANDOM}};
  miss_0_except_1_REG = _RAND_879[0:0];
  _RAND_880 = {1{`RANDOM}};
  miss_0_hit_1_latch_bit = _RAND_880[0:0];
  _RAND_881 = {1{`RANDOM}};
  miss_0_miss_1_latch_bit = _RAND_881[0:0];
  _RAND_882 = {1{`RANDOM}};
  only_0_miss_latch_bit = _RAND_882[0:0];
  _RAND_883 = {1{`RANDOM}};
  hit_0_miss_1_latch_bit = _RAND_883[0:0];
  _RAND_884 = {1{`RANDOM}};
  miss_0_except_1_latch_bit = _RAND_884[0:0];
  _RAND_885 = {1{`RANDOM}};
  only_0_hit_latch_bit = _RAND_885[0:0];
  _RAND_886 = {1{`RANDOM}};
  hit_0_hit_1_latch_bit = _RAND_886[0:0];
  _RAND_887 = {16{`RANDOM}};
  reservedRefillData_0_r = _RAND_887[511:0];
  _RAND_888 = {16{`RANDOM}};
  reservedRefillData_1_r = _RAND_888[511:0];
  _RAND_889 = {1{`RANDOM}};
  REG_8 = _RAND_889[0:0];
  _RAND_890 = {2{`RANDOM}};
  io_errors_0_paddr_REG_2 = _RAND_890[35:0];
  _RAND_891 = {1{`RANDOM}};
  REG_9 = _RAND_891[0:0];
  _RAND_892 = {2{`RANDOM}};
  io_errors_1_paddr_REG_2 = _RAND_892[35:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    missSwitchBit = 1'h0;
  end
  if (reset) begin
    s2_valid = 1'h0;
  end
  if (reset) begin
    miss_0_s2_0_latch_bit = 1'h0;
  end
  if (reset) begin
    missStateQueue_0 = 3'h0;
  end
  if (reset) begin
    miss_1_s2_0_latch_bit = 1'h0;
  end
  if (reset) begin
    missStateQueue_1 = 3'h0;
  end
  if (reset) begin
    miss_0_s2_1_latch_bit = 1'h0;
  end
  if (reset) begin
    miss_1_s2_1_latch_bit = 1'h0;
  end
  if (reset) begin
    wait_state = 4'h0;
  end
  if (reset) begin
    hit_0_except_1_latch_bit = 1'h0;
  end
  if (reset) begin
    except_0_latch_bit = 1'h0;
  end
  if (reset) begin
    tlb_need_back_valid = 1'h0;
  end
  if (reset) begin
    tlb_already_recv_0 = 1'h0;
  end
  if (reset) begin
    tlb_ready_recv_REG = 1'h0;
  end
  if (reset) begin
    s1_valid = 1'h0;
  end
  if (reset) begin
    tlb_need_back_valid_1 = 1'h0;
  end
  if (reset) begin
    tlb_already_recv_1 = 1'h0;
  end
  if (reset) begin
    tlb_ready_recv_REG_1 = 1'h0;
  end
  if (reset) begin
    state_vec__0 = 7'h0;
  end
  if (reset) begin
    state_vec__1 = 7'h0;
  end
  if (reset) begin
    state_vec__2 = 7'h0;
  end
  if (reset) begin
    state_vec__3 = 7'h0;
  end
  if (reset) begin
    state_vec__4 = 7'h0;
  end
  if (reset) begin
    state_vec__5 = 7'h0;
  end
  if (reset) begin
    state_vec__6 = 7'h0;
  end
  if (reset) begin
    state_vec__7 = 7'h0;
  end
  if (reset) begin
    state_vec__8 = 7'h0;
  end
  if (reset) begin
    state_vec__9 = 7'h0;
  end
  if (reset) begin
    state_vec__10 = 7'h0;
  end
  if (reset) begin
    state_vec__11 = 7'h0;
  end
  if (reset) begin
    state_vec__12 = 7'h0;
  end
  if (reset) begin
    state_vec__13 = 7'h0;
  end
  if (reset) begin
    state_vec__14 = 7'h0;
  end
  if (reset) begin
    state_vec__15 = 7'h0;
  end
  if (reset) begin
    state_vec__16 = 7'h0;
  end
  if (reset) begin
    state_vec__17 = 7'h0;
  end
  if (reset) begin
    state_vec__18 = 7'h0;
  end
  if (reset) begin
    state_vec__19 = 7'h0;
  end
  if (reset) begin
    state_vec__20 = 7'h0;
  end
  if (reset) begin
    state_vec__21 = 7'h0;
  end
  if (reset) begin
    state_vec__22 = 7'h0;
  end
  if (reset) begin
    state_vec__23 = 7'h0;
  end
  if (reset) begin
    state_vec__24 = 7'h0;
  end
  if (reset) begin
    state_vec__25 = 7'h0;
  end
  if (reset) begin
    state_vec__26 = 7'h0;
  end
  if (reset) begin
    state_vec__27 = 7'h0;
  end
  if (reset) begin
    state_vec__28 = 7'h0;
  end
  if (reset) begin
    state_vec__29 = 7'h0;
  end
  if (reset) begin
    state_vec__30 = 7'h0;
  end
  if (reset) begin
    state_vec__31 = 7'h0;
  end
  if (reset) begin
    state_vec_1_0 = 7'h0;
  end
  if (reset) begin
    state_vec_1_1 = 7'h0;
  end
  if (reset) begin
    state_vec_1_2 = 7'h0;
  end
  if (reset) begin
    state_vec_1_3 = 7'h0;
  end
  if (reset) begin
    state_vec_1_4 = 7'h0;
  end
  if (reset) begin
    state_vec_1_5 = 7'h0;
  end
  if (reset) begin
    state_vec_1_6 = 7'h0;
  end
  if (reset) begin
    state_vec_1_7 = 7'h0;
  end
  if (reset) begin
    state_vec_1_8 = 7'h0;
  end
  if (reset) begin
    state_vec_1_9 = 7'h0;
  end
  if (reset) begin
    state_vec_1_10 = 7'h0;
  end
  if (reset) begin
    state_vec_1_11 = 7'h0;
  end
  if (reset) begin
    state_vec_1_12 = 7'h0;
  end
  if (reset) begin
    state_vec_1_13 = 7'h0;
  end
  if (reset) begin
    state_vec_1_14 = 7'h0;
  end
  if (reset) begin
    state_vec_1_15 = 7'h0;
  end
  if (reset) begin
    state_vec_1_16 = 7'h0;
  end
  if (reset) begin
    state_vec_1_17 = 7'h0;
  end
  if (reset) begin
    state_vec_1_18 = 7'h0;
  end
  if (reset) begin
    state_vec_1_19 = 7'h0;
  end
  if (reset) begin
    state_vec_1_20 = 7'h0;
  end
  if (reset) begin
    state_vec_1_21 = 7'h0;
  end
  if (reset) begin
    state_vec_1_22 = 7'h0;
  end
  if (reset) begin
    state_vec_1_23 = 7'h0;
  end
  if (reset) begin
    state_vec_1_24 = 7'h0;
  end
  if (reset) begin
    state_vec_1_25 = 7'h0;
  end
  if (reset) begin
    state_vec_1_26 = 7'h0;
  end
  if (reset) begin
    state_vec_1_27 = 7'h0;
  end
  if (reset) begin
    state_vec_1_28 = 7'h0;
  end
  if (reset) begin
    state_vec_1_29 = 7'h0;
  end
  if (reset) begin
    state_vec_1_30 = 7'h0;
  end
  if (reset) begin
    state_vec_1_31 = 7'h0;
  end
  if (reset) begin
    s2_tlb_need_back_valid = 1'h0;
  end
  if (reset) begin
    s2_tlb_need_back_valid_1 = 1'h0;
  end
  if (reset) begin
    missSlot_0_m_vSetIdx = 6'h0;
  end
  if (reset) begin
    missSlot_0_m_pTag = 24'h0;
  end
  if (reset) begin
    missSlot_0_m_data = 512'h0;
  end
  if (reset) begin
    missSlot_0_m_corrupt = 1'h0;
  end
  if (reset) begin
    missSlot_1_m_vSetIdx = 6'h0;
  end
  if (reset) begin
    missSlot_1_m_pTag = 24'h0;
  end
  if (reset) begin
    missSlot_1_m_data = 512'h0;
  end
  if (reset) begin
    missSlot_1_m_corrupt = 1'h0;
  end
  if (reset) begin
    miss_0_hit_1_latch_bit = 1'h0;
  end
  if (reset) begin
    miss_0_miss_1_latch_bit = 1'h0;
  end
  if (reset) begin
    only_0_miss_latch_bit = 1'h0;
  end
  if (reset) begin
    hit_0_miss_1_latch_bit = 1'h0;
  end
  if (reset) begin
    miss_0_except_1_latch_bit = 1'h0;
  end
  if (reset) begin
    only_0_hit_latch_bit = 1'h0;
  end
  if (reset) begin
    hit_0_hit_1_latch_bit = 1'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule

