module CLZ_5(
  input  [107:0] io_in,
  output [6:0]   io_out
);
  wire [6:0] _io_out_T_108 = io_in[1] ? 7'h6a : 7'h6b; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_109 = io_in[2] ? 7'h69 : _io_out_T_108; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_110 = io_in[3] ? 7'h68 : _io_out_T_109; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_111 = io_in[4] ? 7'h67 : _io_out_T_110; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_112 = io_in[5] ? 7'h66 : _io_out_T_111; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_113 = io_in[6] ? 7'h65 : _io_out_T_112; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_114 = io_in[7] ? 7'h64 : _io_out_T_113; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_115 = io_in[8] ? 7'h63 : _io_out_T_114; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_116 = io_in[9] ? 7'h62 : _io_out_T_115; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_117 = io_in[10] ? 7'h61 : _io_out_T_116; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_118 = io_in[11] ? 7'h60 : _io_out_T_117; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_119 = io_in[12] ? 7'h5f : _io_out_T_118; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_120 = io_in[13] ? 7'h5e : _io_out_T_119; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_121 = io_in[14] ? 7'h5d : _io_out_T_120; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_122 = io_in[15] ? 7'h5c : _io_out_T_121; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_123 = io_in[16] ? 7'h5b : _io_out_T_122; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_124 = io_in[17] ? 7'h5a : _io_out_T_123; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_125 = io_in[18] ? 7'h59 : _io_out_T_124; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_126 = io_in[19] ? 7'h58 : _io_out_T_125; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_127 = io_in[20] ? 7'h57 : _io_out_T_126; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_128 = io_in[21] ? 7'h56 : _io_out_T_127; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_129 = io_in[22] ? 7'h55 : _io_out_T_128; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_130 = io_in[23] ? 7'h54 : _io_out_T_129; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_131 = io_in[24] ? 7'h53 : _io_out_T_130; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_132 = io_in[25] ? 7'h52 : _io_out_T_131; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_133 = io_in[26] ? 7'h51 : _io_out_T_132; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_134 = io_in[27] ? 7'h50 : _io_out_T_133; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_135 = io_in[28] ? 7'h4f : _io_out_T_134; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_136 = io_in[29] ? 7'h4e : _io_out_T_135; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_137 = io_in[30] ? 7'h4d : _io_out_T_136; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_138 = io_in[31] ? 7'h4c : _io_out_T_137; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_139 = io_in[32] ? 7'h4b : _io_out_T_138; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_140 = io_in[33] ? 7'h4a : _io_out_T_139; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_141 = io_in[34] ? 7'h49 : _io_out_T_140; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_142 = io_in[35] ? 7'h48 : _io_out_T_141; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_143 = io_in[36] ? 7'h47 : _io_out_T_142; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_144 = io_in[37] ? 7'h46 : _io_out_T_143; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_145 = io_in[38] ? 7'h45 : _io_out_T_144; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_146 = io_in[39] ? 7'h44 : _io_out_T_145; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_147 = io_in[40] ? 7'h43 : _io_out_T_146; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_148 = io_in[41] ? 7'h42 : _io_out_T_147; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_149 = io_in[42] ? 7'h41 : _io_out_T_148; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_150 = io_in[43] ? 7'h40 : _io_out_T_149; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_151 = io_in[44] ? 7'h3f : _io_out_T_150; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_152 = io_in[45] ? 7'h3e : _io_out_T_151; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_153 = io_in[46] ? 7'h3d : _io_out_T_152; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_154 = io_in[47] ? 7'h3c : _io_out_T_153; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_155 = io_in[48] ? 7'h3b : _io_out_T_154; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_156 = io_in[49] ? 7'h3a : _io_out_T_155; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_157 = io_in[50] ? 7'h39 : _io_out_T_156; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_158 = io_in[51] ? 7'h38 : _io_out_T_157; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_159 = io_in[52] ? 7'h37 : _io_out_T_158; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_160 = io_in[53] ? 7'h36 : _io_out_T_159; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_161 = io_in[54] ? 7'h35 : _io_out_T_160; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_162 = io_in[55] ? 7'h34 : _io_out_T_161; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_163 = io_in[56] ? 7'h33 : _io_out_T_162; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_164 = io_in[57] ? 7'h32 : _io_out_T_163; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_165 = io_in[58] ? 7'h31 : _io_out_T_164; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_166 = io_in[59] ? 7'h30 : _io_out_T_165; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_167 = io_in[60] ? 7'h2f : _io_out_T_166; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_168 = io_in[61] ? 7'h2e : _io_out_T_167; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_169 = io_in[62] ? 7'h2d : _io_out_T_168; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_170 = io_in[63] ? 7'h2c : _io_out_T_169; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_171 = io_in[64] ? 7'h2b : _io_out_T_170; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_172 = io_in[65] ? 7'h2a : _io_out_T_171; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_173 = io_in[66] ? 7'h29 : _io_out_T_172; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_174 = io_in[67] ? 7'h28 : _io_out_T_173; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_175 = io_in[68] ? 7'h27 : _io_out_T_174; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_176 = io_in[69] ? 7'h26 : _io_out_T_175; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_177 = io_in[70] ? 7'h25 : _io_out_T_176; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_178 = io_in[71] ? 7'h24 : _io_out_T_177; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_179 = io_in[72] ? 7'h23 : _io_out_T_178; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_180 = io_in[73] ? 7'h22 : _io_out_T_179; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_181 = io_in[74] ? 7'h21 : _io_out_T_180; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_182 = io_in[75] ? 7'h20 : _io_out_T_181; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_183 = io_in[76] ? 7'h1f : _io_out_T_182; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_184 = io_in[77] ? 7'h1e : _io_out_T_183; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_185 = io_in[78] ? 7'h1d : _io_out_T_184; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_186 = io_in[79] ? 7'h1c : _io_out_T_185; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_187 = io_in[80] ? 7'h1b : _io_out_T_186; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_188 = io_in[81] ? 7'h1a : _io_out_T_187; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_189 = io_in[82] ? 7'h19 : _io_out_T_188; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_190 = io_in[83] ? 7'h18 : _io_out_T_189; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_191 = io_in[84] ? 7'h17 : _io_out_T_190; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_192 = io_in[85] ? 7'h16 : _io_out_T_191; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_193 = io_in[86] ? 7'h15 : _io_out_T_192; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_194 = io_in[87] ? 7'h14 : _io_out_T_193; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_195 = io_in[88] ? 7'h13 : _io_out_T_194; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_196 = io_in[89] ? 7'h12 : _io_out_T_195; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_197 = io_in[90] ? 7'h11 : _io_out_T_196; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_198 = io_in[91] ? 7'h10 : _io_out_T_197; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_199 = io_in[92] ? 7'hf : _io_out_T_198; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_200 = io_in[93] ? 7'he : _io_out_T_199; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_201 = io_in[94] ? 7'hd : _io_out_T_200; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_202 = io_in[95] ? 7'hc : _io_out_T_201; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_203 = io_in[96] ? 7'hb : _io_out_T_202; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_204 = io_in[97] ? 7'ha : _io_out_T_203; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_205 = io_in[98] ? 7'h9 : _io_out_T_204; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_206 = io_in[99] ? 7'h8 : _io_out_T_205; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_207 = io_in[100] ? 7'h7 : _io_out_T_206; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_208 = io_in[101] ? 7'h6 : _io_out_T_207; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_209 = io_in[102] ? 7'h5 : _io_out_T_208; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_210 = io_in[103] ? 7'h4 : _io_out_T_209; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_211 = io_in[104] ? 7'h3 : _io_out_T_210; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_212 = io_in[105] ? 7'h2 : _io_out_T_211; // @[Mux.scala 47:70]
  wire [6:0] _io_out_T_213 = io_in[106] ? 7'h1 : _io_out_T_212; // @[Mux.scala 47:70]
  assign io_out = io_in[107] ? 7'h0 : _io_out_T_213; // @[Mux.scala 47:70]
endmodule

