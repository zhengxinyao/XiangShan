module DelayN_46(
  input  [35:0] io_in,
  output [35:0] io_out
);
  assign io_out = io_in; // @[Hold.scala 92:10]
endmodule

