module bosc_CtrlBlock(
  input         clock,
  input         reset,
  input  [7:0]  io_hartId,
  output        io_cpu_halt,
  output        io_frontend_cfVec_0_ready,
  input         io_frontend_cfVec_0_valid,
  input  [31:0] io_frontend_cfVec_0_bits_instr,
  input  [9:0]  io_frontend_cfVec_0_bits_foldpc,
  input         io_frontend_cfVec_0_bits_exceptionVec_1,
  input         io_frontend_cfVec_0_bits_exceptionVec_12,
  input         io_frontend_cfVec_0_bits_trigger_frontendHit_0,
  input         io_frontend_cfVec_0_bits_trigger_frontendHit_1,
  input         io_frontend_cfVec_0_bits_trigger_frontendHit_2,
  input         io_frontend_cfVec_0_bits_trigger_frontendHit_3,
  input         io_frontend_cfVec_0_bits_trigger_backendEn_0,
  input         io_frontend_cfVec_0_bits_trigger_backendEn_1,
  input         io_frontend_cfVec_0_bits_pd_isRVC,
  input  [1:0]  io_frontend_cfVec_0_bits_pd_brType,
  input         io_frontend_cfVec_0_bits_pd_isCall,
  input         io_frontend_cfVec_0_bits_pd_isRet,
  input         io_frontend_cfVec_0_bits_pred_taken,
  input         io_frontend_cfVec_0_bits_crossPageIPFFix,
  input         io_frontend_cfVec_0_bits_ftqPtr_flag,
  input  [2:0]  io_frontend_cfVec_0_bits_ftqPtr_value,
  input  [2:0]  io_frontend_cfVec_0_bits_ftqOffset,
  output        io_frontend_cfVec_1_ready,
  input         io_frontend_cfVec_1_valid,
  input  [31:0] io_frontend_cfVec_1_bits_instr,
  input  [9:0]  io_frontend_cfVec_1_bits_foldpc,
  input         io_frontend_cfVec_1_bits_exceptionVec_1,
  input         io_frontend_cfVec_1_bits_exceptionVec_12,
  input         io_frontend_cfVec_1_bits_trigger_frontendHit_0,
  input         io_frontend_cfVec_1_bits_trigger_frontendHit_1,
  input         io_frontend_cfVec_1_bits_trigger_frontendHit_2,
  input         io_frontend_cfVec_1_bits_trigger_frontendHit_3,
  input         io_frontend_cfVec_1_bits_trigger_backendEn_0,
  input         io_frontend_cfVec_1_bits_trigger_backendEn_1,
  input         io_frontend_cfVec_1_bits_pd_isRVC,
  input  [1:0]  io_frontend_cfVec_1_bits_pd_brType,
  input         io_frontend_cfVec_1_bits_pd_isCall,
  input         io_frontend_cfVec_1_bits_pd_isRet,
  input         io_frontend_cfVec_1_bits_pred_taken,
  input         io_frontend_cfVec_1_bits_crossPageIPFFix,
  input         io_frontend_cfVec_1_bits_ftqPtr_flag,
  input  [2:0]  io_frontend_cfVec_1_bits_ftqPtr_value,
  input  [2:0]  io_frontend_cfVec_1_bits_ftqOffset,
  input         io_frontend_fromFtq_pc_mem_wen,
  input  [2:0]  io_frontend_fromFtq_pc_mem_waddr,
  input  [38:0] io_frontend_fromFtq_pc_mem_wdata_startAddr,
  input  [38:0] io_frontend_fromFtq_pc_mem_wdata_nextLineAddr,
  input         io_frontend_fromFtq_pc_mem_wdata_isNextMask_0,
  input         io_frontend_fromFtq_pc_mem_wdata_isNextMask_1,
  input         io_frontend_fromFtq_pc_mem_wdata_isNextMask_2,
  input         io_frontend_fromFtq_pc_mem_wdata_isNextMask_3,
  input         io_frontend_fromFtq_pc_mem_wdata_isNextMask_4,
  input         io_frontend_fromFtq_pc_mem_wdata_isNextMask_5,
  input         io_frontend_fromFtq_pc_mem_wdata_isNextMask_6,
  input         io_frontend_fromFtq_pc_mem_wdata_isNextMask_7,
  input  [38:0] io_frontend_fromFtq_newest_entry_target,
  input         io_frontend_fromFtq_newest_entry_ptr_flag,
  input  [2:0]  io_frontend_fromFtq_newest_entry_ptr_value,
  output        io_frontend_toFtq_rob_commits_0_valid,
  output [2:0]  io_frontend_toFtq_rob_commits_0_bits_commitType,
  output        io_frontend_toFtq_rob_commits_0_bits_ftqIdx_flag,
  output [2:0]  io_frontend_toFtq_rob_commits_0_bits_ftqIdx_value,
  output [2:0]  io_frontend_toFtq_rob_commits_0_bits_ftqOffset,
  output        io_frontend_toFtq_rob_commits_1_valid,
  output [2:0]  io_frontend_toFtq_rob_commits_1_bits_commitType,
  output        io_frontend_toFtq_rob_commits_1_bits_ftqIdx_flag,
  output [2:0]  io_frontend_toFtq_rob_commits_1_bits_ftqIdx_value,
  output [2:0]  io_frontend_toFtq_rob_commits_1_bits_ftqOffset,
  output        io_frontend_toFtq_redirect_valid,
  output        io_frontend_toFtq_redirect_bits_ftqIdx_flag,
  output [2:0]  io_frontend_toFtq_redirect_bits_ftqIdx_value,
  output [2:0]  io_frontend_toFtq_redirect_bits_ftqOffset,
  output        io_frontend_toFtq_redirect_bits_level,
  output [38:0] io_frontend_toFtq_redirect_bits_cfiUpdate_pc,
  output        io_frontend_toFtq_redirect_bits_cfiUpdate_pd_isRVC,
  output [1:0]  io_frontend_toFtq_redirect_bits_cfiUpdate_pd_brType,
  output        io_frontend_toFtq_redirect_bits_cfiUpdate_pd_isCall,
  output        io_frontend_toFtq_redirect_bits_cfiUpdate_pd_isRet,
  output [38:0] io_frontend_toFtq_redirect_bits_cfiUpdate_target,
  output        io_frontend_toFtq_redirect_bits_cfiUpdate_taken,
  output        io_frontend_toFtq_redirect_bits_cfiUpdate_isMisPred,
  output        io_allocPregs_0_isInt,
  output        io_allocPregs_0_isFp,
  output [5:0]  io_allocPregs_0_preg,
  output        io_allocPregs_1_isInt,
  output        io_allocPregs_1_isFp,
  output [5:0]  io_allocPregs_1_preg,
  output        io_dispatch_0_valid,
  output [9:0]  io_dispatch_0_bits_cf_foldpc,
  output        io_dispatch_0_bits_cf_trigger_backendEn_0,
  output        io_dispatch_0_bits_cf_trigger_backendEn_1,
  output        io_dispatch_0_bits_cf_pd_isRVC,
  output [1:0]  io_dispatch_0_bits_cf_pd_brType,
  output        io_dispatch_0_bits_cf_pd_isCall,
  output        io_dispatch_0_bits_cf_pd_isRet,
  output        io_dispatch_0_bits_cf_pred_taken,
  output        io_dispatch_0_bits_cf_storeSetHit,
  output        io_dispatch_0_bits_cf_waitForRobIdx_flag,
  output [4:0]  io_dispatch_0_bits_cf_waitForRobIdx_value,
  output        io_dispatch_0_bits_cf_loadWaitBit,
  output        io_dispatch_0_bits_cf_loadWaitStrict,
  output [4:0]  io_dispatch_0_bits_cf_ssid,
  output        io_dispatch_0_bits_cf_ftqPtr_flag,
  output [2:0]  io_dispatch_0_bits_cf_ftqPtr_value,
  output [2:0]  io_dispatch_0_bits_cf_ftqOffset,
  output [1:0]  io_dispatch_0_bits_ctrl_srcType_0,
  output [1:0]  io_dispatch_0_bits_ctrl_srcType_1,
  output [3:0]  io_dispatch_0_bits_ctrl_fuType,
  output [6:0]  io_dispatch_0_bits_ctrl_fuOpType,
  output        io_dispatch_0_bits_ctrl_rfWen,
  output        io_dispatch_0_bits_ctrl_fpWen,
  output [3:0]  io_dispatch_0_bits_ctrl_selImm,
  output [19:0] io_dispatch_0_bits_ctrl_imm,
  output        io_dispatch_0_bits_ctrl_fpu_isAddSub,
  output        io_dispatch_0_bits_ctrl_fpu_typeTagIn,
  output        io_dispatch_0_bits_ctrl_fpu_typeTagOut,
  output        io_dispatch_0_bits_ctrl_fpu_fromInt,
  output        io_dispatch_0_bits_ctrl_fpu_wflags,
  output        io_dispatch_0_bits_ctrl_fpu_fpWen,
  output [1:0]  io_dispatch_0_bits_ctrl_fpu_fmaCmd,
  output        io_dispatch_0_bits_ctrl_fpu_div,
  output        io_dispatch_0_bits_ctrl_fpu_sqrt,
  output        io_dispatch_0_bits_ctrl_fpu_fcvt,
  output [1:0]  io_dispatch_0_bits_ctrl_fpu_typ,
  output [1:0]  io_dispatch_0_bits_ctrl_fpu_fmt,
  output        io_dispatch_0_bits_ctrl_fpu_ren3,
  output [2:0]  io_dispatch_0_bits_ctrl_fpu_rm,
  output [5:0]  io_dispatch_0_bits_psrc_0,
  output [5:0]  io_dispatch_0_bits_psrc_1,
  output [5:0]  io_dispatch_0_bits_pdest,
  output        io_dispatch_0_bits_robIdx_flag,
  output [4:0]  io_dispatch_0_bits_robIdx_value,
  output        io_dispatch_0_bits_lqIdx_flag,
  output [3:0]  io_dispatch_0_bits_lqIdx_value,
  output        io_dispatch_0_bits_sqIdx_flag,
  output [3:0]  io_dispatch_0_bits_sqIdx_value,
  output        io_dispatch_1_valid,
  output [9:0]  io_dispatch_1_bits_cf_foldpc,
  output        io_dispatch_1_bits_cf_trigger_backendEn_0,
  output        io_dispatch_1_bits_cf_trigger_backendEn_1,
  output        io_dispatch_1_bits_cf_pd_isRVC,
  output [1:0]  io_dispatch_1_bits_cf_pd_brType,
  output        io_dispatch_1_bits_cf_pd_isCall,
  output        io_dispatch_1_bits_cf_pd_isRet,
  output        io_dispatch_1_bits_cf_pred_taken,
  output        io_dispatch_1_bits_cf_storeSetHit,
  output        io_dispatch_1_bits_cf_waitForRobIdx_flag,
  output [4:0]  io_dispatch_1_bits_cf_waitForRobIdx_value,
  output        io_dispatch_1_bits_cf_loadWaitBit,
  output        io_dispatch_1_bits_cf_loadWaitStrict,
  output [4:0]  io_dispatch_1_bits_cf_ssid,
  output        io_dispatch_1_bits_cf_ftqPtr_flag,
  output [2:0]  io_dispatch_1_bits_cf_ftqPtr_value,
  output [2:0]  io_dispatch_1_bits_cf_ftqOffset,
  output [1:0]  io_dispatch_1_bits_ctrl_srcType_0,
  output [1:0]  io_dispatch_1_bits_ctrl_srcType_1,
  output [3:0]  io_dispatch_1_bits_ctrl_fuType,
  output [6:0]  io_dispatch_1_bits_ctrl_fuOpType,
  output        io_dispatch_1_bits_ctrl_rfWen,
  output        io_dispatch_1_bits_ctrl_fpWen,
  output [3:0]  io_dispatch_1_bits_ctrl_selImm,
  output [19:0] io_dispatch_1_bits_ctrl_imm,
  output [5:0]  io_dispatch_1_bits_psrc_0,
  output [5:0]  io_dispatch_1_bits_psrc_1,
  output [5:0]  io_dispatch_1_bits_pdest,
  output        io_dispatch_1_bits_robIdx_flag,
  output [4:0]  io_dispatch_1_bits_robIdx_value,
  output        io_dispatch_1_bits_lqIdx_flag,
  output [3:0]  io_dispatch_1_bits_lqIdx_value,
  output        io_dispatch_1_bits_sqIdx_flag,
  output [3:0]  io_dispatch_1_bits_sqIdx_value,
  output        io_dispatch_4_valid,
  output [9:0]  io_dispatch_4_bits_cf_foldpc,
  output        io_dispatch_4_bits_cf_trigger_backendEn_0,
  output        io_dispatch_4_bits_cf_trigger_backendEn_1,
  output        io_dispatch_4_bits_cf_pd_isRVC,
  output [1:0]  io_dispatch_4_bits_cf_pd_brType,
  output        io_dispatch_4_bits_cf_pd_isCall,
  output        io_dispatch_4_bits_cf_pd_isRet,
  output        io_dispatch_4_bits_cf_pred_taken,
  output        io_dispatch_4_bits_cf_storeSetHit,
  output        io_dispatch_4_bits_cf_waitForRobIdx_flag,
  output [4:0]  io_dispatch_4_bits_cf_waitForRobIdx_value,
  output        io_dispatch_4_bits_cf_loadWaitBit,
  output        io_dispatch_4_bits_cf_loadWaitStrict,
  output [4:0]  io_dispatch_4_bits_cf_ssid,
  output        io_dispatch_4_bits_cf_ftqPtr_flag,
  output [2:0]  io_dispatch_4_bits_cf_ftqPtr_value,
  output [2:0]  io_dispatch_4_bits_cf_ftqOffset,
  output [1:0]  io_dispatch_4_bits_ctrl_srcType_0,
  output [1:0]  io_dispatch_4_bits_ctrl_srcType_1,
  output [3:0]  io_dispatch_4_bits_ctrl_fuType,
  output [6:0]  io_dispatch_4_bits_ctrl_fuOpType,
  output        io_dispatch_4_bits_ctrl_rfWen,
  output        io_dispatch_4_bits_ctrl_fpWen,
  output        io_dispatch_4_bits_ctrl_flushPipe,
  output [19:0] io_dispatch_4_bits_ctrl_imm,
  output        io_dispatch_4_bits_ctrl_replayInst,
  output [5:0]  io_dispatch_4_bits_psrc_0,
  output [5:0]  io_dispatch_4_bits_psrc_1,
  output [5:0]  io_dispatch_4_bits_pdest,
  output        io_dispatch_4_bits_robIdx_flag,
  output [4:0]  io_dispatch_4_bits_robIdx_value,
  output        io_dispatch_5_valid,
  output [9:0]  io_dispatch_5_bits_cf_foldpc,
  output        io_dispatch_5_bits_cf_trigger_backendEn_0,
  output        io_dispatch_5_bits_cf_trigger_backendEn_1,
  output        io_dispatch_5_bits_cf_pd_isRVC,
  output [1:0]  io_dispatch_5_bits_cf_pd_brType,
  output        io_dispatch_5_bits_cf_pd_isCall,
  output        io_dispatch_5_bits_cf_pd_isRet,
  output        io_dispatch_5_bits_cf_pred_taken,
  output        io_dispatch_5_bits_cf_storeSetHit,
  output        io_dispatch_5_bits_cf_waitForRobIdx_flag,
  output [4:0]  io_dispatch_5_bits_cf_waitForRobIdx_value,
  output        io_dispatch_5_bits_cf_loadWaitBit,
  output        io_dispatch_5_bits_cf_loadWaitStrict,
  output [4:0]  io_dispatch_5_bits_cf_ssid,
  output        io_dispatch_5_bits_cf_ftqPtr_flag,
  output [2:0]  io_dispatch_5_bits_cf_ftqPtr_value,
  output [2:0]  io_dispatch_5_bits_cf_ftqOffset,
  output [1:0]  io_dispatch_5_bits_ctrl_srcType_0,
  output [1:0]  io_dispatch_5_bits_ctrl_srcType_1,
  output [3:0]  io_dispatch_5_bits_ctrl_fuType,
  output [6:0]  io_dispatch_5_bits_ctrl_fuOpType,
  output        io_dispatch_5_bits_ctrl_rfWen,
  output        io_dispatch_5_bits_ctrl_fpWen,
  output        io_dispatch_5_bits_ctrl_flushPipe,
  output [19:0] io_dispatch_5_bits_ctrl_imm,
  output        io_dispatch_5_bits_ctrl_replayInst,
  output [5:0]  io_dispatch_5_bits_psrc_0,
  output [5:0]  io_dispatch_5_bits_psrc_1,
  output [5:0]  io_dispatch_5_bits_pdest,
  output        io_dispatch_5_bits_robIdx_flag,
  output [4:0]  io_dispatch_5_bits_robIdx_value,
  output        io_dispatch_6_valid,
  output [9:0]  io_dispatch_6_bits_cf_foldpc,
  output        io_dispatch_6_bits_cf_trigger_backendEn_0,
  output        io_dispatch_6_bits_cf_trigger_backendEn_1,
  output        io_dispatch_6_bits_cf_pd_isRVC,
  output [1:0]  io_dispatch_6_bits_cf_pd_brType,
  output        io_dispatch_6_bits_cf_pd_isCall,
  output        io_dispatch_6_bits_cf_pd_isRet,
  output        io_dispatch_6_bits_cf_pred_taken,
  output        io_dispatch_6_bits_cf_storeSetHit,
  output        io_dispatch_6_bits_cf_waitForRobIdx_flag,
  output [4:0]  io_dispatch_6_bits_cf_waitForRobIdx_value,
  output        io_dispatch_6_bits_cf_loadWaitBit,
  output        io_dispatch_6_bits_cf_loadWaitStrict,
  output [4:0]  io_dispatch_6_bits_cf_ssid,
  output        io_dispatch_6_bits_cf_ftqPtr_flag,
  output [2:0]  io_dispatch_6_bits_cf_ftqPtr_value,
  output [2:0]  io_dispatch_6_bits_cf_ftqOffset,
  output [1:0]  io_dispatch_6_bits_ctrl_srcType_0,
  output [1:0]  io_dispatch_6_bits_ctrl_srcType_1,
  output [3:0]  io_dispatch_6_bits_ctrl_fuType,
  output [6:0]  io_dispatch_6_bits_ctrl_fuOpType,
  output        io_dispatch_6_bits_ctrl_rfWen,
  output        io_dispatch_6_bits_ctrl_fpWen,
  output        io_dispatch_6_bits_ctrl_flushPipe,
  output [19:0] io_dispatch_6_bits_ctrl_imm,
  output        io_dispatch_6_bits_ctrl_replayInst,
  output [5:0]  io_dispatch_6_bits_psrc_0,
  output [5:0]  io_dispatch_6_bits_psrc_1,
  output [5:0]  io_dispatch_6_bits_pdest,
  output        io_dispatch_6_bits_robIdx_flag,
  output [4:0]  io_dispatch_6_bits_robIdx_value,
  output        io_dispatch_7_valid,
  output [9:0]  io_dispatch_7_bits_cf_foldpc,
  output        io_dispatch_7_bits_cf_trigger_backendEn_0,
  output        io_dispatch_7_bits_cf_trigger_backendEn_1,
  output        io_dispatch_7_bits_cf_pd_isRVC,
  output [1:0]  io_dispatch_7_bits_cf_pd_brType,
  output        io_dispatch_7_bits_cf_pd_isCall,
  output        io_dispatch_7_bits_cf_pd_isRet,
  output        io_dispatch_7_bits_cf_pred_taken,
  output        io_dispatch_7_bits_cf_storeSetHit,
  output        io_dispatch_7_bits_cf_waitForRobIdx_flag,
  output [4:0]  io_dispatch_7_bits_cf_waitForRobIdx_value,
  output        io_dispatch_7_bits_cf_loadWaitBit,
  output        io_dispatch_7_bits_cf_loadWaitStrict,
  output [4:0]  io_dispatch_7_bits_cf_ssid,
  output        io_dispatch_7_bits_cf_ftqPtr_flag,
  output [2:0]  io_dispatch_7_bits_cf_ftqPtr_value,
  output [2:0]  io_dispatch_7_bits_cf_ftqOffset,
  output [1:0]  io_dispatch_7_bits_ctrl_srcType_0,
  output [1:0]  io_dispatch_7_bits_ctrl_srcType_1,
  output [3:0]  io_dispatch_7_bits_ctrl_fuType,
  output [6:0]  io_dispatch_7_bits_ctrl_fuOpType,
  output        io_dispatch_7_bits_ctrl_rfWen,
  output        io_dispatch_7_bits_ctrl_fpWen,
  output        io_dispatch_7_bits_ctrl_flushPipe,
  output [19:0] io_dispatch_7_bits_ctrl_imm,
  output        io_dispatch_7_bits_ctrl_replayInst,
  output [5:0]  io_dispatch_7_bits_psrc_0,
  output [5:0]  io_dispatch_7_bits_psrc_1,
  output [5:0]  io_dispatch_7_bits_pdest,
  output        io_dispatch_7_bits_robIdx_flag,
  output [4:0]  io_dispatch_7_bits_robIdx_value,
  output        io_dispatch_8_valid,
  output        io_dispatch_8_bits_cf_pd_isRVC,
  output [1:0]  io_dispatch_8_bits_cf_pd_brType,
  output        io_dispatch_8_bits_cf_pd_isCall,
  output        io_dispatch_8_bits_cf_pd_isRet,
  output        io_dispatch_8_bits_cf_pred_taken,
  output        io_dispatch_8_bits_cf_ftqPtr_flag,
  output [2:0]  io_dispatch_8_bits_cf_ftqPtr_value,
  output [2:0]  io_dispatch_8_bits_cf_ftqOffset,
  output [1:0]  io_dispatch_8_bits_ctrl_srcType_0,
  output [1:0]  io_dispatch_8_bits_ctrl_srcType_1,
  output [1:0]  io_dispatch_8_bits_ctrl_srcType_2,
  output [3:0]  io_dispatch_8_bits_ctrl_fuType,
  output [6:0]  io_dispatch_8_bits_ctrl_fuOpType,
  output        io_dispatch_8_bits_ctrl_rfWen,
  output        io_dispatch_8_bits_ctrl_fpWen,
  output [19:0] io_dispatch_8_bits_ctrl_imm,
  output        io_dispatch_8_bits_ctrl_fpu_isAddSub,
  output        io_dispatch_8_bits_ctrl_fpu_typeTagIn,
  output        io_dispatch_8_bits_ctrl_fpu_typeTagOut,
  output        io_dispatch_8_bits_ctrl_fpu_fromInt,
  output        io_dispatch_8_bits_ctrl_fpu_wflags,
  output        io_dispatch_8_bits_ctrl_fpu_fpWen,
  output [1:0]  io_dispatch_8_bits_ctrl_fpu_fmaCmd,
  output        io_dispatch_8_bits_ctrl_fpu_div,
  output        io_dispatch_8_bits_ctrl_fpu_sqrt,
  output        io_dispatch_8_bits_ctrl_fpu_fcvt,
  output [1:0]  io_dispatch_8_bits_ctrl_fpu_typ,
  output [1:0]  io_dispatch_8_bits_ctrl_fpu_fmt,
  output        io_dispatch_8_bits_ctrl_fpu_ren3,
  output [2:0]  io_dispatch_8_bits_ctrl_fpu_rm,
  output [5:0]  io_dispatch_8_bits_psrc_0,
  output [5:0]  io_dispatch_8_bits_psrc_1,
  output [5:0]  io_dispatch_8_bits_psrc_2,
  output [5:0]  io_dispatch_8_bits_pdest,
  output        io_dispatch_8_bits_robIdx_flag,
  output [4:0]  io_dispatch_8_bits_robIdx_value,
  input         io_rsReady_0,
  input         io_rsReady_1,
  input         io_rsReady_2,
  input         io_rsReady_3,
  input         io_rsReady_4,
  input         io_rsReady_5,
  input         io_rsReady_6,
  input         io_rsReady_7,
  input         io_rsReady_8,
  output [1:0]  io_enqLsq_needAlloc_0,
  output [1:0]  io_enqLsq_needAlloc_1,
  output [1:0]  io_enqLsq_needAlloc_2,
  output [1:0]  io_enqLsq_needAlloc_3,
  output        io_enqLsq_req_0_valid,
  output        io_enqLsq_req_0_bits_cf_trigger_backendEn_0,
  output        io_enqLsq_req_0_bits_cf_trigger_backendEn_1,
  output [6:0]  io_enqLsq_req_0_bits_ctrl_fuOpType,
  output        io_enqLsq_req_0_bits_ctrl_rfWen,
  output        io_enqLsq_req_0_bits_ctrl_fpWen,
  output        io_enqLsq_req_0_bits_ctrl_flushPipe,
  output        io_enqLsq_req_0_bits_ctrl_replayInst,
  output [5:0]  io_enqLsq_req_0_bits_pdest,
  output        io_enqLsq_req_0_bits_robIdx_flag,
  output [4:0]  io_enqLsq_req_0_bits_robIdx_value,
  output [3:0]  io_enqLsq_req_0_bits_lqIdx_value,
  output [3:0]  io_enqLsq_req_0_bits_sqIdx_value,
  output        io_enqLsq_req_1_valid,
  output        io_enqLsq_req_1_bits_cf_trigger_backendEn_0,
  output        io_enqLsq_req_1_bits_cf_trigger_backendEn_1,
  output [6:0]  io_enqLsq_req_1_bits_ctrl_fuOpType,
  output        io_enqLsq_req_1_bits_ctrl_rfWen,
  output        io_enqLsq_req_1_bits_ctrl_fpWen,
  output        io_enqLsq_req_1_bits_ctrl_flushPipe,
  output        io_enqLsq_req_1_bits_ctrl_replayInst,
  output [5:0]  io_enqLsq_req_1_bits_pdest,
  output        io_enqLsq_req_1_bits_robIdx_flag,
  output [4:0]  io_enqLsq_req_1_bits_robIdx_value,
  output [3:0]  io_enqLsq_req_1_bits_lqIdx_value,
  output [3:0]  io_enqLsq_req_1_bits_sqIdx_value,
  output        io_enqLsq_req_2_valid,
  output        io_enqLsq_req_2_bits_cf_trigger_backendEn_0,
  output        io_enqLsq_req_2_bits_cf_trigger_backendEn_1,
  output [6:0]  io_enqLsq_req_2_bits_ctrl_fuOpType,
  output        io_enqLsq_req_2_bits_ctrl_rfWen,
  output        io_enqLsq_req_2_bits_ctrl_fpWen,
  output        io_enqLsq_req_2_bits_ctrl_flushPipe,
  output        io_enqLsq_req_2_bits_ctrl_replayInst,
  output [5:0]  io_enqLsq_req_2_bits_pdest,
  output        io_enqLsq_req_2_bits_robIdx_flag,
  output [4:0]  io_enqLsq_req_2_bits_robIdx_value,
  output [3:0]  io_enqLsq_req_2_bits_lqIdx_value,
  output [3:0]  io_enqLsq_req_2_bits_sqIdx_value,
  output        io_enqLsq_req_3_valid,
  output        io_enqLsq_req_3_bits_cf_trigger_backendEn_0,
  output        io_enqLsq_req_3_bits_cf_trigger_backendEn_1,
  output [6:0]  io_enqLsq_req_3_bits_ctrl_fuOpType,
  output        io_enqLsq_req_3_bits_ctrl_rfWen,
  output        io_enqLsq_req_3_bits_ctrl_fpWen,
  output        io_enqLsq_req_3_bits_ctrl_flushPipe,
  output        io_enqLsq_req_3_bits_ctrl_replayInst,
  output [5:0]  io_enqLsq_req_3_bits_pdest,
  output        io_enqLsq_req_3_bits_robIdx_flag,
  output [4:0]  io_enqLsq_req_3_bits_robIdx_value,
  output [3:0]  io_enqLsq_req_3_bits_lqIdx_value,
  output [3:0]  io_enqLsq_req_3_bits_sqIdx_value,
  input  [4:0]  io_lqCancelCnt,
  input  [3:0]  io_sqCancelCnt,
  input  [1:0]  io_lqDeq,
  input  [1:0]  io_sqDeq,
  input         io_exuRedirect_0_valid,
  input         io_exuRedirect_0_bits_uop_cf_pd_isRVC,
  input  [1:0]  io_exuRedirect_0_bits_uop_cf_pd_brType,
  input         io_exuRedirect_0_bits_uop_cf_pd_isCall,
  input         io_exuRedirect_0_bits_uop_cf_pd_isRet,
  input  [19:0] io_exuRedirect_0_bits_uop_ctrl_imm,
  input         io_exuRedirect_0_bits_uop_robIdx_flag,
  input  [4:0]  io_exuRedirect_0_bits_uop_robIdx_value,
  input         io_exuRedirect_0_bits_redirectValid,
  input         io_exuRedirect_0_bits_redirect_robIdx_flag,
  input  [4:0]  io_exuRedirect_0_bits_redirect_robIdx_value,
  input         io_exuRedirect_0_bits_redirect_ftqIdx_flag,
  input  [2:0]  io_exuRedirect_0_bits_redirect_ftqIdx_value,
  input  [2:0]  io_exuRedirect_0_bits_redirect_ftqOffset,
  input  [38:0] io_exuRedirect_0_bits_redirect_cfiUpdate_target,
  input         io_exuRedirect_0_bits_redirect_cfiUpdate_isMisPred,
  input         io_exuRedirect_1_valid,
  input         io_exuRedirect_1_bits_uop_cf_pd_isRVC,
  input  [1:0]  io_exuRedirect_1_bits_uop_cf_pd_brType,
  input         io_exuRedirect_1_bits_uop_cf_pd_isCall,
  input         io_exuRedirect_1_bits_uop_cf_pd_isRet,
  input  [19:0] io_exuRedirect_1_bits_uop_ctrl_imm,
  input         io_exuRedirect_1_bits_uop_robIdx_flag,
  input  [4:0]  io_exuRedirect_1_bits_uop_robIdx_value,
  input         io_exuRedirect_1_bits_redirectValid,
  input         io_exuRedirect_1_bits_redirect_robIdx_flag,
  input  [4:0]  io_exuRedirect_1_bits_redirect_robIdx_value,
  input         io_exuRedirect_1_bits_redirect_ftqIdx_flag,
  input  [2:0]  io_exuRedirect_1_bits_redirect_ftqIdx_value,
  input  [2:0]  io_exuRedirect_1_bits_redirect_ftqOffset,
  input         io_exuRedirect_1_bits_redirect_cfiUpdate_taken,
  input         io_exuRedirect_1_bits_redirect_cfiUpdate_isMisPred,
  input         io_exuRedirect_2_valid,
  input         io_exuRedirect_2_bits_uop_cf_pd_isRVC,
  input  [1:0]  io_exuRedirect_2_bits_uop_cf_pd_brType,
  input         io_exuRedirect_2_bits_uop_cf_pd_isCall,
  input         io_exuRedirect_2_bits_uop_cf_pd_isRet,
  input  [19:0] io_exuRedirect_2_bits_uop_ctrl_imm,
  input         io_exuRedirect_2_bits_uop_robIdx_flag,
  input  [4:0]  io_exuRedirect_2_bits_uop_robIdx_value,
  input         io_exuRedirect_2_bits_redirectValid,
  input         io_exuRedirect_2_bits_redirect_robIdx_flag,
  input  [4:0]  io_exuRedirect_2_bits_redirect_robIdx_value,
  input         io_exuRedirect_2_bits_redirect_ftqIdx_flag,
  input  [2:0]  io_exuRedirect_2_bits_redirect_ftqIdx_value,
  input  [2:0]  io_exuRedirect_2_bits_redirect_ftqOffset,
  input         io_exuRedirect_2_bits_redirect_cfiUpdate_taken,
  input         io_exuRedirect_2_bits_redirect_cfiUpdate_isMisPred,
  input         io_stIn_0_valid,
  input         io_stIn_0_bits_uop_cf_storeSetHit,
  input  [4:0]  io_stIn_0_bits_uop_cf_ssid,
  input  [4:0]  io_stIn_0_bits_uop_robIdx_value,
  input         io_stIn_1_valid,
  input         io_stIn_1_bits_uop_cf_storeSetHit,
  input  [4:0]  io_stIn_1_bits_uop_cf_ssid,
  input  [4:0]  io_stIn_1_bits_uop_robIdx_value,
  input         io_memoryViolation_valid,
  input         io_memoryViolation_bits_robIdx_flag,
  input  [4:0]  io_memoryViolation_bits_robIdx_value,
  input         io_memoryViolation_bits_ftqIdx_flag,
  input  [2:0]  io_memoryViolation_bits_ftqIdx_value,
  input  [2:0]  io_memoryViolation_bits_ftqOffset,
  input  [2:0]  io_memoryViolation_bits_stFtqIdx_value,
  input  [2:0]  io_memoryViolation_bits_stFtqOffset,
  output [38:0] io_jumpPc,
  output [38:0] io_jalr_target,
  input         io_robio_toCSR_intrBitSet,
  input  [38:0] io_robio_toCSR_trapTarget,
  input         io_robio_toCSR_isXRet,
  input         io_robio_toCSR_wfiEvent,
  output        io_robio_toCSR_fflags_valid,
  output [4:0]  io_robio_toCSR_fflags_bits,
  output        io_robio_toCSR_dirty_fs,
  output [2:0]  io_robio_toCSR_perfinfo_retiredInstr,
  output        io_robio_exception_valid,
  output [38:0] io_robio_exception_bits_uop_cf_pc,
  output        io_robio_exception_bits_uop_cf_exceptionVec_0,
  output        io_robio_exception_bits_uop_cf_exceptionVec_1,
  output        io_robio_exception_bits_uop_cf_exceptionVec_2,
  output        io_robio_exception_bits_uop_cf_exceptionVec_3,
  output        io_robio_exception_bits_uop_cf_exceptionVec_4,
  output        io_robio_exception_bits_uop_cf_exceptionVec_5,
  output        io_robio_exception_bits_uop_cf_exceptionVec_6,
  output        io_robio_exception_bits_uop_cf_exceptionVec_7,
  output        io_robio_exception_bits_uop_cf_exceptionVec_8,
  output        io_robio_exception_bits_uop_cf_exceptionVec_9,
  output        io_robio_exception_bits_uop_cf_exceptionVec_11,
  output        io_robio_exception_bits_uop_cf_exceptionVec_12,
  output        io_robio_exception_bits_uop_cf_exceptionVec_13,
  output        io_robio_exception_bits_uop_cf_exceptionVec_15,
  output        io_robio_exception_bits_uop_cf_trigger_frontendHit_0,
  output        io_robio_exception_bits_uop_cf_trigger_frontendHit_1,
  output        io_robio_exception_bits_uop_cf_trigger_frontendHit_2,
  output        io_robio_exception_bits_uop_cf_trigger_frontendHit_3,
  output        io_robio_exception_bits_uop_cf_trigger_backendHit_0,
  output        io_robio_exception_bits_uop_cf_trigger_backendHit_1,
  output        io_robio_exception_bits_uop_cf_trigger_backendHit_2,
  output        io_robio_exception_bits_uop_cf_trigger_backendHit_3,
  output        io_robio_exception_bits_uop_cf_trigger_backendHit_4,
  output        io_robio_exception_bits_uop_cf_trigger_backendHit_5,
  output        io_robio_exception_bits_uop_cf_crossPageIPFFix,
  output [2:0]  io_robio_exception_bits_uop_ctrl_commitType,
  output        io_robio_exception_bits_uop_ctrl_singleStep,
  output        io_robio_exception_bits_isInterrupt,
  output [1:0]  io_robio_lsq_scommit,
  output        io_robio_lsq_pendingld,
  output        io_robio_lsq_pendingst,
  output        io_robio_lsq_commit,
  input         io_robio_lsq_isMMIO_0,
  input         io_robio_lsq_isMMIO_1,
  input  [4:0]  io_robio_lsq_uop_0_robIdx_value,
  input  [4:0]  io_robio_lsq_uop_1_robIdx_value,
  input         io_csrCtrl_lvpred_disable,
  input         io_csrCtrl_no_spec_load,
  input         io_csrCtrl_storeset_wait_store,
  input  [4:0]  io_csrCtrl_lvpred_timeout,
  input         io_csrCtrl_fusion_enable,
  input         io_csrCtrl_wfi_enable,
  input         io_csrCtrl_svinval_enable,
  input         io_csrCtrl_distribute_csr_wvalid,
  input  [11:0] io_csrCtrl_distribute_csr_waddr,
  input  [63:0] io_csrCtrl_distribute_csr_wdata,
  input         io_csrCtrl_singlestep,
  input         io_writeback_1_0_valid,
  input         io_writeback_1_0_bits_uop_robIdx_flag,
  input  [4:0]  io_writeback_1_0_bits_uop_robIdx_value,
  input         io_writeback_1_0_bits_redirectValid,
  input         io_writeback_1_0_bits_redirect_cfiUpdate_isMisPred,
  input         io_writeback_1_1_valid,
  input         io_writeback_1_1_bits_uop_robIdx_flag,
  input  [4:0]  io_writeback_1_1_bits_uop_robIdx_value,
  input         io_writeback_1_1_bits_redirectValid,
  input         io_writeback_1_1_bits_redirect_cfiUpdate_isMisPred,
  input         io_writeback_1_2_valid,
  input         io_writeback_1_2_bits_uop_cf_exceptionVec_4,
  input         io_writeback_1_2_bits_uop_cf_exceptionVec_5,
  input         io_writeback_1_2_bits_uop_cf_exceptionVec_13,
  input         io_writeback_1_2_bits_uop_cf_trigger_backendHit_0,
  input         io_writeback_1_2_bits_uop_cf_trigger_backendHit_1,
  input         io_writeback_1_2_bits_uop_cf_trigger_backendHit_2,
  input         io_writeback_1_2_bits_uop_cf_trigger_backendHit_3,
  input         io_writeback_1_2_bits_uop_cf_trigger_backendHit_4,
  input         io_writeback_1_2_bits_uop_cf_trigger_backendHit_5,
  input         io_writeback_1_2_bits_uop_ctrl_flushPipe,
  input         io_writeback_1_2_bits_uop_ctrl_replayInst,
  input         io_writeback_1_2_bits_uop_robIdx_flag,
  input  [4:0]  io_writeback_1_2_bits_uop_robIdx_value,
  input         io_writeback_1_2_bits_debug_isMMIO,
  input         io_writeback_1_3_valid,
  input         io_writeback_1_3_bits_uop_cf_exceptionVec_4,
  input         io_writeback_1_3_bits_uop_cf_exceptionVec_5,
  input         io_writeback_1_3_bits_uop_cf_exceptionVec_13,
  input         io_writeback_1_3_bits_uop_cf_trigger_backendHit_0,
  input         io_writeback_1_3_bits_uop_cf_trigger_backendHit_1,
  input         io_writeback_1_3_bits_uop_cf_trigger_backendHit_2,
  input         io_writeback_1_3_bits_uop_cf_trigger_backendHit_3,
  input         io_writeback_1_3_bits_uop_cf_trigger_backendHit_4,
  input         io_writeback_1_3_bits_uop_cf_trigger_backendHit_5,
  input         io_writeback_1_3_bits_uop_ctrl_flushPipe,
  input         io_writeback_1_3_bits_uop_ctrl_replayInst,
  input         io_writeback_1_3_bits_uop_robIdx_flag,
  input  [4:0]  io_writeback_1_3_bits_uop_robIdx_value,
  input         io_writeback_1_3_bits_debug_isMMIO,
  input         io_writeback_1_4_valid,
  input         io_writeback_1_4_bits_uop_cf_exceptionVec_2,
  input         io_writeback_1_4_bits_uop_cf_exceptionVec_3,
  input         io_writeback_1_4_bits_uop_cf_exceptionVec_8,
  input         io_writeback_1_4_bits_uop_cf_exceptionVec_9,
  input         io_writeback_1_4_bits_uop_cf_exceptionVec_11,
  input         io_writeback_1_4_bits_uop_ctrl_flushPipe,
  input         io_writeback_1_4_bits_uop_robIdx_flag,
  input  [4:0]  io_writeback_1_4_bits_uop_robIdx_value,
  input         io_writeback_1_4_bits_redirectValid,
  input         io_writeback_1_4_bits_redirect_cfiUpdate_isMisPred,
  input         io_writeback_1_4_bits_debug_isPerfCnt,
  input         io_writeback_1_5_valid,
  input         io_writeback_1_5_bits_uop_cf_trigger_backendHit_0,
  input         io_writeback_1_5_bits_uop_cf_trigger_backendHit_1,
  input         io_writeback_1_5_bits_uop_cf_trigger_backendHit_2,
  input         io_writeback_1_5_bits_uop_cf_trigger_backendHit_3,
  input         io_writeback_1_5_bits_uop_cf_trigger_backendHit_4,
  input         io_writeback_1_5_bits_uop_cf_trigger_backendHit_5,
  input         io_writeback_1_5_bits_uop_robIdx_flag,
  input  [4:0]  io_writeback_1_5_bits_uop_robIdx_value,
  input         io_writeback_1_6_valid,
  input         io_writeback_1_6_bits_uop_cf_exceptionVec_2,
  input         io_writeback_1_6_bits_uop_cf_exceptionVec_3,
  input         io_writeback_1_6_bits_uop_cf_exceptionVec_8,
  input         io_writeback_1_6_bits_uop_cf_exceptionVec_9,
  input         io_writeback_1_6_bits_uop_cf_exceptionVec_11,
  input         io_writeback_1_6_bits_uop_ctrl_flushPipe,
  input         io_writeback_1_6_bits_uop_robIdx_flag,
  input  [4:0]  io_writeback_1_6_bits_uop_robIdx_value,
  input         io_writeback_1_6_bits_redirectValid,
  input         io_writeback_1_6_bits_redirect_cfiUpdate_isMisPred,
  input         io_writeback_1_6_bits_debug_isPerfCnt,
  input         io_writeback_1_7_valid,
  input         io_writeback_1_7_bits_uop_cf_exceptionVec_4,
  input         io_writeback_1_7_bits_uop_cf_exceptionVec_5,
  input         io_writeback_1_7_bits_uop_cf_exceptionVec_6,
  input         io_writeback_1_7_bits_uop_cf_exceptionVec_7,
  input         io_writeback_1_7_bits_uop_cf_exceptionVec_13,
  input         io_writeback_1_7_bits_uop_cf_exceptionVec_15,
  input         io_writeback_1_7_bits_uop_cf_trigger_backendHit_0,
  input         io_writeback_1_7_bits_uop_cf_trigger_backendHit_1,
  input         io_writeback_1_7_bits_uop_cf_trigger_backendHit_2,
  input         io_writeback_1_7_bits_uop_cf_trigger_backendHit_3,
  input         io_writeback_1_7_bits_uop_cf_trigger_backendHit_4,
  input         io_writeback_1_7_bits_uop_cf_trigger_backendHit_5,
  input         io_writeback_1_7_bits_uop_robIdx_flag,
  input  [4:0]  io_writeback_1_7_bits_uop_robIdx_value,
  input         io_writeback_1_7_bits_redirectValid,
  input         io_writeback_1_7_bits_redirect_cfiUpdate_isMisPred,
  input         io_writeback_1_7_bits_debug_isMMIO,
  input         io_writeback_1_7_bits_debug_isPerfCnt,
  input         io_writeback_1_8_valid,
  input         io_writeback_1_8_bits_uop_cf_exceptionVec_4,
  input         io_writeback_1_8_bits_uop_cf_exceptionVec_5,
  input         io_writeback_1_8_bits_uop_cf_exceptionVec_6,
  input         io_writeback_1_8_bits_uop_cf_exceptionVec_7,
  input         io_writeback_1_8_bits_uop_cf_exceptionVec_13,
  input         io_writeback_1_8_bits_uop_cf_exceptionVec_15,
  input         io_writeback_1_8_bits_uop_cf_trigger_backendHit_0,
  input         io_writeback_1_8_bits_uop_cf_trigger_backendHit_1,
  input         io_writeback_1_8_bits_uop_cf_trigger_backendHit_2,
  input         io_writeback_1_8_bits_uop_cf_trigger_backendHit_3,
  input         io_writeback_1_8_bits_uop_cf_trigger_backendHit_4,
  input         io_writeback_1_8_bits_uop_cf_trigger_backendHit_5,
  input         io_writeback_1_8_bits_uop_robIdx_flag,
  input  [4:0]  io_writeback_1_8_bits_uop_robIdx_value,
  input         io_writeback_1_8_bits_redirectValid,
  input         io_writeback_1_8_bits_redirect_cfiUpdate_isMisPred,
  input         io_writeback_1_8_bits_debug_isMMIO,
  input         io_writeback_1_8_bits_debug_isPerfCnt,
  input         io_writeback_1_9_valid,
  input         io_writeback_1_9_bits_uop_robIdx_flag,
  input  [4:0]  io_writeback_1_9_bits_uop_robIdx_value,
  input         io_writeback_1_10_valid,
  input         io_writeback_1_10_bits_uop_robIdx_flag,
  input  [4:0]  io_writeback_1_10_bits_uop_robIdx_value,
  input         io_writeback_0_3_valid,
  input         io_writeback_0_3_bits_uop_cf_exceptionVec_2,
  input         io_writeback_0_3_bits_uop_cf_exceptionVec_3,
  input         io_writeback_0_3_bits_uop_cf_exceptionVec_8,
  input         io_writeback_0_3_bits_uop_cf_exceptionVec_9,
  input         io_writeback_0_3_bits_uop_cf_exceptionVec_11,
  input         io_writeback_0_3_bits_uop_ctrl_flushPipe,
  input         io_writeback_0_3_bits_uop_robIdx_flag,
  input  [4:0]  io_writeback_0_3_bits_uop_robIdx_value,
  input  [4:0]  io_writeback_0_3_bits_fflags,
  input         io_writeback_0_4_valid,
  input         io_writeback_0_4_bits_uop_robIdx_flag,
  input  [4:0]  io_writeback_0_4_bits_uop_robIdx_value,
  input  [4:0]  io_writeback_0_4_bits_fflags,
  input         io_writeback_0_5_valid,
  input         io_writeback_0_5_bits_uop_robIdx_flag,
  input  [4:0]  io_writeback_0_5_bits_uop_robIdx_value,
  input  [4:0]  io_writeback_0_5_bits_fflags,
  input         io_writeback_0_6_valid,
  input         io_writeback_0_6_bits_uop_cf_exceptionVec_4,
  input         io_writeback_0_6_bits_uop_cf_exceptionVec_5,
  input         io_writeback_0_6_bits_uop_cf_exceptionVec_13,
  input         io_writeback_0_6_bits_uop_cf_trigger_backendHit_0,
  input         io_writeback_0_6_bits_uop_cf_trigger_backendHit_1,
  input         io_writeback_0_6_bits_uop_cf_trigger_backendHit_2,
  input         io_writeback_0_6_bits_uop_cf_trigger_backendHit_3,
  input         io_writeback_0_6_bits_uop_cf_trigger_backendHit_4,
  input         io_writeback_0_6_bits_uop_cf_trigger_backendHit_5,
  input         io_writeback_0_6_bits_uop_ctrl_flushPipe,
  input         io_writeback_0_6_bits_uop_ctrl_replayInst,
  input         io_writeback_0_6_bits_uop_robIdx_flag,
  input  [4:0]  io_writeback_0_6_bits_uop_robIdx_value,
  input         io_writeback_0_7_valid,
  input         io_writeback_0_7_bits_uop_cf_exceptionVec_4,
  input         io_writeback_0_7_bits_uop_cf_exceptionVec_5,
  input         io_writeback_0_7_bits_uop_cf_exceptionVec_13,
  input         io_writeback_0_7_bits_uop_cf_trigger_backendHit_0,
  input         io_writeback_0_7_bits_uop_cf_trigger_backendHit_1,
  input         io_writeback_0_7_bits_uop_cf_trigger_backendHit_2,
  input         io_writeback_0_7_bits_uop_cf_trigger_backendHit_3,
  input         io_writeback_0_7_bits_uop_cf_trigger_backendHit_4,
  input         io_writeback_0_7_bits_uop_cf_trigger_backendHit_5,
  input         io_writeback_0_7_bits_uop_ctrl_flushPipe,
  input         io_writeback_0_7_bits_uop_ctrl_replayInst,
  input         io_writeback_0_7_bits_uop_robIdx_flag,
  input  [4:0]  io_writeback_0_7_bits_uop_robIdx_value,
  input         io_writeback_0_8_valid,
  input         io_writeback_0_8_bits_uop_cf_exceptionVec_4,
  input         io_writeback_0_8_bits_uop_cf_exceptionVec_5,
  input         io_writeback_0_8_bits_uop_cf_exceptionVec_6,
  input         io_writeback_0_8_bits_uop_cf_exceptionVec_7,
  input         io_writeback_0_8_bits_uop_cf_exceptionVec_13,
  input         io_writeback_0_8_bits_uop_cf_exceptionVec_15,
  input         io_writeback_0_8_bits_uop_cf_trigger_backendHit_0,
  input         io_writeback_0_8_bits_uop_cf_trigger_backendHit_1,
  input         io_writeback_0_8_bits_uop_cf_trigger_backendHit_2,
  input         io_writeback_0_8_bits_uop_cf_trigger_backendHit_3,
  input         io_writeback_0_8_bits_uop_cf_trigger_backendHit_4,
  input         io_writeback_0_8_bits_uop_cf_trigger_backendHit_5,
  input         io_writeback_0_8_bits_uop_robIdx_flag,
  input  [4:0]  io_writeback_0_8_bits_uop_robIdx_value,
  input         io_writeback_0_9_valid,
  input         io_writeback_0_9_bits_uop_cf_exceptionVec_6,
  input         io_writeback_0_9_bits_uop_cf_exceptionVec_7,
  input         io_writeback_0_9_bits_uop_cf_exceptionVec_15,
  input         io_writeback_0_9_bits_uop_cf_trigger_backendHit_0,
  input         io_writeback_0_9_bits_uop_cf_trigger_backendHit_1,
  input         io_writeback_0_9_bits_uop_cf_trigger_backendHit_4,
  input         io_writeback_0_9_bits_uop_robIdx_flag,
  input  [4:0]  io_writeback_0_9_bits_uop_robIdx_value,
  output        io_redirect_valid,
  output        io_redirect_bits_robIdx_flag,
  output [4:0]  io_redirect_bits_robIdx_value,
  output        io_redirect_bits_level,
  output [5:0]  io_debug_int_rat_0,
  output [5:0]  io_debug_int_rat_1,
  output [5:0]  io_debug_int_rat_2,
  output [5:0]  io_debug_int_rat_3,
  output [5:0]  io_debug_int_rat_4,
  output [5:0]  io_debug_int_rat_5,
  output [5:0]  io_debug_int_rat_6,
  output [5:0]  io_debug_int_rat_7,
  output [5:0]  io_debug_int_rat_8,
  output [5:0]  io_debug_int_rat_9,
  output [5:0]  io_debug_int_rat_10,
  output [5:0]  io_debug_int_rat_11,
  output [5:0]  io_debug_int_rat_12,
  output [5:0]  io_debug_int_rat_13,
  output [5:0]  io_debug_int_rat_14,
  output [5:0]  io_debug_int_rat_15,
  output [5:0]  io_debug_int_rat_16,
  output [5:0]  io_debug_int_rat_17,
  output [5:0]  io_debug_int_rat_18,
  output [5:0]  io_debug_int_rat_19,
  output [5:0]  io_debug_int_rat_20,
  output [5:0]  io_debug_int_rat_21,
  output [5:0]  io_debug_int_rat_22,
  output [5:0]  io_debug_int_rat_23,
  output [5:0]  io_debug_int_rat_24,
  output [5:0]  io_debug_int_rat_25,
  output [5:0]  io_debug_int_rat_26,
  output [5:0]  io_debug_int_rat_27,
  output [5:0]  io_debug_int_rat_28,
  output [5:0]  io_debug_int_rat_29,
  output [5:0]  io_debug_int_rat_30,
  output [5:0]  io_debug_int_rat_31,
  output [5:0]  io_debug_fp_rat_0,
  output [5:0]  io_debug_fp_rat_1,
  output [5:0]  io_debug_fp_rat_2,
  output [5:0]  io_debug_fp_rat_3,
  output [5:0]  io_debug_fp_rat_4,
  output [5:0]  io_debug_fp_rat_5,
  output [5:0]  io_debug_fp_rat_6,
  output [5:0]  io_debug_fp_rat_7,
  output [5:0]  io_debug_fp_rat_8,
  output [5:0]  io_debug_fp_rat_9,
  output [5:0]  io_debug_fp_rat_10,
  output [5:0]  io_debug_fp_rat_11,
  output [5:0]  io_debug_fp_rat_12,
  output [5:0]  io_debug_fp_rat_13,
  output [5:0]  io_debug_fp_rat_14,
  output [5:0]  io_debug_fp_rat_15,
  output [5:0]  io_debug_fp_rat_16,
  output [5:0]  io_debug_fp_rat_17,
  output [5:0]  io_debug_fp_rat_18,
  output [5:0]  io_debug_fp_rat_19,
  output [5:0]  io_debug_fp_rat_20,
  output [5:0]  io_debug_fp_rat_21,
  output [5:0]  io_debug_fp_rat_22,
  output [5:0]  io_debug_fp_rat_23,
  output [5:0]  io_debug_fp_rat_24,
  output [5:0]  io_debug_fp_rat_25,
  output [5:0]  io_debug_fp_rat_26,
  output [5:0]  io_debug_fp_rat_27,
  output [5:0]  io_debug_fp_rat_28,
  output [5:0]  io_debug_fp_rat_29,
  output [5:0]  io_debug_fp_rat_30,
  output [5:0]  io_debug_fp_rat_31,
  input  [5:0]  perfinfo_perfEventsRs_0_value,
  input  [5:0]  perfinfo_perfEventsRs_1_value,
  input  [5:0]  perfinfo_perfEventsRs_2_value,
  input  [5:0]  perfinfo_perfEventsRs_3_value,
  input  [5:0]  perfinfo_perfEventsRs_4_value,
  input  [5:0]  perfinfo_perfEventsRs_5_value,
  input  [5:0]  perfinfo_perfEventsRs_6_value,
  input  [5:0]  perfinfo_perfEventsRs_7_value,
  input  [5:0]  perfinfo_perfEventsEu0_0_value,
  input  [5:0]  perfinfo_perfEventsEu0_1_value,
  input  [5:0]  perfinfo_perfEventsEu0_2_value,
  input  [5:0]  perfinfo_perfEventsEu0_3_value,
  input  [5:0]  perfinfo_perfEventsEu0_4_value,
  input  [5:0]  perfinfo_perfEventsEu0_5_value,
  input  [5:0]  perfinfo_perfEventsEu1_0_value,
  input  [5:0]  perfinfo_perfEventsEu1_1_value,
  input  [5:0]  perfinfo_perfEventsEu1_2_value,
  input  [5:0]  perfinfo_perfEventsEu1_3_value,
  input  [5:0]  perfinfo_perfEventsEu1_4_value,
  input  [5:0]  perfinfo_perfEventsEu1_5_value,
  output [5:0]  io_perf_0_value,
  output [5:0]  io_perf_1_value,
  output [5:0]  io_perf_2_value,
  output [5:0]  io_perf_3_value,
  output [5:0]  io_perf_4_value,
  output [5:0]  io_perf_5_value,
  output [5:0]  io_perf_6_value,
  output [5:0]  io_perf_7_value
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [63:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [63:0] _RAND_87;
  reg [63:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [63:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [63:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
`endif // RANDOMIZE_REG_INIT
  wire  rob_clock; // @[CtrlBlock.scala 173:23]
  wire  rob_reset; // @[CtrlBlock.scala 173:23]
  wire [7:0] rob_io_hartId; // @[CtrlBlock.scala 173:23]
  wire  rob_io_redirect_valid; // @[CtrlBlock.scala 173:23]
  wire  rob_io_redirect_bits_robIdx_flag; // @[CtrlBlock.scala 173:23]
  wire [4:0] rob_io_redirect_bits_robIdx_value; // @[CtrlBlock.scala 173:23]
  wire  rob_io_redirect_bits_level; // @[CtrlBlock.scala 173:23]
  wire  rob_io_enq_canAccept; // @[CtrlBlock.scala 173:23]
  wire  rob_io_enq_isEmpty; // @[CtrlBlock.scala 173:23]
  wire  rob_io_enq_needAlloc_0; // @[CtrlBlock.scala 173:23]
  wire  rob_io_enq_req_0_valid; // @[CtrlBlock.scala 173:23]
  wire  rob_io_enq_req_0_bits_cf_exceptionVec_1; // @[CtrlBlock.scala 173:23]
  wire  rob_io_enq_req_0_bits_cf_exceptionVec_2; // @[CtrlBlock.scala 173:23]
  wire  rob_io_enq_req_0_bits_cf_exceptionVec_12; // @[CtrlBlock.scala 173:23]
  wire  rob_io_enq_req_0_bits_cf_trigger_frontendHit_0; // @[CtrlBlock.scala 173:23]
  wire  rob_io_enq_req_0_bits_cf_trigger_frontendHit_1; // @[CtrlBlock.scala 173:23]
  wire  rob_io_enq_req_0_bits_cf_trigger_frontendHit_2; // @[CtrlBlock.scala 173:23]
  wire  rob_io_enq_req_0_bits_cf_trigger_frontendHit_3; // @[CtrlBlock.scala 173:23]
  wire  rob_io_enq_req_0_bits_cf_pd_isRVC; // @[CtrlBlock.scala 173:23]
  wire  rob_io_enq_req_0_bits_cf_crossPageIPFFix; // @[CtrlBlock.scala 173:23]
  wire  rob_io_enq_req_0_bits_cf_loadWaitBit; // @[CtrlBlock.scala 173:23]
  wire  rob_io_enq_req_0_bits_cf_ftqPtr_flag; // @[CtrlBlock.scala 173:23]
  wire [2:0] rob_io_enq_req_0_bits_cf_ftqPtr_value; // @[CtrlBlock.scala 173:23]
  wire [2:0] rob_io_enq_req_0_bits_cf_ftqOffset; // @[CtrlBlock.scala 173:23]
  wire [4:0] rob_io_enq_req_0_bits_ctrl_ldest; // @[CtrlBlock.scala 173:23]
  wire [3:0] rob_io_enq_req_0_bits_ctrl_fuType; // @[CtrlBlock.scala 173:23]
  wire [6:0] rob_io_enq_req_0_bits_ctrl_fuOpType; // @[CtrlBlock.scala 173:23]
  wire  rob_io_enq_req_0_bits_ctrl_rfWen; // @[CtrlBlock.scala 173:23]
  wire  rob_io_enq_req_0_bits_ctrl_fpWen; // @[CtrlBlock.scala 173:23]
  wire  rob_io_enq_req_0_bits_ctrl_isXSTrap; // @[CtrlBlock.scala 173:23]
  wire  rob_io_enq_req_0_bits_ctrl_noSpecExec; // @[CtrlBlock.scala 173:23]
  wire  rob_io_enq_req_0_bits_ctrl_blockBackward; // @[CtrlBlock.scala 173:23]
  wire  rob_io_enq_req_0_bits_ctrl_flushPipe; // @[CtrlBlock.scala 173:23]
  wire [2:0] rob_io_enq_req_0_bits_ctrl_commitType; // @[CtrlBlock.scala 173:23]
  wire  rob_io_enq_req_0_bits_ctrl_fpu_wflags; // @[CtrlBlock.scala 173:23]
  wire  rob_io_enq_req_0_bits_ctrl_isMove; // @[CtrlBlock.scala 173:23]
  wire  rob_io_enq_req_0_bits_ctrl_singleStep; // @[CtrlBlock.scala 173:23]
  wire [5:0] rob_io_enq_req_0_bits_pdest; // @[CtrlBlock.scala 173:23]
  wire [5:0] rob_io_enq_req_0_bits_old_pdest; // @[CtrlBlock.scala 173:23]
  wire  rob_io_enq_req_0_bits_robIdx_flag; // @[CtrlBlock.scala 173:23]
  wire [4:0] rob_io_enq_req_0_bits_robIdx_value; // @[CtrlBlock.scala 173:23]
  wire  rob_io_enq_req_0_bits_eliminatedMove; // @[CtrlBlock.scala 173:23]
  wire  rob_io_enq_req_1_valid; // @[CtrlBlock.scala 173:23]
  wire  rob_io_enq_req_1_bits_cf_exceptionVec_1; // @[CtrlBlock.scala 173:23]
  wire  rob_io_enq_req_1_bits_cf_exceptionVec_2; // @[CtrlBlock.scala 173:23]
  wire  rob_io_enq_req_1_bits_cf_exceptionVec_12; // @[CtrlBlock.scala 173:23]
  wire  rob_io_enq_req_1_bits_cf_trigger_frontendHit_0; // @[CtrlBlock.scala 173:23]
  wire  rob_io_enq_req_1_bits_cf_trigger_frontendHit_1; // @[CtrlBlock.scala 173:23]
  wire  rob_io_enq_req_1_bits_cf_trigger_frontendHit_2; // @[CtrlBlock.scala 173:23]
  wire  rob_io_enq_req_1_bits_cf_trigger_frontendHit_3; // @[CtrlBlock.scala 173:23]
  wire  rob_io_enq_req_1_bits_cf_pd_isRVC; // @[CtrlBlock.scala 173:23]
  wire  rob_io_enq_req_1_bits_cf_crossPageIPFFix; // @[CtrlBlock.scala 173:23]
  wire  rob_io_enq_req_1_bits_cf_loadWaitBit; // @[CtrlBlock.scala 173:23]
  wire  rob_io_enq_req_1_bits_cf_ftqPtr_flag; // @[CtrlBlock.scala 173:23]
  wire [2:0] rob_io_enq_req_1_bits_cf_ftqPtr_value; // @[CtrlBlock.scala 173:23]
  wire [2:0] rob_io_enq_req_1_bits_cf_ftqOffset; // @[CtrlBlock.scala 173:23]
  wire [4:0] rob_io_enq_req_1_bits_ctrl_ldest; // @[CtrlBlock.scala 173:23]
  wire [3:0] rob_io_enq_req_1_bits_ctrl_fuType; // @[CtrlBlock.scala 173:23]
  wire [6:0] rob_io_enq_req_1_bits_ctrl_fuOpType; // @[CtrlBlock.scala 173:23]
  wire  rob_io_enq_req_1_bits_ctrl_rfWen; // @[CtrlBlock.scala 173:23]
  wire  rob_io_enq_req_1_bits_ctrl_fpWen; // @[CtrlBlock.scala 173:23]
  wire  rob_io_enq_req_1_bits_ctrl_isXSTrap; // @[CtrlBlock.scala 173:23]
  wire  rob_io_enq_req_1_bits_ctrl_noSpecExec; // @[CtrlBlock.scala 173:23]
  wire  rob_io_enq_req_1_bits_ctrl_blockBackward; // @[CtrlBlock.scala 173:23]
  wire  rob_io_enq_req_1_bits_ctrl_flushPipe; // @[CtrlBlock.scala 173:23]
  wire [2:0] rob_io_enq_req_1_bits_ctrl_commitType; // @[CtrlBlock.scala 173:23]
  wire  rob_io_enq_req_1_bits_ctrl_fpu_wflags; // @[CtrlBlock.scala 173:23]
  wire  rob_io_enq_req_1_bits_ctrl_isMove; // @[CtrlBlock.scala 173:23]
  wire  rob_io_enq_req_1_bits_ctrl_singleStep; // @[CtrlBlock.scala 173:23]
  wire [5:0] rob_io_enq_req_1_bits_pdest; // @[CtrlBlock.scala 173:23]
  wire [5:0] rob_io_enq_req_1_bits_old_pdest; // @[CtrlBlock.scala 173:23]
  wire  rob_io_enq_req_1_bits_robIdx_flag; // @[CtrlBlock.scala 173:23]
  wire [4:0] rob_io_enq_req_1_bits_robIdx_value; // @[CtrlBlock.scala 173:23]
  wire  rob_io_enq_req_1_bits_eliminatedMove; // @[CtrlBlock.scala 173:23]
  wire  rob_io_flushOut_valid; // @[CtrlBlock.scala 173:23]
  wire  rob_io_flushOut_bits_robIdx_flag; // @[CtrlBlock.scala 173:23]
  wire [4:0] rob_io_flushOut_bits_robIdx_value; // @[CtrlBlock.scala 173:23]
  wire  rob_io_flushOut_bits_ftqIdx_flag; // @[CtrlBlock.scala 173:23]
  wire [2:0] rob_io_flushOut_bits_ftqIdx_value; // @[CtrlBlock.scala 173:23]
  wire [2:0] rob_io_flushOut_bits_ftqOffset; // @[CtrlBlock.scala 173:23]
  wire  rob_io_flushOut_bits_level; // @[CtrlBlock.scala 173:23]
  wire  rob_io_exception_valid; // @[CtrlBlock.scala 173:23]
  wire  rob_io_exception_bits_uop_cf_exceptionVec_0; // @[CtrlBlock.scala 173:23]
  wire  rob_io_exception_bits_uop_cf_exceptionVec_1; // @[CtrlBlock.scala 173:23]
  wire  rob_io_exception_bits_uop_cf_exceptionVec_2; // @[CtrlBlock.scala 173:23]
  wire  rob_io_exception_bits_uop_cf_exceptionVec_3; // @[CtrlBlock.scala 173:23]
  wire  rob_io_exception_bits_uop_cf_exceptionVec_4; // @[CtrlBlock.scala 173:23]
  wire  rob_io_exception_bits_uop_cf_exceptionVec_5; // @[CtrlBlock.scala 173:23]
  wire  rob_io_exception_bits_uop_cf_exceptionVec_6; // @[CtrlBlock.scala 173:23]
  wire  rob_io_exception_bits_uop_cf_exceptionVec_7; // @[CtrlBlock.scala 173:23]
  wire  rob_io_exception_bits_uop_cf_exceptionVec_8; // @[CtrlBlock.scala 173:23]
  wire  rob_io_exception_bits_uop_cf_exceptionVec_9; // @[CtrlBlock.scala 173:23]
  wire  rob_io_exception_bits_uop_cf_exceptionVec_11; // @[CtrlBlock.scala 173:23]
  wire  rob_io_exception_bits_uop_cf_exceptionVec_12; // @[CtrlBlock.scala 173:23]
  wire  rob_io_exception_bits_uop_cf_exceptionVec_13; // @[CtrlBlock.scala 173:23]
  wire  rob_io_exception_bits_uop_cf_exceptionVec_15; // @[CtrlBlock.scala 173:23]
  wire  rob_io_exception_bits_uop_cf_trigger_frontendHit_0; // @[CtrlBlock.scala 173:23]
  wire  rob_io_exception_bits_uop_cf_trigger_frontendHit_1; // @[CtrlBlock.scala 173:23]
  wire  rob_io_exception_bits_uop_cf_trigger_frontendHit_2; // @[CtrlBlock.scala 173:23]
  wire  rob_io_exception_bits_uop_cf_trigger_frontendHit_3; // @[CtrlBlock.scala 173:23]
  wire  rob_io_exception_bits_uop_cf_trigger_backendHit_0; // @[CtrlBlock.scala 173:23]
  wire  rob_io_exception_bits_uop_cf_trigger_backendHit_1; // @[CtrlBlock.scala 173:23]
  wire  rob_io_exception_bits_uop_cf_trigger_backendHit_2; // @[CtrlBlock.scala 173:23]
  wire  rob_io_exception_bits_uop_cf_trigger_backendHit_3; // @[CtrlBlock.scala 173:23]
  wire  rob_io_exception_bits_uop_cf_trigger_backendHit_4; // @[CtrlBlock.scala 173:23]
  wire  rob_io_exception_bits_uop_cf_trigger_backendHit_5; // @[CtrlBlock.scala 173:23]
  wire  rob_io_exception_bits_uop_cf_crossPageIPFFix; // @[CtrlBlock.scala 173:23]
  wire [2:0] rob_io_exception_bits_uop_ctrl_commitType; // @[CtrlBlock.scala 173:23]
  wire  rob_io_exception_bits_uop_ctrl_singleStep; // @[CtrlBlock.scala 173:23]
  wire  rob_io_exception_bits_isInterrupt; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_0_valid; // @[CtrlBlock.scala 173:23]
  wire [4:0] rob_io_writeback_1_0_bits_uop_robIdx_value; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_0_bits_redirectValid; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_0_bits_redirect_cfiUpdate_isMisPred; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_1_valid; // @[CtrlBlock.scala 173:23]
  wire [4:0] rob_io_writeback_1_1_bits_uop_robIdx_value; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_1_bits_redirectValid; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_1_bits_redirect_cfiUpdate_isMisPred; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_2_valid; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_2_bits_uop_cf_exceptionVec_4; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_2_bits_uop_cf_exceptionVec_5; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_2_bits_uop_cf_exceptionVec_13; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_2_bits_uop_cf_trigger_backendHit_0; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_2_bits_uop_cf_trigger_backendHit_1; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_2_bits_uop_cf_trigger_backendHit_2; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_2_bits_uop_cf_trigger_backendHit_3; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_2_bits_uop_cf_trigger_backendHit_4; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_2_bits_uop_cf_trigger_backendHit_5; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_2_bits_uop_ctrl_flushPipe; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_2_bits_uop_ctrl_replayInst; // @[CtrlBlock.scala 173:23]
  wire [4:0] rob_io_writeback_1_2_bits_uop_robIdx_value; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_2_bits_debug_isMMIO; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_3_valid; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_3_bits_uop_cf_exceptionVec_4; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_3_bits_uop_cf_exceptionVec_5; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_3_bits_uop_cf_exceptionVec_13; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_3_bits_uop_cf_trigger_backendHit_0; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_3_bits_uop_cf_trigger_backendHit_1; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_3_bits_uop_cf_trigger_backendHit_2; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_3_bits_uop_cf_trigger_backendHit_3; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_3_bits_uop_cf_trigger_backendHit_4; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_3_bits_uop_cf_trigger_backendHit_5; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_3_bits_uop_ctrl_flushPipe; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_3_bits_uop_ctrl_replayInst; // @[CtrlBlock.scala 173:23]
  wire [4:0] rob_io_writeback_1_3_bits_uop_robIdx_value; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_3_bits_debug_isMMIO; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_4_valid; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_4_bits_uop_cf_exceptionVec_2; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_4_bits_uop_cf_exceptionVec_3; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_4_bits_uop_cf_exceptionVec_8; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_4_bits_uop_cf_exceptionVec_9; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_4_bits_uop_cf_exceptionVec_11; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_4_bits_uop_ctrl_flushPipe; // @[CtrlBlock.scala 173:23]
  wire [4:0] rob_io_writeback_1_4_bits_uop_robIdx_value; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_4_bits_redirectValid; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_4_bits_redirect_cfiUpdate_isMisPred; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_4_bits_debug_isPerfCnt; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_5_valid; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_5_bits_uop_cf_trigger_backendHit_0; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_5_bits_uop_cf_trigger_backendHit_1; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_5_bits_uop_cf_trigger_backendHit_2; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_5_bits_uop_cf_trigger_backendHit_3; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_5_bits_uop_cf_trigger_backendHit_4; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_5_bits_uop_cf_trigger_backendHit_5; // @[CtrlBlock.scala 173:23]
  wire [4:0] rob_io_writeback_1_5_bits_uop_robIdx_value; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_6_valid; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_6_bits_uop_cf_exceptionVec_2; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_6_bits_uop_cf_exceptionVec_3; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_6_bits_uop_cf_exceptionVec_8; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_6_bits_uop_cf_exceptionVec_9; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_6_bits_uop_cf_exceptionVec_11; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_6_bits_uop_ctrl_flushPipe; // @[CtrlBlock.scala 173:23]
  wire [4:0] rob_io_writeback_1_6_bits_uop_robIdx_value; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_6_bits_redirectValid; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_6_bits_redirect_cfiUpdate_isMisPred; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_6_bits_debug_isPerfCnt; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_7_valid; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_7_bits_uop_cf_exceptionVec_4; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_7_bits_uop_cf_exceptionVec_5; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_7_bits_uop_cf_exceptionVec_6; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_7_bits_uop_cf_exceptionVec_7; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_7_bits_uop_cf_exceptionVec_13; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_7_bits_uop_cf_exceptionVec_15; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_7_bits_uop_cf_trigger_backendHit_0; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_7_bits_uop_cf_trigger_backendHit_1; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_7_bits_uop_cf_trigger_backendHit_2; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_7_bits_uop_cf_trigger_backendHit_3; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_7_bits_uop_cf_trigger_backendHit_4; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_7_bits_uop_cf_trigger_backendHit_5; // @[CtrlBlock.scala 173:23]
  wire [4:0] rob_io_writeback_1_7_bits_uop_robIdx_value; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_7_bits_redirectValid; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_7_bits_redirect_cfiUpdate_isMisPred; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_7_bits_debug_isMMIO; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_7_bits_debug_isPerfCnt; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_8_valid; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_8_bits_uop_cf_exceptionVec_4; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_8_bits_uop_cf_exceptionVec_5; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_8_bits_uop_cf_exceptionVec_6; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_8_bits_uop_cf_exceptionVec_7; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_8_bits_uop_cf_exceptionVec_13; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_8_bits_uop_cf_exceptionVec_15; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_8_bits_uop_cf_trigger_backendHit_0; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_8_bits_uop_cf_trigger_backendHit_1; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_8_bits_uop_cf_trigger_backendHit_2; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_8_bits_uop_cf_trigger_backendHit_3; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_8_bits_uop_cf_trigger_backendHit_4; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_8_bits_uop_cf_trigger_backendHit_5; // @[CtrlBlock.scala 173:23]
  wire [4:0] rob_io_writeback_1_8_bits_uop_robIdx_value; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_8_bits_redirectValid; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_8_bits_redirect_cfiUpdate_isMisPred; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_8_bits_debug_isMMIO; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_8_bits_debug_isPerfCnt; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_9_valid; // @[CtrlBlock.scala 173:23]
  wire [4:0] rob_io_writeback_1_9_bits_uop_robIdx_value; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_1_10_valid; // @[CtrlBlock.scala 173:23]
  wire [4:0] rob_io_writeback_1_10_bits_uop_robIdx_value; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_0_3_valid; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_0_3_bits_uop_cf_exceptionVec_2; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_0_3_bits_uop_cf_exceptionVec_3; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_0_3_bits_uop_cf_exceptionVec_8; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_0_3_bits_uop_cf_exceptionVec_9; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_0_3_bits_uop_cf_exceptionVec_11; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_0_3_bits_uop_ctrl_flushPipe; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_0_3_bits_uop_robIdx_flag; // @[CtrlBlock.scala 173:23]
  wire [4:0] rob_io_writeback_0_3_bits_uop_robIdx_value; // @[CtrlBlock.scala 173:23]
  wire [4:0] rob_io_writeback_0_3_bits_fflags; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_0_4_valid; // @[CtrlBlock.scala 173:23]
  wire [4:0] rob_io_writeback_0_4_bits_uop_robIdx_value; // @[CtrlBlock.scala 173:23]
  wire [4:0] rob_io_writeback_0_4_bits_fflags; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_0_5_valid; // @[CtrlBlock.scala 173:23]
  wire [4:0] rob_io_writeback_0_5_bits_uop_robIdx_value; // @[CtrlBlock.scala 173:23]
  wire [4:0] rob_io_writeback_0_5_bits_fflags; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_0_6_valid; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_0_6_bits_uop_cf_exceptionVec_4; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_0_6_bits_uop_cf_exceptionVec_5; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_0_6_bits_uop_cf_exceptionVec_13; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_0_6_bits_uop_cf_trigger_backendHit_0; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_0_6_bits_uop_cf_trigger_backendHit_1; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_0_6_bits_uop_cf_trigger_backendHit_2; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_0_6_bits_uop_cf_trigger_backendHit_3; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_0_6_bits_uop_cf_trigger_backendHit_4; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_0_6_bits_uop_cf_trigger_backendHit_5; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_0_6_bits_uop_ctrl_flushPipe; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_0_6_bits_uop_ctrl_replayInst; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_0_6_bits_uop_robIdx_flag; // @[CtrlBlock.scala 173:23]
  wire [4:0] rob_io_writeback_0_6_bits_uop_robIdx_value; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_0_7_valid; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_0_7_bits_uop_cf_exceptionVec_4; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_0_7_bits_uop_cf_exceptionVec_5; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_0_7_bits_uop_cf_exceptionVec_13; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_0_7_bits_uop_cf_trigger_backendHit_0; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_0_7_bits_uop_cf_trigger_backendHit_1; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_0_7_bits_uop_cf_trigger_backendHit_2; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_0_7_bits_uop_cf_trigger_backendHit_3; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_0_7_bits_uop_cf_trigger_backendHit_4; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_0_7_bits_uop_cf_trigger_backendHit_5; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_0_7_bits_uop_ctrl_flushPipe; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_0_7_bits_uop_ctrl_replayInst; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_0_7_bits_uop_robIdx_flag; // @[CtrlBlock.scala 173:23]
  wire [4:0] rob_io_writeback_0_7_bits_uop_robIdx_value; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_0_8_valid; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_0_8_bits_uop_cf_exceptionVec_4; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_0_8_bits_uop_cf_exceptionVec_5; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_0_8_bits_uop_cf_exceptionVec_6; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_0_8_bits_uop_cf_exceptionVec_7; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_0_8_bits_uop_cf_exceptionVec_13; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_0_8_bits_uop_cf_exceptionVec_15; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_0_8_bits_uop_cf_trigger_backendHit_0; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_0_8_bits_uop_cf_trigger_backendHit_1; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_0_8_bits_uop_cf_trigger_backendHit_2; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_0_8_bits_uop_cf_trigger_backendHit_3; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_0_8_bits_uop_cf_trigger_backendHit_4; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_0_8_bits_uop_cf_trigger_backendHit_5; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_0_8_bits_uop_robIdx_flag; // @[CtrlBlock.scala 173:23]
  wire [4:0] rob_io_writeback_0_8_bits_uop_robIdx_value; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_0_9_valid; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_0_9_bits_uop_cf_exceptionVec_6; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_0_9_bits_uop_cf_exceptionVec_7; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_0_9_bits_uop_cf_exceptionVec_15; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_0_9_bits_uop_cf_trigger_backendHit_0; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_0_9_bits_uop_cf_trigger_backendHit_1; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_0_9_bits_uop_cf_trigger_backendHit_4; // @[CtrlBlock.scala 173:23]
  wire  rob_io_writeback_0_9_bits_uop_robIdx_flag; // @[CtrlBlock.scala 173:23]
  wire [4:0] rob_io_writeback_0_9_bits_uop_robIdx_value; // @[CtrlBlock.scala 173:23]
  wire  rob_io_commits_isCommit; // @[CtrlBlock.scala 173:23]
  wire  rob_io_commits_commitValid_0; // @[CtrlBlock.scala 173:23]
  wire  rob_io_commits_commitValid_1; // @[CtrlBlock.scala 173:23]
  wire  rob_io_commits_isWalk; // @[CtrlBlock.scala 173:23]
  wire  rob_io_commits_walkValid_0; // @[CtrlBlock.scala 173:23]
  wire  rob_io_commits_walkValid_1; // @[CtrlBlock.scala 173:23]
  wire [4:0] rob_io_commits_info_0_ldest; // @[CtrlBlock.scala 173:23]
  wire  rob_io_commits_info_0_rfWen; // @[CtrlBlock.scala 173:23]
  wire  rob_io_commits_info_0_fpWen; // @[CtrlBlock.scala 173:23]
  wire  rob_io_commits_info_0_wflags; // @[CtrlBlock.scala 173:23]
  wire [2:0] rob_io_commits_info_0_commitType; // @[CtrlBlock.scala 173:23]
  wire [5:0] rob_io_commits_info_0_pdest; // @[CtrlBlock.scala 173:23]
  wire [5:0] rob_io_commits_info_0_old_pdest; // @[CtrlBlock.scala 173:23]
  wire  rob_io_commits_info_0_ftqIdx_flag; // @[CtrlBlock.scala 173:23]
  wire [2:0] rob_io_commits_info_0_ftqIdx_value; // @[CtrlBlock.scala 173:23]
  wire [2:0] rob_io_commits_info_0_ftqOffset; // @[CtrlBlock.scala 173:23]
  wire  rob_io_commits_info_0_isMove; // @[CtrlBlock.scala 173:23]
  wire [4:0] rob_io_commits_info_1_ldest; // @[CtrlBlock.scala 173:23]
  wire  rob_io_commits_info_1_rfWen; // @[CtrlBlock.scala 173:23]
  wire  rob_io_commits_info_1_fpWen; // @[CtrlBlock.scala 173:23]
  wire  rob_io_commits_info_1_wflags; // @[CtrlBlock.scala 173:23]
  wire [2:0] rob_io_commits_info_1_commitType; // @[CtrlBlock.scala 173:23]
  wire [5:0] rob_io_commits_info_1_pdest; // @[CtrlBlock.scala 173:23]
  wire [5:0] rob_io_commits_info_1_old_pdest; // @[CtrlBlock.scala 173:23]
  wire  rob_io_commits_info_1_ftqIdx_flag; // @[CtrlBlock.scala 173:23]
  wire [2:0] rob_io_commits_info_1_ftqIdx_value; // @[CtrlBlock.scala 173:23]
  wire [2:0] rob_io_commits_info_1_ftqOffset; // @[CtrlBlock.scala 173:23]
  wire  rob_io_commits_info_1_isMove; // @[CtrlBlock.scala 173:23]
  wire [1:0] rob_io_lsq_scommit; // @[CtrlBlock.scala 173:23]
  wire  rob_io_lsq_pendingld; // @[CtrlBlock.scala 173:23]
  wire  rob_io_lsq_pendingst; // @[CtrlBlock.scala 173:23]
  wire  rob_io_lsq_commit; // @[CtrlBlock.scala 173:23]
  wire  rob_io_lsq_isMMIO_0; // @[CtrlBlock.scala 173:23]
  wire  rob_io_lsq_isMMIO_1; // @[CtrlBlock.scala 173:23]
  wire [4:0] rob_io_lsq_uop_0_robIdx_value; // @[CtrlBlock.scala 173:23]
  wire [4:0] rob_io_lsq_uop_1_robIdx_value; // @[CtrlBlock.scala 173:23]
  wire  rob_io_csr_intrBitSet; // @[CtrlBlock.scala 173:23]
  wire  rob_io_csr_wfiEvent; // @[CtrlBlock.scala 173:23]
  wire  rob_io_csr_fflags_valid; // @[CtrlBlock.scala 173:23]
  wire [4:0] rob_io_csr_fflags_bits; // @[CtrlBlock.scala 173:23]
  wire  rob_io_csr_dirty_fs; // @[CtrlBlock.scala 173:23]
  wire [2:0] rob_io_csr_perfinfo_retiredInstr; // @[CtrlBlock.scala 173:23]
  wire  rob_io_cpu_halt; // @[CtrlBlock.scala 173:23]
  wire  rob_io_wfi_enable; // @[CtrlBlock.scala 173:23]
  wire [5:0] rob_io_perf_0_value; // @[CtrlBlock.scala 173:23]
  wire [5:0] rob_io_perf_1_value; // @[CtrlBlock.scala 173:23]
  wire [5:0] rob_io_perf_2_value; // @[CtrlBlock.scala 173:23]
  wire [5:0] rob_io_perf_3_value; // @[CtrlBlock.scala 173:23]
  wire [5:0] rob_io_perf_4_value; // @[CtrlBlock.scala 173:23]
  wire [5:0] rob_io_perf_5_value; // @[CtrlBlock.scala 173:23]
  wire [5:0] rob_io_perf_6_value; // @[CtrlBlock.scala 173:23]
  wire [5:0] rob_io_perf_7_value; // @[CtrlBlock.scala 173:23]
  wire [5:0] rob_io_perf_8_value; // @[CtrlBlock.scala 173:23]
  wire [5:0] rob_io_perf_9_value; // @[CtrlBlock.scala 173:23]
  wire [5:0] rob_io_perf_10_value; // @[CtrlBlock.scala 173:23]
  wire [5:0] rob_io_perf_11_value; // @[CtrlBlock.scala 173:23]
  wire [5:0] rob_io_perf_12_value; // @[CtrlBlock.scala 173:23]
  wire [5:0] rob_io_perf_13_value; // @[CtrlBlock.scala 173:23]
  wire [5:0] rob_io_perf_14_value; // @[CtrlBlock.scala 173:23]
  wire [5:0] rob_io_perf_15_value; // @[CtrlBlock.scala 173:23]
  wire [5:0] rob_io_perf_16_value; // @[CtrlBlock.scala 173:23]
  wire [5:0] rob_io_perf_17_value; // @[CtrlBlock.scala 173:23]
  wire  dispatch2_io_in_0_ready; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_io_in_1_ready; // @[CtrlBlock.scala 181:51]
  wire [3:0] dispatch2_io_in_1_bits_ctrl_fuType; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_io_out_0_ready; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_io_out_1_ready; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_clock; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_reset; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_redirect_valid; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_redirect_bits_robIdx_flag; // @[CtrlBlock.scala 181:51]
  wire [4:0] dispatch2_1_io_redirect_bits_robIdx_value; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_redirect_bits_level; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_in_0_ready; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_in_0_valid; // @[CtrlBlock.scala 181:51]
  wire [9:0] dispatch2_1_io_in_0_bits_cf_foldpc; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_in_0_bits_cf_trigger_backendEn_0; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_in_0_bits_cf_trigger_backendEn_1; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_in_0_bits_cf_pd_isRVC; // @[CtrlBlock.scala 181:51]
  wire [1:0] dispatch2_1_io_in_0_bits_cf_pd_brType; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_in_0_bits_cf_pd_isCall; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_in_0_bits_cf_pd_isRet; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_in_0_bits_cf_pred_taken; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_in_0_bits_cf_storeSetHit; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_in_0_bits_cf_waitForRobIdx_flag; // @[CtrlBlock.scala 181:51]
  wire [4:0] dispatch2_1_io_in_0_bits_cf_waitForRobIdx_value; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_in_0_bits_cf_loadWaitBit; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_in_0_bits_cf_loadWaitStrict; // @[CtrlBlock.scala 181:51]
  wire [4:0] dispatch2_1_io_in_0_bits_cf_ssid; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_in_0_bits_cf_ftqPtr_flag; // @[CtrlBlock.scala 181:51]
  wire [2:0] dispatch2_1_io_in_0_bits_cf_ftqPtr_value; // @[CtrlBlock.scala 181:51]
  wire [2:0] dispatch2_1_io_in_0_bits_cf_ftqOffset; // @[CtrlBlock.scala 181:51]
  wire [1:0] dispatch2_1_io_in_0_bits_ctrl_srcType_0; // @[CtrlBlock.scala 181:51]
  wire [1:0] dispatch2_1_io_in_0_bits_ctrl_srcType_1; // @[CtrlBlock.scala 181:51]
  wire [3:0] dispatch2_1_io_in_0_bits_ctrl_fuType; // @[CtrlBlock.scala 181:51]
  wire [6:0] dispatch2_1_io_in_0_bits_ctrl_fuOpType; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_in_0_bits_ctrl_rfWen; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_in_0_bits_ctrl_fpWen; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_in_0_bits_ctrl_flushPipe; // @[CtrlBlock.scala 181:51]
  wire [19:0] dispatch2_1_io_in_0_bits_ctrl_imm; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_in_0_bits_ctrl_replayInst; // @[CtrlBlock.scala 181:51]
  wire [5:0] dispatch2_1_io_in_0_bits_psrc_0; // @[CtrlBlock.scala 181:51]
  wire [5:0] dispatch2_1_io_in_0_bits_psrc_1; // @[CtrlBlock.scala 181:51]
  wire [5:0] dispatch2_1_io_in_0_bits_pdest; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_in_0_bits_robIdx_flag; // @[CtrlBlock.scala 181:51]
  wire [4:0] dispatch2_1_io_in_0_bits_robIdx_value; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_in_1_ready; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_in_1_valid; // @[CtrlBlock.scala 181:51]
  wire [9:0] dispatch2_1_io_in_1_bits_cf_foldpc; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_in_1_bits_cf_trigger_backendEn_0; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_in_1_bits_cf_trigger_backendEn_1; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_in_1_bits_cf_pd_isRVC; // @[CtrlBlock.scala 181:51]
  wire [1:0] dispatch2_1_io_in_1_bits_cf_pd_brType; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_in_1_bits_cf_pd_isCall; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_in_1_bits_cf_pd_isRet; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_in_1_bits_cf_pred_taken; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_in_1_bits_cf_storeSetHit; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_in_1_bits_cf_waitForRobIdx_flag; // @[CtrlBlock.scala 181:51]
  wire [4:0] dispatch2_1_io_in_1_bits_cf_waitForRobIdx_value; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_in_1_bits_cf_loadWaitBit; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_in_1_bits_cf_loadWaitStrict; // @[CtrlBlock.scala 181:51]
  wire [4:0] dispatch2_1_io_in_1_bits_cf_ssid; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_in_1_bits_cf_ftqPtr_flag; // @[CtrlBlock.scala 181:51]
  wire [2:0] dispatch2_1_io_in_1_bits_cf_ftqPtr_value; // @[CtrlBlock.scala 181:51]
  wire [2:0] dispatch2_1_io_in_1_bits_cf_ftqOffset; // @[CtrlBlock.scala 181:51]
  wire [1:0] dispatch2_1_io_in_1_bits_ctrl_srcType_0; // @[CtrlBlock.scala 181:51]
  wire [1:0] dispatch2_1_io_in_1_bits_ctrl_srcType_1; // @[CtrlBlock.scala 181:51]
  wire [3:0] dispatch2_1_io_in_1_bits_ctrl_fuType; // @[CtrlBlock.scala 181:51]
  wire [6:0] dispatch2_1_io_in_1_bits_ctrl_fuOpType; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_in_1_bits_ctrl_rfWen; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_in_1_bits_ctrl_fpWen; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_in_1_bits_ctrl_flushPipe; // @[CtrlBlock.scala 181:51]
  wire [19:0] dispatch2_1_io_in_1_bits_ctrl_imm; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_in_1_bits_ctrl_replayInst; // @[CtrlBlock.scala 181:51]
  wire [5:0] dispatch2_1_io_in_1_bits_psrc_0; // @[CtrlBlock.scala 181:51]
  wire [5:0] dispatch2_1_io_in_1_bits_psrc_1; // @[CtrlBlock.scala 181:51]
  wire [5:0] dispatch2_1_io_in_1_bits_pdest; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_in_1_bits_robIdx_flag; // @[CtrlBlock.scala 181:51]
  wire [4:0] dispatch2_1_io_in_1_bits_robIdx_value; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_in_2_ready; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_in_2_valid; // @[CtrlBlock.scala 181:51]
  wire [9:0] dispatch2_1_io_in_2_bits_cf_foldpc; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_in_2_bits_cf_trigger_backendEn_0; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_in_2_bits_cf_trigger_backendEn_1; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_in_2_bits_cf_pd_isRVC; // @[CtrlBlock.scala 181:51]
  wire [1:0] dispatch2_1_io_in_2_bits_cf_pd_brType; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_in_2_bits_cf_pd_isCall; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_in_2_bits_cf_pd_isRet; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_in_2_bits_cf_pred_taken; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_in_2_bits_cf_storeSetHit; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_in_2_bits_cf_waitForRobIdx_flag; // @[CtrlBlock.scala 181:51]
  wire [4:0] dispatch2_1_io_in_2_bits_cf_waitForRobIdx_value; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_in_2_bits_cf_loadWaitBit; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_in_2_bits_cf_loadWaitStrict; // @[CtrlBlock.scala 181:51]
  wire [4:0] dispatch2_1_io_in_2_bits_cf_ssid; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_in_2_bits_cf_ftqPtr_flag; // @[CtrlBlock.scala 181:51]
  wire [2:0] dispatch2_1_io_in_2_bits_cf_ftqPtr_value; // @[CtrlBlock.scala 181:51]
  wire [2:0] dispatch2_1_io_in_2_bits_cf_ftqOffset; // @[CtrlBlock.scala 181:51]
  wire [1:0] dispatch2_1_io_in_2_bits_ctrl_srcType_0; // @[CtrlBlock.scala 181:51]
  wire [1:0] dispatch2_1_io_in_2_bits_ctrl_srcType_1; // @[CtrlBlock.scala 181:51]
  wire [3:0] dispatch2_1_io_in_2_bits_ctrl_fuType; // @[CtrlBlock.scala 181:51]
  wire [6:0] dispatch2_1_io_in_2_bits_ctrl_fuOpType; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_in_2_bits_ctrl_rfWen; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_in_2_bits_ctrl_fpWen; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_in_2_bits_ctrl_flushPipe; // @[CtrlBlock.scala 181:51]
  wire [19:0] dispatch2_1_io_in_2_bits_ctrl_imm; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_in_2_bits_ctrl_replayInst; // @[CtrlBlock.scala 181:51]
  wire [5:0] dispatch2_1_io_in_2_bits_psrc_0; // @[CtrlBlock.scala 181:51]
  wire [5:0] dispatch2_1_io_in_2_bits_psrc_1; // @[CtrlBlock.scala 181:51]
  wire [5:0] dispatch2_1_io_in_2_bits_pdest; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_in_2_bits_robIdx_flag; // @[CtrlBlock.scala 181:51]
  wire [4:0] dispatch2_1_io_in_2_bits_robIdx_value; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_in_3_ready; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_in_3_valid; // @[CtrlBlock.scala 181:51]
  wire [9:0] dispatch2_1_io_in_3_bits_cf_foldpc; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_in_3_bits_cf_trigger_backendEn_0; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_in_3_bits_cf_trigger_backendEn_1; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_in_3_bits_cf_pd_isRVC; // @[CtrlBlock.scala 181:51]
  wire [1:0] dispatch2_1_io_in_3_bits_cf_pd_brType; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_in_3_bits_cf_pd_isCall; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_in_3_bits_cf_pd_isRet; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_in_3_bits_cf_pred_taken; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_in_3_bits_cf_storeSetHit; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_in_3_bits_cf_waitForRobIdx_flag; // @[CtrlBlock.scala 181:51]
  wire [4:0] dispatch2_1_io_in_3_bits_cf_waitForRobIdx_value; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_in_3_bits_cf_loadWaitBit; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_in_3_bits_cf_loadWaitStrict; // @[CtrlBlock.scala 181:51]
  wire [4:0] dispatch2_1_io_in_3_bits_cf_ssid; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_in_3_bits_cf_ftqPtr_flag; // @[CtrlBlock.scala 181:51]
  wire [2:0] dispatch2_1_io_in_3_bits_cf_ftqPtr_value; // @[CtrlBlock.scala 181:51]
  wire [2:0] dispatch2_1_io_in_3_bits_cf_ftqOffset; // @[CtrlBlock.scala 181:51]
  wire [1:0] dispatch2_1_io_in_3_bits_ctrl_srcType_0; // @[CtrlBlock.scala 181:51]
  wire [1:0] dispatch2_1_io_in_3_bits_ctrl_srcType_1; // @[CtrlBlock.scala 181:51]
  wire [3:0] dispatch2_1_io_in_3_bits_ctrl_fuType; // @[CtrlBlock.scala 181:51]
  wire [6:0] dispatch2_1_io_in_3_bits_ctrl_fuOpType; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_in_3_bits_ctrl_rfWen; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_in_3_bits_ctrl_fpWen; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_in_3_bits_ctrl_flushPipe; // @[CtrlBlock.scala 181:51]
  wire [19:0] dispatch2_1_io_in_3_bits_ctrl_imm; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_in_3_bits_ctrl_replayInst; // @[CtrlBlock.scala 181:51]
  wire [5:0] dispatch2_1_io_in_3_bits_psrc_0; // @[CtrlBlock.scala 181:51]
  wire [5:0] dispatch2_1_io_in_3_bits_psrc_1; // @[CtrlBlock.scala 181:51]
  wire [5:0] dispatch2_1_io_in_3_bits_pdest; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_in_3_bits_robIdx_flag; // @[CtrlBlock.scala 181:51]
  wire [4:0] dispatch2_1_io_in_3_bits_robIdx_value; // @[CtrlBlock.scala 181:51]
  wire [5:0] dispatch2_1_io_readIntState_0_req; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_readIntState_0_resp; // @[CtrlBlock.scala 181:51]
  wire [5:0] dispatch2_1_io_readIntState_1_req; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_readIntState_1_resp; // @[CtrlBlock.scala 181:51]
  wire [5:0] dispatch2_1_io_readIntState_2_req; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_readIntState_2_resp; // @[CtrlBlock.scala 181:51]
  wire [5:0] dispatch2_1_io_readIntState_3_req; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_readIntState_3_resp; // @[CtrlBlock.scala 181:51]
  wire [5:0] dispatch2_1_io_readIntState_4_req; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_readIntState_4_resp; // @[CtrlBlock.scala 181:51]
  wire [5:0] dispatch2_1_io_readIntState_5_req; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_readIntState_5_resp; // @[CtrlBlock.scala 181:51]
  wire [5:0] dispatch2_1_io_readFpState_0_req; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_readFpState_0_resp; // @[CtrlBlock.scala 181:51]
  wire [5:0] dispatch2_1_io_readFpState_1_req; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_readFpState_1_resp; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_0_ready; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_0_valid; // @[CtrlBlock.scala 181:51]
  wire [9:0] dispatch2_1_io_out_0_bits_cf_foldpc; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_0_bits_cf_trigger_backendEn_0; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_0_bits_cf_trigger_backendEn_1; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_0_bits_cf_pd_isRVC; // @[CtrlBlock.scala 181:51]
  wire [1:0] dispatch2_1_io_out_0_bits_cf_pd_brType; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_0_bits_cf_pd_isCall; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_0_bits_cf_pd_isRet; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_0_bits_cf_pred_taken; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_0_bits_cf_storeSetHit; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_0_bits_cf_waitForRobIdx_flag; // @[CtrlBlock.scala 181:51]
  wire [4:0] dispatch2_1_io_out_0_bits_cf_waitForRobIdx_value; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_0_bits_cf_loadWaitBit; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_0_bits_cf_loadWaitStrict; // @[CtrlBlock.scala 181:51]
  wire [4:0] dispatch2_1_io_out_0_bits_cf_ssid; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_0_bits_cf_ftqPtr_flag; // @[CtrlBlock.scala 181:51]
  wire [2:0] dispatch2_1_io_out_0_bits_cf_ftqPtr_value; // @[CtrlBlock.scala 181:51]
  wire [2:0] dispatch2_1_io_out_0_bits_cf_ftqOffset; // @[CtrlBlock.scala 181:51]
  wire [1:0] dispatch2_1_io_out_0_bits_ctrl_srcType_0; // @[CtrlBlock.scala 181:51]
  wire [3:0] dispatch2_1_io_out_0_bits_ctrl_fuType; // @[CtrlBlock.scala 181:51]
  wire [6:0] dispatch2_1_io_out_0_bits_ctrl_fuOpType; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_0_bits_ctrl_rfWen; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_0_bits_ctrl_fpWen; // @[CtrlBlock.scala 181:51]
  wire [19:0] dispatch2_1_io_out_0_bits_ctrl_imm; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_0_bits_srcState_0; // @[CtrlBlock.scala 181:51]
  wire [5:0] dispatch2_1_io_out_0_bits_psrc_0; // @[CtrlBlock.scala 181:51]
  wire [5:0] dispatch2_1_io_out_0_bits_psrc_1; // @[CtrlBlock.scala 181:51]
  wire [5:0] dispatch2_1_io_out_0_bits_pdest; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_0_bits_robIdx_flag; // @[CtrlBlock.scala 181:51]
  wire [4:0] dispatch2_1_io_out_0_bits_robIdx_value; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_0_bits_lqIdx_flag; // @[CtrlBlock.scala 181:51]
  wire [3:0] dispatch2_1_io_out_0_bits_lqIdx_value; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_0_bits_sqIdx_flag; // @[CtrlBlock.scala 181:51]
  wire [3:0] dispatch2_1_io_out_0_bits_sqIdx_value; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_1_ready; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_1_valid; // @[CtrlBlock.scala 181:51]
  wire [9:0] dispatch2_1_io_out_1_bits_cf_foldpc; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_1_bits_cf_trigger_backendEn_0; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_1_bits_cf_trigger_backendEn_1; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_1_bits_cf_pd_isRVC; // @[CtrlBlock.scala 181:51]
  wire [1:0] dispatch2_1_io_out_1_bits_cf_pd_brType; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_1_bits_cf_pd_isCall; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_1_bits_cf_pd_isRet; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_1_bits_cf_pred_taken; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_1_bits_cf_storeSetHit; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_1_bits_cf_waitForRobIdx_flag; // @[CtrlBlock.scala 181:51]
  wire [4:0] dispatch2_1_io_out_1_bits_cf_waitForRobIdx_value; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_1_bits_cf_loadWaitBit; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_1_bits_cf_loadWaitStrict; // @[CtrlBlock.scala 181:51]
  wire [4:0] dispatch2_1_io_out_1_bits_cf_ssid; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_1_bits_cf_ftqPtr_flag; // @[CtrlBlock.scala 181:51]
  wire [2:0] dispatch2_1_io_out_1_bits_cf_ftqPtr_value; // @[CtrlBlock.scala 181:51]
  wire [2:0] dispatch2_1_io_out_1_bits_cf_ftqOffset; // @[CtrlBlock.scala 181:51]
  wire [1:0] dispatch2_1_io_out_1_bits_ctrl_srcType_0; // @[CtrlBlock.scala 181:51]
  wire [3:0] dispatch2_1_io_out_1_bits_ctrl_fuType; // @[CtrlBlock.scala 181:51]
  wire [6:0] dispatch2_1_io_out_1_bits_ctrl_fuOpType; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_1_bits_ctrl_rfWen; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_1_bits_ctrl_fpWen; // @[CtrlBlock.scala 181:51]
  wire [19:0] dispatch2_1_io_out_1_bits_ctrl_imm; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_1_bits_srcState_0; // @[CtrlBlock.scala 181:51]
  wire [5:0] dispatch2_1_io_out_1_bits_psrc_0; // @[CtrlBlock.scala 181:51]
  wire [5:0] dispatch2_1_io_out_1_bits_psrc_1; // @[CtrlBlock.scala 181:51]
  wire [5:0] dispatch2_1_io_out_1_bits_pdest; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_1_bits_robIdx_flag; // @[CtrlBlock.scala 181:51]
  wire [4:0] dispatch2_1_io_out_1_bits_robIdx_value; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_1_bits_lqIdx_flag; // @[CtrlBlock.scala 181:51]
  wire [3:0] dispatch2_1_io_out_1_bits_lqIdx_value; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_1_bits_sqIdx_flag; // @[CtrlBlock.scala 181:51]
  wire [3:0] dispatch2_1_io_out_1_bits_sqIdx_value; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_2_ready; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_2_valid; // @[CtrlBlock.scala 181:51]
  wire [9:0] dispatch2_1_io_out_2_bits_cf_foldpc; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_2_bits_cf_trigger_backendEn_0; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_2_bits_cf_trigger_backendEn_1; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_2_bits_cf_pd_isRVC; // @[CtrlBlock.scala 181:51]
  wire [1:0] dispatch2_1_io_out_2_bits_cf_pd_brType; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_2_bits_cf_pd_isCall; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_2_bits_cf_pd_isRet; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_2_bits_cf_pred_taken; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_2_bits_cf_storeSetHit; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_2_bits_cf_waitForRobIdx_flag; // @[CtrlBlock.scala 181:51]
  wire [4:0] dispatch2_1_io_out_2_bits_cf_waitForRobIdx_value; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_2_bits_cf_loadWaitBit; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_2_bits_cf_loadWaitStrict; // @[CtrlBlock.scala 181:51]
  wire [4:0] dispatch2_1_io_out_2_bits_cf_ssid; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_2_bits_cf_ftqPtr_flag; // @[CtrlBlock.scala 181:51]
  wire [2:0] dispatch2_1_io_out_2_bits_cf_ftqPtr_value; // @[CtrlBlock.scala 181:51]
  wire [2:0] dispatch2_1_io_out_2_bits_cf_ftqOffset; // @[CtrlBlock.scala 181:51]
  wire [1:0] dispatch2_1_io_out_2_bits_ctrl_srcType_0; // @[CtrlBlock.scala 181:51]
  wire [3:0] dispatch2_1_io_out_2_bits_ctrl_fuType; // @[CtrlBlock.scala 181:51]
  wire [6:0] dispatch2_1_io_out_2_bits_ctrl_fuOpType; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_2_bits_ctrl_rfWen; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_2_bits_ctrl_fpWen; // @[CtrlBlock.scala 181:51]
  wire [19:0] dispatch2_1_io_out_2_bits_ctrl_imm; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_2_bits_srcState_0; // @[CtrlBlock.scala 181:51]
  wire [5:0] dispatch2_1_io_out_2_bits_psrc_0; // @[CtrlBlock.scala 181:51]
  wire [5:0] dispatch2_1_io_out_2_bits_pdest; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_2_bits_robIdx_flag; // @[CtrlBlock.scala 181:51]
  wire [4:0] dispatch2_1_io_out_2_bits_robIdx_value; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_2_bits_lqIdx_flag; // @[CtrlBlock.scala 181:51]
  wire [3:0] dispatch2_1_io_out_2_bits_lqIdx_value; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_2_bits_sqIdx_flag; // @[CtrlBlock.scala 181:51]
  wire [3:0] dispatch2_1_io_out_2_bits_sqIdx_value; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_3_ready; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_3_valid; // @[CtrlBlock.scala 181:51]
  wire [9:0] dispatch2_1_io_out_3_bits_cf_foldpc; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_3_bits_cf_trigger_backendEn_0; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_3_bits_cf_trigger_backendEn_1; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_3_bits_cf_pd_isRVC; // @[CtrlBlock.scala 181:51]
  wire [1:0] dispatch2_1_io_out_3_bits_cf_pd_brType; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_3_bits_cf_pd_isCall; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_3_bits_cf_pd_isRet; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_3_bits_cf_pred_taken; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_3_bits_cf_storeSetHit; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_3_bits_cf_waitForRobIdx_flag; // @[CtrlBlock.scala 181:51]
  wire [4:0] dispatch2_1_io_out_3_bits_cf_waitForRobIdx_value; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_3_bits_cf_loadWaitBit; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_3_bits_cf_loadWaitStrict; // @[CtrlBlock.scala 181:51]
  wire [4:0] dispatch2_1_io_out_3_bits_cf_ssid; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_3_bits_cf_ftqPtr_flag; // @[CtrlBlock.scala 181:51]
  wire [2:0] dispatch2_1_io_out_3_bits_cf_ftqPtr_value; // @[CtrlBlock.scala 181:51]
  wire [2:0] dispatch2_1_io_out_3_bits_cf_ftqOffset; // @[CtrlBlock.scala 181:51]
  wire [1:0] dispatch2_1_io_out_3_bits_ctrl_srcType_0; // @[CtrlBlock.scala 181:51]
  wire [3:0] dispatch2_1_io_out_3_bits_ctrl_fuType; // @[CtrlBlock.scala 181:51]
  wire [6:0] dispatch2_1_io_out_3_bits_ctrl_fuOpType; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_3_bits_ctrl_rfWen; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_3_bits_ctrl_fpWen; // @[CtrlBlock.scala 181:51]
  wire [19:0] dispatch2_1_io_out_3_bits_ctrl_imm; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_3_bits_srcState_0; // @[CtrlBlock.scala 181:51]
  wire [5:0] dispatch2_1_io_out_3_bits_psrc_0; // @[CtrlBlock.scala 181:51]
  wire [5:0] dispatch2_1_io_out_3_bits_pdest; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_3_bits_robIdx_flag; // @[CtrlBlock.scala 181:51]
  wire [4:0] dispatch2_1_io_out_3_bits_robIdx_value; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_3_bits_lqIdx_flag; // @[CtrlBlock.scala 181:51]
  wire [3:0] dispatch2_1_io_out_3_bits_lqIdx_value; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_3_bits_sqIdx_flag; // @[CtrlBlock.scala 181:51]
  wire [3:0] dispatch2_1_io_out_3_bits_sqIdx_value; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_4_ready; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_4_valid; // @[CtrlBlock.scala 181:51]
  wire [9:0] dispatch2_1_io_out_4_bits_cf_foldpc; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_4_bits_cf_trigger_backendEn_0; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_4_bits_cf_trigger_backendEn_1; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_4_bits_cf_pd_isRVC; // @[CtrlBlock.scala 181:51]
  wire [1:0] dispatch2_1_io_out_4_bits_cf_pd_brType; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_4_bits_cf_pd_isCall; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_4_bits_cf_pd_isRet; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_4_bits_cf_pred_taken; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_4_bits_cf_storeSetHit; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_4_bits_cf_waitForRobIdx_flag; // @[CtrlBlock.scala 181:51]
  wire [4:0] dispatch2_1_io_out_4_bits_cf_waitForRobIdx_value; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_4_bits_cf_loadWaitBit; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_4_bits_cf_loadWaitStrict; // @[CtrlBlock.scala 181:51]
  wire [4:0] dispatch2_1_io_out_4_bits_cf_ssid; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_4_bits_cf_ftqPtr_flag; // @[CtrlBlock.scala 181:51]
  wire [2:0] dispatch2_1_io_out_4_bits_cf_ftqPtr_value; // @[CtrlBlock.scala 181:51]
  wire [2:0] dispatch2_1_io_out_4_bits_cf_ftqOffset; // @[CtrlBlock.scala 181:51]
  wire [1:0] dispatch2_1_io_out_4_bits_ctrl_srcType_0; // @[CtrlBlock.scala 181:51]
  wire [3:0] dispatch2_1_io_out_4_bits_ctrl_fuType; // @[CtrlBlock.scala 181:51]
  wire [6:0] dispatch2_1_io_out_4_bits_ctrl_fuOpType; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_4_bits_ctrl_rfWen; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_4_bits_ctrl_fpWen; // @[CtrlBlock.scala 181:51]
  wire [19:0] dispatch2_1_io_out_4_bits_ctrl_imm; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_4_bits_srcState_0; // @[CtrlBlock.scala 181:51]
  wire [5:0] dispatch2_1_io_out_4_bits_psrc_0; // @[CtrlBlock.scala 181:51]
  wire [5:0] dispatch2_1_io_out_4_bits_pdest; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_4_bits_robIdx_flag; // @[CtrlBlock.scala 181:51]
  wire [4:0] dispatch2_1_io_out_4_bits_robIdx_value; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_4_bits_lqIdx_flag; // @[CtrlBlock.scala 181:51]
  wire [3:0] dispatch2_1_io_out_4_bits_lqIdx_value; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_4_bits_sqIdx_flag; // @[CtrlBlock.scala 181:51]
  wire [3:0] dispatch2_1_io_out_4_bits_sqIdx_value; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_5_ready; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_5_valid; // @[CtrlBlock.scala 181:51]
  wire [9:0] dispatch2_1_io_out_5_bits_cf_foldpc; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_5_bits_cf_trigger_backendEn_0; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_5_bits_cf_trigger_backendEn_1; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_5_bits_cf_pd_isRVC; // @[CtrlBlock.scala 181:51]
  wire [1:0] dispatch2_1_io_out_5_bits_cf_pd_brType; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_5_bits_cf_pd_isCall; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_5_bits_cf_pd_isRet; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_5_bits_cf_pred_taken; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_5_bits_cf_storeSetHit; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_5_bits_cf_waitForRobIdx_flag; // @[CtrlBlock.scala 181:51]
  wire [4:0] dispatch2_1_io_out_5_bits_cf_waitForRobIdx_value; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_5_bits_cf_loadWaitBit; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_5_bits_cf_loadWaitStrict; // @[CtrlBlock.scala 181:51]
  wire [4:0] dispatch2_1_io_out_5_bits_cf_ssid; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_5_bits_cf_ftqPtr_flag; // @[CtrlBlock.scala 181:51]
  wire [2:0] dispatch2_1_io_out_5_bits_cf_ftqPtr_value; // @[CtrlBlock.scala 181:51]
  wire [2:0] dispatch2_1_io_out_5_bits_cf_ftqOffset; // @[CtrlBlock.scala 181:51]
  wire [1:0] dispatch2_1_io_out_5_bits_ctrl_srcType_0; // @[CtrlBlock.scala 181:51]
  wire [3:0] dispatch2_1_io_out_5_bits_ctrl_fuType; // @[CtrlBlock.scala 181:51]
  wire [6:0] dispatch2_1_io_out_5_bits_ctrl_fuOpType; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_5_bits_ctrl_rfWen; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_5_bits_ctrl_fpWen; // @[CtrlBlock.scala 181:51]
  wire [19:0] dispatch2_1_io_out_5_bits_ctrl_imm; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_5_bits_srcState_0; // @[CtrlBlock.scala 181:51]
  wire [5:0] dispatch2_1_io_out_5_bits_psrc_0; // @[CtrlBlock.scala 181:51]
  wire [5:0] dispatch2_1_io_out_5_bits_pdest; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_5_bits_robIdx_flag; // @[CtrlBlock.scala 181:51]
  wire [4:0] dispatch2_1_io_out_5_bits_robIdx_value; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_5_bits_lqIdx_flag; // @[CtrlBlock.scala 181:51]
  wire [3:0] dispatch2_1_io_out_5_bits_lqIdx_value; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_out_5_bits_sqIdx_flag; // @[CtrlBlock.scala 181:51]
  wire [3:0] dispatch2_1_io_out_5_bits_sqIdx_value; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_enqLsq_canAccept; // @[CtrlBlock.scala 181:51]
  wire [1:0] dispatch2_1_io_enqLsq_needAlloc_0; // @[CtrlBlock.scala 181:51]
  wire [1:0] dispatch2_1_io_enqLsq_needAlloc_1; // @[CtrlBlock.scala 181:51]
  wire [1:0] dispatch2_1_io_enqLsq_needAlloc_2; // @[CtrlBlock.scala 181:51]
  wire [1:0] dispatch2_1_io_enqLsq_needAlloc_3; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_enqLsq_req_0_valid; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_enqLsq_req_0_bits_cf_trigger_backendEn_0; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_enqLsq_req_0_bits_cf_trigger_backendEn_1; // @[CtrlBlock.scala 181:51]
  wire [6:0] dispatch2_1_io_enqLsq_req_0_bits_ctrl_fuOpType; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_enqLsq_req_0_bits_ctrl_rfWen; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_enqLsq_req_0_bits_ctrl_fpWen; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_enqLsq_req_0_bits_ctrl_flushPipe; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_enqLsq_req_0_bits_ctrl_replayInst; // @[CtrlBlock.scala 181:51]
  wire [5:0] dispatch2_1_io_enqLsq_req_0_bits_pdest; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_enqLsq_req_0_bits_robIdx_flag; // @[CtrlBlock.scala 181:51]
  wire [4:0] dispatch2_1_io_enqLsq_req_0_bits_robIdx_value; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_enqLsq_req_1_valid; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_enqLsq_req_1_bits_cf_trigger_backendEn_0; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_enqLsq_req_1_bits_cf_trigger_backendEn_1; // @[CtrlBlock.scala 181:51]
  wire [6:0] dispatch2_1_io_enqLsq_req_1_bits_ctrl_fuOpType; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_enqLsq_req_1_bits_ctrl_rfWen; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_enqLsq_req_1_bits_ctrl_fpWen; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_enqLsq_req_1_bits_ctrl_flushPipe; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_enqLsq_req_1_bits_ctrl_replayInst; // @[CtrlBlock.scala 181:51]
  wire [5:0] dispatch2_1_io_enqLsq_req_1_bits_pdest; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_enqLsq_req_1_bits_robIdx_flag; // @[CtrlBlock.scala 181:51]
  wire [4:0] dispatch2_1_io_enqLsq_req_1_bits_robIdx_value; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_enqLsq_req_2_valid; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_enqLsq_req_2_bits_cf_trigger_backendEn_0; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_enqLsq_req_2_bits_cf_trigger_backendEn_1; // @[CtrlBlock.scala 181:51]
  wire [6:0] dispatch2_1_io_enqLsq_req_2_bits_ctrl_fuOpType; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_enqLsq_req_2_bits_ctrl_rfWen; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_enqLsq_req_2_bits_ctrl_fpWen; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_enqLsq_req_2_bits_ctrl_flushPipe; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_enqLsq_req_2_bits_ctrl_replayInst; // @[CtrlBlock.scala 181:51]
  wire [5:0] dispatch2_1_io_enqLsq_req_2_bits_pdest; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_enqLsq_req_2_bits_robIdx_flag; // @[CtrlBlock.scala 181:51]
  wire [4:0] dispatch2_1_io_enqLsq_req_2_bits_robIdx_value; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_enqLsq_req_3_valid; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_enqLsq_req_3_bits_cf_trigger_backendEn_0; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_enqLsq_req_3_bits_cf_trigger_backendEn_1; // @[CtrlBlock.scala 181:51]
  wire [6:0] dispatch2_1_io_enqLsq_req_3_bits_ctrl_fuOpType; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_enqLsq_req_3_bits_ctrl_rfWen; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_enqLsq_req_3_bits_ctrl_fpWen; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_enqLsq_req_3_bits_ctrl_flushPipe; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_enqLsq_req_3_bits_ctrl_replayInst; // @[CtrlBlock.scala 181:51]
  wire [5:0] dispatch2_1_io_enqLsq_req_3_bits_pdest; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_enqLsq_req_3_bits_robIdx_flag; // @[CtrlBlock.scala 181:51]
  wire [4:0] dispatch2_1_io_enqLsq_req_3_bits_robIdx_value; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_enqLsq_resp_0_lqIdx_flag; // @[CtrlBlock.scala 181:51]
  wire [3:0] dispatch2_1_io_enqLsq_resp_0_lqIdx_value; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_enqLsq_resp_0_sqIdx_flag; // @[CtrlBlock.scala 181:51]
  wire [3:0] dispatch2_1_io_enqLsq_resp_0_sqIdx_value; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_enqLsq_resp_1_lqIdx_flag; // @[CtrlBlock.scala 181:51]
  wire [3:0] dispatch2_1_io_enqLsq_resp_1_lqIdx_value; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_enqLsq_resp_1_sqIdx_flag; // @[CtrlBlock.scala 181:51]
  wire [3:0] dispatch2_1_io_enqLsq_resp_1_sqIdx_value; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_enqLsq_resp_2_lqIdx_flag; // @[CtrlBlock.scala 181:51]
  wire [3:0] dispatch2_1_io_enqLsq_resp_2_lqIdx_value; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_enqLsq_resp_2_sqIdx_flag; // @[CtrlBlock.scala 181:51]
  wire [3:0] dispatch2_1_io_enqLsq_resp_2_sqIdx_value; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_enqLsq_resp_3_lqIdx_flag; // @[CtrlBlock.scala 181:51]
  wire [3:0] dispatch2_1_io_enqLsq_resp_3_lqIdx_value; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_1_io_enqLsq_resp_3_sqIdx_flag; // @[CtrlBlock.scala 181:51]
  wire [3:0] dispatch2_1_io_enqLsq_resp_3_sqIdx_value; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_2_io_in_0_ready; // @[CtrlBlock.scala 181:51]
  wire  dispatch2_2_io_out_0_ready; // @[CtrlBlock.scala 181:51]
  wire  decode_clock; // @[CtrlBlock.scala 263:22]
  wire  decode_io_in_0_ready; // @[CtrlBlock.scala 263:22]
  wire  decode_io_in_0_valid; // @[CtrlBlock.scala 263:22]
  wire [31:0] decode_io_in_0_bits_instr; // @[CtrlBlock.scala 263:22]
  wire [9:0] decode_io_in_0_bits_foldpc; // @[CtrlBlock.scala 263:22]
  wire  decode_io_in_0_bits_exceptionVec_1; // @[CtrlBlock.scala 263:22]
  wire  decode_io_in_0_bits_exceptionVec_12; // @[CtrlBlock.scala 263:22]
  wire  decode_io_in_0_bits_trigger_frontendHit_0; // @[CtrlBlock.scala 263:22]
  wire  decode_io_in_0_bits_trigger_frontendHit_1; // @[CtrlBlock.scala 263:22]
  wire  decode_io_in_0_bits_trigger_frontendHit_2; // @[CtrlBlock.scala 263:22]
  wire  decode_io_in_0_bits_trigger_frontendHit_3; // @[CtrlBlock.scala 263:22]
  wire  decode_io_in_0_bits_trigger_backendEn_0; // @[CtrlBlock.scala 263:22]
  wire  decode_io_in_0_bits_trigger_backendEn_1; // @[CtrlBlock.scala 263:22]
  wire  decode_io_in_0_bits_pd_isRVC; // @[CtrlBlock.scala 263:22]
  wire [1:0] decode_io_in_0_bits_pd_brType; // @[CtrlBlock.scala 263:22]
  wire  decode_io_in_0_bits_pd_isCall; // @[CtrlBlock.scala 263:22]
  wire  decode_io_in_0_bits_pd_isRet; // @[CtrlBlock.scala 263:22]
  wire  decode_io_in_0_bits_pred_taken; // @[CtrlBlock.scala 263:22]
  wire  decode_io_in_0_bits_crossPageIPFFix; // @[CtrlBlock.scala 263:22]
  wire  decode_io_in_0_bits_ftqPtr_flag; // @[CtrlBlock.scala 263:22]
  wire [2:0] decode_io_in_0_bits_ftqPtr_value; // @[CtrlBlock.scala 263:22]
  wire [2:0] decode_io_in_0_bits_ftqOffset; // @[CtrlBlock.scala 263:22]
  wire  decode_io_in_1_ready; // @[CtrlBlock.scala 263:22]
  wire  decode_io_in_1_valid; // @[CtrlBlock.scala 263:22]
  wire [31:0] decode_io_in_1_bits_instr; // @[CtrlBlock.scala 263:22]
  wire [9:0] decode_io_in_1_bits_foldpc; // @[CtrlBlock.scala 263:22]
  wire  decode_io_in_1_bits_exceptionVec_1; // @[CtrlBlock.scala 263:22]
  wire  decode_io_in_1_bits_exceptionVec_12; // @[CtrlBlock.scala 263:22]
  wire  decode_io_in_1_bits_trigger_frontendHit_0; // @[CtrlBlock.scala 263:22]
  wire  decode_io_in_1_bits_trigger_frontendHit_1; // @[CtrlBlock.scala 263:22]
  wire  decode_io_in_1_bits_trigger_frontendHit_2; // @[CtrlBlock.scala 263:22]
  wire  decode_io_in_1_bits_trigger_frontendHit_3; // @[CtrlBlock.scala 263:22]
  wire  decode_io_in_1_bits_trigger_backendEn_0; // @[CtrlBlock.scala 263:22]
  wire  decode_io_in_1_bits_trigger_backendEn_1; // @[CtrlBlock.scala 263:22]
  wire  decode_io_in_1_bits_pd_isRVC; // @[CtrlBlock.scala 263:22]
  wire [1:0] decode_io_in_1_bits_pd_brType; // @[CtrlBlock.scala 263:22]
  wire  decode_io_in_1_bits_pd_isCall; // @[CtrlBlock.scala 263:22]
  wire  decode_io_in_1_bits_pd_isRet; // @[CtrlBlock.scala 263:22]
  wire  decode_io_in_1_bits_pred_taken; // @[CtrlBlock.scala 263:22]
  wire  decode_io_in_1_bits_crossPageIPFFix; // @[CtrlBlock.scala 263:22]
  wire  decode_io_in_1_bits_ftqPtr_flag; // @[CtrlBlock.scala 263:22]
  wire [2:0] decode_io_in_1_bits_ftqPtr_value; // @[CtrlBlock.scala 263:22]
  wire [2:0] decode_io_in_1_bits_ftqOffset; // @[CtrlBlock.scala 263:22]
  wire  decode_io_out_0_ready; // @[CtrlBlock.scala 263:22]
  wire  decode_io_out_0_valid; // @[CtrlBlock.scala 263:22]
  wire [9:0] decode_io_out_0_bits_cf_foldpc; // @[CtrlBlock.scala 263:22]
  wire  decode_io_out_0_bits_cf_exceptionVec_1; // @[CtrlBlock.scala 263:22]
  wire  decode_io_out_0_bits_cf_exceptionVec_2; // @[CtrlBlock.scala 263:22]
  wire  decode_io_out_0_bits_cf_exceptionVec_12; // @[CtrlBlock.scala 263:22]
  wire  decode_io_out_0_bits_cf_trigger_frontendHit_0; // @[CtrlBlock.scala 263:22]
  wire  decode_io_out_0_bits_cf_trigger_frontendHit_1; // @[CtrlBlock.scala 263:22]
  wire  decode_io_out_0_bits_cf_trigger_frontendHit_2; // @[CtrlBlock.scala 263:22]
  wire  decode_io_out_0_bits_cf_trigger_frontendHit_3; // @[CtrlBlock.scala 263:22]
  wire  decode_io_out_0_bits_cf_trigger_backendEn_0; // @[CtrlBlock.scala 263:22]
  wire  decode_io_out_0_bits_cf_trigger_backendEn_1; // @[CtrlBlock.scala 263:22]
  wire  decode_io_out_0_bits_cf_pd_isRVC; // @[CtrlBlock.scala 263:22]
  wire [1:0] decode_io_out_0_bits_cf_pd_brType; // @[CtrlBlock.scala 263:22]
  wire  decode_io_out_0_bits_cf_pd_isCall; // @[CtrlBlock.scala 263:22]
  wire  decode_io_out_0_bits_cf_pd_isRet; // @[CtrlBlock.scala 263:22]
  wire  decode_io_out_0_bits_cf_pred_taken; // @[CtrlBlock.scala 263:22]
  wire  decode_io_out_0_bits_cf_crossPageIPFFix; // @[CtrlBlock.scala 263:22]
  wire  decode_io_out_0_bits_cf_ftqPtr_flag; // @[CtrlBlock.scala 263:22]
  wire [2:0] decode_io_out_0_bits_cf_ftqPtr_value; // @[CtrlBlock.scala 263:22]
  wire [2:0] decode_io_out_0_bits_cf_ftqOffset; // @[CtrlBlock.scala 263:22]
  wire [1:0] decode_io_out_0_bits_ctrl_srcType_0; // @[CtrlBlock.scala 263:22]
  wire [1:0] decode_io_out_0_bits_ctrl_srcType_1; // @[CtrlBlock.scala 263:22]
  wire [1:0] decode_io_out_0_bits_ctrl_srcType_2; // @[CtrlBlock.scala 263:22]
  wire [4:0] decode_io_out_0_bits_ctrl_lsrc_0; // @[CtrlBlock.scala 263:22]
  wire [4:0] decode_io_out_0_bits_ctrl_lsrc_1; // @[CtrlBlock.scala 263:22]
  wire [4:0] decode_io_out_0_bits_ctrl_ldest; // @[CtrlBlock.scala 263:22]
  wire [3:0] decode_io_out_0_bits_ctrl_fuType; // @[CtrlBlock.scala 263:22]
  wire [6:0] decode_io_out_0_bits_ctrl_fuOpType; // @[CtrlBlock.scala 263:22]
  wire  decode_io_out_0_bits_ctrl_rfWen; // @[CtrlBlock.scala 263:22]
  wire  decode_io_out_0_bits_ctrl_fpWen; // @[CtrlBlock.scala 263:22]
  wire  decode_io_out_0_bits_ctrl_isXSTrap; // @[CtrlBlock.scala 263:22]
  wire  decode_io_out_0_bits_ctrl_noSpecExec; // @[CtrlBlock.scala 263:22]
  wire  decode_io_out_0_bits_ctrl_blockBackward; // @[CtrlBlock.scala 263:22]
  wire  decode_io_out_0_bits_ctrl_flushPipe; // @[CtrlBlock.scala 263:22]
  wire [3:0] decode_io_out_0_bits_ctrl_selImm; // @[CtrlBlock.scala 263:22]
  wire [19:0] decode_io_out_0_bits_ctrl_imm; // @[CtrlBlock.scala 263:22]
  wire  decode_io_out_0_bits_ctrl_fpu_isAddSub; // @[CtrlBlock.scala 263:22]
  wire  decode_io_out_0_bits_ctrl_fpu_typeTagIn; // @[CtrlBlock.scala 263:22]
  wire  decode_io_out_0_bits_ctrl_fpu_typeTagOut; // @[CtrlBlock.scala 263:22]
  wire  decode_io_out_0_bits_ctrl_fpu_fromInt; // @[CtrlBlock.scala 263:22]
  wire  decode_io_out_0_bits_ctrl_fpu_wflags; // @[CtrlBlock.scala 263:22]
  wire  decode_io_out_0_bits_ctrl_fpu_fpWen; // @[CtrlBlock.scala 263:22]
  wire [1:0] decode_io_out_0_bits_ctrl_fpu_fmaCmd; // @[CtrlBlock.scala 263:22]
  wire  decode_io_out_0_bits_ctrl_fpu_div; // @[CtrlBlock.scala 263:22]
  wire  decode_io_out_0_bits_ctrl_fpu_sqrt; // @[CtrlBlock.scala 263:22]
  wire  decode_io_out_0_bits_ctrl_fpu_fcvt; // @[CtrlBlock.scala 263:22]
  wire [1:0] decode_io_out_0_bits_ctrl_fpu_typ; // @[CtrlBlock.scala 263:22]
  wire [1:0] decode_io_out_0_bits_ctrl_fpu_fmt; // @[CtrlBlock.scala 263:22]
  wire  decode_io_out_0_bits_ctrl_fpu_ren3; // @[CtrlBlock.scala 263:22]
  wire [2:0] decode_io_out_0_bits_ctrl_fpu_rm; // @[CtrlBlock.scala 263:22]
  wire  decode_io_out_0_bits_ctrl_isMove; // @[CtrlBlock.scala 263:22]
  wire  decode_io_out_1_ready; // @[CtrlBlock.scala 263:22]
  wire  decode_io_out_1_valid; // @[CtrlBlock.scala 263:22]
  wire [9:0] decode_io_out_1_bits_cf_foldpc; // @[CtrlBlock.scala 263:22]
  wire  decode_io_out_1_bits_cf_exceptionVec_1; // @[CtrlBlock.scala 263:22]
  wire  decode_io_out_1_bits_cf_exceptionVec_2; // @[CtrlBlock.scala 263:22]
  wire  decode_io_out_1_bits_cf_exceptionVec_12; // @[CtrlBlock.scala 263:22]
  wire  decode_io_out_1_bits_cf_trigger_frontendHit_0; // @[CtrlBlock.scala 263:22]
  wire  decode_io_out_1_bits_cf_trigger_frontendHit_1; // @[CtrlBlock.scala 263:22]
  wire  decode_io_out_1_bits_cf_trigger_frontendHit_2; // @[CtrlBlock.scala 263:22]
  wire  decode_io_out_1_bits_cf_trigger_frontendHit_3; // @[CtrlBlock.scala 263:22]
  wire  decode_io_out_1_bits_cf_trigger_backendEn_0; // @[CtrlBlock.scala 263:22]
  wire  decode_io_out_1_bits_cf_trigger_backendEn_1; // @[CtrlBlock.scala 263:22]
  wire  decode_io_out_1_bits_cf_pd_isRVC; // @[CtrlBlock.scala 263:22]
  wire [1:0] decode_io_out_1_bits_cf_pd_brType; // @[CtrlBlock.scala 263:22]
  wire  decode_io_out_1_bits_cf_pd_isCall; // @[CtrlBlock.scala 263:22]
  wire  decode_io_out_1_bits_cf_pd_isRet; // @[CtrlBlock.scala 263:22]
  wire  decode_io_out_1_bits_cf_pred_taken; // @[CtrlBlock.scala 263:22]
  wire  decode_io_out_1_bits_cf_crossPageIPFFix; // @[CtrlBlock.scala 263:22]
  wire  decode_io_out_1_bits_cf_ftqPtr_flag; // @[CtrlBlock.scala 263:22]
  wire [2:0] decode_io_out_1_bits_cf_ftqPtr_value; // @[CtrlBlock.scala 263:22]
  wire [2:0] decode_io_out_1_bits_cf_ftqOffset; // @[CtrlBlock.scala 263:22]
  wire [1:0] decode_io_out_1_bits_ctrl_srcType_0; // @[CtrlBlock.scala 263:22]
  wire [1:0] decode_io_out_1_bits_ctrl_srcType_1; // @[CtrlBlock.scala 263:22]
  wire [1:0] decode_io_out_1_bits_ctrl_srcType_2; // @[CtrlBlock.scala 263:22]
  wire [4:0] decode_io_out_1_bits_ctrl_lsrc_0; // @[CtrlBlock.scala 263:22]
  wire [4:0] decode_io_out_1_bits_ctrl_lsrc_1; // @[CtrlBlock.scala 263:22]
  wire [4:0] decode_io_out_1_bits_ctrl_lsrc_2; // @[CtrlBlock.scala 263:22]
  wire [4:0] decode_io_out_1_bits_ctrl_ldest; // @[CtrlBlock.scala 263:22]
  wire [3:0] decode_io_out_1_bits_ctrl_fuType; // @[CtrlBlock.scala 263:22]
  wire [6:0] decode_io_out_1_bits_ctrl_fuOpType; // @[CtrlBlock.scala 263:22]
  wire  decode_io_out_1_bits_ctrl_rfWen; // @[CtrlBlock.scala 263:22]
  wire  decode_io_out_1_bits_ctrl_fpWen; // @[CtrlBlock.scala 263:22]
  wire  decode_io_out_1_bits_ctrl_isXSTrap; // @[CtrlBlock.scala 263:22]
  wire  decode_io_out_1_bits_ctrl_noSpecExec; // @[CtrlBlock.scala 263:22]
  wire  decode_io_out_1_bits_ctrl_blockBackward; // @[CtrlBlock.scala 263:22]
  wire  decode_io_out_1_bits_ctrl_flushPipe; // @[CtrlBlock.scala 263:22]
  wire [3:0] decode_io_out_1_bits_ctrl_selImm; // @[CtrlBlock.scala 263:22]
  wire [19:0] decode_io_out_1_bits_ctrl_imm; // @[CtrlBlock.scala 263:22]
  wire  decode_io_out_1_bits_ctrl_fpu_isAddSub; // @[CtrlBlock.scala 263:22]
  wire  decode_io_out_1_bits_ctrl_fpu_typeTagIn; // @[CtrlBlock.scala 263:22]
  wire  decode_io_out_1_bits_ctrl_fpu_typeTagOut; // @[CtrlBlock.scala 263:22]
  wire  decode_io_out_1_bits_ctrl_fpu_fromInt; // @[CtrlBlock.scala 263:22]
  wire  decode_io_out_1_bits_ctrl_fpu_wflags; // @[CtrlBlock.scala 263:22]
  wire  decode_io_out_1_bits_ctrl_fpu_fpWen; // @[CtrlBlock.scala 263:22]
  wire [1:0] decode_io_out_1_bits_ctrl_fpu_fmaCmd; // @[CtrlBlock.scala 263:22]
  wire  decode_io_out_1_bits_ctrl_fpu_div; // @[CtrlBlock.scala 263:22]
  wire  decode_io_out_1_bits_ctrl_fpu_sqrt; // @[CtrlBlock.scala 263:22]
  wire  decode_io_out_1_bits_ctrl_fpu_fcvt; // @[CtrlBlock.scala 263:22]
  wire [1:0] decode_io_out_1_bits_ctrl_fpu_typ; // @[CtrlBlock.scala 263:22]
  wire [1:0] decode_io_out_1_bits_ctrl_fpu_fmt; // @[CtrlBlock.scala 263:22]
  wire  decode_io_out_1_bits_ctrl_fpu_ren3; // @[CtrlBlock.scala 263:22]
  wire [2:0] decode_io_out_1_bits_ctrl_fpu_rm; // @[CtrlBlock.scala 263:22]
  wire  decode_io_out_1_bits_ctrl_isMove; // @[CtrlBlock.scala 263:22]
  wire  decode_io_intRat_0_0_hold; // @[CtrlBlock.scala 263:22]
  wire [4:0] decode_io_intRat_0_0_addr; // @[CtrlBlock.scala 263:22]
  wire  decode_io_intRat_0_1_hold; // @[CtrlBlock.scala 263:22]
  wire [4:0] decode_io_intRat_0_1_addr; // @[CtrlBlock.scala 263:22]
  wire  decode_io_intRat_0_2_hold; // @[CtrlBlock.scala 263:22]
  wire [4:0] decode_io_intRat_0_2_addr; // @[CtrlBlock.scala 263:22]
  wire  decode_io_intRat_1_0_hold; // @[CtrlBlock.scala 263:22]
  wire [4:0] decode_io_intRat_1_0_addr; // @[CtrlBlock.scala 263:22]
  wire  decode_io_intRat_1_1_hold; // @[CtrlBlock.scala 263:22]
  wire [4:0] decode_io_intRat_1_1_addr; // @[CtrlBlock.scala 263:22]
  wire  decode_io_intRat_1_2_hold; // @[CtrlBlock.scala 263:22]
  wire [4:0] decode_io_intRat_1_2_addr; // @[CtrlBlock.scala 263:22]
  wire  decode_io_fpRat_0_0_hold; // @[CtrlBlock.scala 263:22]
  wire [4:0] decode_io_fpRat_0_0_addr; // @[CtrlBlock.scala 263:22]
  wire  decode_io_fpRat_0_1_hold; // @[CtrlBlock.scala 263:22]
  wire [4:0] decode_io_fpRat_0_1_addr; // @[CtrlBlock.scala 263:22]
  wire  decode_io_fpRat_0_2_hold; // @[CtrlBlock.scala 263:22]
  wire [4:0] decode_io_fpRat_0_2_addr; // @[CtrlBlock.scala 263:22]
  wire  decode_io_fpRat_0_3_hold; // @[CtrlBlock.scala 263:22]
  wire [4:0] decode_io_fpRat_0_3_addr; // @[CtrlBlock.scala 263:22]
  wire  decode_io_fpRat_1_0_hold; // @[CtrlBlock.scala 263:22]
  wire [4:0] decode_io_fpRat_1_0_addr; // @[CtrlBlock.scala 263:22]
  wire  decode_io_fpRat_1_1_hold; // @[CtrlBlock.scala 263:22]
  wire [4:0] decode_io_fpRat_1_1_addr; // @[CtrlBlock.scala 263:22]
  wire  decode_io_fpRat_1_2_hold; // @[CtrlBlock.scala 263:22]
  wire [4:0] decode_io_fpRat_1_2_addr; // @[CtrlBlock.scala 263:22]
  wire  decode_io_fpRat_1_3_hold; // @[CtrlBlock.scala 263:22]
  wire [4:0] decode_io_fpRat_1_3_addr; // @[CtrlBlock.scala 263:22]
  wire  decode_io_csrCtrl_fusion_enable; // @[CtrlBlock.scala 263:22]
  wire  decode_io_csrCtrl_wfi_enable; // @[CtrlBlock.scala 263:22]
  wire  decode_io_csrCtrl_svinval_enable; // @[CtrlBlock.scala 263:22]
  wire  decode_io_csrCtrl_singlestep; // @[CtrlBlock.scala 263:22]
  wire  decode_io_fusion_0; // @[CtrlBlock.scala 263:22]
  wire [5:0] decode_io_perf_0_value; // @[CtrlBlock.scala 263:22]
  wire [5:0] decode_io_perf_1_value; // @[CtrlBlock.scala 263:22]
  wire [5:0] decode_io_perf_2_value; // @[CtrlBlock.scala 263:22]
  wire [5:0] decode_io_perf_3_value; // @[CtrlBlock.scala 263:22]
  wire  fusionDecoder_clock; // @[CtrlBlock.scala 264:29]
  wire  fusionDecoder_reset; // @[CtrlBlock.scala 264:29]
  wire  fusionDecoder_io_in_0_valid; // @[CtrlBlock.scala 264:29]
  wire [31:0] fusionDecoder_io_in_0_bits; // @[CtrlBlock.scala 264:29]
  wire  fusionDecoder_io_in_1_valid; // @[CtrlBlock.scala 264:29]
  wire [31:0] fusionDecoder_io_in_1_bits; // @[CtrlBlock.scala 264:29]
  wire  fusionDecoder_io_inReady_0; // @[CtrlBlock.scala 264:29]
  wire [6:0] fusionDecoder_io_dec_0_fuOpType; // @[CtrlBlock.scala 264:29]
  wire  fusionDecoder_io_out_0_valid; // @[CtrlBlock.scala 264:29]
  wire  fusionDecoder_io_out_0_bits_fuType_valid; // @[CtrlBlock.scala 264:29]
  wire  fusionDecoder_io_out_0_bits_fuOpType_valid; // @[CtrlBlock.scala 264:29]
  wire [6:0] fusionDecoder_io_out_0_bits_fuOpType_bits; // @[CtrlBlock.scala 264:29]
  wire  fusionDecoder_io_out_0_bits_lsrc2_valid; // @[CtrlBlock.scala 264:29]
  wire [4:0] fusionDecoder_io_out_0_bits_lsrc2_bits; // @[CtrlBlock.scala 264:29]
  wire  fusionDecoder_io_out_0_bits_src2Type_valid; // @[CtrlBlock.scala 264:29]
  wire  fusionDecoder_io_info_0_rs2FromRs1; // @[CtrlBlock.scala 264:29]
  wire  fusionDecoder_io_info_0_rs2FromRs2; // @[CtrlBlock.scala 264:29]
  wire  fusionDecoder_io_info_0_rs2FromZero; // @[CtrlBlock.scala 264:29]
  wire  fusionDecoder_io_clear_0; // @[CtrlBlock.scala 264:29]
  wire  fusionDecoder_io_clear_1; // @[CtrlBlock.scala 264:29]
  wire  rat_clock; // @[CtrlBlock.scala 265:19]
  wire  rat_reset; // @[CtrlBlock.scala 265:19]
  wire  rat_io_redirect; // @[CtrlBlock.scala 265:19]
  wire  rat_io_robCommits_isCommit; // @[CtrlBlock.scala 265:19]
  wire  rat_io_robCommits_commitValid_0; // @[CtrlBlock.scala 265:19]
  wire  rat_io_robCommits_commitValid_1; // @[CtrlBlock.scala 265:19]
  wire  rat_io_robCommits_isWalk; // @[CtrlBlock.scala 265:19]
  wire  rat_io_robCommits_walkValid_0; // @[CtrlBlock.scala 265:19]
  wire  rat_io_robCommits_walkValid_1; // @[CtrlBlock.scala 265:19]
  wire [4:0] rat_io_robCommits_info_0_ldest; // @[CtrlBlock.scala 265:19]
  wire  rat_io_robCommits_info_0_rfWen; // @[CtrlBlock.scala 265:19]
  wire  rat_io_robCommits_info_0_fpWen; // @[CtrlBlock.scala 265:19]
  wire [5:0] rat_io_robCommits_info_0_pdest; // @[CtrlBlock.scala 265:19]
  wire [4:0] rat_io_robCommits_info_1_ldest; // @[CtrlBlock.scala 265:19]
  wire  rat_io_robCommits_info_1_rfWen; // @[CtrlBlock.scala 265:19]
  wire  rat_io_robCommits_info_1_fpWen; // @[CtrlBlock.scala 265:19]
  wire [5:0] rat_io_robCommits_info_1_pdest; // @[CtrlBlock.scala 265:19]
  wire  rat_io_intReadPorts_0_0_hold; // @[CtrlBlock.scala 265:19]
  wire [4:0] rat_io_intReadPorts_0_0_addr; // @[CtrlBlock.scala 265:19]
  wire [5:0] rat_io_intReadPorts_0_0_data; // @[CtrlBlock.scala 265:19]
  wire  rat_io_intReadPorts_0_1_hold; // @[CtrlBlock.scala 265:19]
  wire [4:0] rat_io_intReadPorts_0_1_addr; // @[CtrlBlock.scala 265:19]
  wire [5:0] rat_io_intReadPorts_0_1_data; // @[CtrlBlock.scala 265:19]
  wire  rat_io_intReadPorts_0_2_hold; // @[CtrlBlock.scala 265:19]
  wire [4:0] rat_io_intReadPorts_0_2_addr; // @[CtrlBlock.scala 265:19]
  wire [5:0] rat_io_intReadPorts_0_2_data; // @[CtrlBlock.scala 265:19]
  wire  rat_io_intReadPorts_1_0_hold; // @[CtrlBlock.scala 265:19]
  wire [4:0] rat_io_intReadPorts_1_0_addr; // @[CtrlBlock.scala 265:19]
  wire [5:0] rat_io_intReadPorts_1_0_data; // @[CtrlBlock.scala 265:19]
  wire  rat_io_intReadPorts_1_1_hold; // @[CtrlBlock.scala 265:19]
  wire [4:0] rat_io_intReadPorts_1_1_addr; // @[CtrlBlock.scala 265:19]
  wire [5:0] rat_io_intReadPorts_1_1_data; // @[CtrlBlock.scala 265:19]
  wire  rat_io_intReadPorts_1_2_hold; // @[CtrlBlock.scala 265:19]
  wire [4:0] rat_io_intReadPorts_1_2_addr; // @[CtrlBlock.scala 265:19]
  wire [5:0] rat_io_intReadPorts_1_2_data; // @[CtrlBlock.scala 265:19]
  wire  rat_io_intRenamePorts_0_wen; // @[CtrlBlock.scala 265:19]
  wire [4:0] rat_io_intRenamePorts_0_addr; // @[CtrlBlock.scala 265:19]
  wire [5:0] rat_io_intRenamePorts_0_data; // @[CtrlBlock.scala 265:19]
  wire  rat_io_intRenamePorts_1_wen; // @[CtrlBlock.scala 265:19]
  wire [4:0] rat_io_intRenamePorts_1_addr; // @[CtrlBlock.scala 265:19]
  wire [5:0] rat_io_intRenamePorts_1_data; // @[CtrlBlock.scala 265:19]
  wire  rat_io_fpReadPorts_0_0_hold; // @[CtrlBlock.scala 265:19]
  wire [4:0] rat_io_fpReadPorts_0_0_addr; // @[CtrlBlock.scala 265:19]
  wire [5:0] rat_io_fpReadPorts_0_0_data; // @[CtrlBlock.scala 265:19]
  wire  rat_io_fpReadPorts_0_1_hold; // @[CtrlBlock.scala 265:19]
  wire [4:0] rat_io_fpReadPorts_0_1_addr; // @[CtrlBlock.scala 265:19]
  wire [5:0] rat_io_fpReadPorts_0_1_data; // @[CtrlBlock.scala 265:19]
  wire  rat_io_fpReadPorts_0_2_hold; // @[CtrlBlock.scala 265:19]
  wire [4:0] rat_io_fpReadPorts_0_2_addr; // @[CtrlBlock.scala 265:19]
  wire [5:0] rat_io_fpReadPorts_0_2_data; // @[CtrlBlock.scala 265:19]
  wire  rat_io_fpReadPorts_0_3_hold; // @[CtrlBlock.scala 265:19]
  wire [4:0] rat_io_fpReadPorts_0_3_addr; // @[CtrlBlock.scala 265:19]
  wire [5:0] rat_io_fpReadPorts_0_3_data; // @[CtrlBlock.scala 265:19]
  wire  rat_io_fpReadPorts_1_0_hold; // @[CtrlBlock.scala 265:19]
  wire [4:0] rat_io_fpReadPorts_1_0_addr; // @[CtrlBlock.scala 265:19]
  wire [5:0] rat_io_fpReadPorts_1_0_data; // @[CtrlBlock.scala 265:19]
  wire  rat_io_fpReadPorts_1_1_hold; // @[CtrlBlock.scala 265:19]
  wire [4:0] rat_io_fpReadPorts_1_1_addr; // @[CtrlBlock.scala 265:19]
  wire [5:0] rat_io_fpReadPorts_1_1_data; // @[CtrlBlock.scala 265:19]
  wire  rat_io_fpReadPorts_1_2_hold; // @[CtrlBlock.scala 265:19]
  wire [4:0] rat_io_fpReadPorts_1_2_addr; // @[CtrlBlock.scala 265:19]
  wire [5:0] rat_io_fpReadPorts_1_2_data; // @[CtrlBlock.scala 265:19]
  wire  rat_io_fpReadPorts_1_3_hold; // @[CtrlBlock.scala 265:19]
  wire [4:0] rat_io_fpReadPorts_1_3_addr; // @[CtrlBlock.scala 265:19]
  wire [5:0] rat_io_fpReadPorts_1_3_data; // @[CtrlBlock.scala 265:19]
  wire  rat_io_fpRenamePorts_0_wen; // @[CtrlBlock.scala 265:19]
  wire [4:0] rat_io_fpRenamePorts_0_addr; // @[CtrlBlock.scala 265:19]
  wire [5:0] rat_io_fpRenamePorts_0_data; // @[CtrlBlock.scala 265:19]
  wire  rat_io_fpRenamePorts_1_wen; // @[CtrlBlock.scala 265:19]
  wire [4:0] rat_io_fpRenamePorts_1_addr; // @[CtrlBlock.scala 265:19]
  wire [5:0] rat_io_fpRenamePorts_1_data; // @[CtrlBlock.scala 265:19]
  wire [5:0] rat_io_debug_int_rat_0; // @[CtrlBlock.scala 265:19]
  wire [5:0] rat_io_debug_int_rat_1; // @[CtrlBlock.scala 265:19]
  wire [5:0] rat_io_debug_int_rat_2; // @[CtrlBlock.scala 265:19]
  wire [5:0] rat_io_debug_int_rat_3; // @[CtrlBlock.scala 265:19]
  wire [5:0] rat_io_debug_int_rat_4; // @[CtrlBlock.scala 265:19]
  wire [5:0] rat_io_debug_int_rat_5; // @[CtrlBlock.scala 265:19]
  wire [5:0] rat_io_debug_int_rat_6; // @[CtrlBlock.scala 265:19]
  wire [5:0] rat_io_debug_int_rat_7; // @[CtrlBlock.scala 265:19]
  wire [5:0] rat_io_debug_int_rat_8; // @[CtrlBlock.scala 265:19]
  wire [5:0] rat_io_debug_int_rat_9; // @[CtrlBlock.scala 265:19]
  wire [5:0] rat_io_debug_int_rat_10; // @[CtrlBlock.scala 265:19]
  wire [5:0] rat_io_debug_int_rat_11; // @[CtrlBlock.scala 265:19]
  wire [5:0] rat_io_debug_int_rat_12; // @[CtrlBlock.scala 265:19]
  wire [5:0] rat_io_debug_int_rat_13; // @[CtrlBlock.scala 265:19]
  wire [5:0] rat_io_debug_int_rat_14; // @[CtrlBlock.scala 265:19]
  wire [5:0] rat_io_debug_int_rat_15; // @[CtrlBlock.scala 265:19]
  wire [5:0] rat_io_debug_int_rat_16; // @[CtrlBlock.scala 265:19]
  wire [5:0] rat_io_debug_int_rat_17; // @[CtrlBlock.scala 265:19]
  wire [5:0] rat_io_debug_int_rat_18; // @[CtrlBlock.scala 265:19]
  wire [5:0] rat_io_debug_int_rat_19; // @[CtrlBlock.scala 265:19]
  wire [5:0] rat_io_debug_int_rat_20; // @[CtrlBlock.scala 265:19]
  wire [5:0] rat_io_debug_int_rat_21; // @[CtrlBlock.scala 265:19]
  wire [5:0] rat_io_debug_int_rat_22; // @[CtrlBlock.scala 265:19]
  wire [5:0] rat_io_debug_int_rat_23; // @[CtrlBlock.scala 265:19]
  wire [5:0] rat_io_debug_int_rat_24; // @[CtrlBlock.scala 265:19]
  wire [5:0] rat_io_debug_int_rat_25; // @[CtrlBlock.scala 265:19]
  wire [5:0] rat_io_debug_int_rat_26; // @[CtrlBlock.scala 265:19]
  wire [5:0] rat_io_debug_int_rat_27; // @[CtrlBlock.scala 265:19]
  wire [5:0] rat_io_debug_int_rat_28; // @[CtrlBlock.scala 265:19]
  wire [5:0] rat_io_debug_int_rat_29; // @[CtrlBlock.scala 265:19]
  wire [5:0] rat_io_debug_int_rat_30; // @[CtrlBlock.scala 265:19]
  wire [5:0] rat_io_debug_int_rat_31; // @[CtrlBlock.scala 265:19]
  wire [5:0] rat_io_debug_fp_rat_0; // @[CtrlBlock.scala 265:19]
  wire [5:0] rat_io_debug_fp_rat_1; // @[CtrlBlock.scala 265:19]
  wire [5:0] rat_io_debug_fp_rat_2; // @[CtrlBlock.scala 265:19]
  wire [5:0] rat_io_debug_fp_rat_3; // @[CtrlBlock.scala 265:19]
  wire [5:0] rat_io_debug_fp_rat_4; // @[CtrlBlock.scala 265:19]
  wire [5:0] rat_io_debug_fp_rat_5; // @[CtrlBlock.scala 265:19]
  wire [5:0] rat_io_debug_fp_rat_6; // @[CtrlBlock.scala 265:19]
  wire [5:0] rat_io_debug_fp_rat_7; // @[CtrlBlock.scala 265:19]
  wire [5:0] rat_io_debug_fp_rat_8; // @[CtrlBlock.scala 265:19]
  wire [5:0] rat_io_debug_fp_rat_9; // @[CtrlBlock.scala 265:19]
  wire [5:0] rat_io_debug_fp_rat_10; // @[CtrlBlock.scala 265:19]
  wire [5:0] rat_io_debug_fp_rat_11; // @[CtrlBlock.scala 265:19]
  wire [5:0] rat_io_debug_fp_rat_12; // @[CtrlBlock.scala 265:19]
  wire [5:0] rat_io_debug_fp_rat_13; // @[CtrlBlock.scala 265:19]
  wire [5:0] rat_io_debug_fp_rat_14; // @[CtrlBlock.scala 265:19]
  wire [5:0] rat_io_debug_fp_rat_15; // @[CtrlBlock.scala 265:19]
  wire [5:0] rat_io_debug_fp_rat_16; // @[CtrlBlock.scala 265:19]
  wire [5:0] rat_io_debug_fp_rat_17; // @[CtrlBlock.scala 265:19]
  wire [5:0] rat_io_debug_fp_rat_18; // @[CtrlBlock.scala 265:19]
  wire [5:0] rat_io_debug_fp_rat_19; // @[CtrlBlock.scala 265:19]
  wire [5:0] rat_io_debug_fp_rat_20; // @[CtrlBlock.scala 265:19]
  wire [5:0] rat_io_debug_fp_rat_21; // @[CtrlBlock.scala 265:19]
  wire [5:0] rat_io_debug_fp_rat_22; // @[CtrlBlock.scala 265:19]
  wire [5:0] rat_io_debug_fp_rat_23; // @[CtrlBlock.scala 265:19]
  wire [5:0] rat_io_debug_fp_rat_24; // @[CtrlBlock.scala 265:19]
  wire [5:0] rat_io_debug_fp_rat_25; // @[CtrlBlock.scala 265:19]
  wire [5:0] rat_io_debug_fp_rat_26; // @[CtrlBlock.scala 265:19]
  wire [5:0] rat_io_debug_fp_rat_27; // @[CtrlBlock.scala 265:19]
  wire [5:0] rat_io_debug_fp_rat_28; // @[CtrlBlock.scala 265:19]
  wire [5:0] rat_io_debug_fp_rat_29; // @[CtrlBlock.scala 265:19]
  wire [5:0] rat_io_debug_fp_rat_30; // @[CtrlBlock.scala 265:19]
  wire [5:0] rat_io_debug_fp_rat_31; // @[CtrlBlock.scala 265:19]
  wire  ssit_clock; // @[CtrlBlock.scala 266:20]
  wire  ssit_reset; // @[CtrlBlock.scala 266:20]
  wire [9:0] ssit_io_raddr_0; // @[CtrlBlock.scala 266:20]
  wire [9:0] ssit_io_raddr_1; // @[CtrlBlock.scala 266:20]
  wire  ssit_io_rdata_0_valid; // @[CtrlBlock.scala 266:20]
  wire [4:0] ssit_io_rdata_0_ssid; // @[CtrlBlock.scala 266:20]
  wire  ssit_io_rdata_0_strict; // @[CtrlBlock.scala 266:20]
  wire  ssit_io_rdata_1_valid; // @[CtrlBlock.scala 266:20]
  wire [4:0] ssit_io_rdata_1_ssid; // @[CtrlBlock.scala 266:20]
  wire  ssit_io_rdata_1_strict; // @[CtrlBlock.scala 266:20]
  wire  ssit_io_update_valid; // @[CtrlBlock.scala 266:20]
  wire [9:0] ssit_io_update_ldpc; // @[CtrlBlock.scala 266:20]
  wire [9:0] ssit_io_update_stpc; // @[CtrlBlock.scala 266:20]
  wire [4:0] ssit_io_csrCtrl_lvpred_timeout; // @[CtrlBlock.scala 266:20]
  wire  rename_clock; // @[CtrlBlock.scala 268:22]
  wire  rename_reset; // @[CtrlBlock.scala 268:22]
  wire  rename_io_redirect_valid; // @[CtrlBlock.scala 268:22]
  wire  rename_io_redirect_bits_robIdx_flag; // @[CtrlBlock.scala 268:22]
  wire [4:0] rename_io_redirect_bits_robIdx_value; // @[CtrlBlock.scala 268:22]
  wire  rename_io_redirect_bits_level; // @[CtrlBlock.scala 268:22]
  wire  rename_io_robCommits_isCommit; // @[CtrlBlock.scala 268:22]
  wire  rename_io_robCommits_commitValid_0; // @[CtrlBlock.scala 268:22]
  wire  rename_io_robCommits_commitValid_1; // @[CtrlBlock.scala 268:22]
  wire  rename_io_robCommits_isWalk; // @[CtrlBlock.scala 268:22]
  wire  rename_io_robCommits_walkValid_0; // @[CtrlBlock.scala 268:22]
  wire  rename_io_robCommits_walkValid_1; // @[CtrlBlock.scala 268:22]
  wire [4:0] rename_io_robCommits_info_0_ldest; // @[CtrlBlock.scala 268:22]
  wire  rename_io_robCommits_info_0_rfWen; // @[CtrlBlock.scala 268:22]
  wire  rename_io_robCommits_info_0_fpWen; // @[CtrlBlock.scala 268:22]
  wire [5:0] rename_io_robCommits_info_0_pdest; // @[CtrlBlock.scala 268:22]
  wire [5:0] rename_io_robCommits_info_0_old_pdest; // @[CtrlBlock.scala 268:22]
  wire  rename_io_robCommits_info_0_isMove; // @[CtrlBlock.scala 268:22]
  wire [4:0] rename_io_robCommits_info_1_ldest; // @[CtrlBlock.scala 268:22]
  wire  rename_io_robCommits_info_1_rfWen; // @[CtrlBlock.scala 268:22]
  wire  rename_io_robCommits_info_1_fpWen; // @[CtrlBlock.scala 268:22]
  wire [5:0] rename_io_robCommits_info_1_pdest; // @[CtrlBlock.scala 268:22]
  wire [5:0] rename_io_robCommits_info_1_old_pdest; // @[CtrlBlock.scala 268:22]
  wire  rename_io_robCommits_info_1_isMove; // @[CtrlBlock.scala 268:22]
  wire  rename_io_in_0_ready; // @[CtrlBlock.scala 268:22]
  wire  rename_io_in_0_valid; // @[CtrlBlock.scala 268:22]
  wire [9:0] rename_io_in_0_bits_cf_foldpc; // @[CtrlBlock.scala 268:22]
  wire  rename_io_in_0_bits_cf_exceptionVec_1; // @[CtrlBlock.scala 268:22]
  wire  rename_io_in_0_bits_cf_exceptionVec_2; // @[CtrlBlock.scala 268:22]
  wire  rename_io_in_0_bits_cf_exceptionVec_12; // @[CtrlBlock.scala 268:22]
  wire  rename_io_in_0_bits_cf_trigger_frontendHit_0; // @[CtrlBlock.scala 268:22]
  wire  rename_io_in_0_bits_cf_trigger_frontendHit_1; // @[CtrlBlock.scala 268:22]
  wire  rename_io_in_0_bits_cf_trigger_frontendHit_2; // @[CtrlBlock.scala 268:22]
  wire  rename_io_in_0_bits_cf_trigger_frontendHit_3; // @[CtrlBlock.scala 268:22]
  wire  rename_io_in_0_bits_cf_trigger_backendEn_0; // @[CtrlBlock.scala 268:22]
  wire  rename_io_in_0_bits_cf_trigger_backendEn_1; // @[CtrlBlock.scala 268:22]
  wire  rename_io_in_0_bits_cf_pd_isRVC; // @[CtrlBlock.scala 268:22]
  wire [1:0] rename_io_in_0_bits_cf_pd_brType; // @[CtrlBlock.scala 268:22]
  wire  rename_io_in_0_bits_cf_pd_isCall; // @[CtrlBlock.scala 268:22]
  wire  rename_io_in_0_bits_cf_pd_isRet; // @[CtrlBlock.scala 268:22]
  wire  rename_io_in_0_bits_cf_pred_taken; // @[CtrlBlock.scala 268:22]
  wire  rename_io_in_0_bits_cf_crossPageIPFFix; // @[CtrlBlock.scala 268:22]
  wire  rename_io_in_0_bits_cf_ftqPtr_flag; // @[CtrlBlock.scala 268:22]
  wire [2:0] rename_io_in_0_bits_cf_ftqPtr_value; // @[CtrlBlock.scala 268:22]
  wire [2:0] rename_io_in_0_bits_cf_ftqOffset; // @[CtrlBlock.scala 268:22]
  wire [1:0] rename_io_in_0_bits_ctrl_srcType_0; // @[CtrlBlock.scala 268:22]
  wire [1:0] rename_io_in_0_bits_ctrl_srcType_1; // @[CtrlBlock.scala 268:22]
  wire [1:0] rename_io_in_0_bits_ctrl_srcType_2; // @[CtrlBlock.scala 268:22]
  wire [4:0] rename_io_in_0_bits_ctrl_lsrc_0; // @[CtrlBlock.scala 268:22]
  wire [4:0] rename_io_in_0_bits_ctrl_lsrc_1; // @[CtrlBlock.scala 268:22]
  wire [4:0] rename_io_in_0_bits_ctrl_ldest; // @[CtrlBlock.scala 268:22]
  wire [3:0] rename_io_in_0_bits_ctrl_fuType; // @[CtrlBlock.scala 268:22]
  wire [6:0] rename_io_in_0_bits_ctrl_fuOpType; // @[CtrlBlock.scala 268:22]
  wire  rename_io_in_0_bits_ctrl_rfWen; // @[CtrlBlock.scala 268:22]
  wire  rename_io_in_0_bits_ctrl_fpWen; // @[CtrlBlock.scala 268:22]
  wire  rename_io_in_0_bits_ctrl_isXSTrap; // @[CtrlBlock.scala 268:22]
  wire  rename_io_in_0_bits_ctrl_noSpecExec; // @[CtrlBlock.scala 268:22]
  wire  rename_io_in_0_bits_ctrl_blockBackward; // @[CtrlBlock.scala 268:22]
  wire  rename_io_in_0_bits_ctrl_flushPipe; // @[CtrlBlock.scala 268:22]
  wire [3:0] rename_io_in_0_bits_ctrl_selImm; // @[CtrlBlock.scala 268:22]
  wire [19:0] rename_io_in_0_bits_ctrl_imm; // @[CtrlBlock.scala 268:22]
  wire [2:0] rename_io_in_0_bits_ctrl_commitType; // @[CtrlBlock.scala 268:22]
  wire  rename_io_in_0_bits_ctrl_fpu_isAddSub; // @[CtrlBlock.scala 268:22]
  wire  rename_io_in_0_bits_ctrl_fpu_typeTagIn; // @[CtrlBlock.scala 268:22]
  wire  rename_io_in_0_bits_ctrl_fpu_typeTagOut; // @[CtrlBlock.scala 268:22]
  wire  rename_io_in_0_bits_ctrl_fpu_fromInt; // @[CtrlBlock.scala 268:22]
  wire  rename_io_in_0_bits_ctrl_fpu_wflags; // @[CtrlBlock.scala 268:22]
  wire  rename_io_in_0_bits_ctrl_fpu_fpWen; // @[CtrlBlock.scala 268:22]
  wire [1:0] rename_io_in_0_bits_ctrl_fpu_fmaCmd; // @[CtrlBlock.scala 268:22]
  wire  rename_io_in_0_bits_ctrl_fpu_div; // @[CtrlBlock.scala 268:22]
  wire  rename_io_in_0_bits_ctrl_fpu_sqrt; // @[CtrlBlock.scala 268:22]
  wire  rename_io_in_0_bits_ctrl_fpu_fcvt; // @[CtrlBlock.scala 268:22]
  wire [1:0] rename_io_in_0_bits_ctrl_fpu_typ; // @[CtrlBlock.scala 268:22]
  wire [1:0] rename_io_in_0_bits_ctrl_fpu_fmt; // @[CtrlBlock.scala 268:22]
  wire  rename_io_in_0_bits_ctrl_fpu_ren3; // @[CtrlBlock.scala 268:22]
  wire [2:0] rename_io_in_0_bits_ctrl_fpu_rm; // @[CtrlBlock.scala 268:22]
  wire  rename_io_in_0_bits_ctrl_isMove; // @[CtrlBlock.scala 268:22]
  wire  rename_io_in_1_ready; // @[CtrlBlock.scala 268:22]
  wire  rename_io_in_1_valid; // @[CtrlBlock.scala 268:22]
  wire [9:0] rename_io_in_1_bits_cf_foldpc; // @[CtrlBlock.scala 268:22]
  wire  rename_io_in_1_bits_cf_exceptionVec_1; // @[CtrlBlock.scala 268:22]
  wire  rename_io_in_1_bits_cf_exceptionVec_2; // @[CtrlBlock.scala 268:22]
  wire  rename_io_in_1_bits_cf_exceptionVec_12; // @[CtrlBlock.scala 268:22]
  wire  rename_io_in_1_bits_cf_trigger_frontendHit_0; // @[CtrlBlock.scala 268:22]
  wire  rename_io_in_1_bits_cf_trigger_frontendHit_1; // @[CtrlBlock.scala 268:22]
  wire  rename_io_in_1_bits_cf_trigger_frontendHit_2; // @[CtrlBlock.scala 268:22]
  wire  rename_io_in_1_bits_cf_trigger_frontendHit_3; // @[CtrlBlock.scala 268:22]
  wire  rename_io_in_1_bits_cf_trigger_backendEn_0; // @[CtrlBlock.scala 268:22]
  wire  rename_io_in_1_bits_cf_trigger_backendEn_1; // @[CtrlBlock.scala 268:22]
  wire  rename_io_in_1_bits_cf_pd_isRVC; // @[CtrlBlock.scala 268:22]
  wire [1:0] rename_io_in_1_bits_cf_pd_brType; // @[CtrlBlock.scala 268:22]
  wire  rename_io_in_1_bits_cf_pd_isCall; // @[CtrlBlock.scala 268:22]
  wire  rename_io_in_1_bits_cf_pd_isRet; // @[CtrlBlock.scala 268:22]
  wire  rename_io_in_1_bits_cf_pred_taken; // @[CtrlBlock.scala 268:22]
  wire  rename_io_in_1_bits_cf_crossPageIPFFix; // @[CtrlBlock.scala 268:22]
  wire  rename_io_in_1_bits_cf_ftqPtr_flag; // @[CtrlBlock.scala 268:22]
  wire [2:0] rename_io_in_1_bits_cf_ftqPtr_value; // @[CtrlBlock.scala 268:22]
  wire [2:0] rename_io_in_1_bits_cf_ftqOffset; // @[CtrlBlock.scala 268:22]
  wire [1:0] rename_io_in_1_bits_ctrl_srcType_0; // @[CtrlBlock.scala 268:22]
  wire [1:0] rename_io_in_1_bits_ctrl_srcType_1; // @[CtrlBlock.scala 268:22]
  wire [1:0] rename_io_in_1_bits_ctrl_srcType_2; // @[CtrlBlock.scala 268:22]
  wire [4:0] rename_io_in_1_bits_ctrl_lsrc_0; // @[CtrlBlock.scala 268:22]
  wire [4:0] rename_io_in_1_bits_ctrl_lsrc_1; // @[CtrlBlock.scala 268:22]
  wire [4:0] rename_io_in_1_bits_ctrl_lsrc_2; // @[CtrlBlock.scala 268:22]
  wire [4:0] rename_io_in_1_bits_ctrl_ldest; // @[CtrlBlock.scala 268:22]
  wire [3:0] rename_io_in_1_bits_ctrl_fuType; // @[CtrlBlock.scala 268:22]
  wire [6:0] rename_io_in_1_bits_ctrl_fuOpType; // @[CtrlBlock.scala 268:22]
  wire  rename_io_in_1_bits_ctrl_rfWen; // @[CtrlBlock.scala 268:22]
  wire  rename_io_in_1_bits_ctrl_fpWen; // @[CtrlBlock.scala 268:22]
  wire  rename_io_in_1_bits_ctrl_isXSTrap; // @[CtrlBlock.scala 268:22]
  wire  rename_io_in_1_bits_ctrl_noSpecExec; // @[CtrlBlock.scala 268:22]
  wire  rename_io_in_1_bits_ctrl_blockBackward; // @[CtrlBlock.scala 268:22]
  wire  rename_io_in_1_bits_ctrl_flushPipe; // @[CtrlBlock.scala 268:22]
  wire [3:0] rename_io_in_1_bits_ctrl_selImm; // @[CtrlBlock.scala 268:22]
  wire [19:0] rename_io_in_1_bits_ctrl_imm; // @[CtrlBlock.scala 268:22]
  wire  rename_io_in_1_bits_ctrl_fpu_isAddSub; // @[CtrlBlock.scala 268:22]
  wire  rename_io_in_1_bits_ctrl_fpu_typeTagIn; // @[CtrlBlock.scala 268:22]
  wire  rename_io_in_1_bits_ctrl_fpu_typeTagOut; // @[CtrlBlock.scala 268:22]
  wire  rename_io_in_1_bits_ctrl_fpu_fromInt; // @[CtrlBlock.scala 268:22]
  wire  rename_io_in_1_bits_ctrl_fpu_wflags; // @[CtrlBlock.scala 268:22]
  wire  rename_io_in_1_bits_ctrl_fpu_fpWen; // @[CtrlBlock.scala 268:22]
  wire [1:0] rename_io_in_1_bits_ctrl_fpu_fmaCmd; // @[CtrlBlock.scala 268:22]
  wire  rename_io_in_1_bits_ctrl_fpu_div; // @[CtrlBlock.scala 268:22]
  wire  rename_io_in_1_bits_ctrl_fpu_sqrt; // @[CtrlBlock.scala 268:22]
  wire  rename_io_in_1_bits_ctrl_fpu_fcvt; // @[CtrlBlock.scala 268:22]
  wire [1:0] rename_io_in_1_bits_ctrl_fpu_typ; // @[CtrlBlock.scala 268:22]
  wire [1:0] rename_io_in_1_bits_ctrl_fpu_fmt; // @[CtrlBlock.scala 268:22]
  wire  rename_io_in_1_bits_ctrl_fpu_ren3; // @[CtrlBlock.scala 268:22]
  wire [2:0] rename_io_in_1_bits_ctrl_fpu_rm; // @[CtrlBlock.scala 268:22]
  wire  rename_io_in_1_bits_ctrl_isMove; // @[CtrlBlock.scala 268:22]
  wire  rename_io_fusionInfo_0_rs2FromRs1; // @[CtrlBlock.scala 268:22]
  wire  rename_io_fusionInfo_0_rs2FromRs2; // @[CtrlBlock.scala 268:22]
  wire  rename_io_fusionInfo_0_rs2FromZero; // @[CtrlBlock.scala 268:22]
  wire  rename_io_ssit_0_valid; // @[CtrlBlock.scala 268:22]
  wire [4:0] rename_io_ssit_0_ssid; // @[CtrlBlock.scala 268:22]
  wire  rename_io_ssit_0_strict; // @[CtrlBlock.scala 268:22]
  wire  rename_io_ssit_1_valid; // @[CtrlBlock.scala 268:22]
  wire [4:0] rename_io_ssit_1_ssid; // @[CtrlBlock.scala 268:22]
  wire  rename_io_ssit_1_strict; // @[CtrlBlock.scala 268:22]
  wire [5:0] rename_io_intReadPorts_0_0; // @[CtrlBlock.scala 268:22]
  wire [5:0] rename_io_intReadPorts_0_1; // @[CtrlBlock.scala 268:22]
  wire [5:0] rename_io_intReadPorts_0_2; // @[CtrlBlock.scala 268:22]
  wire [5:0] rename_io_intReadPorts_1_0; // @[CtrlBlock.scala 268:22]
  wire [5:0] rename_io_intReadPorts_1_1; // @[CtrlBlock.scala 268:22]
  wire [5:0] rename_io_intReadPorts_1_2; // @[CtrlBlock.scala 268:22]
  wire [5:0] rename_io_fpReadPorts_0_0; // @[CtrlBlock.scala 268:22]
  wire [5:0] rename_io_fpReadPorts_0_1; // @[CtrlBlock.scala 268:22]
  wire [5:0] rename_io_fpReadPorts_0_2; // @[CtrlBlock.scala 268:22]
  wire [5:0] rename_io_fpReadPorts_0_3; // @[CtrlBlock.scala 268:22]
  wire [5:0] rename_io_fpReadPorts_1_0; // @[CtrlBlock.scala 268:22]
  wire [5:0] rename_io_fpReadPorts_1_1; // @[CtrlBlock.scala 268:22]
  wire [5:0] rename_io_fpReadPorts_1_2; // @[CtrlBlock.scala 268:22]
  wire [5:0] rename_io_fpReadPorts_1_3; // @[CtrlBlock.scala 268:22]
  wire  rename_io_intRenamePorts_0_wen; // @[CtrlBlock.scala 268:22]
  wire [4:0] rename_io_intRenamePorts_0_addr; // @[CtrlBlock.scala 268:22]
  wire [5:0] rename_io_intRenamePorts_0_data; // @[CtrlBlock.scala 268:22]
  wire  rename_io_intRenamePorts_1_wen; // @[CtrlBlock.scala 268:22]
  wire [4:0] rename_io_intRenamePorts_1_addr; // @[CtrlBlock.scala 268:22]
  wire [5:0] rename_io_intRenamePorts_1_data; // @[CtrlBlock.scala 268:22]
  wire  rename_io_fpRenamePorts_0_wen; // @[CtrlBlock.scala 268:22]
  wire [4:0] rename_io_fpRenamePorts_0_addr; // @[CtrlBlock.scala 268:22]
  wire [5:0] rename_io_fpRenamePorts_0_data; // @[CtrlBlock.scala 268:22]
  wire  rename_io_fpRenamePorts_1_wen; // @[CtrlBlock.scala 268:22]
  wire [4:0] rename_io_fpRenamePorts_1_addr; // @[CtrlBlock.scala 268:22]
  wire [5:0] rename_io_fpRenamePorts_1_data; // @[CtrlBlock.scala 268:22]
  wire  rename_io_out_0_ready; // @[CtrlBlock.scala 268:22]
  wire  rename_io_out_0_valid; // @[CtrlBlock.scala 268:22]
  wire [9:0] rename_io_out_0_bits_cf_foldpc; // @[CtrlBlock.scala 268:22]
  wire  rename_io_out_0_bits_cf_exceptionVec_1; // @[CtrlBlock.scala 268:22]
  wire  rename_io_out_0_bits_cf_exceptionVec_2; // @[CtrlBlock.scala 268:22]
  wire  rename_io_out_0_bits_cf_exceptionVec_12; // @[CtrlBlock.scala 268:22]
  wire  rename_io_out_0_bits_cf_trigger_frontendHit_0; // @[CtrlBlock.scala 268:22]
  wire  rename_io_out_0_bits_cf_trigger_frontendHit_1; // @[CtrlBlock.scala 268:22]
  wire  rename_io_out_0_bits_cf_trigger_frontendHit_2; // @[CtrlBlock.scala 268:22]
  wire  rename_io_out_0_bits_cf_trigger_frontendHit_3; // @[CtrlBlock.scala 268:22]
  wire  rename_io_out_0_bits_cf_trigger_backendEn_0; // @[CtrlBlock.scala 268:22]
  wire  rename_io_out_0_bits_cf_trigger_backendEn_1; // @[CtrlBlock.scala 268:22]
  wire  rename_io_out_0_bits_cf_pd_isRVC; // @[CtrlBlock.scala 268:22]
  wire [1:0] rename_io_out_0_bits_cf_pd_brType; // @[CtrlBlock.scala 268:22]
  wire  rename_io_out_0_bits_cf_pd_isCall; // @[CtrlBlock.scala 268:22]
  wire  rename_io_out_0_bits_cf_pd_isRet; // @[CtrlBlock.scala 268:22]
  wire  rename_io_out_0_bits_cf_pred_taken; // @[CtrlBlock.scala 268:22]
  wire  rename_io_out_0_bits_cf_crossPageIPFFix; // @[CtrlBlock.scala 268:22]
  wire  rename_io_out_0_bits_cf_storeSetHit; // @[CtrlBlock.scala 268:22]
  wire  rename_io_out_0_bits_cf_loadWaitStrict; // @[CtrlBlock.scala 268:22]
  wire [4:0] rename_io_out_0_bits_cf_ssid; // @[CtrlBlock.scala 268:22]
  wire  rename_io_out_0_bits_cf_ftqPtr_flag; // @[CtrlBlock.scala 268:22]
  wire [2:0] rename_io_out_0_bits_cf_ftqPtr_value; // @[CtrlBlock.scala 268:22]
  wire [2:0] rename_io_out_0_bits_cf_ftqOffset; // @[CtrlBlock.scala 268:22]
  wire [1:0] rename_io_out_0_bits_ctrl_srcType_0; // @[CtrlBlock.scala 268:22]
  wire [1:0] rename_io_out_0_bits_ctrl_srcType_1; // @[CtrlBlock.scala 268:22]
  wire [1:0] rename_io_out_0_bits_ctrl_srcType_2; // @[CtrlBlock.scala 268:22]
  wire [4:0] rename_io_out_0_bits_ctrl_ldest; // @[CtrlBlock.scala 268:22]
  wire [3:0] rename_io_out_0_bits_ctrl_fuType; // @[CtrlBlock.scala 268:22]
  wire [6:0] rename_io_out_0_bits_ctrl_fuOpType; // @[CtrlBlock.scala 268:22]
  wire  rename_io_out_0_bits_ctrl_rfWen; // @[CtrlBlock.scala 268:22]
  wire  rename_io_out_0_bits_ctrl_fpWen; // @[CtrlBlock.scala 268:22]
  wire  rename_io_out_0_bits_ctrl_isXSTrap; // @[CtrlBlock.scala 268:22]
  wire  rename_io_out_0_bits_ctrl_noSpecExec; // @[CtrlBlock.scala 268:22]
  wire  rename_io_out_0_bits_ctrl_blockBackward; // @[CtrlBlock.scala 268:22]
  wire  rename_io_out_0_bits_ctrl_flushPipe; // @[CtrlBlock.scala 268:22]
  wire [3:0] rename_io_out_0_bits_ctrl_selImm; // @[CtrlBlock.scala 268:22]
  wire [19:0] rename_io_out_0_bits_ctrl_imm; // @[CtrlBlock.scala 268:22]
  wire [2:0] rename_io_out_0_bits_ctrl_commitType; // @[CtrlBlock.scala 268:22]
  wire  rename_io_out_0_bits_ctrl_fpu_isAddSub; // @[CtrlBlock.scala 268:22]
  wire  rename_io_out_0_bits_ctrl_fpu_typeTagIn; // @[CtrlBlock.scala 268:22]
  wire  rename_io_out_0_bits_ctrl_fpu_typeTagOut; // @[CtrlBlock.scala 268:22]
  wire  rename_io_out_0_bits_ctrl_fpu_fromInt; // @[CtrlBlock.scala 268:22]
  wire  rename_io_out_0_bits_ctrl_fpu_wflags; // @[CtrlBlock.scala 268:22]
  wire  rename_io_out_0_bits_ctrl_fpu_fpWen; // @[CtrlBlock.scala 268:22]
  wire [1:0] rename_io_out_0_bits_ctrl_fpu_fmaCmd; // @[CtrlBlock.scala 268:22]
  wire  rename_io_out_0_bits_ctrl_fpu_div; // @[CtrlBlock.scala 268:22]
  wire  rename_io_out_0_bits_ctrl_fpu_sqrt; // @[CtrlBlock.scala 268:22]
  wire  rename_io_out_0_bits_ctrl_fpu_fcvt; // @[CtrlBlock.scala 268:22]
  wire [1:0] rename_io_out_0_bits_ctrl_fpu_typ; // @[CtrlBlock.scala 268:22]
  wire [1:0] rename_io_out_0_bits_ctrl_fpu_fmt; // @[CtrlBlock.scala 268:22]
  wire  rename_io_out_0_bits_ctrl_fpu_ren3; // @[CtrlBlock.scala 268:22]
  wire [2:0] rename_io_out_0_bits_ctrl_fpu_rm; // @[CtrlBlock.scala 268:22]
  wire  rename_io_out_0_bits_ctrl_isMove; // @[CtrlBlock.scala 268:22]
  wire [5:0] rename_io_out_0_bits_psrc_0; // @[CtrlBlock.scala 268:22]
  wire [5:0] rename_io_out_0_bits_psrc_1; // @[CtrlBlock.scala 268:22]
  wire [5:0] rename_io_out_0_bits_psrc_2; // @[CtrlBlock.scala 268:22]
  wire [5:0] rename_io_out_0_bits_pdest; // @[CtrlBlock.scala 268:22]
  wire [5:0] rename_io_out_0_bits_old_pdest; // @[CtrlBlock.scala 268:22]
  wire  rename_io_out_0_bits_robIdx_flag; // @[CtrlBlock.scala 268:22]
  wire [4:0] rename_io_out_0_bits_robIdx_value; // @[CtrlBlock.scala 268:22]
  wire  rename_io_out_0_bits_eliminatedMove; // @[CtrlBlock.scala 268:22]
  wire  rename_io_out_1_valid; // @[CtrlBlock.scala 268:22]
  wire [9:0] rename_io_out_1_bits_cf_foldpc; // @[CtrlBlock.scala 268:22]
  wire  rename_io_out_1_bits_cf_exceptionVec_1; // @[CtrlBlock.scala 268:22]
  wire  rename_io_out_1_bits_cf_exceptionVec_2; // @[CtrlBlock.scala 268:22]
  wire  rename_io_out_1_bits_cf_exceptionVec_12; // @[CtrlBlock.scala 268:22]
  wire  rename_io_out_1_bits_cf_trigger_frontendHit_0; // @[CtrlBlock.scala 268:22]
  wire  rename_io_out_1_bits_cf_trigger_frontendHit_1; // @[CtrlBlock.scala 268:22]
  wire  rename_io_out_1_bits_cf_trigger_frontendHit_2; // @[CtrlBlock.scala 268:22]
  wire  rename_io_out_1_bits_cf_trigger_frontendHit_3; // @[CtrlBlock.scala 268:22]
  wire  rename_io_out_1_bits_cf_trigger_backendEn_0; // @[CtrlBlock.scala 268:22]
  wire  rename_io_out_1_bits_cf_trigger_backendEn_1; // @[CtrlBlock.scala 268:22]
  wire  rename_io_out_1_bits_cf_pd_isRVC; // @[CtrlBlock.scala 268:22]
  wire [1:0] rename_io_out_1_bits_cf_pd_brType; // @[CtrlBlock.scala 268:22]
  wire  rename_io_out_1_bits_cf_pd_isCall; // @[CtrlBlock.scala 268:22]
  wire  rename_io_out_1_bits_cf_pd_isRet; // @[CtrlBlock.scala 268:22]
  wire  rename_io_out_1_bits_cf_pred_taken; // @[CtrlBlock.scala 268:22]
  wire  rename_io_out_1_bits_cf_crossPageIPFFix; // @[CtrlBlock.scala 268:22]
  wire  rename_io_out_1_bits_cf_storeSetHit; // @[CtrlBlock.scala 268:22]
  wire  rename_io_out_1_bits_cf_loadWaitStrict; // @[CtrlBlock.scala 268:22]
  wire [4:0] rename_io_out_1_bits_cf_ssid; // @[CtrlBlock.scala 268:22]
  wire  rename_io_out_1_bits_cf_ftqPtr_flag; // @[CtrlBlock.scala 268:22]
  wire [2:0] rename_io_out_1_bits_cf_ftqPtr_value; // @[CtrlBlock.scala 268:22]
  wire [2:0] rename_io_out_1_bits_cf_ftqOffset; // @[CtrlBlock.scala 268:22]
  wire [1:0] rename_io_out_1_bits_ctrl_srcType_0; // @[CtrlBlock.scala 268:22]
  wire [1:0] rename_io_out_1_bits_ctrl_srcType_1; // @[CtrlBlock.scala 268:22]
  wire [1:0] rename_io_out_1_bits_ctrl_srcType_2; // @[CtrlBlock.scala 268:22]
  wire [4:0] rename_io_out_1_bits_ctrl_ldest; // @[CtrlBlock.scala 268:22]
  wire [3:0] rename_io_out_1_bits_ctrl_fuType; // @[CtrlBlock.scala 268:22]
  wire [6:0] rename_io_out_1_bits_ctrl_fuOpType; // @[CtrlBlock.scala 268:22]
  wire  rename_io_out_1_bits_ctrl_rfWen; // @[CtrlBlock.scala 268:22]
  wire  rename_io_out_1_bits_ctrl_fpWen; // @[CtrlBlock.scala 268:22]
  wire  rename_io_out_1_bits_ctrl_isXSTrap; // @[CtrlBlock.scala 268:22]
  wire  rename_io_out_1_bits_ctrl_noSpecExec; // @[CtrlBlock.scala 268:22]
  wire  rename_io_out_1_bits_ctrl_blockBackward; // @[CtrlBlock.scala 268:22]
  wire  rename_io_out_1_bits_ctrl_flushPipe; // @[CtrlBlock.scala 268:22]
  wire [3:0] rename_io_out_1_bits_ctrl_selImm; // @[CtrlBlock.scala 268:22]
  wire [19:0] rename_io_out_1_bits_ctrl_imm; // @[CtrlBlock.scala 268:22]
  wire  rename_io_out_1_bits_ctrl_fpu_isAddSub; // @[CtrlBlock.scala 268:22]
  wire  rename_io_out_1_bits_ctrl_fpu_typeTagIn; // @[CtrlBlock.scala 268:22]
  wire  rename_io_out_1_bits_ctrl_fpu_typeTagOut; // @[CtrlBlock.scala 268:22]
  wire  rename_io_out_1_bits_ctrl_fpu_fromInt; // @[CtrlBlock.scala 268:22]
  wire  rename_io_out_1_bits_ctrl_fpu_wflags; // @[CtrlBlock.scala 268:22]
  wire  rename_io_out_1_bits_ctrl_fpu_fpWen; // @[CtrlBlock.scala 268:22]
  wire [1:0] rename_io_out_1_bits_ctrl_fpu_fmaCmd; // @[CtrlBlock.scala 268:22]
  wire  rename_io_out_1_bits_ctrl_fpu_div; // @[CtrlBlock.scala 268:22]
  wire  rename_io_out_1_bits_ctrl_fpu_sqrt; // @[CtrlBlock.scala 268:22]
  wire  rename_io_out_1_bits_ctrl_fpu_fcvt; // @[CtrlBlock.scala 268:22]
  wire [1:0] rename_io_out_1_bits_ctrl_fpu_typ; // @[CtrlBlock.scala 268:22]
  wire [1:0] rename_io_out_1_bits_ctrl_fpu_fmt; // @[CtrlBlock.scala 268:22]
  wire  rename_io_out_1_bits_ctrl_fpu_ren3; // @[CtrlBlock.scala 268:22]
  wire [2:0] rename_io_out_1_bits_ctrl_fpu_rm; // @[CtrlBlock.scala 268:22]
  wire  rename_io_out_1_bits_ctrl_isMove; // @[CtrlBlock.scala 268:22]
  wire [5:0] rename_io_out_1_bits_psrc_0; // @[CtrlBlock.scala 268:22]
  wire [5:0] rename_io_out_1_bits_psrc_1; // @[CtrlBlock.scala 268:22]
  wire [5:0] rename_io_out_1_bits_psrc_2; // @[CtrlBlock.scala 268:22]
  wire [5:0] rename_io_out_1_bits_pdest; // @[CtrlBlock.scala 268:22]
  wire [5:0] rename_io_out_1_bits_old_pdest; // @[CtrlBlock.scala 268:22]
  wire  rename_io_out_1_bits_robIdx_flag; // @[CtrlBlock.scala 268:22]
  wire [4:0] rename_io_out_1_bits_robIdx_value; // @[CtrlBlock.scala 268:22]
  wire  rename_io_out_1_bits_eliminatedMove; // @[CtrlBlock.scala 268:22]
  wire [5:0] rename_io_perf_0_value; // @[CtrlBlock.scala 268:22]
  wire [5:0] rename_io_perf_1_value; // @[CtrlBlock.scala 268:22]
  wire [5:0] rename_io_perf_2_value; // @[CtrlBlock.scala 268:22]
  wire [5:0] rename_io_perf_3_value; // @[CtrlBlock.scala 268:22]
  wire [5:0] rename_io_perf_4_value; // @[CtrlBlock.scala 268:22]
  wire [5:0] rename_io_perf_5_value; // @[CtrlBlock.scala 268:22]
  wire [5:0] rename_io_perf_6_value; // @[CtrlBlock.scala 268:22]
  wire [5:0] rename_io_perf_7_value; // @[CtrlBlock.scala 268:22]
  wire [5:0] rename_io_perf_8_value; // @[CtrlBlock.scala 268:22]
  wire [5:0] rename_io_perf_9_value; // @[CtrlBlock.scala 268:22]
  wire [5:0] rename_io_perf_10_value; // @[CtrlBlock.scala 268:22]
  wire [5:0] rename_io_perf_11_value; // @[CtrlBlock.scala 268:22]
  wire [5:0] rename_io_perf_12_value; // @[CtrlBlock.scala 268:22]
  wire [5:0] rename_io_perf_13_value; // @[CtrlBlock.scala 268:22]
  wire  dispatch_clock; // @[CtrlBlock.scala 269:24]
  wire  dispatch_reset; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_fromRename_0_ready; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_fromRename_0_valid; // @[CtrlBlock.scala 269:24]
  wire [9:0] dispatch_io_fromRename_0_bits_cf_foldpc; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_fromRename_0_bits_cf_exceptionVec_1; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_fromRename_0_bits_cf_exceptionVec_2; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_fromRename_0_bits_cf_exceptionVec_12; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_fromRename_0_bits_cf_trigger_frontendHit_0; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_fromRename_0_bits_cf_trigger_frontendHit_1; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_fromRename_0_bits_cf_trigger_frontendHit_2; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_fromRename_0_bits_cf_trigger_frontendHit_3; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_fromRename_0_bits_cf_trigger_backendEn_0; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_fromRename_0_bits_cf_trigger_backendEn_1; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_fromRename_0_bits_cf_pd_isRVC; // @[CtrlBlock.scala 269:24]
  wire [1:0] dispatch_io_fromRename_0_bits_cf_pd_brType; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_fromRename_0_bits_cf_pd_isCall; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_fromRename_0_bits_cf_pd_isRet; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_fromRename_0_bits_cf_pred_taken; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_fromRename_0_bits_cf_crossPageIPFFix; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_fromRename_0_bits_cf_storeSetHit; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_fromRename_0_bits_cf_loadWaitStrict; // @[CtrlBlock.scala 269:24]
  wire [4:0] dispatch_io_fromRename_0_bits_cf_ssid; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_fromRename_0_bits_cf_ftqPtr_flag; // @[CtrlBlock.scala 269:24]
  wire [2:0] dispatch_io_fromRename_0_bits_cf_ftqPtr_value; // @[CtrlBlock.scala 269:24]
  wire [2:0] dispatch_io_fromRename_0_bits_cf_ftqOffset; // @[CtrlBlock.scala 269:24]
  wire [1:0] dispatch_io_fromRename_0_bits_ctrl_srcType_0; // @[CtrlBlock.scala 269:24]
  wire [1:0] dispatch_io_fromRename_0_bits_ctrl_srcType_1; // @[CtrlBlock.scala 269:24]
  wire [1:0] dispatch_io_fromRename_0_bits_ctrl_srcType_2; // @[CtrlBlock.scala 269:24]
  wire [4:0] dispatch_io_fromRename_0_bits_ctrl_ldest; // @[CtrlBlock.scala 269:24]
  wire [3:0] dispatch_io_fromRename_0_bits_ctrl_fuType; // @[CtrlBlock.scala 269:24]
  wire [6:0] dispatch_io_fromRename_0_bits_ctrl_fuOpType; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_fromRename_0_bits_ctrl_rfWen; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_fromRename_0_bits_ctrl_fpWen; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_fromRename_0_bits_ctrl_isXSTrap; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_fromRename_0_bits_ctrl_noSpecExec; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_fromRename_0_bits_ctrl_blockBackward; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_fromRename_0_bits_ctrl_flushPipe; // @[CtrlBlock.scala 269:24]
  wire [3:0] dispatch_io_fromRename_0_bits_ctrl_selImm; // @[CtrlBlock.scala 269:24]
  wire [19:0] dispatch_io_fromRename_0_bits_ctrl_imm; // @[CtrlBlock.scala 269:24]
  wire [2:0] dispatch_io_fromRename_0_bits_ctrl_commitType; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_fromRename_0_bits_ctrl_fpu_isAddSub; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_fromRename_0_bits_ctrl_fpu_typeTagIn; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_fromRename_0_bits_ctrl_fpu_typeTagOut; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_fromRename_0_bits_ctrl_fpu_fromInt; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_fromRename_0_bits_ctrl_fpu_wflags; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_fromRename_0_bits_ctrl_fpu_fpWen; // @[CtrlBlock.scala 269:24]
  wire [1:0] dispatch_io_fromRename_0_bits_ctrl_fpu_fmaCmd; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_fromRename_0_bits_ctrl_fpu_div; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_fromRename_0_bits_ctrl_fpu_sqrt; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_fromRename_0_bits_ctrl_fpu_fcvt; // @[CtrlBlock.scala 269:24]
  wire [1:0] dispatch_io_fromRename_0_bits_ctrl_fpu_typ; // @[CtrlBlock.scala 269:24]
  wire [1:0] dispatch_io_fromRename_0_bits_ctrl_fpu_fmt; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_fromRename_0_bits_ctrl_fpu_ren3; // @[CtrlBlock.scala 269:24]
  wire [2:0] dispatch_io_fromRename_0_bits_ctrl_fpu_rm; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_fromRename_0_bits_ctrl_isMove; // @[CtrlBlock.scala 269:24]
  wire [5:0] dispatch_io_fromRename_0_bits_psrc_0; // @[CtrlBlock.scala 269:24]
  wire [5:0] dispatch_io_fromRename_0_bits_psrc_1; // @[CtrlBlock.scala 269:24]
  wire [5:0] dispatch_io_fromRename_0_bits_psrc_2; // @[CtrlBlock.scala 269:24]
  wire [5:0] dispatch_io_fromRename_0_bits_pdest; // @[CtrlBlock.scala 269:24]
  wire [5:0] dispatch_io_fromRename_0_bits_old_pdest; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_fromRename_0_bits_robIdx_flag; // @[CtrlBlock.scala 269:24]
  wire [4:0] dispatch_io_fromRename_0_bits_robIdx_value; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_fromRename_0_bits_eliminatedMove; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_fromRename_1_ready; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_fromRename_1_valid; // @[CtrlBlock.scala 269:24]
  wire [9:0] dispatch_io_fromRename_1_bits_cf_foldpc; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_fromRename_1_bits_cf_exceptionVec_1; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_fromRename_1_bits_cf_exceptionVec_2; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_fromRename_1_bits_cf_exceptionVec_12; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_fromRename_1_bits_cf_trigger_frontendHit_0; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_fromRename_1_bits_cf_trigger_frontendHit_1; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_fromRename_1_bits_cf_trigger_frontendHit_2; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_fromRename_1_bits_cf_trigger_frontendHit_3; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_fromRename_1_bits_cf_trigger_backendEn_0; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_fromRename_1_bits_cf_trigger_backendEn_1; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_fromRename_1_bits_cf_pd_isRVC; // @[CtrlBlock.scala 269:24]
  wire [1:0] dispatch_io_fromRename_1_bits_cf_pd_brType; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_fromRename_1_bits_cf_pd_isCall; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_fromRename_1_bits_cf_pd_isRet; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_fromRename_1_bits_cf_pred_taken; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_fromRename_1_bits_cf_crossPageIPFFix; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_fromRename_1_bits_cf_storeSetHit; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_fromRename_1_bits_cf_loadWaitStrict; // @[CtrlBlock.scala 269:24]
  wire [4:0] dispatch_io_fromRename_1_bits_cf_ssid; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_fromRename_1_bits_cf_ftqPtr_flag; // @[CtrlBlock.scala 269:24]
  wire [2:0] dispatch_io_fromRename_1_bits_cf_ftqPtr_value; // @[CtrlBlock.scala 269:24]
  wire [2:0] dispatch_io_fromRename_1_bits_cf_ftqOffset; // @[CtrlBlock.scala 269:24]
  wire [1:0] dispatch_io_fromRename_1_bits_ctrl_srcType_0; // @[CtrlBlock.scala 269:24]
  wire [1:0] dispatch_io_fromRename_1_bits_ctrl_srcType_1; // @[CtrlBlock.scala 269:24]
  wire [1:0] dispatch_io_fromRename_1_bits_ctrl_srcType_2; // @[CtrlBlock.scala 269:24]
  wire [4:0] dispatch_io_fromRename_1_bits_ctrl_ldest; // @[CtrlBlock.scala 269:24]
  wire [3:0] dispatch_io_fromRename_1_bits_ctrl_fuType; // @[CtrlBlock.scala 269:24]
  wire [6:0] dispatch_io_fromRename_1_bits_ctrl_fuOpType; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_fromRename_1_bits_ctrl_rfWen; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_fromRename_1_bits_ctrl_fpWen; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_fromRename_1_bits_ctrl_isXSTrap; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_fromRename_1_bits_ctrl_noSpecExec; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_fromRename_1_bits_ctrl_blockBackward; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_fromRename_1_bits_ctrl_flushPipe; // @[CtrlBlock.scala 269:24]
  wire [3:0] dispatch_io_fromRename_1_bits_ctrl_selImm; // @[CtrlBlock.scala 269:24]
  wire [19:0] dispatch_io_fromRename_1_bits_ctrl_imm; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_fromRename_1_bits_ctrl_fpu_isAddSub; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_fromRename_1_bits_ctrl_fpu_typeTagIn; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_fromRename_1_bits_ctrl_fpu_typeTagOut; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_fromRename_1_bits_ctrl_fpu_fromInt; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_fromRename_1_bits_ctrl_fpu_wflags; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_fromRename_1_bits_ctrl_fpu_fpWen; // @[CtrlBlock.scala 269:24]
  wire [1:0] dispatch_io_fromRename_1_bits_ctrl_fpu_fmaCmd; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_fromRename_1_bits_ctrl_fpu_div; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_fromRename_1_bits_ctrl_fpu_sqrt; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_fromRename_1_bits_ctrl_fpu_fcvt; // @[CtrlBlock.scala 269:24]
  wire [1:0] dispatch_io_fromRename_1_bits_ctrl_fpu_typ; // @[CtrlBlock.scala 269:24]
  wire [1:0] dispatch_io_fromRename_1_bits_ctrl_fpu_fmt; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_fromRename_1_bits_ctrl_fpu_ren3; // @[CtrlBlock.scala 269:24]
  wire [2:0] dispatch_io_fromRename_1_bits_ctrl_fpu_rm; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_fromRename_1_bits_ctrl_isMove; // @[CtrlBlock.scala 269:24]
  wire [5:0] dispatch_io_fromRename_1_bits_psrc_0; // @[CtrlBlock.scala 269:24]
  wire [5:0] dispatch_io_fromRename_1_bits_psrc_1; // @[CtrlBlock.scala 269:24]
  wire [5:0] dispatch_io_fromRename_1_bits_psrc_2; // @[CtrlBlock.scala 269:24]
  wire [5:0] dispatch_io_fromRename_1_bits_pdest; // @[CtrlBlock.scala 269:24]
  wire [5:0] dispatch_io_fromRename_1_bits_old_pdest; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_fromRename_1_bits_robIdx_flag; // @[CtrlBlock.scala 269:24]
  wire [4:0] dispatch_io_fromRename_1_bits_robIdx_value; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_fromRename_1_bits_eliminatedMove; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_recv_0; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_recv_1; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_enqRob_canAccept; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_enqRob_isEmpty; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_enqRob_needAlloc_0; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_enqRob_req_0_valid; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_enqRob_req_0_bits_cf_exceptionVec_1; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_enqRob_req_0_bits_cf_exceptionVec_2; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_enqRob_req_0_bits_cf_exceptionVec_12; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_enqRob_req_0_bits_cf_trigger_frontendHit_0; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_enqRob_req_0_bits_cf_trigger_frontendHit_1; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_enqRob_req_0_bits_cf_trigger_frontendHit_2; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_enqRob_req_0_bits_cf_trigger_frontendHit_3; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_enqRob_req_0_bits_cf_pd_isRVC; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_enqRob_req_0_bits_cf_crossPageIPFFix; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_enqRob_req_0_bits_cf_loadWaitBit; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_enqRob_req_0_bits_cf_ftqPtr_flag; // @[CtrlBlock.scala 269:24]
  wire [2:0] dispatch_io_enqRob_req_0_bits_cf_ftqPtr_value; // @[CtrlBlock.scala 269:24]
  wire [2:0] dispatch_io_enqRob_req_0_bits_cf_ftqOffset; // @[CtrlBlock.scala 269:24]
  wire [4:0] dispatch_io_enqRob_req_0_bits_ctrl_ldest; // @[CtrlBlock.scala 269:24]
  wire [3:0] dispatch_io_enqRob_req_0_bits_ctrl_fuType; // @[CtrlBlock.scala 269:24]
  wire [6:0] dispatch_io_enqRob_req_0_bits_ctrl_fuOpType; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_enqRob_req_0_bits_ctrl_rfWen; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_enqRob_req_0_bits_ctrl_fpWen; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_enqRob_req_0_bits_ctrl_isXSTrap; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_enqRob_req_0_bits_ctrl_noSpecExec; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_enqRob_req_0_bits_ctrl_blockBackward; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_enqRob_req_0_bits_ctrl_flushPipe; // @[CtrlBlock.scala 269:24]
  wire [2:0] dispatch_io_enqRob_req_0_bits_ctrl_commitType; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_enqRob_req_0_bits_ctrl_fpu_wflags; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_enqRob_req_0_bits_ctrl_isMove; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_enqRob_req_0_bits_ctrl_singleStep; // @[CtrlBlock.scala 269:24]
  wire [5:0] dispatch_io_enqRob_req_0_bits_pdest; // @[CtrlBlock.scala 269:24]
  wire [5:0] dispatch_io_enqRob_req_0_bits_old_pdest; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_enqRob_req_0_bits_robIdx_flag; // @[CtrlBlock.scala 269:24]
  wire [4:0] dispatch_io_enqRob_req_0_bits_robIdx_value; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_enqRob_req_0_bits_eliminatedMove; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_enqRob_req_1_valid; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_enqRob_req_1_bits_cf_exceptionVec_1; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_enqRob_req_1_bits_cf_exceptionVec_2; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_enqRob_req_1_bits_cf_exceptionVec_12; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_enqRob_req_1_bits_cf_trigger_frontendHit_0; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_enqRob_req_1_bits_cf_trigger_frontendHit_1; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_enqRob_req_1_bits_cf_trigger_frontendHit_2; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_enqRob_req_1_bits_cf_trigger_frontendHit_3; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_enqRob_req_1_bits_cf_pd_isRVC; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_enqRob_req_1_bits_cf_crossPageIPFFix; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_enqRob_req_1_bits_cf_loadWaitBit; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_enqRob_req_1_bits_cf_ftqPtr_flag; // @[CtrlBlock.scala 269:24]
  wire [2:0] dispatch_io_enqRob_req_1_bits_cf_ftqPtr_value; // @[CtrlBlock.scala 269:24]
  wire [2:0] dispatch_io_enqRob_req_1_bits_cf_ftqOffset; // @[CtrlBlock.scala 269:24]
  wire [4:0] dispatch_io_enqRob_req_1_bits_ctrl_ldest; // @[CtrlBlock.scala 269:24]
  wire [3:0] dispatch_io_enqRob_req_1_bits_ctrl_fuType; // @[CtrlBlock.scala 269:24]
  wire [6:0] dispatch_io_enqRob_req_1_bits_ctrl_fuOpType; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_enqRob_req_1_bits_ctrl_rfWen; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_enqRob_req_1_bits_ctrl_fpWen; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_enqRob_req_1_bits_ctrl_isXSTrap; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_enqRob_req_1_bits_ctrl_noSpecExec; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_enqRob_req_1_bits_ctrl_blockBackward; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_enqRob_req_1_bits_ctrl_flushPipe; // @[CtrlBlock.scala 269:24]
  wire [2:0] dispatch_io_enqRob_req_1_bits_ctrl_commitType; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_enqRob_req_1_bits_ctrl_fpu_wflags; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_enqRob_req_1_bits_ctrl_isMove; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_enqRob_req_1_bits_ctrl_singleStep; // @[CtrlBlock.scala 269:24]
  wire [5:0] dispatch_io_enqRob_req_1_bits_pdest; // @[CtrlBlock.scala 269:24]
  wire [5:0] dispatch_io_enqRob_req_1_bits_old_pdest; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_enqRob_req_1_bits_robIdx_flag; // @[CtrlBlock.scala 269:24]
  wire [4:0] dispatch_io_enqRob_req_1_bits_robIdx_value; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_enqRob_req_1_bits_eliminatedMove; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_allocPregs_0_isInt; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_allocPregs_0_isFp; // @[CtrlBlock.scala 269:24]
  wire [5:0] dispatch_io_allocPregs_0_preg; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_allocPregs_1_isInt; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_allocPregs_1_isFp; // @[CtrlBlock.scala 269:24]
  wire [5:0] dispatch_io_allocPregs_1_preg; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toIntDq_canAccept; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toIntDq_needAlloc_0; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toIntDq_needAlloc_1; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toIntDq_req_0_valid; // @[CtrlBlock.scala 269:24]
  wire [9:0] dispatch_io_toIntDq_req_0_bits_cf_foldpc; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toIntDq_req_0_bits_cf_trigger_backendEn_0; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toIntDq_req_0_bits_cf_trigger_backendEn_1; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toIntDq_req_0_bits_cf_pd_isRVC; // @[CtrlBlock.scala 269:24]
  wire [1:0] dispatch_io_toIntDq_req_0_bits_cf_pd_brType; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toIntDq_req_0_bits_cf_pd_isCall; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toIntDq_req_0_bits_cf_pd_isRet; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toIntDq_req_0_bits_cf_pred_taken; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toIntDq_req_0_bits_cf_storeSetHit; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toIntDq_req_0_bits_cf_waitForRobIdx_flag; // @[CtrlBlock.scala 269:24]
  wire [4:0] dispatch_io_toIntDq_req_0_bits_cf_waitForRobIdx_value; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toIntDq_req_0_bits_cf_loadWaitBit; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toIntDq_req_0_bits_cf_loadWaitStrict; // @[CtrlBlock.scala 269:24]
  wire [4:0] dispatch_io_toIntDq_req_0_bits_cf_ssid; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toIntDq_req_0_bits_cf_ftqPtr_flag; // @[CtrlBlock.scala 269:24]
  wire [2:0] dispatch_io_toIntDq_req_0_bits_cf_ftqPtr_value; // @[CtrlBlock.scala 269:24]
  wire [2:0] dispatch_io_toIntDq_req_0_bits_cf_ftqOffset; // @[CtrlBlock.scala 269:24]
  wire [1:0] dispatch_io_toIntDq_req_0_bits_ctrl_srcType_0; // @[CtrlBlock.scala 269:24]
  wire [1:0] dispatch_io_toIntDq_req_0_bits_ctrl_srcType_1; // @[CtrlBlock.scala 269:24]
  wire [1:0] dispatch_io_toIntDq_req_0_bits_ctrl_srcType_2; // @[CtrlBlock.scala 269:24]
  wire [3:0] dispatch_io_toIntDq_req_0_bits_ctrl_fuType; // @[CtrlBlock.scala 269:24]
  wire [6:0] dispatch_io_toIntDq_req_0_bits_ctrl_fuOpType; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toIntDq_req_0_bits_ctrl_rfWen; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toIntDq_req_0_bits_ctrl_fpWen; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toIntDq_req_0_bits_ctrl_flushPipe; // @[CtrlBlock.scala 269:24]
  wire [3:0] dispatch_io_toIntDq_req_0_bits_ctrl_selImm; // @[CtrlBlock.scala 269:24]
  wire [19:0] dispatch_io_toIntDq_req_0_bits_ctrl_imm; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toIntDq_req_0_bits_ctrl_fpu_isAddSub; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toIntDq_req_0_bits_ctrl_fpu_typeTagIn; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toIntDq_req_0_bits_ctrl_fpu_typeTagOut; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toIntDq_req_0_bits_ctrl_fpu_fromInt; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toIntDq_req_0_bits_ctrl_fpu_wflags; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toIntDq_req_0_bits_ctrl_fpu_fpWen; // @[CtrlBlock.scala 269:24]
  wire [1:0] dispatch_io_toIntDq_req_0_bits_ctrl_fpu_fmaCmd; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toIntDq_req_0_bits_ctrl_fpu_div; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toIntDq_req_0_bits_ctrl_fpu_sqrt; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toIntDq_req_0_bits_ctrl_fpu_fcvt; // @[CtrlBlock.scala 269:24]
  wire [1:0] dispatch_io_toIntDq_req_0_bits_ctrl_fpu_typ; // @[CtrlBlock.scala 269:24]
  wire [1:0] dispatch_io_toIntDq_req_0_bits_ctrl_fpu_fmt; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toIntDq_req_0_bits_ctrl_fpu_ren3; // @[CtrlBlock.scala 269:24]
  wire [2:0] dispatch_io_toIntDq_req_0_bits_ctrl_fpu_rm; // @[CtrlBlock.scala 269:24]
  wire [5:0] dispatch_io_toIntDq_req_0_bits_psrc_0; // @[CtrlBlock.scala 269:24]
  wire [5:0] dispatch_io_toIntDq_req_0_bits_psrc_1; // @[CtrlBlock.scala 269:24]
  wire [5:0] dispatch_io_toIntDq_req_0_bits_psrc_2; // @[CtrlBlock.scala 269:24]
  wire [5:0] dispatch_io_toIntDq_req_0_bits_pdest; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toIntDq_req_0_bits_robIdx_flag; // @[CtrlBlock.scala 269:24]
  wire [4:0] dispatch_io_toIntDq_req_0_bits_robIdx_value; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toIntDq_req_1_valid; // @[CtrlBlock.scala 269:24]
  wire [9:0] dispatch_io_toIntDq_req_1_bits_cf_foldpc; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toIntDq_req_1_bits_cf_trigger_backendEn_0; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toIntDq_req_1_bits_cf_trigger_backendEn_1; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toIntDq_req_1_bits_cf_pd_isRVC; // @[CtrlBlock.scala 269:24]
  wire [1:0] dispatch_io_toIntDq_req_1_bits_cf_pd_brType; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toIntDq_req_1_bits_cf_pd_isCall; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toIntDq_req_1_bits_cf_pd_isRet; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toIntDq_req_1_bits_cf_pred_taken; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toIntDq_req_1_bits_cf_storeSetHit; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toIntDq_req_1_bits_cf_waitForRobIdx_flag; // @[CtrlBlock.scala 269:24]
  wire [4:0] dispatch_io_toIntDq_req_1_bits_cf_waitForRobIdx_value; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toIntDq_req_1_bits_cf_loadWaitBit; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toIntDq_req_1_bits_cf_loadWaitStrict; // @[CtrlBlock.scala 269:24]
  wire [4:0] dispatch_io_toIntDq_req_1_bits_cf_ssid; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toIntDq_req_1_bits_cf_ftqPtr_flag; // @[CtrlBlock.scala 269:24]
  wire [2:0] dispatch_io_toIntDq_req_1_bits_cf_ftqPtr_value; // @[CtrlBlock.scala 269:24]
  wire [2:0] dispatch_io_toIntDq_req_1_bits_cf_ftqOffset; // @[CtrlBlock.scala 269:24]
  wire [1:0] dispatch_io_toIntDq_req_1_bits_ctrl_srcType_0; // @[CtrlBlock.scala 269:24]
  wire [1:0] dispatch_io_toIntDq_req_1_bits_ctrl_srcType_1; // @[CtrlBlock.scala 269:24]
  wire [1:0] dispatch_io_toIntDq_req_1_bits_ctrl_srcType_2; // @[CtrlBlock.scala 269:24]
  wire [3:0] dispatch_io_toIntDq_req_1_bits_ctrl_fuType; // @[CtrlBlock.scala 269:24]
  wire [6:0] dispatch_io_toIntDq_req_1_bits_ctrl_fuOpType; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toIntDq_req_1_bits_ctrl_rfWen; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toIntDq_req_1_bits_ctrl_fpWen; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toIntDq_req_1_bits_ctrl_flushPipe; // @[CtrlBlock.scala 269:24]
  wire [3:0] dispatch_io_toIntDq_req_1_bits_ctrl_selImm; // @[CtrlBlock.scala 269:24]
  wire [19:0] dispatch_io_toIntDq_req_1_bits_ctrl_imm; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toIntDq_req_1_bits_ctrl_fpu_isAddSub; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toIntDq_req_1_bits_ctrl_fpu_typeTagIn; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toIntDq_req_1_bits_ctrl_fpu_typeTagOut; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toIntDq_req_1_bits_ctrl_fpu_fromInt; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toIntDq_req_1_bits_ctrl_fpu_wflags; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toIntDq_req_1_bits_ctrl_fpu_fpWen; // @[CtrlBlock.scala 269:24]
  wire [1:0] dispatch_io_toIntDq_req_1_bits_ctrl_fpu_fmaCmd; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toIntDq_req_1_bits_ctrl_fpu_div; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toIntDq_req_1_bits_ctrl_fpu_sqrt; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toIntDq_req_1_bits_ctrl_fpu_fcvt; // @[CtrlBlock.scala 269:24]
  wire [1:0] dispatch_io_toIntDq_req_1_bits_ctrl_fpu_typ; // @[CtrlBlock.scala 269:24]
  wire [1:0] dispatch_io_toIntDq_req_1_bits_ctrl_fpu_fmt; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toIntDq_req_1_bits_ctrl_fpu_ren3; // @[CtrlBlock.scala 269:24]
  wire [2:0] dispatch_io_toIntDq_req_1_bits_ctrl_fpu_rm; // @[CtrlBlock.scala 269:24]
  wire [5:0] dispatch_io_toIntDq_req_1_bits_psrc_0; // @[CtrlBlock.scala 269:24]
  wire [5:0] dispatch_io_toIntDq_req_1_bits_psrc_1; // @[CtrlBlock.scala 269:24]
  wire [5:0] dispatch_io_toIntDq_req_1_bits_psrc_2; // @[CtrlBlock.scala 269:24]
  wire [5:0] dispatch_io_toIntDq_req_1_bits_pdest; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toIntDq_req_1_bits_robIdx_flag; // @[CtrlBlock.scala 269:24]
  wire [4:0] dispatch_io_toIntDq_req_1_bits_robIdx_value; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toFpDq_canAccept; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toFpDq_needAlloc_0; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toFpDq_needAlloc_1; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toFpDq_req_0_valid; // @[CtrlBlock.scala 269:24]
  wire [9:0] dispatch_io_toFpDq_req_0_bits_cf_foldpc; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toFpDq_req_0_bits_cf_trigger_backendEn_0; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toFpDq_req_0_bits_cf_trigger_backendEn_1; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toFpDq_req_0_bits_cf_pd_isRVC; // @[CtrlBlock.scala 269:24]
  wire [1:0] dispatch_io_toFpDq_req_0_bits_cf_pd_brType; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toFpDq_req_0_bits_cf_pd_isCall; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toFpDq_req_0_bits_cf_pd_isRet; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toFpDq_req_0_bits_cf_pred_taken; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toFpDq_req_0_bits_cf_storeSetHit; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toFpDq_req_0_bits_cf_waitForRobIdx_flag; // @[CtrlBlock.scala 269:24]
  wire [4:0] dispatch_io_toFpDq_req_0_bits_cf_waitForRobIdx_value; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toFpDq_req_0_bits_cf_loadWaitBit; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toFpDq_req_0_bits_cf_loadWaitStrict; // @[CtrlBlock.scala 269:24]
  wire [4:0] dispatch_io_toFpDq_req_0_bits_cf_ssid; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toFpDq_req_0_bits_cf_ftqPtr_flag; // @[CtrlBlock.scala 269:24]
  wire [2:0] dispatch_io_toFpDq_req_0_bits_cf_ftqPtr_value; // @[CtrlBlock.scala 269:24]
  wire [2:0] dispatch_io_toFpDq_req_0_bits_cf_ftqOffset; // @[CtrlBlock.scala 269:24]
  wire [1:0] dispatch_io_toFpDq_req_0_bits_ctrl_srcType_0; // @[CtrlBlock.scala 269:24]
  wire [1:0] dispatch_io_toFpDq_req_0_bits_ctrl_srcType_1; // @[CtrlBlock.scala 269:24]
  wire [1:0] dispatch_io_toFpDq_req_0_bits_ctrl_srcType_2; // @[CtrlBlock.scala 269:24]
  wire [3:0] dispatch_io_toFpDq_req_0_bits_ctrl_fuType; // @[CtrlBlock.scala 269:24]
  wire [6:0] dispatch_io_toFpDq_req_0_bits_ctrl_fuOpType; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toFpDq_req_0_bits_ctrl_rfWen; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toFpDq_req_0_bits_ctrl_fpWen; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toFpDq_req_0_bits_ctrl_flushPipe; // @[CtrlBlock.scala 269:24]
  wire [3:0] dispatch_io_toFpDq_req_0_bits_ctrl_selImm; // @[CtrlBlock.scala 269:24]
  wire [19:0] dispatch_io_toFpDq_req_0_bits_ctrl_imm; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toFpDq_req_0_bits_ctrl_fpu_isAddSub; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toFpDq_req_0_bits_ctrl_fpu_typeTagIn; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toFpDq_req_0_bits_ctrl_fpu_typeTagOut; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toFpDq_req_0_bits_ctrl_fpu_fromInt; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toFpDq_req_0_bits_ctrl_fpu_wflags; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toFpDq_req_0_bits_ctrl_fpu_fpWen; // @[CtrlBlock.scala 269:24]
  wire [1:0] dispatch_io_toFpDq_req_0_bits_ctrl_fpu_fmaCmd; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toFpDq_req_0_bits_ctrl_fpu_div; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toFpDq_req_0_bits_ctrl_fpu_sqrt; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toFpDq_req_0_bits_ctrl_fpu_fcvt; // @[CtrlBlock.scala 269:24]
  wire [1:0] dispatch_io_toFpDq_req_0_bits_ctrl_fpu_typ; // @[CtrlBlock.scala 269:24]
  wire [1:0] dispatch_io_toFpDq_req_0_bits_ctrl_fpu_fmt; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toFpDq_req_0_bits_ctrl_fpu_ren3; // @[CtrlBlock.scala 269:24]
  wire [2:0] dispatch_io_toFpDq_req_0_bits_ctrl_fpu_rm; // @[CtrlBlock.scala 269:24]
  wire [5:0] dispatch_io_toFpDq_req_0_bits_psrc_0; // @[CtrlBlock.scala 269:24]
  wire [5:0] dispatch_io_toFpDq_req_0_bits_psrc_1; // @[CtrlBlock.scala 269:24]
  wire [5:0] dispatch_io_toFpDq_req_0_bits_psrc_2; // @[CtrlBlock.scala 269:24]
  wire [5:0] dispatch_io_toFpDq_req_0_bits_pdest; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toFpDq_req_0_bits_robIdx_flag; // @[CtrlBlock.scala 269:24]
  wire [4:0] dispatch_io_toFpDq_req_0_bits_robIdx_value; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toFpDq_req_1_valid; // @[CtrlBlock.scala 269:24]
  wire [9:0] dispatch_io_toFpDq_req_1_bits_cf_foldpc; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toFpDq_req_1_bits_cf_trigger_backendEn_0; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toFpDq_req_1_bits_cf_trigger_backendEn_1; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toFpDq_req_1_bits_cf_pd_isRVC; // @[CtrlBlock.scala 269:24]
  wire [1:0] dispatch_io_toFpDq_req_1_bits_cf_pd_brType; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toFpDq_req_1_bits_cf_pd_isCall; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toFpDq_req_1_bits_cf_pd_isRet; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toFpDq_req_1_bits_cf_pred_taken; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toFpDq_req_1_bits_cf_storeSetHit; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toFpDq_req_1_bits_cf_waitForRobIdx_flag; // @[CtrlBlock.scala 269:24]
  wire [4:0] dispatch_io_toFpDq_req_1_bits_cf_waitForRobIdx_value; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toFpDq_req_1_bits_cf_loadWaitBit; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toFpDq_req_1_bits_cf_loadWaitStrict; // @[CtrlBlock.scala 269:24]
  wire [4:0] dispatch_io_toFpDq_req_1_bits_cf_ssid; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toFpDq_req_1_bits_cf_ftqPtr_flag; // @[CtrlBlock.scala 269:24]
  wire [2:0] dispatch_io_toFpDq_req_1_bits_cf_ftqPtr_value; // @[CtrlBlock.scala 269:24]
  wire [2:0] dispatch_io_toFpDq_req_1_bits_cf_ftqOffset; // @[CtrlBlock.scala 269:24]
  wire [1:0] dispatch_io_toFpDq_req_1_bits_ctrl_srcType_0; // @[CtrlBlock.scala 269:24]
  wire [1:0] dispatch_io_toFpDq_req_1_bits_ctrl_srcType_1; // @[CtrlBlock.scala 269:24]
  wire [1:0] dispatch_io_toFpDq_req_1_bits_ctrl_srcType_2; // @[CtrlBlock.scala 269:24]
  wire [3:0] dispatch_io_toFpDq_req_1_bits_ctrl_fuType; // @[CtrlBlock.scala 269:24]
  wire [6:0] dispatch_io_toFpDq_req_1_bits_ctrl_fuOpType; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toFpDq_req_1_bits_ctrl_rfWen; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toFpDq_req_1_bits_ctrl_fpWen; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toFpDq_req_1_bits_ctrl_flushPipe; // @[CtrlBlock.scala 269:24]
  wire [3:0] dispatch_io_toFpDq_req_1_bits_ctrl_selImm; // @[CtrlBlock.scala 269:24]
  wire [19:0] dispatch_io_toFpDq_req_1_bits_ctrl_imm; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toFpDq_req_1_bits_ctrl_fpu_isAddSub; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toFpDq_req_1_bits_ctrl_fpu_typeTagIn; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toFpDq_req_1_bits_ctrl_fpu_typeTagOut; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toFpDq_req_1_bits_ctrl_fpu_fromInt; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toFpDq_req_1_bits_ctrl_fpu_wflags; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toFpDq_req_1_bits_ctrl_fpu_fpWen; // @[CtrlBlock.scala 269:24]
  wire [1:0] dispatch_io_toFpDq_req_1_bits_ctrl_fpu_fmaCmd; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toFpDq_req_1_bits_ctrl_fpu_div; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toFpDq_req_1_bits_ctrl_fpu_sqrt; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toFpDq_req_1_bits_ctrl_fpu_fcvt; // @[CtrlBlock.scala 269:24]
  wire [1:0] dispatch_io_toFpDq_req_1_bits_ctrl_fpu_typ; // @[CtrlBlock.scala 269:24]
  wire [1:0] dispatch_io_toFpDq_req_1_bits_ctrl_fpu_fmt; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toFpDq_req_1_bits_ctrl_fpu_ren3; // @[CtrlBlock.scala 269:24]
  wire [2:0] dispatch_io_toFpDq_req_1_bits_ctrl_fpu_rm; // @[CtrlBlock.scala 269:24]
  wire [5:0] dispatch_io_toFpDq_req_1_bits_psrc_0; // @[CtrlBlock.scala 269:24]
  wire [5:0] dispatch_io_toFpDq_req_1_bits_psrc_1; // @[CtrlBlock.scala 269:24]
  wire [5:0] dispatch_io_toFpDq_req_1_bits_psrc_2; // @[CtrlBlock.scala 269:24]
  wire [5:0] dispatch_io_toFpDq_req_1_bits_pdest; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toFpDq_req_1_bits_robIdx_flag; // @[CtrlBlock.scala 269:24]
  wire [4:0] dispatch_io_toFpDq_req_1_bits_robIdx_value; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toLsDq_canAccept; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toLsDq_needAlloc_0; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toLsDq_needAlloc_1; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toLsDq_req_0_valid; // @[CtrlBlock.scala 269:24]
  wire [9:0] dispatch_io_toLsDq_req_0_bits_cf_foldpc; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toLsDq_req_0_bits_cf_trigger_backendEn_0; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toLsDq_req_0_bits_cf_trigger_backendEn_1; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toLsDq_req_0_bits_cf_pd_isRVC; // @[CtrlBlock.scala 269:24]
  wire [1:0] dispatch_io_toLsDq_req_0_bits_cf_pd_brType; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toLsDq_req_0_bits_cf_pd_isCall; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toLsDq_req_0_bits_cf_pd_isRet; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toLsDq_req_0_bits_cf_pred_taken; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toLsDq_req_0_bits_cf_storeSetHit; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toLsDq_req_0_bits_cf_waitForRobIdx_flag; // @[CtrlBlock.scala 269:24]
  wire [4:0] dispatch_io_toLsDq_req_0_bits_cf_waitForRobIdx_value; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toLsDq_req_0_bits_cf_loadWaitBit; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toLsDq_req_0_bits_cf_loadWaitStrict; // @[CtrlBlock.scala 269:24]
  wire [4:0] dispatch_io_toLsDq_req_0_bits_cf_ssid; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toLsDq_req_0_bits_cf_ftqPtr_flag; // @[CtrlBlock.scala 269:24]
  wire [2:0] dispatch_io_toLsDq_req_0_bits_cf_ftqPtr_value; // @[CtrlBlock.scala 269:24]
  wire [2:0] dispatch_io_toLsDq_req_0_bits_cf_ftqOffset; // @[CtrlBlock.scala 269:24]
  wire [1:0] dispatch_io_toLsDq_req_0_bits_ctrl_srcType_0; // @[CtrlBlock.scala 269:24]
  wire [1:0] dispatch_io_toLsDq_req_0_bits_ctrl_srcType_1; // @[CtrlBlock.scala 269:24]
  wire [1:0] dispatch_io_toLsDq_req_0_bits_ctrl_srcType_2; // @[CtrlBlock.scala 269:24]
  wire [3:0] dispatch_io_toLsDq_req_0_bits_ctrl_fuType; // @[CtrlBlock.scala 269:24]
  wire [6:0] dispatch_io_toLsDq_req_0_bits_ctrl_fuOpType; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toLsDq_req_0_bits_ctrl_rfWen; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toLsDq_req_0_bits_ctrl_fpWen; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toLsDq_req_0_bits_ctrl_flushPipe; // @[CtrlBlock.scala 269:24]
  wire [3:0] dispatch_io_toLsDq_req_0_bits_ctrl_selImm; // @[CtrlBlock.scala 269:24]
  wire [19:0] dispatch_io_toLsDq_req_0_bits_ctrl_imm; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toLsDq_req_0_bits_ctrl_fpu_isAddSub; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toLsDq_req_0_bits_ctrl_fpu_typeTagIn; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toLsDq_req_0_bits_ctrl_fpu_typeTagOut; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toLsDq_req_0_bits_ctrl_fpu_fromInt; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toLsDq_req_0_bits_ctrl_fpu_wflags; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toLsDq_req_0_bits_ctrl_fpu_fpWen; // @[CtrlBlock.scala 269:24]
  wire [1:0] dispatch_io_toLsDq_req_0_bits_ctrl_fpu_fmaCmd; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toLsDq_req_0_bits_ctrl_fpu_div; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toLsDq_req_0_bits_ctrl_fpu_sqrt; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toLsDq_req_0_bits_ctrl_fpu_fcvt; // @[CtrlBlock.scala 269:24]
  wire [1:0] dispatch_io_toLsDq_req_0_bits_ctrl_fpu_typ; // @[CtrlBlock.scala 269:24]
  wire [1:0] dispatch_io_toLsDq_req_0_bits_ctrl_fpu_fmt; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toLsDq_req_0_bits_ctrl_fpu_ren3; // @[CtrlBlock.scala 269:24]
  wire [2:0] dispatch_io_toLsDq_req_0_bits_ctrl_fpu_rm; // @[CtrlBlock.scala 269:24]
  wire [5:0] dispatch_io_toLsDq_req_0_bits_psrc_0; // @[CtrlBlock.scala 269:24]
  wire [5:0] dispatch_io_toLsDq_req_0_bits_psrc_1; // @[CtrlBlock.scala 269:24]
  wire [5:0] dispatch_io_toLsDq_req_0_bits_psrc_2; // @[CtrlBlock.scala 269:24]
  wire [5:0] dispatch_io_toLsDq_req_0_bits_pdest; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toLsDq_req_0_bits_robIdx_flag; // @[CtrlBlock.scala 269:24]
  wire [4:0] dispatch_io_toLsDq_req_0_bits_robIdx_value; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toLsDq_req_1_valid; // @[CtrlBlock.scala 269:24]
  wire [9:0] dispatch_io_toLsDq_req_1_bits_cf_foldpc; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toLsDq_req_1_bits_cf_trigger_backendEn_0; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toLsDq_req_1_bits_cf_trigger_backendEn_1; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toLsDq_req_1_bits_cf_pd_isRVC; // @[CtrlBlock.scala 269:24]
  wire [1:0] dispatch_io_toLsDq_req_1_bits_cf_pd_brType; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toLsDq_req_1_bits_cf_pd_isCall; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toLsDq_req_1_bits_cf_pd_isRet; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toLsDq_req_1_bits_cf_pred_taken; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toLsDq_req_1_bits_cf_storeSetHit; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toLsDq_req_1_bits_cf_waitForRobIdx_flag; // @[CtrlBlock.scala 269:24]
  wire [4:0] dispatch_io_toLsDq_req_1_bits_cf_waitForRobIdx_value; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toLsDq_req_1_bits_cf_loadWaitBit; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toLsDq_req_1_bits_cf_loadWaitStrict; // @[CtrlBlock.scala 269:24]
  wire [4:0] dispatch_io_toLsDq_req_1_bits_cf_ssid; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toLsDq_req_1_bits_cf_ftqPtr_flag; // @[CtrlBlock.scala 269:24]
  wire [2:0] dispatch_io_toLsDq_req_1_bits_cf_ftqPtr_value; // @[CtrlBlock.scala 269:24]
  wire [2:0] dispatch_io_toLsDq_req_1_bits_cf_ftqOffset; // @[CtrlBlock.scala 269:24]
  wire [1:0] dispatch_io_toLsDq_req_1_bits_ctrl_srcType_0; // @[CtrlBlock.scala 269:24]
  wire [1:0] dispatch_io_toLsDq_req_1_bits_ctrl_srcType_1; // @[CtrlBlock.scala 269:24]
  wire [1:0] dispatch_io_toLsDq_req_1_bits_ctrl_srcType_2; // @[CtrlBlock.scala 269:24]
  wire [3:0] dispatch_io_toLsDq_req_1_bits_ctrl_fuType; // @[CtrlBlock.scala 269:24]
  wire [6:0] dispatch_io_toLsDq_req_1_bits_ctrl_fuOpType; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toLsDq_req_1_bits_ctrl_rfWen; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toLsDq_req_1_bits_ctrl_fpWen; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toLsDq_req_1_bits_ctrl_flushPipe; // @[CtrlBlock.scala 269:24]
  wire [3:0] dispatch_io_toLsDq_req_1_bits_ctrl_selImm; // @[CtrlBlock.scala 269:24]
  wire [19:0] dispatch_io_toLsDq_req_1_bits_ctrl_imm; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toLsDq_req_1_bits_ctrl_fpu_isAddSub; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toLsDq_req_1_bits_ctrl_fpu_typeTagIn; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toLsDq_req_1_bits_ctrl_fpu_typeTagOut; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toLsDq_req_1_bits_ctrl_fpu_fromInt; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toLsDq_req_1_bits_ctrl_fpu_wflags; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toLsDq_req_1_bits_ctrl_fpu_fpWen; // @[CtrlBlock.scala 269:24]
  wire [1:0] dispatch_io_toLsDq_req_1_bits_ctrl_fpu_fmaCmd; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toLsDq_req_1_bits_ctrl_fpu_div; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toLsDq_req_1_bits_ctrl_fpu_sqrt; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toLsDq_req_1_bits_ctrl_fpu_fcvt; // @[CtrlBlock.scala 269:24]
  wire [1:0] dispatch_io_toLsDq_req_1_bits_ctrl_fpu_typ; // @[CtrlBlock.scala 269:24]
  wire [1:0] dispatch_io_toLsDq_req_1_bits_ctrl_fpu_fmt; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toLsDq_req_1_bits_ctrl_fpu_ren3; // @[CtrlBlock.scala 269:24]
  wire [2:0] dispatch_io_toLsDq_req_1_bits_ctrl_fpu_rm; // @[CtrlBlock.scala 269:24]
  wire [5:0] dispatch_io_toLsDq_req_1_bits_psrc_0; // @[CtrlBlock.scala 269:24]
  wire [5:0] dispatch_io_toLsDq_req_1_bits_psrc_1; // @[CtrlBlock.scala 269:24]
  wire [5:0] dispatch_io_toLsDq_req_1_bits_psrc_2; // @[CtrlBlock.scala 269:24]
  wire [5:0] dispatch_io_toLsDq_req_1_bits_pdest; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_toLsDq_req_1_bits_robIdx_flag; // @[CtrlBlock.scala 269:24]
  wire [4:0] dispatch_io_toLsDq_req_1_bits_robIdx_value; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_redirect_valid; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_singleStep; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_lfst_req_0_valid; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_lfst_req_0_bits_isstore; // @[CtrlBlock.scala 269:24]
  wire [4:0] dispatch_io_lfst_req_0_bits_ssid; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_lfst_req_0_bits_robIdx_flag; // @[CtrlBlock.scala 269:24]
  wire [4:0] dispatch_io_lfst_req_0_bits_robIdx_value; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_lfst_req_1_valid; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_lfst_req_1_bits_isstore; // @[CtrlBlock.scala 269:24]
  wire [4:0] dispatch_io_lfst_req_1_bits_ssid; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_lfst_req_1_bits_robIdx_flag; // @[CtrlBlock.scala 269:24]
  wire [4:0] dispatch_io_lfst_req_1_bits_robIdx_value; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_lfst_resp_0_bits_shouldWait; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_lfst_resp_0_bits_robIdx_flag; // @[CtrlBlock.scala 269:24]
  wire [4:0] dispatch_io_lfst_resp_0_bits_robIdx_value; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_lfst_resp_1_bits_shouldWait; // @[CtrlBlock.scala 269:24]
  wire  dispatch_io_lfst_resp_1_bits_robIdx_flag; // @[CtrlBlock.scala 269:24]
  wire [4:0] dispatch_io_lfst_resp_1_bits_robIdx_value; // @[CtrlBlock.scala 269:24]
  wire [5:0] dispatch_io_perf_0_value; // @[CtrlBlock.scala 269:24]
  wire [5:0] dispatch_io_perf_1_value; // @[CtrlBlock.scala 269:24]
  wire [5:0] dispatch_io_perf_2_value; // @[CtrlBlock.scala 269:24]
  wire [5:0] dispatch_io_perf_3_value; // @[CtrlBlock.scala 269:24]
  wire [5:0] dispatch_io_perf_5_value; // @[CtrlBlock.scala 269:24]
  wire [5:0] dispatch_io_perf_6_value; // @[CtrlBlock.scala 269:24]
  wire [5:0] dispatch_io_perf_7_value; // @[CtrlBlock.scala 269:24]
  wire [5:0] dispatch_io_perf_8_value; // @[CtrlBlock.scala 269:24]
  wire  intDq_clock; // @[CtrlBlock.scala 270:21]
  wire  intDq_reset; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_enq_canAccept; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_enq_needAlloc_0; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_enq_needAlloc_1; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_enq_req_0_valid; // @[CtrlBlock.scala 270:21]
  wire [9:0] intDq_io_enq_req_0_bits_cf_foldpc; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_enq_req_0_bits_cf_trigger_backendEn_0; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_enq_req_0_bits_cf_trigger_backendEn_1; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_enq_req_0_bits_cf_pd_isRVC; // @[CtrlBlock.scala 270:21]
  wire [1:0] intDq_io_enq_req_0_bits_cf_pd_brType; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_enq_req_0_bits_cf_pd_isCall; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_enq_req_0_bits_cf_pd_isRet; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_enq_req_0_bits_cf_pred_taken; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_enq_req_0_bits_cf_storeSetHit; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_enq_req_0_bits_cf_waitForRobIdx_flag; // @[CtrlBlock.scala 270:21]
  wire [4:0] intDq_io_enq_req_0_bits_cf_waitForRobIdx_value; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_enq_req_0_bits_cf_loadWaitBit; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_enq_req_0_bits_cf_loadWaitStrict; // @[CtrlBlock.scala 270:21]
  wire [4:0] intDq_io_enq_req_0_bits_cf_ssid; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_enq_req_0_bits_cf_ftqPtr_flag; // @[CtrlBlock.scala 270:21]
  wire [2:0] intDq_io_enq_req_0_bits_cf_ftqPtr_value; // @[CtrlBlock.scala 270:21]
  wire [2:0] intDq_io_enq_req_0_bits_cf_ftqOffset; // @[CtrlBlock.scala 270:21]
  wire [1:0] intDq_io_enq_req_0_bits_ctrl_srcType_0; // @[CtrlBlock.scala 270:21]
  wire [1:0] intDq_io_enq_req_0_bits_ctrl_srcType_1; // @[CtrlBlock.scala 270:21]
  wire [1:0] intDq_io_enq_req_0_bits_ctrl_srcType_2; // @[CtrlBlock.scala 270:21]
  wire [3:0] intDq_io_enq_req_0_bits_ctrl_fuType; // @[CtrlBlock.scala 270:21]
  wire [6:0] intDq_io_enq_req_0_bits_ctrl_fuOpType; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_enq_req_0_bits_ctrl_rfWen; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_enq_req_0_bits_ctrl_fpWen; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_enq_req_0_bits_ctrl_flushPipe; // @[CtrlBlock.scala 270:21]
  wire [3:0] intDq_io_enq_req_0_bits_ctrl_selImm; // @[CtrlBlock.scala 270:21]
  wire [19:0] intDq_io_enq_req_0_bits_ctrl_imm; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_enq_req_0_bits_ctrl_fpu_isAddSub; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_enq_req_0_bits_ctrl_fpu_typeTagIn; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_enq_req_0_bits_ctrl_fpu_typeTagOut; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_enq_req_0_bits_ctrl_fpu_fromInt; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_enq_req_0_bits_ctrl_fpu_wflags; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_enq_req_0_bits_ctrl_fpu_fpWen; // @[CtrlBlock.scala 270:21]
  wire [1:0] intDq_io_enq_req_0_bits_ctrl_fpu_fmaCmd; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_enq_req_0_bits_ctrl_fpu_div; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_enq_req_0_bits_ctrl_fpu_sqrt; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_enq_req_0_bits_ctrl_fpu_fcvt; // @[CtrlBlock.scala 270:21]
  wire [1:0] intDq_io_enq_req_0_bits_ctrl_fpu_typ; // @[CtrlBlock.scala 270:21]
  wire [1:0] intDq_io_enq_req_0_bits_ctrl_fpu_fmt; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_enq_req_0_bits_ctrl_fpu_ren3; // @[CtrlBlock.scala 270:21]
  wire [2:0] intDq_io_enq_req_0_bits_ctrl_fpu_rm; // @[CtrlBlock.scala 270:21]
  wire [5:0] intDq_io_enq_req_0_bits_psrc_0; // @[CtrlBlock.scala 270:21]
  wire [5:0] intDq_io_enq_req_0_bits_psrc_1; // @[CtrlBlock.scala 270:21]
  wire [5:0] intDq_io_enq_req_0_bits_psrc_2; // @[CtrlBlock.scala 270:21]
  wire [5:0] intDq_io_enq_req_0_bits_pdest; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_enq_req_0_bits_robIdx_flag; // @[CtrlBlock.scala 270:21]
  wire [4:0] intDq_io_enq_req_0_bits_robIdx_value; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_enq_req_1_valid; // @[CtrlBlock.scala 270:21]
  wire [9:0] intDq_io_enq_req_1_bits_cf_foldpc; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_enq_req_1_bits_cf_trigger_backendEn_0; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_enq_req_1_bits_cf_trigger_backendEn_1; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_enq_req_1_bits_cf_pd_isRVC; // @[CtrlBlock.scala 270:21]
  wire [1:0] intDq_io_enq_req_1_bits_cf_pd_brType; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_enq_req_1_bits_cf_pd_isCall; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_enq_req_1_bits_cf_pd_isRet; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_enq_req_1_bits_cf_pred_taken; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_enq_req_1_bits_cf_storeSetHit; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_enq_req_1_bits_cf_waitForRobIdx_flag; // @[CtrlBlock.scala 270:21]
  wire [4:0] intDq_io_enq_req_1_bits_cf_waitForRobIdx_value; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_enq_req_1_bits_cf_loadWaitBit; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_enq_req_1_bits_cf_loadWaitStrict; // @[CtrlBlock.scala 270:21]
  wire [4:0] intDq_io_enq_req_1_bits_cf_ssid; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_enq_req_1_bits_cf_ftqPtr_flag; // @[CtrlBlock.scala 270:21]
  wire [2:0] intDq_io_enq_req_1_bits_cf_ftqPtr_value; // @[CtrlBlock.scala 270:21]
  wire [2:0] intDq_io_enq_req_1_bits_cf_ftqOffset; // @[CtrlBlock.scala 270:21]
  wire [1:0] intDq_io_enq_req_1_bits_ctrl_srcType_0; // @[CtrlBlock.scala 270:21]
  wire [1:0] intDq_io_enq_req_1_bits_ctrl_srcType_1; // @[CtrlBlock.scala 270:21]
  wire [1:0] intDq_io_enq_req_1_bits_ctrl_srcType_2; // @[CtrlBlock.scala 270:21]
  wire [3:0] intDq_io_enq_req_1_bits_ctrl_fuType; // @[CtrlBlock.scala 270:21]
  wire [6:0] intDq_io_enq_req_1_bits_ctrl_fuOpType; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_enq_req_1_bits_ctrl_rfWen; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_enq_req_1_bits_ctrl_fpWen; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_enq_req_1_bits_ctrl_flushPipe; // @[CtrlBlock.scala 270:21]
  wire [3:0] intDq_io_enq_req_1_bits_ctrl_selImm; // @[CtrlBlock.scala 270:21]
  wire [19:0] intDq_io_enq_req_1_bits_ctrl_imm; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_enq_req_1_bits_ctrl_fpu_isAddSub; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_enq_req_1_bits_ctrl_fpu_typeTagIn; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_enq_req_1_bits_ctrl_fpu_typeTagOut; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_enq_req_1_bits_ctrl_fpu_fromInt; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_enq_req_1_bits_ctrl_fpu_wflags; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_enq_req_1_bits_ctrl_fpu_fpWen; // @[CtrlBlock.scala 270:21]
  wire [1:0] intDq_io_enq_req_1_bits_ctrl_fpu_fmaCmd; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_enq_req_1_bits_ctrl_fpu_div; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_enq_req_1_bits_ctrl_fpu_sqrt; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_enq_req_1_bits_ctrl_fpu_fcvt; // @[CtrlBlock.scala 270:21]
  wire [1:0] intDq_io_enq_req_1_bits_ctrl_fpu_typ; // @[CtrlBlock.scala 270:21]
  wire [1:0] intDq_io_enq_req_1_bits_ctrl_fpu_fmt; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_enq_req_1_bits_ctrl_fpu_ren3; // @[CtrlBlock.scala 270:21]
  wire [2:0] intDq_io_enq_req_1_bits_ctrl_fpu_rm; // @[CtrlBlock.scala 270:21]
  wire [5:0] intDq_io_enq_req_1_bits_psrc_0; // @[CtrlBlock.scala 270:21]
  wire [5:0] intDq_io_enq_req_1_bits_psrc_1; // @[CtrlBlock.scala 270:21]
  wire [5:0] intDq_io_enq_req_1_bits_psrc_2; // @[CtrlBlock.scala 270:21]
  wire [5:0] intDq_io_enq_req_1_bits_pdest; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_enq_req_1_bits_robIdx_flag; // @[CtrlBlock.scala 270:21]
  wire [4:0] intDq_io_enq_req_1_bits_robIdx_value; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deq_0_ready; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deq_0_valid; // @[CtrlBlock.scala 270:21]
  wire [9:0] intDq_io_deq_0_bits_cf_foldpc; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deq_0_bits_cf_trigger_backendEn_0; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deq_0_bits_cf_trigger_backendEn_1; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deq_0_bits_cf_pd_isRVC; // @[CtrlBlock.scala 270:21]
  wire [1:0] intDq_io_deq_0_bits_cf_pd_brType; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deq_0_bits_cf_pd_isCall; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deq_0_bits_cf_pd_isRet; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deq_0_bits_cf_pred_taken; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deq_0_bits_cf_storeSetHit; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deq_0_bits_cf_waitForRobIdx_flag; // @[CtrlBlock.scala 270:21]
  wire [4:0] intDq_io_deq_0_bits_cf_waitForRobIdx_value; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deq_0_bits_cf_loadWaitBit; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deq_0_bits_cf_loadWaitStrict; // @[CtrlBlock.scala 270:21]
  wire [4:0] intDq_io_deq_0_bits_cf_ssid; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deq_0_bits_cf_ftqPtr_flag; // @[CtrlBlock.scala 270:21]
  wire [2:0] intDq_io_deq_0_bits_cf_ftqPtr_value; // @[CtrlBlock.scala 270:21]
  wire [2:0] intDq_io_deq_0_bits_cf_ftqOffset; // @[CtrlBlock.scala 270:21]
  wire [1:0] intDq_io_deq_0_bits_ctrl_srcType_0; // @[CtrlBlock.scala 270:21]
  wire [1:0] intDq_io_deq_0_bits_ctrl_srcType_1; // @[CtrlBlock.scala 270:21]
  wire [1:0] intDq_io_deq_0_bits_ctrl_srcType_2; // @[CtrlBlock.scala 270:21]
  wire [3:0] intDq_io_deq_0_bits_ctrl_fuType; // @[CtrlBlock.scala 270:21]
  wire [6:0] intDq_io_deq_0_bits_ctrl_fuOpType; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deq_0_bits_ctrl_rfWen; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deq_0_bits_ctrl_fpWen; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deq_0_bits_ctrl_flushPipe; // @[CtrlBlock.scala 270:21]
  wire [3:0] intDq_io_deq_0_bits_ctrl_selImm; // @[CtrlBlock.scala 270:21]
  wire [19:0] intDq_io_deq_0_bits_ctrl_imm; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deq_0_bits_ctrl_fpu_isAddSub; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deq_0_bits_ctrl_fpu_typeTagIn; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deq_0_bits_ctrl_fpu_typeTagOut; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deq_0_bits_ctrl_fpu_fromInt; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deq_0_bits_ctrl_fpu_wflags; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deq_0_bits_ctrl_fpu_fpWen; // @[CtrlBlock.scala 270:21]
  wire [1:0] intDq_io_deq_0_bits_ctrl_fpu_fmaCmd; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deq_0_bits_ctrl_fpu_div; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deq_0_bits_ctrl_fpu_sqrt; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deq_0_bits_ctrl_fpu_fcvt; // @[CtrlBlock.scala 270:21]
  wire [1:0] intDq_io_deq_0_bits_ctrl_fpu_typ; // @[CtrlBlock.scala 270:21]
  wire [1:0] intDq_io_deq_0_bits_ctrl_fpu_fmt; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deq_0_bits_ctrl_fpu_ren3; // @[CtrlBlock.scala 270:21]
  wire [2:0] intDq_io_deq_0_bits_ctrl_fpu_rm; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deq_0_bits_ctrl_replayInst; // @[CtrlBlock.scala 270:21]
  wire [5:0] intDq_io_deq_0_bits_psrc_0; // @[CtrlBlock.scala 270:21]
  wire [5:0] intDq_io_deq_0_bits_psrc_1; // @[CtrlBlock.scala 270:21]
  wire [5:0] intDq_io_deq_0_bits_psrc_2; // @[CtrlBlock.scala 270:21]
  wire [5:0] intDq_io_deq_0_bits_pdest; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deq_0_bits_robIdx_flag; // @[CtrlBlock.scala 270:21]
  wire [4:0] intDq_io_deq_0_bits_robIdx_value; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deq_0_bits_lqIdx_flag; // @[CtrlBlock.scala 270:21]
  wire [3:0] intDq_io_deq_0_bits_lqIdx_value; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deq_0_bits_sqIdx_flag; // @[CtrlBlock.scala 270:21]
  wire [3:0] intDq_io_deq_0_bits_sqIdx_value; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deq_1_ready; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deq_1_valid; // @[CtrlBlock.scala 270:21]
  wire [9:0] intDq_io_deq_1_bits_cf_foldpc; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deq_1_bits_cf_trigger_backendEn_0; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deq_1_bits_cf_trigger_backendEn_1; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deq_1_bits_cf_pd_isRVC; // @[CtrlBlock.scala 270:21]
  wire [1:0] intDq_io_deq_1_bits_cf_pd_brType; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deq_1_bits_cf_pd_isCall; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deq_1_bits_cf_pd_isRet; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deq_1_bits_cf_pred_taken; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deq_1_bits_cf_storeSetHit; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deq_1_bits_cf_waitForRobIdx_flag; // @[CtrlBlock.scala 270:21]
  wire [4:0] intDq_io_deq_1_bits_cf_waitForRobIdx_value; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deq_1_bits_cf_loadWaitBit; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deq_1_bits_cf_loadWaitStrict; // @[CtrlBlock.scala 270:21]
  wire [4:0] intDq_io_deq_1_bits_cf_ssid; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deq_1_bits_cf_ftqPtr_flag; // @[CtrlBlock.scala 270:21]
  wire [2:0] intDq_io_deq_1_bits_cf_ftqPtr_value; // @[CtrlBlock.scala 270:21]
  wire [2:0] intDq_io_deq_1_bits_cf_ftqOffset; // @[CtrlBlock.scala 270:21]
  wire [1:0] intDq_io_deq_1_bits_ctrl_srcType_0; // @[CtrlBlock.scala 270:21]
  wire [1:0] intDq_io_deq_1_bits_ctrl_srcType_1; // @[CtrlBlock.scala 270:21]
  wire [3:0] intDq_io_deq_1_bits_ctrl_fuType; // @[CtrlBlock.scala 270:21]
  wire [6:0] intDq_io_deq_1_bits_ctrl_fuOpType; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deq_1_bits_ctrl_rfWen; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deq_1_bits_ctrl_fpWen; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deq_1_bits_ctrl_flushPipe; // @[CtrlBlock.scala 270:21]
  wire [3:0] intDq_io_deq_1_bits_ctrl_selImm; // @[CtrlBlock.scala 270:21]
  wire [19:0] intDq_io_deq_1_bits_ctrl_imm; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deq_1_bits_ctrl_replayInst; // @[CtrlBlock.scala 270:21]
  wire [5:0] intDq_io_deq_1_bits_psrc_0; // @[CtrlBlock.scala 270:21]
  wire [5:0] intDq_io_deq_1_bits_psrc_1; // @[CtrlBlock.scala 270:21]
  wire [5:0] intDq_io_deq_1_bits_pdest; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deq_1_bits_robIdx_flag; // @[CtrlBlock.scala 270:21]
  wire [4:0] intDq_io_deq_1_bits_robIdx_value; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deq_1_bits_lqIdx_flag; // @[CtrlBlock.scala 270:21]
  wire [3:0] intDq_io_deq_1_bits_lqIdx_value; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deq_1_bits_sqIdx_flag; // @[CtrlBlock.scala 270:21]
  wire [3:0] intDq_io_deq_1_bits_sqIdx_value; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deq_2_ready; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deq_2_valid; // @[CtrlBlock.scala 270:21]
  wire [9:0] intDq_io_deq_2_bits_cf_foldpc; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deq_2_bits_cf_trigger_backendEn_0; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deq_2_bits_cf_trigger_backendEn_1; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deq_2_bits_cf_pd_isRVC; // @[CtrlBlock.scala 270:21]
  wire [1:0] intDq_io_deq_2_bits_cf_pd_brType; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deq_2_bits_cf_pd_isCall; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deq_2_bits_cf_pd_isRet; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deq_2_bits_cf_pred_taken; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deq_2_bits_cf_storeSetHit; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deq_2_bits_cf_waitForRobIdx_flag; // @[CtrlBlock.scala 270:21]
  wire [4:0] intDq_io_deq_2_bits_cf_waitForRobIdx_value; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deq_2_bits_cf_loadWaitBit; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deq_2_bits_cf_loadWaitStrict; // @[CtrlBlock.scala 270:21]
  wire [4:0] intDq_io_deq_2_bits_cf_ssid; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deq_2_bits_cf_ftqPtr_flag; // @[CtrlBlock.scala 270:21]
  wire [2:0] intDq_io_deq_2_bits_cf_ftqPtr_value; // @[CtrlBlock.scala 270:21]
  wire [2:0] intDq_io_deq_2_bits_cf_ftqOffset; // @[CtrlBlock.scala 270:21]
  wire [1:0] intDq_io_deq_2_bits_ctrl_srcType_0; // @[CtrlBlock.scala 270:21]
  wire [1:0] intDq_io_deq_2_bits_ctrl_srcType_1; // @[CtrlBlock.scala 270:21]
  wire [3:0] intDq_io_deq_2_bits_ctrl_fuType; // @[CtrlBlock.scala 270:21]
  wire [6:0] intDq_io_deq_2_bits_ctrl_fuOpType; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deq_2_bits_ctrl_rfWen; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deq_2_bits_ctrl_fpWen; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deq_2_bits_ctrl_flushPipe; // @[CtrlBlock.scala 270:21]
  wire [19:0] intDq_io_deq_2_bits_ctrl_imm; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deq_2_bits_ctrl_replayInst; // @[CtrlBlock.scala 270:21]
  wire [5:0] intDq_io_deq_2_bits_psrc_0; // @[CtrlBlock.scala 270:21]
  wire [5:0] intDq_io_deq_2_bits_psrc_1; // @[CtrlBlock.scala 270:21]
  wire [5:0] intDq_io_deq_2_bits_pdest; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deq_2_bits_robIdx_flag; // @[CtrlBlock.scala 270:21]
  wire [4:0] intDq_io_deq_2_bits_robIdx_value; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deq_3_ready; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deq_3_valid; // @[CtrlBlock.scala 270:21]
  wire [9:0] intDq_io_deq_3_bits_cf_foldpc; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deq_3_bits_cf_trigger_backendEn_0; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deq_3_bits_cf_trigger_backendEn_1; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deq_3_bits_cf_pd_isRVC; // @[CtrlBlock.scala 270:21]
  wire [1:0] intDq_io_deq_3_bits_cf_pd_brType; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deq_3_bits_cf_pd_isCall; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deq_3_bits_cf_pd_isRet; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deq_3_bits_cf_pred_taken; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deq_3_bits_cf_storeSetHit; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deq_3_bits_cf_waitForRobIdx_flag; // @[CtrlBlock.scala 270:21]
  wire [4:0] intDq_io_deq_3_bits_cf_waitForRobIdx_value; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deq_3_bits_cf_loadWaitBit; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deq_3_bits_cf_loadWaitStrict; // @[CtrlBlock.scala 270:21]
  wire [4:0] intDq_io_deq_3_bits_cf_ssid; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deq_3_bits_cf_ftqPtr_flag; // @[CtrlBlock.scala 270:21]
  wire [2:0] intDq_io_deq_3_bits_cf_ftqPtr_value; // @[CtrlBlock.scala 270:21]
  wire [2:0] intDq_io_deq_3_bits_cf_ftqOffset; // @[CtrlBlock.scala 270:21]
  wire [1:0] intDq_io_deq_3_bits_ctrl_srcType_0; // @[CtrlBlock.scala 270:21]
  wire [1:0] intDq_io_deq_3_bits_ctrl_srcType_1; // @[CtrlBlock.scala 270:21]
  wire [3:0] intDq_io_deq_3_bits_ctrl_fuType; // @[CtrlBlock.scala 270:21]
  wire [6:0] intDq_io_deq_3_bits_ctrl_fuOpType; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deq_3_bits_ctrl_rfWen; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deq_3_bits_ctrl_fpWen; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deq_3_bits_ctrl_flushPipe; // @[CtrlBlock.scala 270:21]
  wire [19:0] intDq_io_deq_3_bits_ctrl_imm; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deq_3_bits_ctrl_replayInst; // @[CtrlBlock.scala 270:21]
  wire [5:0] intDq_io_deq_3_bits_psrc_0; // @[CtrlBlock.scala 270:21]
  wire [5:0] intDq_io_deq_3_bits_psrc_1; // @[CtrlBlock.scala 270:21]
  wire [5:0] intDq_io_deq_3_bits_pdest; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deq_3_bits_robIdx_flag; // @[CtrlBlock.scala 270:21]
  wire [4:0] intDq_io_deq_3_bits_robIdx_value; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_redirect_valid; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_redirect_bits_robIdx_flag; // @[CtrlBlock.scala 270:21]
  wire [4:0] intDq_io_redirect_bits_robIdx_value; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_redirect_bits_level; // @[CtrlBlock.scala 270:21]
  wire [2:0] intDq_io_deqNext_0_cf_ftqPtr_value; // @[CtrlBlock.scala 270:21]
  wire [2:0] intDq_io_deqNext_0_cf_ftqOffset; // @[CtrlBlock.scala 270:21]
  wire [1:0] intDq_io_deqNext_0_ctrl_srcType_0; // @[CtrlBlock.scala 270:21]
  wire [1:0] intDq_io_deqNext_0_ctrl_srcType_1; // @[CtrlBlock.scala 270:21]
  wire [1:0] intDq_io_deqNext_0_ctrl_srcType_2; // @[CtrlBlock.scala 270:21]
  wire [3:0] intDq_io_deqNext_0_ctrl_fuType; // @[CtrlBlock.scala 270:21]
  wire [6:0] intDq_io_deqNext_0_ctrl_fuOpType; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deqNext_0_ctrl_rfWen; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deqNext_0_ctrl_fpWen; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deqNext_0_ctrl_flushPipe; // @[CtrlBlock.scala 270:21]
  wire [3:0] intDq_io_deqNext_0_ctrl_selImm; // @[CtrlBlock.scala 270:21]
  wire [19:0] intDq_io_deqNext_0_ctrl_imm; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deqNext_0_ctrl_replayInst; // @[CtrlBlock.scala 270:21]
  wire [5:0] intDq_io_deqNext_0_psrc_0; // @[CtrlBlock.scala 270:21]
  wire [5:0] intDq_io_deqNext_0_psrc_1; // @[CtrlBlock.scala 270:21]
  wire [5:0] intDq_io_deqNext_0_psrc_2; // @[CtrlBlock.scala 270:21]
  wire [5:0] intDq_io_deqNext_0_pdest; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deqNext_0_robIdx_flag; // @[CtrlBlock.scala 270:21]
  wire [4:0] intDq_io_deqNext_0_robIdx_value; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deqNext_0_lqIdx_flag; // @[CtrlBlock.scala 270:21]
  wire [3:0] intDq_io_deqNext_0_lqIdx_value; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deqNext_0_sqIdx_flag; // @[CtrlBlock.scala 270:21]
  wire [3:0] intDq_io_deqNext_0_sqIdx_value; // @[CtrlBlock.scala 270:21]
  wire [2:0] intDq_io_deqNext_1_cf_ftqPtr_value; // @[CtrlBlock.scala 270:21]
  wire [2:0] intDq_io_deqNext_1_cf_ftqOffset; // @[CtrlBlock.scala 270:21]
  wire [1:0] intDq_io_deqNext_1_ctrl_srcType_0; // @[CtrlBlock.scala 270:21]
  wire [1:0] intDq_io_deqNext_1_ctrl_srcType_1; // @[CtrlBlock.scala 270:21]
  wire [1:0] intDq_io_deqNext_1_ctrl_srcType_2; // @[CtrlBlock.scala 270:21]
  wire [3:0] intDq_io_deqNext_1_ctrl_fuType; // @[CtrlBlock.scala 270:21]
  wire [6:0] intDq_io_deqNext_1_ctrl_fuOpType; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deqNext_1_ctrl_rfWen; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deqNext_1_ctrl_fpWen; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deqNext_1_ctrl_flushPipe; // @[CtrlBlock.scala 270:21]
  wire [3:0] intDq_io_deqNext_1_ctrl_selImm; // @[CtrlBlock.scala 270:21]
  wire [19:0] intDq_io_deqNext_1_ctrl_imm; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deqNext_1_ctrl_replayInst; // @[CtrlBlock.scala 270:21]
  wire [5:0] intDq_io_deqNext_1_psrc_0; // @[CtrlBlock.scala 270:21]
  wire [5:0] intDq_io_deqNext_1_psrc_1; // @[CtrlBlock.scala 270:21]
  wire [5:0] intDq_io_deqNext_1_psrc_2; // @[CtrlBlock.scala 270:21]
  wire [5:0] intDq_io_deqNext_1_pdest; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deqNext_1_robIdx_flag; // @[CtrlBlock.scala 270:21]
  wire [4:0] intDq_io_deqNext_1_robIdx_value; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deqNext_1_lqIdx_flag; // @[CtrlBlock.scala 270:21]
  wire [3:0] intDq_io_deqNext_1_lqIdx_value; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deqNext_1_sqIdx_flag; // @[CtrlBlock.scala 270:21]
  wire [3:0] intDq_io_deqNext_1_sqIdx_value; // @[CtrlBlock.scala 270:21]
  wire [2:0] intDq_io_deqNext_2_cf_ftqPtr_value; // @[CtrlBlock.scala 270:21]
  wire [2:0] intDq_io_deqNext_2_cf_ftqOffset; // @[CtrlBlock.scala 270:21]
  wire [1:0] intDq_io_deqNext_2_ctrl_srcType_0; // @[CtrlBlock.scala 270:21]
  wire [1:0] intDq_io_deqNext_2_ctrl_srcType_1; // @[CtrlBlock.scala 270:21]
  wire [1:0] intDq_io_deqNext_2_ctrl_srcType_2; // @[CtrlBlock.scala 270:21]
  wire [3:0] intDq_io_deqNext_2_ctrl_fuType; // @[CtrlBlock.scala 270:21]
  wire [6:0] intDq_io_deqNext_2_ctrl_fuOpType; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deqNext_2_ctrl_rfWen; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deqNext_2_ctrl_fpWen; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deqNext_2_ctrl_flushPipe; // @[CtrlBlock.scala 270:21]
  wire [3:0] intDq_io_deqNext_2_ctrl_selImm; // @[CtrlBlock.scala 270:21]
  wire [19:0] intDq_io_deqNext_2_ctrl_imm; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deqNext_2_ctrl_replayInst; // @[CtrlBlock.scala 270:21]
  wire [5:0] intDq_io_deqNext_2_psrc_0; // @[CtrlBlock.scala 270:21]
  wire [5:0] intDq_io_deqNext_2_psrc_1; // @[CtrlBlock.scala 270:21]
  wire [5:0] intDq_io_deqNext_2_psrc_2; // @[CtrlBlock.scala 270:21]
  wire [5:0] intDq_io_deqNext_2_pdest; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deqNext_2_robIdx_flag; // @[CtrlBlock.scala 270:21]
  wire [4:0] intDq_io_deqNext_2_robIdx_value; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deqNext_2_lqIdx_flag; // @[CtrlBlock.scala 270:21]
  wire [3:0] intDq_io_deqNext_2_lqIdx_value; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deqNext_2_sqIdx_flag; // @[CtrlBlock.scala 270:21]
  wire [3:0] intDq_io_deqNext_2_sqIdx_value; // @[CtrlBlock.scala 270:21]
  wire [2:0] intDq_io_deqNext_3_cf_ftqPtr_value; // @[CtrlBlock.scala 270:21]
  wire [2:0] intDq_io_deqNext_3_cf_ftqOffset; // @[CtrlBlock.scala 270:21]
  wire [1:0] intDq_io_deqNext_3_ctrl_srcType_0; // @[CtrlBlock.scala 270:21]
  wire [1:0] intDq_io_deqNext_3_ctrl_srcType_1; // @[CtrlBlock.scala 270:21]
  wire [1:0] intDq_io_deqNext_3_ctrl_srcType_2; // @[CtrlBlock.scala 270:21]
  wire [3:0] intDq_io_deqNext_3_ctrl_fuType; // @[CtrlBlock.scala 270:21]
  wire [6:0] intDq_io_deqNext_3_ctrl_fuOpType; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deqNext_3_ctrl_rfWen; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deqNext_3_ctrl_fpWen; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deqNext_3_ctrl_flushPipe; // @[CtrlBlock.scala 270:21]
  wire [3:0] intDq_io_deqNext_3_ctrl_selImm; // @[CtrlBlock.scala 270:21]
  wire [19:0] intDq_io_deqNext_3_ctrl_imm; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deqNext_3_ctrl_replayInst; // @[CtrlBlock.scala 270:21]
  wire [5:0] intDq_io_deqNext_3_psrc_0; // @[CtrlBlock.scala 270:21]
  wire [5:0] intDq_io_deqNext_3_psrc_1; // @[CtrlBlock.scala 270:21]
  wire [5:0] intDq_io_deqNext_3_psrc_2; // @[CtrlBlock.scala 270:21]
  wire [5:0] intDq_io_deqNext_3_pdest; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deqNext_3_robIdx_flag; // @[CtrlBlock.scala 270:21]
  wire [4:0] intDq_io_deqNext_3_robIdx_value; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deqNext_3_lqIdx_flag; // @[CtrlBlock.scala 270:21]
  wire [3:0] intDq_io_deqNext_3_lqIdx_value; // @[CtrlBlock.scala 270:21]
  wire  intDq_io_deqNext_3_sqIdx_flag; // @[CtrlBlock.scala 270:21]
  wire [3:0] intDq_io_deqNext_3_sqIdx_value; // @[CtrlBlock.scala 270:21]
  wire [5:0] intDq_io_perf_0_value; // @[CtrlBlock.scala 270:21]
  wire [5:0] intDq_io_perf_1_value; // @[CtrlBlock.scala 270:21]
  wire [5:0] intDq_io_perf_2_value; // @[CtrlBlock.scala 270:21]
  wire [5:0] intDq_io_perf_3_value; // @[CtrlBlock.scala 270:21]
  wire [5:0] intDq_io_perf_4_value; // @[CtrlBlock.scala 270:21]
  wire [5:0] intDq_io_perf_5_value; // @[CtrlBlock.scala 270:21]
  wire [5:0] intDq_io_perf_6_value; // @[CtrlBlock.scala 270:21]
  wire [5:0] intDq_io_perf_7_value; // @[CtrlBlock.scala 270:21]
  wire  fpDq_clock; // @[CtrlBlock.scala 271:20]
  wire  fpDq_reset; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_enq_canAccept; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_enq_needAlloc_0; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_enq_needAlloc_1; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_enq_req_0_valid; // @[CtrlBlock.scala 271:20]
  wire [9:0] fpDq_io_enq_req_0_bits_cf_foldpc; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_enq_req_0_bits_cf_trigger_backendEn_0; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_enq_req_0_bits_cf_trigger_backendEn_1; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_enq_req_0_bits_cf_pd_isRVC; // @[CtrlBlock.scala 271:20]
  wire [1:0] fpDq_io_enq_req_0_bits_cf_pd_brType; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_enq_req_0_bits_cf_pd_isCall; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_enq_req_0_bits_cf_pd_isRet; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_enq_req_0_bits_cf_pred_taken; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_enq_req_0_bits_cf_storeSetHit; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_enq_req_0_bits_cf_waitForRobIdx_flag; // @[CtrlBlock.scala 271:20]
  wire [4:0] fpDq_io_enq_req_0_bits_cf_waitForRobIdx_value; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_enq_req_0_bits_cf_loadWaitBit; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_enq_req_0_bits_cf_loadWaitStrict; // @[CtrlBlock.scala 271:20]
  wire [4:0] fpDq_io_enq_req_0_bits_cf_ssid; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_enq_req_0_bits_cf_ftqPtr_flag; // @[CtrlBlock.scala 271:20]
  wire [2:0] fpDq_io_enq_req_0_bits_cf_ftqPtr_value; // @[CtrlBlock.scala 271:20]
  wire [2:0] fpDq_io_enq_req_0_bits_cf_ftqOffset; // @[CtrlBlock.scala 271:20]
  wire [1:0] fpDq_io_enq_req_0_bits_ctrl_srcType_0; // @[CtrlBlock.scala 271:20]
  wire [1:0] fpDq_io_enq_req_0_bits_ctrl_srcType_1; // @[CtrlBlock.scala 271:20]
  wire [1:0] fpDq_io_enq_req_0_bits_ctrl_srcType_2; // @[CtrlBlock.scala 271:20]
  wire [3:0] fpDq_io_enq_req_0_bits_ctrl_fuType; // @[CtrlBlock.scala 271:20]
  wire [6:0] fpDq_io_enq_req_0_bits_ctrl_fuOpType; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_enq_req_0_bits_ctrl_rfWen; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_enq_req_0_bits_ctrl_fpWen; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_enq_req_0_bits_ctrl_flushPipe; // @[CtrlBlock.scala 271:20]
  wire [3:0] fpDq_io_enq_req_0_bits_ctrl_selImm; // @[CtrlBlock.scala 271:20]
  wire [19:0] fpDq_io_enq_req_0_bits_ctrl_imm; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_enq_req_0_bits_ctrl_fpu_isAddSub; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_enq_req_0_bits_ctrl_fpu_typeTagIn; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_enq_req_0_bits_ctrl_fpu_typeTagOut; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_enq_req_0_bits_ctrl_fpu_fromInt; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_enq_req_0_bits_ctrl_fpu_wflags; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_enq_req_0_bits_ctrl_fpu_fpWen; // @[CtrlBlock.scala 271:20]
  wire [1:0] fpDq_io_enq_req_0_bits_ctrl_fpu_fmaCmd; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_enq_req_0_bits_ctrl_fpu_div; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_enq_req_0_bits_ctrl_fpu_sqrt; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_enq_req_0_bits_ctrl_fpu_fcvt; // @[CtrlBlock.scala 271:20]
  wire [1:0] fpDq_io_enq_req_0_bits_ctrl_fpu_typ; // @[CtrlBlock.scala 271:20]
  wire [1:0] fpDq_io_enq_req_0_bits_ctrl_fpu_fmt; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_enq_req_0_bits_ctrl_fpu_ren3; // @[CtrlBlock.scala 271:20]
  wire [2:0] fpDq_io_enq_req_0_bits_ctrl_fpu_rm; // @[CtrlBlock.scala 271:20]
  wire [5:0] fpDq_io_enq_req_0_bits_psrc_0; // @[CtrlBlock.scala 271:20]
  wire [5:0] fpDq_io_enq_req_0_bits_psrc_1; // @[CtrlBlock.scala 271:20]
  wire [5:0] fpDq_io_enq_req_0_bits_psrc_2; // @[CtrlBlock.scala 271:20]
  wire [5:0] fpDq_io_enq_req_0_bits_pdest; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_enq_req_0_bits_robIdx_flag; // @[CtrlBlock.scala 271:20]
  wire [4:0] fpDq_io_enq_req_0_bits_robIdx_value; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_enq_req_1_valid; // @[CtrlBlock.scala 271:20]
  wire [9:0] fpDq_io_enq_req_1_bits_cf_foldpc; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_enq_req_1_bits_cf_trigger_backendEn_0; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_enq_req_1_bits_cf_trigger_backendEn_1; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_enq_req_1_bits_cf_pd_isRVC; // @[CtrlBlock.scala 271:20]
  wire [1:0] fpDq_io_enq_req_1_bits_cf_pd_brType; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_enq_req_1_bits_cf_pd_isCall; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_enq_req_1_bits_cf_pd_isRet; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_enq_req_1_bits_cf_pred_taken; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_enq_req_1_bits_cf_storeSetHit; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_enq_req_1_bits_cf_waitForRobIdx_flag; // @[CtrlBlock.scala 271:20]
  wire [4:0] fpDq_io_enq_req_1_bits_cf_waitForRobIdx_value; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_enq_req_1_bits_cf_loadWaitBit; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_enq_req_1_bits_cf_loadWaitStrict; // @[CtrlBlock.scala 271:20]
  wire [4:0] fpDq_io_enq_req_1_bits_cf_ssid; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_enq_req_1_bits_cf_ftqPtr_flag; // @[CtrlBlock.scala 271:20]
  wire [2:0] fpDq_io_enq_req_1_bits_cf_ftqPtr_value; // @[CtrlBlock.scala 271:20]
  wire [2:0] fpDq_io_enq_req_1_bits_cf_ftqOffset; // @[CtrlBlock.scala 271:20]
  wire [1:0] fpDq_io_enq_req_1_bits_ctrl_srcType_0; // @[CtrlBlock.scala 271:20]
  wire [1:0] fpDq_io_enq_req_1_bits_ctrl_srcType_1; // @[CtrlBlock.scala 271:20]
  wire [1:0] fpDq_io_enq_req_1_bits_ctrl_srcType_2; // @[CtrlBlock.scala 271:20]
  wire [3:0] fpDq_io_enq_req_1_bits_ctrl_fuType; // @[CtrlBlock.scala 271:20]
  wire [6:0] fpDq_io_enq_req_1_bits_ctrl_fuOpType; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_enq_req_1_bits_ctrl_rfWen; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_enq_req_1_bits_ctrl_fpWen; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_enq_req_1_bits_ctrl_flushPipe; // @[CtrlBlock.scala 271:20]
  wire [3:0] fpDq_io_enq_req_1_bits_ctrl_selImm; // @[CtrlBlock.scala 271:20]
  wire [19:0] fpDq_io_enq_req_1_bits_ctrl_imm; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_enq_req_1_bits_ctrl_fpu_isAddSub; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_enq_req_1_bits_ctrl_fpu_typeTagIn; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_enq_req_1_bits_ctrl_fpu_typeTagOut; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_enq_req_1_bits_ctrl_fpu_fromInt; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_enq_req_1_bits_ctrl_fpu_wflags; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_enq_req_1_bits_ctrl_fpu_fpWen; // @[CtrlBlock.scala 271:20]
  wire [1:0] fpDq_io_enq_req_1_bits_ctrl_fpu_fmaCmd; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_enq_req_1_bits_ctrl_fpu_div; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_enq_req_1_bits_ctrl_fpu_sqrt; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_enq_req_1_bits_ctrl_fpu_fcvt; // @[CtrlBlock.scala 271:20]
  wire [1:0] fpDq_io_enq_req_1_bits_ctrl_fpu_typ; // @[CtrlBlock.scala 271:20]
  wire [1:0] fpDq_io_enq_req_1_bits_ctrl_fpu_fmt; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_enq_req_1_bits_ctrl_fpu_ren3; // @[CtrlBlock.scala 271:20]
  wire [2:0] fpDq_io_enq_req_1_bits_ctrl_fpu_rm; // @[CtrlBlock.scala 271:20]
  wire [5:0] fpDq_io_enq_req_1_bits_psrc_0; // @[CtrlBlock.scala 271:20]
  wire [5:0] fpDq_io_enq_req_1_bits_psrc_1; // @[CtrlBlock.scala 271:20]
  wire [5:0] fpDq_io_enq_req_1_bits_psrc_2; // @[CtrlBlock.scala 271:20]
  wire [5:0] fpDq_io_enq_req_1_bits_pdest; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_enq_req_1_bits_robIdx_flag; // @[CtrlBlock.scala 271:20]
  wire [4:0] fpDq_io_enq_req_1_bits_robIdx_value; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deq_0_ready; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deq_0_valid; // @[CtrlBlock.scala 271:20]
  wire [9:0] fpDq_io_deq_0_bits_cf_foldpc; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deq_0_bits_cf_trigger_backendEn_0; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deq_0_bits_cf_trigger_backendEn_1; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deq_0_bits_cf_pd_isRVC; // @[CtrlBlock.scala 271:20]
  wire [1:0] fpDq_io_deq_0_bits_cf_pd_brType; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deq_0_bits_cf_pd_isCall; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deq_0_bits_cf_pd_isRet; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deq_0_bits_cf_pred_taken; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deq_0_bits_cf_storeSetHit; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deq_0_bits_cf_waitForRobIdx_flag; // @[CtrlBlock.scala 271:20]
  wire [4:0] fpDq_io_deq_0_bits_cf_waitForRobIdx_value; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deq_0_bits_cf_loadWaitBit; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deq_0_bits_cf_loadWaitStrict; // @[CtrlBlock.scala 271:20]
  wire [4:0] fpDq_io_deq_0_bits_cf_ssid; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deq_0_bits_cf_ftqPtr_flag; // @[CtrlBlock.scala 271:20]
  wire [2:0] fpDq_io_deq_0_bits_cf_ftqPtr_value; // @[CtrlBlock.scala 271:20]
  wire [2:0] fpDq_io_deq_0_bits_cf_ftqOffset; // @[CtrlBlock.scala 271:20]
  wire [1:0] fpDq_io_deq_0_bits_ctrl_srcType_0; // @[CtrlBlock.scala 271:20]
  wire [1:0] fpDq_io_deq_0_bits_ctrl_srcType_1; // @[CtrlBlock.scala 271:20]
  wire [1:0] fpDq_io_deq_0_bits_ctrl_srcType_2; // @[CtrlBlock.scala 271:20]
  wire [3:0] fpDq_io_deq_0_bits_ctrl_fuType; // @[CtrlBlock.scala 271:20]
  wire [6:0] fpDq_io_deq_0_bits_ctrl_fuOpType; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deq_0_bits_ctrl_rfWen; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deq_0_bits_ctrl_fpWen; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deq_0_bits_ctrl_flushPipe; // @[CtrlBlock.scala 271:20]
  wire [3:0] fpDq_io_deq_0_bits_ctrl_selImm; // @[CtrlBlock.scala 271:20]
  wire [19:0] fpDq_io_deq_0_bits_ctrl_imm; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deq_0_bits_ctrl_fpu_isAddSub; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deq_0_bits_ctrl_fpu_typeTagIn; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deq_0_bits_ctrl_fpu_typeTagOut; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deq_0_bits_ctrl_fpu_fromInt; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deq_0_bits_ctrl_fpu_wflags; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deq_0_bits_ctrl_fpu_fpWen; // @[CtrlBlock.scala 271:20]
  wire [1:0] fpDq_io_deq_0_bits_ctrl_fpu_fmaCmd; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deq_0_bits_ctrl_fpu_div; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deq_0_bits_ctrl_fpu_sqrt; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deq_0_bits_ctrl_fpu_fcvt; // @[CtrlBlock.scala 271:20]
  wire [1:0] fpDq_io_deq_0_bits_ctrl_fpu_typ; // @[CtrlBlock.scala 271:20]
  wire [1:0] fpDq_io_deq_0_bits_ctrl_fpu_fmt; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deq_0_bits_ctrl_fpu_ren3; // @[CtrlBlock.scala 271:20]
  wire [2:0] fpDq_io_deq_0_bits_ctrl_fpu_rm; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deq_0_bits_ctrl_replayInst; // @[CtrlBlock.scala 271:20]
  wire [5:0] fpDq_io_deq_0_bits_psrc_0; // @[CtrlBlock.scala 271:20]
  wire [5:0] fpDq_io_deq_0_bits_psrc_1; // @[CtrlBlock.scala 271:20]
  wire [5:0] fpDq_io_deq_0_bits_psrc_2; // @[CtrlBlock.scala 271:20]
  wire [5:0] fpDq_io_deq_0_bits_pdest; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deq_0_bits_robIdx_flag; // @[CtrlBlock.scala 271:20]
  wire [4:0] fpDq_io_deq_0_bits_robIdx_value; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deq_0_bits_lqIdx_flag; // @[CtrlBlock.scala 271:20]
  wire [3:0] fpDq_io_deq_0_bits_lqIdx_value; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deq_0_bits_sqIdx_flag; // @[CtrlBlock.scala 271:20]
  wire [3:0] fpDq_io_deq_0_bits_sqIdx_value; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deq_1_ready; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deq_1_valid; // @[CtrlBlock.scala 271:20]
  wire [9:0] fpDq_io_deq_1_bits_cf_foldpc; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deq_1_bits_cf_trigger_backendEn_0; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deq_1_bits_cf_trigger_backendEn_1; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deq_1_bits_cf_pd_isRVC; // @[CtrlBlock.scala 271:20]
  wire [1:0] fpDq_io_deq_1_bits_cf_pd_brType; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deq_1_bits_cf_pd_isCall; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deq_1_bits_cf_pd_isRet; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deq_1_bits_cf_pred_taken; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deq_1_bits_cf_storeSetHit; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deq_1_bits_cf_waitForRobIdx_flag; // @[CtrlBlock.scala 271:20]
  wire [4:0] fpDq_io_deq_1_bits_cf_waitForRobIdx_value; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deq_1_bits_cf_loadWaitBit; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deq_1_bits_cf_loadWaitStrict; // @[CtrlBlock.scala 271:20]
  wire [4:0] fpDq_io_deq_1_bits_cf_ssid; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deq_1_bits_cf_ftqPtr_flag; // @[CtrlBlock.scala 271:20]
  wire [2:0] fpDq_io_deq_1_bits_cf_ftqPtr_value; // @[CtrlBlock.scala 271:20]
  wire [2:0] fpDq_io_deq_1_bits_cf_ftqOffset; // @[CtrlBlock.scala 271:20]
  wire [1:0] fpDq_io_deq_1_bits_ctrl_srcType_0; // @[CtrlBlock.scala 271:20]
  wire [1:0] fpDq_io_deq_1_bits_ctrl_srcType_1; // @[CtrlBlock.scala 271:20]
  wire [3:0] fpDq_io_deq_1_bits_ctrl_fuType; // @[CtrlBlock.scala 271:20]
  wire [6:0] fpDq_io_deq_1_bits_ctrl_fuOpType; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deq_1_bits_ctrl_rfWen; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deq_1_bits_ctrl_fpWen; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deq_1_bits_ctrl_flushPipe; // @[CtrlBlock.scala 271:20]
  wire [3:0] fpDq_io_deq_1_bits_ctrl_selImm; // @[CtrlBlock.scala 271:20]
  wire [19:0] fpDq_io_deq_1_bits_ctrl_imm; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deq_1_bits_ctrl_replayInst; // @[CtrlBlock.scala 271:20]
  wire [5:0] fpDq_io_deq_1_bits_psrc_0; // @[CtrlBlock.scala 271:20]
  wire [5:0] fpDq_io_deq_1_bits_psrc_1; // @[CtrlBlock.scala 271:20]
  wire [5:0] fpDq_io_deq_1_bits_pdest; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deq_1_bits_robIdx_flag; // @[CtrlBlock.scala 271:20]
  wire [4:0] fpDq_io_deq_1_bits_robIdx_value; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deq_1_bits_lqIdx_flag; // @[CtrlBlock.scala 271:20]
  wire [3:0] fpDq_io_deq_1_bits_lqIdx_value; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deq_1_bits_sqIdx_flag; // @[CtrlBlock.scala 271:20]
  wire [3:0] fpDq_io_deq_1_bits_sqIdx_value; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deq_2_ready; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deq_2_valid; // @[CtrlBlock.scala 271:20]
  wire [9:0] fpDq_io_deq_2_bits_cf_foldpc; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deq_2_bits_cf_trigger_backendEn_0; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deq_2_bits_cf_trigger_backendEn_1; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deq_2_bits_cf_pd_isRVC; // @[CtrlBlock.scala 271:20]
  wire [1:0] fpDq_io_deq_2_bits_cf_pd_brType; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deq_2_bits_cf_pd_isCall; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deq_2_bits_cf_pd_isRet; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deq_2_bits_cf_pred_taken; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deq_2_bits_cf_storeSetHit; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deq_2_bits_cf_waitForRobIdx_flag; // @[CtrlBlock.scala 271:20]
  wire [4:0] fpDq_io_deq_2_bits_cf_waitForRobIdx_value; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deq_2_bits_cf_loadWaitBit; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deq_2_bits_cf_loadWaitStrict; // @[CtrlBlock.scala 271:20]
  wire [4:0] fpDq_io_deq_2_bits_cf_ssid; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deq_2_bits_cf_ftqPtr_flag; // @[CtrlBlock.scala 271:20]
  wire [2:0] fpDq_io_deq_2_bits_cf_ftqPtr_value; // @[CtrlBlock.scala 271:20]
  wire [2:0] fpDq_io_deq_2_bits_cf_ftqOffset; // @[CtrlBlock.scala 271:20]
  wire [1:0] fpDq_io_deq_2_bits_ctrl_srcType_0; // @[CtrlBlock.scala 271:20]
  wire [1:0] fpDq_io_deq_2_bits_ctrl_srcType_1; // @[CtrlBlock.scala 271:20]
  wire [3:0] fpDq_io_deq_2_bits_ctrl_fuType; // @[CtrlBlock.scala 271:20]
  wire [6:0] fpDq_io_deq_2_bits_ctrl_fuOpType; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deq_2_bits_ctrl_rfWen; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deq_2_bits_ctrl_fpWen; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deq_2_bits_ctrl_flushPipe; // @[CtrlBlock.scala 271:20]
  wire [19:0] fpDq_io_deq_2_bits_ctrl_imm; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deq_2_bits_ctrl_replayInst; // @[CtrlBlock.scala 271:20]
  wire [5:0] fpDq_io_deq_2_bits_psrc_0; // @[CtrlBlock.scala 271:20]
  wire [5:0] fpDq_io_deq_2_bits_psrc_1; // @[CtrlBlock.scala 271:20]
  wire [5:0] fpDq_io_deq_2_bits_pdest; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deq_2_bits_robIdx_flag; // @[CtrlBlock.scala 271:20]
  wire [4:0] fpDq_io_deq_2_bits_robIdx_value; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deq_3_ready; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deq_3_valid; // @[CtrlBlock.scala 271:20]
  wire [9:0] fpDq_io_deq_3_bits_cf_foldpc; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deq_3_bits_cf_trigger_backendEn_0; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deq_3_bits_cf_trigger_backendEn_1; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deq_3_bits_cf_pd_isRVC; // @[CtrlBlock.scala 271:20]
  wire [1:0] fpDq_io_deq_3_bits_cf_pd_brType; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deq_3_bits_cf_pd_isCall; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deq_3_bits_cf_pd_isRet; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deq_3_bits_cf_pred_taken; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deq_3_bits_cf_storeSetHit; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deq_3_bits_cf_waitForRobIdx_flag; // @[CtrlBlock.scala 271:20]
  wire [4:0] fpDq_io_deq_3_bits_cf_waitForRobIdx_value; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deq_3_bits_cf_loadWaitBit; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deq_3_bits_cf_loadWaitStrict; // @[CtrlBlock.scala 271:20]
  wire [4:0] fpDq_io_deq_3_bits_cf_ssid; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deq_3_bits_cf_ftqPtr_flag; // @[CtrlBlock.scala 271:20]
  wire [2:0] fpDq_io_deq_3_bits_cf_ftqPtr_value; // @[CtrlBlock.scala 271:20]
  wire [2:0] fpDq_io_deq_3_bits_cf_ftqOffset; // @[CtrlBlock.scala 271:20]
  wire [1:0] fpDq_io_deq_3_bits_ctrl_srcType_0; // @[CtrlBlock.scala 271:20]
  wire [1:0] fpDq_io_deq_3_bits_ctrl_srcType_1; // @[CtrlBlock.scala 271:20]
  wire [3:0] fpDq_io_deq_3_bits_ctrl_fuType; // @[CtrlBlock.scala 271:20]
  wire [6:0] fpDq_io_deq_3_bits_ctrl_fuOpType; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deq_3_bits_ctrl_rfWen; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deq_3_bits_ctrl_fpWen; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deq_3_bits_ctrl_flushPipe; // @[CtrlBlock.scala 271:20]
  wire [19:0] fpDq_io_deq_3_bits_ctrl_imm; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deq_3_bits_ctrl_replayInst; // @[CtrlBlock.scala 271:20]
  wire [5:0] fpDq_io_deq_3_bits_psrc_0; // @[CtrlBlock.scala 271:20]
  wire [5:0] fpDq_io_deq_3_bits_psrc_1; // @[CtrlBlock.scala 271:20]
  wire [5:0] fpDq_io_deq_3_bits_pdest; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deq_3_bits_robIdx_flag; // @[CtrlBlock.scala 271:20]
  wire [4:0] fpDq_io_deq_3_bits_robIdx_value; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_redirect_valid; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_redirect_bits_robIdx_flag; // @[CtrlBlock.scala 271:20]
  wire [4:0] fpDq_io_redirect_bits_robIdx_value; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_redirect_bits_level; // @[CtrlBlock.scala 271:20]
  wire [2:0] fpDq_io_deqNext_0_cf_ftqPtr_value; // @[CtrlBlock.scala 271:20]
  wire [2:0] fpDq_io_deqNext_0_cf_ftqOffset; // @[CtrlBlock.scala 271:20]
  wire [1:0] fpDq_io_deqNext_0_ctrl_srcType_0; // @[CtrlBlock.scala 271:20]
  wire [1:0] fpDq_io_deqNext_0_ctrl_srcType_1; // @[CtrlBlock.scala 271:20]
  wire [1:0] fpDq_io_deqNext_0_ctrl_srcType_2; // @[CtrlBlock.scala 271:20]
  wire [3:0] fpDq_io_deqNext_0_ctrl_fuType; // @[CtrlBlock.scala 271:20]
  wire [6:0] fpDq_io_deqNext_0_ctrl_fuOpType; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deqNext_0_ctrl_rfWen; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deqNext_0_ctrl_fpWen; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deqNext_0_ctrl_flushPipe; // @[CtrlBlock.scala 271:20]
  wire [3:0] fpDq_io_deqNext_0_ctrl_selImm; // @[CtrlBlock.scala 271:20]
  wire [19:0] fpDq_io_deqNext_0_ctrl_imm; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deqNext_0_ctrl_replayInst; // @[CtrlBlock.scala 271:20]
  wire [5:0] fpDq_io_deqNext_0_psrc_0; // @[CtrlBlock.scala 271:20]
  wire [5:0] fpDq_io_deqNext_0_psrc_1; // @[CtrlBlock.scala 271:20]
  wire [5:0] fpDq_io_deqNext_0_psrc_2; // @[CtrlBlock.scala 271:20]
  wire [5:0] fpDq_io_deqNext_0_pdest; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deqNext_0_robIdx_flag; // @[CtrlBlock.scala 271:20]
  wire [4:0] fpDq_io_deqNext_0_robIdx_value; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deqNext_0_lqIdx_flag; // @[CtrlBlock.scala 271:20]
  wire [3:0] fpDq_io_deqNext_0_lqIdx_value; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deqNext_0_sqIdx_flag; // @[CtrlBlock.scala 271:20]
  wire [3:0] fpDq_io_deqNext_0_sqIdx_value; // @[CtrlBlock.scala 271:20]
  wire [2:0] fpDq_io_deqNext_1_cf_ftqPtr_value; // @[CtrlBlock.scala 271:20]
  wire [2:0] fpDq_io_deqNext_1_cf_ftqOffset; // @[CtrlBlock.scala 271:20]
  wire [1:0] fpDq_io_deqNext_1_ctrl_srcType_0; // @[CtrlBlock.scala 271:20]
  wire [1:0] fpDq_io_deqNext_1_ctrl_srcType_1; // @[CtrlBlock.scala 271:20]
  wire [1:0] fpDq_io_deqNext_1_ctrl_srcType_2; // @[CtrlBlock.scala 271:20]
  wire [3:0] fpDq_io_deqNext_1_ctrl_fuType; // @[CtrlBlock.scala 271:20]
  wire [6:0] fpDq_io_deqNext_1_ctrl_fuOpType; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deqNext_1_ctrl_rfWen; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deqNext_1_ctrl_fpWen; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deqNext_1_ctrl_flushPipe; // @[CtrlBlock.scala 271:20]
  wire [3:0] fpDq_io_deqNext_1_ctrl_selImm; // @[CtrlBlock.scala 271:20]
  wire [19:0] fpDq_io_deqNext_1_ctrl_imm; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deqNext_1_ctrl_replayInst; // @[CtrlBlock.scala 271:20]
  wire [5:0] fpDq_io_deqNext_1_psrc_0; // @[CtrlBlock.scala 271:20]
  wire [5:0] fpDq_io_deqNext_1_psrc_1; // @[CtrlBlock.scala 271:20]
  wire [5:0] fpDq_io_deqNext_1_psrc_2; // @[CtrlBlock.scala 271:20]
  wire [5:0] fpDq_io_deqNext_1_pdest; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deqNext_1_robIdx_flag; // @[CtrlBlock.scala 271:20]
  wire [4:0] fpDq_io_deqNext_1_robIdx_value; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deqNext_1_lqIdx_flag; // @[CtrlBlock.scala 271:20]
  wire [3:0] fpDq_io_deqNext_1_lqIdx_value; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deqNext_1_sqIdx_flag; // @[CtrlBlock.scala 271:20]
  wire [3:0] fpDq_io_deqNext_1_sqIdx_value; // @[CtrlBlock.scala 271:20]
  wire [2:0] fpDq_io_deqNext_2_cf_ftqPtr_value; // @[CtrlBlock.scala 271:20]
  wire [2:0] fpDq_io_deqNext_2_cf_ftqOffset; // @[CtrlBlock.scala 271:20]
  wire [1:0] fpDq_io_deqNext_2_ctrl_srcType_0; // @[CtrlBlock.scala 271:20]
  wire [1:0] fpDq_io_deqNext_2_ctrl_srcType_1; // @[CtrlBlock.scala 271:20]
  wire [1:0] fpDq_io_deqNext_2_ctrl_srcType_2; // @[CtrlBlock.scala 271:20]
  wire [3:0] fpDq_io_deqNext_2_ctrl_fuType; // @[CtrlBlock.scala 271:20]
  wire [6:0] fpDq_io_deqNext_2_ctrl_fuOpType; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deqNext_2_ctrl_rfWen; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deqNext_2_ctrl_fpWen; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deqNext_2_ctrl_flushPipe; // @[CtrlBlock.scala 271:20]
  wire [3:0] fpDq_io_deqNext_2_ctrl_selImm; // @[CtrlBlock.scala 271:20]
  wire [19:0] fpDq_io_deqNext_2_ctrl_imm; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deqNext_2_ctrl_replayInst; // @[CtrlBlock.scala 271:20]
  wire [5:0] fpDq_io_deqNext_2_psrc_0; // @[CtrlBlock.scala 271:20]
  wire [5:0] fpDq_io_deqNext_2_psrc_1; // @[CtrlBlock.scala 271:20]
  wire [5:0] fpDq_io_deqNext_2_psrc_2; // @[CtrlBlock.scala 271:20]
  wire [5:0] fpDq_io_deqNext_2_pdest; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deqNext_2_robIdx_flag; // @[CtrlBlock.scala 271:20]
  wire [4:0] fpDq_io_deqNext_2_robIdx_value; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deqNext_2_lqIdx_flag; // @[CtrlBlock.scala 271:20]
  wire [3:0] fpDq_io_deqNext_2_lqIdx_value; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deqNext_2_sqIdx_flag; // @[CtrlBlock.scala 271:20]
  wire [3:0] fpDq_io_deqNext_2_sqIdx_value; // @[CtrlBlock.scala 271:20]
  wire [2:0] fpDq_io_deqNext_3_cf_ftqPtr_value; // @[CtrlBlock.scala 271:20]
  wire [2:0] fpDq_io_deqNext_3_cf_ftqOffset; // @[CtrlBlock.scala 271:20]
  wire [1:0] fpDq_io_deqNext_3_ctrl_srcType_0; // @[CtrlBlock.scala 271:20]
  wire [1:0] fpDq_io_deqNext_3_ctrl_srcType_1; // @[CtrlBlock.scala 271:20]
  wire [1:0] fpDq_io_deqNext_3_ctrl_srcType_2; // @[CtrlBlock.scala 271:20]
  wire [3:0] fpDq_io_deqNext_3_ctrl_fuType; // @[CtrlBlock.scala 271:20]
  wire [6:0] fpDq_io_deqNext_3_ctrl_fuOpType; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deqNext_3_ctrl_rfWen; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deqNext_3_ctrl_fpWen; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deqNext_3_ctrl_flushPipe; // @[CtrlBlock.scala 271:20]
  wire [3:0] fpDq_io_deqNext_3_ctrl_selImm; // @[CtrlBlock.scala 271:20]
  wire [19:0] fpDq_io_deqNext_3_ctrl_imm; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deqNext_3_ctrl_replayInst; // @[CtrlBlock.scala 271:20]
  wire [5:0] fpDq_io_deqNext_3_psrc_0; // @[CtrlBlock.scala 271:20]
  wire [5:0] fpDq_io_deqNext_3_psrc_1; // @[CtrlBlock.scala 271:20]
  wire [5:0] fpDq_io_deqNext_3_psrc_2; // @[CtrlBlock.scala 271:20]
  wire [5:0] fpDq_io_deqNext_3_pdest; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deqNext_3_robIdx_flag; // @[CtrlBlock.scala 271:20]
  wire [4:0] fpDq_io_deqNext_3_robIdx_value; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deqNext_3_lqIdx_flag; // @[CtrlBlock.scala 271:20]
  wire [3:0] fpDq_io_deqNext_3_lqIdx_value; // @[CtrlBlock.scala 271:20]
  wire  fpDq_io_deqNext_3_sqIdx_flag; // @[CtrlBlock.scala 271:20]
  wire [3:0] fpDq_io_deqNext_3_sqIdx_value; // @[CtrlBlock.scala 271:20]
  wire [5:0] fpDq_io_perf_0_value; // @[CtrlBlock.scala 271:20]
  wire [5:0] fpDq_io_perf_1_value; // @[CtrlBlock.scala 271:20]
  wire [5:0] fpDq_io_perf_2_value; // @[CtrlBlock.scala 271:20]
  wire [5:0] fpDq_io_perf_3_value; // @[CtrlBlock.scala 271:20]
  wire [5:0] fpDq_io_perf_4_value; // @[CtrlBlock.scala 271:20]
  wire [5:0] fpDq_io_perf_5_value; // @[CtrlBlock.scala 271:20]
  wire [5:0] fpDq_io_perf_6_value; // @[CtrlBlock.scala 271:20]
  wire [5:0] fpDq_io_perf_7_value; // @[CtrlBlock.scala 271:20]
  wire  lsDq_clock; // @[CtrlBlock.scala 272:20]
  wire  lsDq_reset; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_enq_canAccept; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_enq_needAlloc_0; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_enq_needAlloc_1; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_enq_req_0_valid; // @[CtrlBlock.scala 272:20]
  wire [9:0] lsDq_io_enq_req_0_bits_cf_foldpc; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_enq_req_0_bits_cf_trigger_backendEn_0; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_enq_req_0_bits_cf_trigger_backendEn_1; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_enq_req_0_bits_cf_pd_isRVC; // @[CtrlBlock.scala 272:20]
  wire [1:0] lsDq_io_enq_req_0_bits_cf_pd_brType; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_enq_req_0_bits_cf_pd_isCall; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_enq_req_0_bits_cf_pd_isRet; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_enq_req_0_bits_cf_pred_taken; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_enq_req_0_bits_cf_storeSetHit; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_enq_req_0_bits_cf_waitForRobIdx_flag; // @[CtrlBlock.scala 272:20]
  wire [4:0] lsDq_io_enq_req_0_bits_cf_waitForRobIdx_value; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_enq_req_0_bits_cf_loadWaitBit; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_enq_req_0_bits_cf_loadWaitStrict; // @[CtrlBlock.scala 272:20]
  wire [4:0] lsDq_io_enq_req_0_bits_cf_ssid; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_enq_req_0_bits_cf_ftqPtr_flag; // @[CtrlBlock.scala 272:20]
  wire [2:0] lsDq_io_enq_req_0_bits_cf_ftqPtr_value; // @[CtrlBlock.scala 272:20]
  wire [2:0] lsDq_io_enq_req_0_bits_cf_ftqOffset; // @[CtrlBlock.scala 272:20]
  wire [1:0] lsDq_io_enq_req_0_bits_ctrl_srcType_0; // @[CtrlBlock.scala 272:20]
  wire [1:0] lsDq_io_enq_req_0_bits_ctrl_srcType_1; // @[CtrlBlock.scala 272:20]
  wire [1:0] lsDq_io_enq_req_0_bits_ctrl_srcType_2; // @[CtrlBlock.scala 272:20]
  wire [3:0] lsDq_io_enq_req_0_bits_ctrl_fuType; // @[CtrlBlock.scala 272:20]
  wire [6:0] lsDq_io_enq_req_0_bits_ctrl_fuOpType; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_enq_req_0_bits_ctrl_rfWen; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_enq_req_0_bits_ctrl_fpWen; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_enq_req_0_bits_ctrl_flushPipe; // @[CtrlBlock.scala 272:20]
  wire [3:0] lsDq_io_enq_req_0_bits_ctrl_selImm; // @[CtrlBlock.scala 272:20]
  wire [19:0] lsDq_io_enq_req_0_bits_ctrl_imm; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_enq_req_0_bits_ctrl_fpu_isAddSub; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_enq_req_0_bits_ctrl_fpu_typeTagIn; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_enq_req_0_bits_ctrl_fpu_typeTagOut; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_enq_req_0_bits_ctrl_fpu_fromInt; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_enq_req_0_bits_ctrl_fpu_wflags; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_enq_req_0_bits_ctrl_fpu_fpWen; // @[CtrlBlock.scala 272:20]
  wire [1:0] lsDq_io_enq_req_0_bits_ctrl_fpu_fmaCmd; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_enq_req_0_bits_ctrl_fpu_div; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_enq_req_0_bits_ctrl_fpu_sqrt; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_enq_req_0_bits_ctrl_fpu_fcvt; // @[CtrlBlock.scala 272:20]
  wire [1:0] lsDq_io_enq_req_0_bits_ctrl_fpu_typ; // @[CtrlBlock.scala 272:20]
  wire [1:0] lsDq_io_enq_req_0_bits_ctrl_fpu_fmt; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_enq_req_0_bits_ctrl_fpu_ren3; // @[CtrlBlock.scala 272:20]
  wire [2:0] lsDq_io_enq_req_0_bits_ctrl_fpu_rm; // @[CtrlBlock.scala 272:20]
  wire [5:0] lsDq_io_enq_req_0_bits_psrc_0; // @[CtrlBlock.scala 272:20]
  wire [5:0] lsDq_io_enq_req_0_bits_psrc_1; // @[CtrlBlock.scala 272:20]
  wire [5:0] lsDq_io_enq_req_0_bits_psrc_2; // @[CtrlBlock.scala 272:20]
  wire [5:0] lsDq_io_enq_req_0_bits_pdest; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_enq_req_0_bits_robIdx_flag; // @[CtrlBlock.scala 272:20]
  wire [4:0] lsDq_io_enq_req_0_bits_robIdx_value; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_enq_req_1_valid; // @[CtrlBlock.scala 272:20]
  wire [9:0] lsDq_io_enq_req_1_bits_cf_foldpc; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_enq_req_1_bits_cf_trigger_backendEn_0; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_enq_req_1_bits_cf_trigger_backendEn_1; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_enq_req_1_bits_cf_pd_isRVC; // @[CtrlBlock.scala 272:20]
  wire [1:0] lsDq_io_enq_req_1_bits_cf_pd_brType; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_enq_req_1_bits_cf_pd_isCall; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_enq_req_1_bits_cf_pd_isRet; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_enq_req_1_bits_cf_pred_taken; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_enq_req_1_bits_cf_storeSetHit; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_enq_req_1_bits_cf_waitForRobIdx_flag; // @[CtrlBlock.scala 272:20]
  wire [4:0] lsDq_io_enq_req_1_bits_cf_waitForRobIdx_value; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_enq_req_1_bits_cf_loadWaitBit; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_enq_req_1_bits_cf_loadWaitStrict; // @[CtrlBlock.scala 272:20]
  wire [4:0] lsDq_io_enq_req_1_bits_cf_ssid; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_enq_req_1_bits_cf_ftqPtr_flag; // @[CtrlBlock.scala 272:20]
  wire [2:0] lsDq_io_enq_req_1_bits_cf_ftqPtr_value; // @[CtrlBlock.scala 272:20]
  wire [2:0] lsDq_io_enq_req_1_bits_cf_ftqOffset; // @[CtrlBlock.scala 272:20]
  wire [1:0] lsDq_io_enq_req_1_bits_ctrl_srcType_0; // @[CtrlBlock.scala 272:20]
  wire [1:0] lsDq_io_enq_req_1_bits_ctrl_srcType_1; // @[CtrlBlock.scala 272:20]
  wire [1:0] lsDq_io_enq_req_1_bits_ctrl_srcType_2; // @[CtrlBlock.scala 272:20]
  wire [3:0] lsDq_io_enq_req_1_bits_ctrl_fuType; // @[CtrlBlock.scala 272:20]
  wire [6:0] lsDq_io_enq_req_1_bits_ctrl_fuOpType; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_enq_req_1_bits_ctrl_rfWen; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_enq_req_1_bits_ctrl_fpWen; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_enq_req_1_bits_ctrl_flushPipe; // @[CtrlBlock.scala 272:20]
  wire [3:0] lsDq_io_enq_req_1_bits_ctrl_selImm; // @[CtrlBlock.scala 272:20]
  wire [19:0] lsDq_io_enq_req_1_bits_ctrl_imm; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_enq_req_1_bits_ctrl_fpu_isAddSub; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_enq_req_1_bits_ctrl_fpu_typeTagIn; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_enq_req_1_bits_ctrl_fpu_typeTagOut; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_enq_req_1_bits_ctrl_fpu_fromInt; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_enq_req_1_bits_ctrl_fpu_wflags; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_enq_req_1_bits_ctrl_fpu_fpWen; // @[CtrlBlock.scala 272:20]
  wire [1:0] lsDq_io_enq_req_1_bits_ctrl_fpu_fmaCmd; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_enq_req_1_bits_ctrl_fpu_div; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_enq_req_1_bits_ctrl_fpu_sqrt; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_enq_req_1_bits_ctrl_fpu_fcvt; // @[CtrlBlock.scala 272:20]
  wire [1:0] lsDq_io_enq_req_1_bits_ctrl_fpu_typ; // @[CtrlBlock.scala 272:20]
  wire [1:0] lsDq_io_enq_req_1_bits_ctrl_fpu_fmt; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_enq_req_1_bits_ctrl_fpu_ren3; // @[CtrlBlock.scala 272:20]
  wire [2:0] lsDq_io_enq_req_1_bits_ctrl_fpu_rm; // @[CtrlBlock.scala 272:20]
  wire [5:0] lsDq_io_enq_req_1_bits_psrc_0; // @[CtrlBlock.scala 272:20]
  wire [5:0] lsDq_io_enq_req_1_bits_psrc_1; // @[CtrlBlock.scala 272:20]
  wire [5:0] lsDq_io_enq_req_1_bits_psrc_2; // @[CtrlBlock.scala 272:20]
  wire [5:0] lsDq_io_enq_req_1_bits_pdest; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_enq_req_1_bits_robIdx_flag; // @[CtrlBlock.scala 272:20]
  wire [4:0] lsDq_io_enq_req_1_bits_robIdx_value; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deq_0_ready; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deq_0_valid; // @[CtrlBlock.scala 272:20]
  wire [9:0] lsDq_io_deq_0_bits_cf_foldpc; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deq_0_bits_cf_trigger_backendEn_0; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deq_0_bits_cf_trigger_backendEn_1; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deq_0_bits_cf_pd_isRVC; // @[CtrlBlock.scala 272:20]
  wire [1:0] lsDq_io_deq_0_bits_cf_pd_brType; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deq_0_bits_cf_pd_isCall; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deq_0_bits_cf_pd_isRet; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deq_0_bits_cf_pred_taken; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deq_0_bits_cf_storeSetHit; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deq_0_bits_cf_waitForRobIdx_flag; // @[CtrlBlock.scala 272:20]
  wire [4:0] lsDq_io_deq_0_bits_cf_waitForRobIdx_value; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deq_0_bits_cf_loadWaitBit; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deq_0_bits_cf_loadWaitStrict; // @[CtrlBlock.scala 272:20]
  wire [4:0] lsDq_io_deq_0_bits_cf_ssid; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deq_0_bits_cf_ftqPtr_flag; // @[CtrlBlock.scala 272:20]
  wire [2:0] lsDq_io_deq_0_bits_cf_ftqPtr_value; // @[CtrlBlock.scala 272:20]
  wire [2:0] lsDq_io_deq_0_bits_cf_ftqOffset; // @[CtrlBlock.scala 272:20]
  wire [1:0] lsDq_io_deq_0_bits_ctrl_srcType_0; // @[CtrlBlock.scala 272:20]
  wire [1:0] lsDq_io_deq_0_bits_ctrl_srcType_1; // @[CtrlBlock.scala 272:20]
  wire [1:0] lsDq_io_deq_0_bits_ctrl_srcType_2; // @[CtrlBlock.scala 272:20]
  wire [3:0] lsDq_io_deq_0_bits_ctrl_fuType; // @[CtrlBlock.scala 272:20]
  wire [6:0] lsDq_io_deq_0_bits_ctrl_fuOpType; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deq_0_bits_ctrl_rfWen; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deq_0_bits_ctrl_fpWen; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deq_0_bits_ctrl_flushPipe; // @[CtrlBlock.scala 272:20]
  wire [3:0] lsDq_io_deq_0_bits_ctrl_selImm; // @[CtrlBlock.scala 272:20]
  wire [19:0] lsDq_io_deq_0_bits_ctrl_imm; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deq_0_bits_ctrl_fpu_isAddSub; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deq_0_bits_ctrl_fpu_typeTagIn; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deq_0_bits_ctrl_fpu_typeTagOut; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deq_0_bits_ctrl_fpu_fromInt; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deq_0_bits_ctrl_fpu_wflags; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deq_0_bits_ctrl_fpu_fpWen; // @[CtrlBlock.scala 272:20]
  wire [1:0] lsDq_io_deq_0_bits_ctrl_fpu_fmaCmd; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deq_0_bits_ctrl_fpu_div; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deq_0_bits_ctrl_fpu_sqrt; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deq_0_bits_ctrl_fpu_fcvt; // @[CtrlBlock.scala 272:20]
  wire [1:0] lsDq_io_deq_0_bits_ctrl_fpu_typ; // @[CtrlBlock.scala 272:20]
  wire [1:0] lsDq_io_deq_0_bits_ctrl_fpu_fmt; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deq_0_bits_ctrl_fpu_ren3; // @[CtrlBlock.scala 272:20]
  wire [2:0] lsDq_io_deq_0_bits_ctrl_fpu_rm; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deq_0_bits_ctrl_replayInst; // @[CtrlBlock.scala 272:20]
  wire [5:0] lsDq_io_deq_0_bits_psrc_0; // @[CtrlBlock.scala 272:20]
  wire [5:0] lsDq_io_deq_0_bits_psrc_1; // @[CtrlBlock.scala 272:20]
  wire [5:0] lsDq_io_deq_0_bits_psrc_2; // @[CtrlBlock.scala 272:20]
  wire [5:0] lsDq_io_deq_0_bits_pdest; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deq_0_bits_robIdx_flag; // @[CtrlBlock.scala 272:20]
  wire [4:0] lsDq_io_deq_0_bits_robIdx_value; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deq_0_bits_lqIdx_flag; // @[CtrlBlock.scala 272:20]
  wire [3:0] lsDq_io_deq_0_bits_lqIdx_value; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deq_0_bits_sqIdx_flag; // @[CtrlBlock.scala 272:20]
  wire [3:0] lsDq_io_deq_0_bits_sqIdx_value; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deq_1_ready; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deq_1_valid; // @[CtrlBlock.scala 272:20]
  wire [9:0] lsDq_io_deq_1_bits_cf_foldpc; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deq_1_bits_cf_trigger_backendEn_0; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deq_1_bits_cf_trigger_backendEn_1; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deq_1_bits_cf_pd_isRVC; // @[CtrlBlock.scala 272:20]
  wire [1:0] lsDq_io_deq_1_bits_cf_pd_brType; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deq_1_bits_cf_pd_isCall; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deq_1_bits_cf_pd_isRet; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deq_1_bits_cf_pred_taken; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deq_1_bits_cf_storeSetHit; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deq_1_bits_cf_waitForRobIdx_flag; // @[CtrlBlock.scala 272:20]
  wire [4:0] lsDq_io_deq_1_bits_cf_waitForRobIdx_value; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deq_1_bits_cf_loadWaitBit; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deq_1_bits_cf_loadWaitStrict; // @[CtrlBlock.scala 272:20]
  wire [4:0] lsDq_io_deq_1_bits_cf_ssid; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deq_1_bits_cf_ftqPtr_flag; // @[CtrlBlock.scala 272:20]
  wire [2:0] lsDq_io_deq_1_bits_cf_ftqPtr_value; // @[CtrlBlock.scala 272:20]
  wire [2:0] lsDq_io_deq_1_bits_cf_ftqOffset; // @[CtrlBlock.scala 272:20]
  wire [1:0] lsDq_io_deq_1_bits_ctrl_srcType_0; // @[CtrlBlock.scala 272:20]
  wire [1:0] lsDq_io_deq_1_bits_ctrl_srcType_1; // @[CtrlBlock.scala 272:20]
  wire [3:0] lsDq_io_deq_1_bits_ctrl_fuType; // @[CtrlBlock.scala 272:20]
  wire [6:0] lsDq_io_deq_1_bits_ctrl_fuOpType; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deq_1_bits_ctrl_rfWen; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deq_1_bits_ctrl_fpWen; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deq_1_bits_ctrl_flushPipe; // @[CtrlBlock.scala 272:20]
  wire [3:0] lsDq_io_deq_1_bits_ctrl_selImm; // @[CtrlBlock.scala 272:20]
  wire [19:0] lsDq_io_deq_1_bits_ctrl_imm; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deq_1_bits_ctrl_replayInst; // @[CtrlBlock.scala 272:20]
  wire [5:0] lsDq_io_deq_1_bits_psrc_0; // @[CtrlBlock.scala 272:20]
  wire [5:0] lsDq_io_deq_1_bits_psrc_1; // @[CtrlBlock.scala 272:20]
  wire [5:0] lsDq_io_deq_1_bits_pdest; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deq_1_bits_robIdx_flag; // @[CtrlBlock.scala 272:20]
  wire [4:0] lsDq_io_deq_1_bits_robIdx_value; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deq_1_bits_lqIdx_flag; // @[CtrlBlock.scala 272:20]
  wire [3:0] lsDq_io_deq_1_bits_lqIdx_value; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deq_1_bits_sqIdx_flag; // @[CtrlBlock.scala 272:20]
  wire [3:0] lsDq_io_deq_1_bits_sqIdx_value; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deq_2_ready; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deq_2_valid; // @[CtrlBlock.scala 272:20]
  wire [9:0] lsDq_io_deq_2_bits_cf_foldpc; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deq_2_bits_cf_trigger_backendEn_0; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deq_2_bits_cf_trigger_backendEn_1; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deq_2_bits_cf_pd_isRVC; // @[CtrlBlock.scala 272:20]
  wire [1:0] lsDq_io_deq_2_bits_cf_pd_brType; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deq_2_bits_cf_pd_isCall; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deq_2_bits_cf_pd_isRet; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deq_2_bits_cf_pred_taken; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deq_2_bits_cf_storeSetHit; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deq_2_bits_cf_waitForRobIdx_flag; // @[CtrlBlock.scala 272:20]
  wire [4:0] lsDq_io_deq_2_bits_cf_waitForRobIdx_value; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deq_2_bits_cf_loadWaitBit; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deq_2_bits_cf_loadWaitStrict; // @[CtrlBlock.scala 272:20]
  wire [4:0] lsDq_io_deq_2_bits_cf_ssid; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deq_2_bits_cf_ftqPtr_flag; // @[CtrlBlock.scala 272:20]
  wire [2:0] lsDq_io_deq_2_bits_cf_ftqPtr_value; // @[CtrlBlock.scala 272:20]
  wire [2:0] lsDq_io_deq_2_bits_cf_ftqOffset; // @[CtrlBlock.scala 272:20]
  wire [1:0] lsDq_io_deq_2_bits_ctrl_srcType_0; // @[CtrlBlock.scala 272:20]
  wire [1:0] lsDq_io_deq_2_bits_ctrl_srcType_1; // @[CtrlBlock.scala 272:20]
  wire [3:0] lsDq_io_deq_2_bits_ctrl_fuType; // @[CtrlBlock.scala 272:20]
  wire [6:0] lsDq_io_deq_2_bits_ctrl_fuOpType; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deq_2_bits_ctrl_rfWen; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deq_2_bits_ctrl_fpWen; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deq_2_bits_ctrl_flushPipe; // @[CtrlBlock.scala 272:20]
  wire [19:0] lsDq_io_deq_2_bits_ctrl_imm; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deq_2_bits_ctrl_replayInst; // @[CtrlBlock.scala 272:20]
  wire [5:0] lsDq_io_deq_2_bits_psrc_0; // @[CtrlBlock.scala 272:20]
  wire [5:0] lsDq_io_deq_2_bits_psrc_1; // @[CtrlBlock.scala 272:20]
  wire [5:0] lsDq_io_deq_2_bits_pdest; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deq_2_bits_robIdx_flag; // @[CtrlBlock.scala 272:20]
  wire [4:0] lsDq_io_deq_2_bits_robIdx_value; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deq_3_ready; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deq_3_valid; // @[CtrlBlock.scala 272:20]
  wire [9:0] lsDq_io_deq_3_bits_cf_foldpc; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deq_3_bits_cf_trigger_backendEn_0; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deq_3_bits_cf_trigger_backendEn_1; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deq_3_bits_cf_pd_isRVC; // @[CtrlBlock.scala 272:20]
  wire [1:0] lsDq_io_deq_3_bits_cf_pd_brType; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deq_3_bits_cf_pd_isCall; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deq_3_bits_cf_pd_isRet; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deq_3_bits_cf_pred_taken; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deq_3_bits_cf_storeSetHit; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deq_3_bits_cf_waitForRobIdx_flag; // @[CtrlBlock.scala 272:20]
  wire [4:0] lsDq_io_deq_3_bits_cf_waitForRobIdx_value; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deq_3_bits_cf_loadWaitBit; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deq_3_bits_cf_loadWaitStrict; // @[CtrlBlock.scala 272:20]
  wire [4:0] lsDq_io_deq_3_bits_cf_ssid; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deq_3_bits_cf_ftqPtr_flag; // @[CtrlBlock.scala 272:20]
  wire [2:0] lsDq_io_deq_3_bits_cf_ftqPtr_value; // @[CtrlBlock.scala 272:20]
  wire [2:0] lsDq_io_deq_3_bits_cf_ftqOffset; // @[CtrlBlock.scala 272:20]
  wire [1:0] lsDq_io_deq_3_bits_ctrl_srcType_0; // @[CtrlBlock.scala 272:20]
  wire [1:0] lsDq_io_deq_3_bits_ctrl_srcType_1; // @[CtrlBlock.scala 272:20]
  wire [3:0] lsDq_io_deq_3_bits_ctrl_fuType; // @[CtrlBlock.scala 272:20]
  wire [6:0] lsDq_io_deq_3_bits_ctrl_fuOpType; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deq_3_bits_ctrl_rfWen; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deq_3_bits_ctrl_fpWen; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deq_3_bits_ctrl_flushPipe; // @[CtrlBlock.scala 272:20]
  wire [19:0] lsDq_io_deq_3_bits_ctrl_imm; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deq_3_bits_ctrl_replayInst; // @[CtrlBlock.scala 272:20]
  wire [5:0] lsDq_io_deq_3_bits_psrc_0; // @[CtrlBlock.scala 272:20]
  wire [5:0] lsDq_io_deq_3_bits_psrc_1; // @[CtrlBlock.scala 272:20]
  wire [5:0] lsDq_io_deq_3_bits_pdest; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deq_3_bits_robIdx_flag; // @[CtrlBlock.scala 272:20]
  wire [4:0] lsDq_io_deq_3_bits_robIdx_value; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_redirect_valid; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_redirect_bits_robIdx_flag; // @[CtrlBlock.scala 272:20]
  wire [4:0] lsDq_io_redirect_bits_robIdx_value; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_redirect_bits_level; // @[CtrlBlock.scala 272:20]
  wire [2:0] lsDq_io_deqNext_0_cf_ftqPtr_value; // @[CtrlBlock.scala 272:20]
  wire [2:0] lsDq_io_deqNext_0_cf_ftqOffset; // @[CtrlBlock.scala 272:20]
  wire [1:0] lsDq_io_deqNext_0_ctrl_srcType_0; // @[CtrlBlock.scala 272:20]
  wire [1:0] lsDq_io_deqNext_0_ctrl_srcType_1; // @[CtrlBlock.scala 272:20]
  wire [1:0] lsDq_io_deqNext_0_ctrl_srcType_2; // @[CtrlBlock.scala 272:20]
  wire [3:0] lsDq_io_deqNext_0_ctrl_fuType; // @[CtrlBlock.scala 272:20]
  wire [6:0] lsDq_io_deqNext_0_ctrl_fuOpType; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deqNext_0_ctrl_rfWen; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deqNext_0_ctrl_fpWen; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deqNext_0_ctrl_flushPipe; // @[CtrlBlock.scala 272:20]
  wire [3:0] lsDq_io_deqNext_0_ctrl_selImm; // @[CtrlBlock.scala 272:20]
  wire [19:0] lsDq_io_deqNext_0_ctrl_imm; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deqNext_0_ctrl_replayInst; // @[CtrlBlock.scala 272:20]
  wire [5:0] lsDq_io_deqNext_0_psrc_0; // @[CtrlBlock.scala 272:20]
  wire [5:0] lsDq_io_deqNext_0_psrc_1; // @[CtrlBlock.scala 272:20]
  wire [5:0] lsDq_io_deqNext_0_psrc_2; // @[CtrlBlock.scala 272:20]
  wire [5:0] lsDq_io_deqNext_0_pdest; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deqNext_0_robIdx_flag; // @[CtrlBlock.scala 272:20]
  wire [4:0] lsDq_io_deqNext_0_robIdx_value; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deqNext_0_lqIdx_flag; // @[CtrlBlock.scala 272:20]
  wire [3:0] lsDq_io_deqNext_0_lqIdx_value; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deqNext_0_sqIdx_flag; // @[CtrlBlock.scala 272:20]
  wire [3:0] lsDq_io_deqNext_0_sqIdx_value; // @[CtrlBlock.scala 272:20]
  wire [2:0] lsDq_io_deqNext_1_cf_ftqPtr_value; // @[CtrlBlock.scala 272:20]
  wire [2:0] lsDq_io_deqNext_1_cf_ftqOffset; // @[CtrlBlock.scala 272:20]
  wire [1:0] lsDq_io_deqNext_1_ctrl_srcType_0; // @[CtrlBlock.scala 272:20]
  wire [1:0] lsDq_io_deqNext_1_ctrl_srcType_1; // @[CtrlBlock.scala 272:20]
  wire [1:0] lsDq_io_deqNext_1_ctrl_srcType_2; // @[CtrlBlock.scala 272:20]
  wire [3:0] lsDq_io_deqNext_1_ctrl_fuType; // @[CtrlBlock.scala 272:20]
  wire [6:0] lsDq_io_deqNext_1_ctrl_fuOpType; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deqNext_1_ctrl_rfWen; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deqNext_1_ctrl_fpWen; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deqNext_1_ctrl_flushPipe; // @[CtrlBlock.scala 272:20]
  wire [3:0] lsDq_io_deqNext_1_ctrl_selImm; // @[CtrlBlock.scala 272:20]
  wire [19:0] lsDq_io_deqNext_1_ctrl_imm; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deqNext_1_ctrl_replayInst; // @[CtrlBlock.scala 272:20]
  wire [5:0] lsDq_io_deqNext_1_psrc_0; // @[CtrlBlock.scala 272:20]
  wire [5:0] lsDq_io_deqNext_1_psrc_1; // @[CtrlBlock.scala 272:20]
  wire [5:0] lsDq_io_deqNext_1_psrc_2; // @[CtrlBlock.scala 272:20]
  wire [5:0] lsDq_io_deqNext_1_pdest; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deqNext_1_robIdx_flag; // @[CtrlBlock.scala 272:20]
  wire [4:0] lsDq_io_deqNext_1_robIdx_value; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deqNext_1_lqIdx_flag; // @[CtrlBlock.scala 272:20]
  wire [3:0] lsDq_io_deqNext_1_lqIdx_value; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deqNext_1_sqIdx_flag; // @[CtrlBlock.scala 272:20]
  wire [3:0] lsDq_io_deqNext_1_sqIdx_value; // @[CtrlBlock.scala 272:20]
  wire [2:0] lsDq_io_deqNext_2_cf_ftqPtr_value; // @[CtrlBlock.scala 272:20]
  wire [2:0] lsDq_io_deqNext_2_cf_ftqOffset; // @[CtrlBlock.scala 272:20]
  wire [1:0] lsDq_io_deqNext_2_ctrl_srcType_0; // @[CtrlBlock.scala 272:20]
  wire [1:0] lsDq_io_deqNext_2_ctrl_srcType_1; // @[CtrlBlock.scala 272:20]
  wire [1:0] lsDq_io_deqNext_2_ctrl_srcType_2; // @[CtrlBlock.scala 272:20]
  wire [3:0] lsDq_io_deqNext_2_ctrl_fuType; // @[CtrlBlock.scala 272:20]
  wire [6:0] lsDq_io_deqNext_2_ctrl_fuOpType; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deqNext_2_ctrl_rfWen; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deqNext_2_ctrl_fpWen; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deqNext_2_ctrl_flushPipe; // @[CtrlBlock.scala 272:20]
  wire [3:0] lsDq_io_deqNext_2_ctrl_selImm; // @[CtrlBlock.scala 272:20]
  wire [19:0] lsDq_io_deqNext_2_ctrl_imm; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deqNext_2_ctrl_replayInst; // @[CtrlBlock.scala 272:20]
  wire [5:0] lsDq_io_deqNext_2_psrc_0; // @[CtrlBlock.scala 272:20]
  wire [5:0] lsDq_io_deqNext_2_psrc_1; // @[CtrlBlock.scala 272:20]
  wire [5:0] lsDq_io_deqNext_2_psrc_2; // @[CtrlBlock.scala 272:20]
  wire [5:0] lsDq_io_deqNext_2_pdest; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deqNext_2_robIdx_flag; // @[CtrlBlock.scala 272:20]
  wire [4:0] lsDq_io_deqNext_2_robIdx_value; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deqNext_2_lqIdx_flag; // @[CtrlBlock.scala 272:20]
  wire [3:0] lsDq_io_deqNext_2_lqIdx_value; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deqNext_2_sqIdx_flag; // @[CtrlBlock.scala 272:20]
  wire [3:0] lsDq_io_deqNext_2_sqIdx_value; // @[CtrlBlock.scala 272:20]
  wire [2:0] lsDq_io_deqNext_3_cf_ftqPtr_value; // @[CtrlBlock.scala 272:20]
  wire [2:0] lsDq_io_deqNext_3_cf_ftqOffset; // @[CtrlBlock.scala 272:20]
  wire [1:0] lsDq_io_deqNext_3_ctrl_srcType_0; // @[CtrlBlock.scala 272:20]
  wire [1:0] lsDq_io_deqNext_3_ctrl_srcType_1; // @[CtrlBlock.scala 272:20]
  wire [1:0] lsDq_io_deqNext_3_ctrl_srcType_2; // @[CtrlBlock.scala 272:20]
  wire [3:0] lsDq_io_deqNext_3_ctrl_fuType; // @[CtrlBlock.scala 272:20]
  wire [6:0] lsDq_io_deqNext_3_ctrl_fuOpType; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deqNext_3_ctrl_rfWen; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deqNext_3_ctrl_fpWen; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deqNext_3_ctrl_flushPipe; // @[CtrlBlock.scala 272:20]
  wire [3:0] lsDq_io_deqNext_3_ctrl_selImm; // @[CtrlBlock.scala 272:20]
  wire [19:0] lsDq_io_deqNext_3_ctrl_imm; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deqNext_3_ctrl_replayInst; // @[CtrlBlock.scala 272:20]
  wire [5:0] lsDq_io_deqNext_3_psrc_0; // @[CtrlBlock.scala 272:20]
  wire [5:0] lsDq_io_deqNext_3_psrc_1; // @[CtrlBlock.scala 272:20]
  wire [5:0] lsDq_io_deqNext_3_psrc_2; // @[CtrlBlock.scala 272:20]
  wire [5:0] lsDq_io_deqNext_3_pdest; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deqNext_3_robIdx_flag; // @[CtrlBlock.scala 272:20]
  wire [4:0] lsDq_io_deqNext_3_robIdx_value; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deqNext_3_lqIdx_flag; // @[CtrlBlock.scala 272:20]
  wire [3:0] lsDq_io_deqNext_3_lqIdx_value; // @[CtrlBlock.scala 272:20]
  wire  lsDq_io_deqNext_3_sqIdx_flag; // @[CtrlBlock.scala 272:20]
  wire [3:0] lsDq_io_deqNext_3_sqIdx_value; // @[CtrlBlock.scala 272:20]
  wire [5:0] lsDq_io_perf_0_value; // @[CtrlBlock.scala 272:20]
  wire [5:0] lsDq_io_perf_1_value; // @[CtrlBlock.scala 272:20]
  wire [5:0] lsDq_io_perf_2_value; // @[CtrlBlock.scala 272:20]
  wire [5:0] lsDq_io_perf_3_value; // @[CtrlBlock.scala 272:20]
  wire [5:0] lsDq_io_perf_4_value; // @[CtrlBlock.scala 272:20]
  wire [5:0] lsDq_io_perf_5_value; // @[CtrlBlock.scala 272:20]
  wire [5:0] lsDq_io_perf_6_value; // @[CtrlBlock.scala 272:20]
  wire [5:0] lsDq_io_perf_7_value; // @[CtrlBlock.scala 272:20]
  wire  redirectGen_clock; // @[CtrlBlock.scala 273:27]
  wire  redirectGen_reset; // @[CtrlBlock.scala 273:27]
  wire  redirectGen_io_exuMispredict_0_valid; // @[CtrlBlock.scala 273:27]
  wire  redirectGen_io_exuMispredict_0_bits_uop_cf_pd_isRVC; // @[CtrlBlock.scala 273:27]
  wire [1:0] redirectGen_io_exuMispredict_0_bits_uop_cf_pd_brType; // @[CtrlBlock.scala 273:27]
  wire  redirectGen_io_exuMispredict_0_bits_uop_cf_pd_isCall; // @[CtrlBlock.scala 273:27]
  wire  redirectGen_io_exuMispredict_0_bits_uop_cf_pd_isRet; // @[CtrlBlock.scala 273:27]
  wire [19:0] redirectGen_io_exuMispredict_0_bits_uop_ctrl_imm; // @[CtrlBlock.scala 273:27]
  wire  redirectGen_io_exuMispredict_0_bits_redirect_robIdx_flag; // @[CtrlBlock.scala 273:27]
  wire [4:0] redirectGen_io_exuMispredict_0_bits_redirect_robIdx_value; // @[CtrlBlock.scala 273:27]
  wire  redirectGen_io_exuMispredict_0_bits_redirect_ftqIdx_flag; // @[CtrlBlock.scala 273:27]
  wire [2:0] redirectGen_io_exuMispredict_0_bits_redirect_ftqIdx_value; // @[CtrlBlock.scala 273:27]
  wire [2:0] redirectGen_io_exuMispredict_0_bits_redirect_ftqOffset; // @[CtrlBlock.scala 273:27]
  wire [38:0] redirectGen_io_exuMispredict_0_bits_redirect_cfiUpdate_target; // @[CtrlBlock.scala 273:27]
  wire  redirectGen_io_exuMispredict_0_bits_redirect_cfiUpdate_isMisPred; // @[CtrlBlock.scala 273:27]
  wire  redirectGen_io_exuMispredict_1_valid; // @[CtrlBlock.scala 273:27]
  wire  redirectGen_io_exuMispredict_1_bits_uop_cf_pd_isRVC; // @[CtrlBlock.scala 273:27]
  wire [1:0] redirectGen_io_exuMispredict_1_bits_uop_cf_pd_brType; // @[CtrlBlock.scala 273:27]
  wire  redirectGen_io_exuMispredict_1_bits_uop_cf_pd_isCall; // @[CtrlBlock.scala 273:27]
  wire  redirectGen_io_exuMispredict_1_bits_uop_cf_pd_isRet; // @[CtrlBlock.scala 273:27]
  wire [19:0] redirectGen_io_exuMispredict_1_bits_uop_ctrl_imm; // @[CtrlBlock.scala 273:27]
  wire  redirectGen_io_exuMispredict_1_bits_redirect_robIdx_flag; // @[CtrlBlock.scala 273:27]
  wire [4:0] redirectGen_io_exuMispredict_1_bits_redirect_robIdx_value; // @[CtrlBlock.scala 273:27]
  wire  redirectGen_io_exuMispredict_1_bits_redirect_ftqIdx_flag; // @[CtrlBlock.scala 273:27]
  wire [2:0] redirectGen_io_exuMispredict_1_bits_redirect_ftqIdx_value; // @[CtrlBlock.scala 273:27]
  wire [2:0] redirectGen_io_exuMispredict_1_bits_redirect_ftqOffset; // @[CtrlBlock.scala 273:27]
  wire  redirectGen_io_exuMispredict_1_bits_redirect_cfiUpdate_taken; // @[CtrlBlock.scala 273:27]
  wire  redirectGen_io_exuMispredict_1_bits_redirect_cfiUpdate_isMisPred; // @[CtrlBlock.scala 273:27]
  wire  redirectGen_io_exuMispredict_2_valid; // @[CtrlBlock.scala 273:27]
  wire  redirectGen_io_exuMispredict_2_bits_uop_cf_pd_isRVC; // @[CtrlBlock.scala 273:27]
  wire [1:0] redirectGen_io_exuMispredict_2_bits_uop_cf_pd_brType; // @[CtrlBlock.scala 273:27]
  wire  redirectGen_io_exuMispredict_2_bits_uop_cf_pd_isCall; // @[CtrlBlock.scala 273:27]
  wire  redirectGen_io_exuMispredict_2_bits_uop_cf_pd_isRet; // @[CtrlBlock.scala 273:27]
  wire [19:0] redirectGen_io_exuMispredict_2_bits_uop_ctrl_imm; // @[CtrlBlock.scala 273:27]
  wire  redirectGen_io_exuMispredict_2_bits_redirect_robIdx_flag; // @[CtrlBlock.scala 273:27]
  wire [4:0] redirectGen_io_exuMispredict_2_bits_redirect_robIdx_value; // @[CtrlBlock.scala 273:27]
  wire  redirectGen_io_exuMispredict_2_bits_redirect_ftqIdx_flag; // @[CtrlBlock.scala 273:27]
  wire [2:0] redirectGen_io_exuMispredict_2_bits_redirect_ftqIdx_value; // @[CtrlBlock.scala 273:27]
  wire [2:0] redirectGen_io_exuMispredict_2_bits_redirect_ftqOffset; // @[CtrlBlock.scala 273:27]
  wire  redirectGen_io_exuMispredict_2_bits_redirect_cfiUpdate_taken; // @[CtrlBlock.scala 273:27]
  wire  redirectGen_io_exuMispredict_2_bits_redirect_cfiUpdate_isMisPred; // @[CtrlBlock.scala 273:27]
  wire  redirectGen_io_loadReplay_valid; // @[CtrlBlock.scala 273:27]
  wire  redirectGen_io_loadReplay_bits_robIdx_flag; // @[CtrlBlock.scala 273:27]
  wire [4:0] redirectGen_io_loadReplay_bits_robIdx_value; // @[CtrlBlock.scala 273:27]
  wire  redirectGen_io_loadReplay_bits_ftqIdx_flag; // @[CtrlBlock.scala 273:27]
  wire [2:0] redirectGen_io_loadReplay_bits_ftqIdx_value; // @[CtrlBlock.scala 273:27]
  wire [2:0] redirectGen_io_loadReplay_bits_ftqOffset; // @[CtrlBlock.scala 273:27]
  wire [2:0] redirectGen_io_loadReplay_bits_stFtqIdx_value; // @[CtrlBlock.scala 273:27]
  wire [2:0] redirectGen_io_loadReplay_bits_stFtqOffset; // @[CtrlBlock.scala 273:27]
  wire  redirectGen_io_flush; // @[CtrlBlock.scala 273:27]
  wire [2:0] redirectGen_io_redirectPcRead_ptr_value; // @[CtrlBlock.scala 273:27]
  wire [2:0] redirectGen_io_redirectPcRead_offset; // @[CtrlBlock.scala 273:27]
  wire [38:0] redirectGen_io_redirectPcRead_data; // @[CtrlBlock.scala 273:27]
  wire  redirectGen_io_stage2Redirect_valid; // @[CtrlBlock.scala 273:27]
  wire  redirectGen_io_stage2Redirect_bits_robIdx_flag; // @[CtrlBlock.scala 273:27]
  wire [4:0] redirectGen_io_stage2Redirect_bits_robIdx_value; // @[CtrlBlock.scala 273:27]
  wire  redirectGen_io_stage2Redirect_bits_ftqIdx_flag; // @[CtrlBlock.scala 273:27]
  wire [2:0] redirectGen_io_stage2Redirect_bits_ftqIdx_value; // @[CtrlBlock.scala 273:27]
  wire [2:0] redirectGen_io_stage2Redirect_bits_ftqOffset; // @[CtrlBlock.scala 273:27]
  wire  redirectGen_io_stage2Redirect_bits_level; // @[CtrlBlock.scala 273:27]
  wire [38:0] redirectGen_io_stage2Redirect_bits_cfiUpdate_pc; // @[CtrlBlock.scala 273:27]
  wire  redirectGen_io_stage2Redirect_bits_cfiUpdate_pd_isRVC; // @[CtrlBlock.scala 273:27]
  wire [1:0] redirectGen_io_stage2Redirect_bits_cfiUpdate_pd_brType; // @[CtrlBlock.scala 273:27]
  wire  redirectGen_io_stage2Redirect_bits_cfiUpdate_pd_isCall; // @[CtrlBlock.scala 273:27]
  wire  redirectGen_io_stage2Redirect_bits_cfiUpdate_pd_isRet; // @[CtrlBlock.scala 273:27]
  wire [38:0] redirectGen_io_stage2Redirect_bits_cfiUpdate_target; // @[CtrlBlock.scala 273:27]
  wire  redirectGen_io_stage2Redirect_bits_cfiUpdate_taken; // @[CtrlBlock.scala 273:27]
  wire  redirectGen_io_stage2Redirect_bits_cfiUpdate_isMisPred; // @[CtrlBlock.scala 273:27]
  wire  redirectGen_io_memPredUpdate_valid; // @[CtrlBlock.scala 273:27]
  wire [9:0] redirectGen_io_memPredUpdate_ldpc; // @[CtrlBlock.scala 273:27]
  wire [9:0] redirectGen_io_memPredUpdate_stpc; // @[CtrlBlock.scala 273:27]
  wire [2:0] redirectGen_io_memPredPcRead_ptr_value; // @[CtrlBlock.scala 273:27]
  wire [2:0] redirectGen_io_memPredPcRead_offset; // @[CtrlBlock.scala 273:27]
  wire [38:0] redirectGen_io_memPredPcRead_data; // @[CtrlBlock.scala 273:27]
  wire  pcMem_clock; // @[CtrlBlock.scala 283:21]
  wire [2:0] pcMem_io_raddr_0; // @[CtrlBlock.scala 283:21]
  wire [2:0] pcMem_io_raddr_2; // @[CtrlBlock.scala 283:21]
  wire [2:0] pcMem_io_raddr_3; // @[CtrlBlock.scala 283:21]
  wire [2:0] pcMem_io_raddr_4; // @[CtrlBlock.scala 283:21]
  wire [2:0] pcMem_io_raddr_7; // @[CtrlBlock.scala 283:21]
  wire [38:0] pcMem_io_rdata_0_startAddr; // @[CtrlBlock.scala 283:21]
  wire [38:0] pcMem_io_rdata_0_nextLineAddr; // @[CtrlBlock.scala 283:21]
  wire  pcMem_io_rdata_0_isNextMask_0; // @[CtrlBlock.scala 283:21]
  wire  pcMem_io_rdata_0_isNextMask_1; // @[CtrlBlock.scala 283:21]
  wire  pcMem_io_rdata_0_isNextMask_2; // @[CtrlBlock.scala 283:21]
  wire  pcMem_io_rdata_0_isNextMask_3; // @[CtrlBlock.scala 283:21]
  wire  pcMem_io_rdata_0_isNextMask_4; // @[CtrlBlock.scala 283:21]
  wire  pcMem_io_rdata_0_isNextMask_5; // @[CtrlBlock.scala 283:21]
  wire  pcMem_io_rdata_0_isNextMask_6; // @[CtrlBlock.scala 283:21]
  wire  pcMem_io_rdata_0_isNextMask_7; // @[CtrlBlock.scala 283:21]
  wire [38:0] pcMem_io_rdata_2_startAddr; // @[CtrlBlock.scala 283:21]
  wire [38:0] pcMem_io_rdata_2_nextLineAddr; // @[CtrlBlock.scala 283:21]
  wire  pcMem_io_rdata_2_isNextMask_0; // @[CtrlBlock.scala 283:21]
  wire  pcMem_io_rdata_2_isNextMask_1; // @[CtrlBlock.scala 283:21]
  wire  pcMem_io_rdata_2_isNextMask_2; // @[CtrlBlock.scala 283:21]
  wire  pcMem_io_rdata_2_isNextMask_3; // @[CtrlBlock.scala 283:21]
  wire  pcMem_io_rdata_2_isNextMask_4; // @[CtrlBlock.scala 283:21]
  wire  pcMem_io_rdata_2_isNextMask_5; // @[CtrlBlock.scala 283:21]
  wire  pcMem_io_rdata_2_isNextMask_6; // @[CtrlBlock.scala 283:21]
  wire  pcMem_io_rdata_2_isNextMask_7; // @[CtrlBlock.scala 283:21]
  wire [38:0] pcMem_io_rdata_3_startAddr; // @[CtrlBlock.scala 283:21]
  wire [38:0] pcMem_io_rdata_3_nextLineAddr; // @[CtrlBlock.scala 283:21]
  wire  pcMem_io_rdata_3_isNextMask_0; // @[CtrlBlock.scala 283:21]
  wire  pcMem_io_rdata_3_isNextMask_1; // @[CtrlBlock.scala 283:21]
  wire  pcMem_io_rdata_3_isNextMask_2; // @[CtrlBlock.scala 283:21]
  wire  pcMem_io_rdata_3_isNextMask_3; // @[CtrlBlock.scala 283:21]
  wire  pcMem_io_rdata_3_isNextMask_4; // @[CtrlBlock.scala 283:21]
  wire  pcMem_io_rdata_3_isNextMask_5; // @[CtrlBlock.scala 283:21]
  wire  pcMem_io_rdata_3_isNextMask_6; // @[CtrlBlock.scala 283:21]
  wire  pcMem_io_rdata_3_isNextMask_7; // @[CtrlBlock.scala 283:21]
  wire [38:0] pcMem_io_rdata_4_startAddr; // @[CtrlBlock.scala 283:21]
  wire [38:0] pcMem_io_rdata_7_startAddr; // @[CtrlBlock.scala 283:21]
  wire [38:0] pcMem_io_rdata_7_nextLineAddr; // @[CtrlBlock.scala 283:21]
  wire  pcMem_io_rdata_7_isNextMask_0; // @[CtrlBlock.scala 283:21]
  wire  pcMem_io_rdata_7_isNextMask_1; // @[CtrlBlock.scala 283:21]
  wire  pcMem_io_rdata_7_isNextMask_2; // @[CtrlBlock.scala 283:21]
  wire  pcMem_io_rdata_7_isNextMask_3; // @[CtrlBlock.scala 283:21]
  wire  pcMem_io_rdata_7_isNextMask_4; // @[CtrlBlock.scala 283:21]
  wire  pcMem_io_rdata_7_isNextMask_5; // @[CtrlBlock.scala 283:21]
  wire  pcMem_io_rdata_7_isNextMask_6; // @[CtrlBlock.scala 283:21]
  wire  pcMem_io_rdata_7_isNextMask_7; // @[CtrlBlock.scala 283:21]
  wire  pcMem_io_wen_0; // @[CtrlBlock.scala 283:21]
  wire [2:0] pcMem_io_waddr_0; // @[CtrlBlock.scala 283:21]
  wire [38:0] pcMem_io_wdata_0_startAddr; // @[CtrlBlock.scala 283:21]
  wire [38:0] pcMem_io_wdata_0_nextLineAddr; // @[CtrlBlock.scala 283:21]
  wire  pcMem_io_wdata_0_isNextMask_0; // @[CtrlBlock.scala 283:21]
  wire  pcMem_io_wdata_0_isNextMask_1; // @[CtrlBlock.scala 283:21]
  wire  pcMem_io_wdata_0_isNextMask_2; // @[CtrlBlock.scala 283:21]
  wire  pcMem_io_wdata_0_isNextMask_3; // @[CtrlBlock.scala 283:21]
  wire  pcMem_io_wdata_0_isNextMask_4; // @[CtrlBlock.scala 283:21]
  wire  pcMem_io_wdata_0_isNextMask_5; // @[CtrlBlock.scala 283:21]
  wire  pcMem_io_wdata_0_isNextMask_6; // @[CtrlBlock.scala 283:21]
  wire  pcMem_io_wdata_0_isNextMask_7; // @[CtrlBlock.scala 283:21]
  wire  frontendFlushValid_delay_clock; // @[Hold.scala 97:23]
  wire  frontendFlushValid_delay_io_in; // @[Hold.scala 97:23]
  wire  frontendFlushValid_delay_io_out; // @[Hold.scala 97:23]
  wire  pc_from_csr_delay_clock; // @[Hold.scala 97:23]
  wire  pc_from_csr_delay_io_in; // @[Hold.scala 97:23]
  wire  pc_from_csr_delay_io_out; // @[Hold.scala 97:23]
  wire  lfst_clock; // @[CtrlBlock.scala 425:20]
  wire  lfst_reset; // @[CtrlBlock.scala 425:20]
  wire  lfst_io_redirect_valid; // @[CtrlBlock.scala 425:20]
  wire  lfst_io_redirect_bits_robIdx_flag; // @[CtrlBlock.scala 425:20]
  wire [4:0] lfst_io_redirect_bits_robIdx_value; // @[CtrlBlock.scala 425:20]
  wire  lfst_io_redirect_bits_level; // @[CtrlBlock.scala 425:20]
  wire  lfst_io_dispatch_req_0_valid; // @[CtrlBlock.scala 425:20]
  wire  lfst_io_dispatch_req_0_bits_isstore; // @[CtrlBlock.scala 425:20]
  wire [4:0] lfst_io_dispatch_req_0_bits_ssid; // @[CtrlBlock.scala 425:20]
  wire  lfst_io_dispatch_req_0_bits_robIdx_flag; // @[CtrlBlock.scala 425:20]
  wire [4:0] lfst_io_dispatch_req_0_bits_robIdx_value; // @[CtrlBlock.scala 425:20]
  wire  lfst_io_dispatch_req_1_valid; // @[CtrlBlock.scala 425:20]
  wire  lfst_io_dispatch_req_1_bits_isstore; // @[CtrlBlock.scala 425:20]
  wire [4:0] lfst_io_dispatch_req_1_bits_ssid; // @[CtrlBlock.scala 425:20]
  wire  lfst_io_dispatch_req_1_bits_robIdx_flag; // @[CtrlBlock.scala 425:20]
  wire [4:0] lfst_io_dispatch_req_1_bits_robIdx_value; // @[CtrlBlock.scala 425:20]
  wire  lfst_io_dispatch_resp_0_bits_shouldWait; // @[CtrlBlock.scala 425:20]
  wire  lfst_io_dispatch_resp_0_bits_robIdx_flag; // @[CtrlBlock.scala 425:20]
  wire [4:0] lfst_io_dispatch_resp_0_bits_robIdx_value; // @[CtrlBlock.scala 425:20]
  wire  lfst_io_dispatch_resp_1_bits_shouldWait; // @[CtrlBlock.scala 425:20]
  wire  lfst_io_dispatch_resp_1_bits_robIdx_flag; // @[CtrlBlock.scala 425:20]
  wire [4:0] lfst_io_dispatch_resp_1_bits_robIdx_value; // @[CtrlBlock.scala 425:20]
  wire  lfst_io_storeIssue_0_valid; // @[CtrlBlock.scala 425:20]
  wire  lfst_io_storeIssue_0_bits_uop_cf_storeSetHit; // @[CtrlBlock.scala 425:20]
  wire [4:0] lfst_io_storeIssue_0_bits_uop_cf_ssid; // @[CtrlBlock.scala 425:20]
  wire [4:0] lfst_io_storeIssue_0_bits_uop_robIdx_value; // @[CtrlBlock.scala 425:20]
  wire  lfst_io_storeIssue_1_valid; // @[CtrlBlock.scala 425:20]
  wire  lfst_io_storeIssue_1_bits_uop_cf_storeSetHit; // @[CtrlBlock.scala 425:20]
  wire [4:0] lfst_io_storeIssue_1_bits_uop_cf_ssid; // @[CtrlBlock.scala 425:20]
  wire [4:0] lfst_io_storeIssue_1_bits_uop_robIdx_value; // @[CtrlBlock.scala 425:20]
  wire  lfst_io_csrCtrl_lvpred_disable; // @[CtrlBlock.scala 425:20]
  wire  lfst_io_csrCtrl_no_spec_load; // @[CtrlBlock.scala 425:20]
  wire  lfst_io_csrCtrl_storeset_wait_store; // @[CtrlBlock.scala 425:20]
  wire  lsqCtrl_clock; // @[CtrlBlock.scala 519:27]
  wire  lsqCtrl_reset; // @[CtrlBlock.scala 519:27]
  wire  lsqCtrl_io_redirect_valid; // @[CtrlBlock.scala 519:27]
  wire  lsqCtrl_io_enq_canAccept; // @[CtrlBlock.scala 519:27]
  wire [1:0] lsqCtrl_io_enq_needAlloc_0; // @[CtrlBlock.scala 519:27]
  wire [1:0] lsqCtrl_io_enq_needAlloc_1; // @[CtrlBlock.scala 519:27]
  wire [1:0] lsqCtrl_io_enq_needAlloc_2; // @[CtrlBlock.scala 519:27]
  wire [1:0] lsqCtrl_io_enq_needAlloc_3; // @[CtrlBlock.scala 519:27]
  wire  lsqCtrl_io_enq_req_0_valid; // @[CtrlBlock.scala 519:27]
  wire  lsqCtrl_io_enq_req_0_bits_cf_trigger_backendEn_0; // @[CtrlBlock.scala 519:27]
  wire  lsqCtrl_io_enq_req_0_bits_cf_trigger_backendEn_1; // @[CtrlBlock.scala 519:27]
  wire [6:0] lsqCtrl_io_enq_req_0_bits_ctrl_fuOpType; // @[CtrlBlock.scala 519:27]
  wire  lsqCtrl_io_enq_req_0_bits_ctrl_rfWen; // @[CtrlBlock.scala 519:27]
  wire  lsqCtrl_io_enq_req_0_bits_ctrl_fpWen; // @[CtrlBlock.scala 519:27]
  wire  lsqCtrl_io_enq_req_0_bits_ctrl_flushPipe; // @[CtrlBlock.scala 519:27]
  wire  lsqCtrl_io_enq_req_0_bits_ctrl_replayInst; // @[CtrlBlock.scala 519:27]
  wire [5:0] lsqCtrl_io_enq_req_0_bits_pdest; // @[CtrlBlock.scala 519:27]
  wire  lsqCtrl_io_enq_req_0_bits_robIdx_flag; // @[CtrlBlock.scala 519:27]
  wire [4:0] lsqCtrl_io_enq_req_0_bits_robIdx_value; // @[CtrlBlock.scala 519:27]
  wire  lsqCtrl_io_enq_req_1_valid; // @[CtrlBlock.scala 519:27]
  wire  lsqCtrl_io_enq_req_1_bits_cf_trigger_backendEn_0; // @[CtrlBlock.scala 519:27]
  wire  lsqCtrl_io_enq_req_1_bits_cf_trigger_backendEn_1; // @[CtrlBlock.scala 519:27]
  wire [6:0] lsqCtrl_io_enq_req_1_bits_ctrl_fuOpType; // @[CtrlBlock.scala 519:27]
  wire  lsqCtrl_io_enq_req_1_bits_ctrl_rfWen; // @[CtrlBlock.scala 519:27]
  wire  lsqCtrl_io_enq_req_1_bits_ctrl_fpWen; // @[CtrlBlock.scala 519:27]
  wire  lsqCtrl_io_enq_req_1_bits_ctrl_flushPipe; // @[CtrlBlock.scala 519:27]
  wire  lsqCtrl_io_enq_req_1_bits_ctrl_replayInst; // @[CtrlBlock.scala 519:27]
  wire [5:0] lsqCtrl_io_enq_req_1_bits_pdest; // @[CtrlBlock.scala 519:27]
  wire  lsqCtrl_io_enq_req_1_bits_robIdx_flag; // @[CtrlBlock.scala 519:27]
  wire [4:0] lsqCtrl_io_enq_req_1_bits_robIdx_value; // @[CtrlBlock.scala 519:27]
  wire  lsqCtrl_io_enq_req_2_valid; // @[CtrlBlock.scala 519:27]
  wire  lsqCtrl_io_enq_req_2_bits_cf_trigger_backendEn_0; // @[CtrlBlock.scala 519:27]
  wire  lsqCtrl_io_enq_req_2_bits_cf_trigger_backendEn_1; // @[CtrlBlock.scala 519:27]
  wire [6:0] lsqCtrl_io_enq_req_2_bits_ctrl_fuOpType; // @[CtrlBlock.scala 519:27]
  wire  lsqCtrl_io_enq_req_2_bits_ctrl_rfWen; // @[CtrlBlock.scala 519:27]
  wire  lsqCtrl_io_enq_req_2_bits_ctrl_fpWen; // @[CtrlBlock.scala 519:27]
  wire  lsqCtrl_io_enq_req_2_bits_ctrl_flushPipe; // @[CtrlBlock.scala 519:27]
  wire  lsqCtrl_io_enq_req_2_bits_ctrl_replayInst; // @[CtrlBlock.scala 519:27]
  wire [5:0] lsqCtrl_io_enq_req_2_bits_pdest; // @[CtrlBlock.scala 519:27]
  wire  lsqCtrl_io_enq_req_2_bits_robIdx_flag; // @[CtrlBlock.scala 519:27]
  wire [4:0] lsqCtrl_io_enq_req_2_bits_robIdx_value; // @[CtrlBlock.scala 519:27]
  wire  lsqCtrl_io_enq_req_3_valid; // @[CtrlBlock.scala 519:27]
  wire  lsqCtrl_io_enq_req_3_bits_cf_trigger_backendEn_0; // @[CtrlBlock.scala 519:27]
  wire  lsqCtrl_io_enq_req_3_bits_cf_trigger_backendEn_1; // @[CtrlBlock.scala 519:27]
  wire [6:0] lsqCtrl_io_enq_req_3_bits_ctrl_fuOpType; // @[CtrlBlock.scala 519:27]
  wire  lsqCtrl_io_enq_req_3_bits_ctrl_rfWen; // @[CtrlBlock.scala 519:27]
  wire  lsqCtrl_io_enq_req_3_bits_ctrl_fpWen; // @[CtrlBlock.scala 519:27]
  wire  lsqCtrl_io_enq_req_3_bits_ctrl_flushPipe; // @[CtrlBlock.scala 519:27]
  wire  lsqCtrl_io_enq_req_3_bits_ctrl_replayInst; // @[CtrlBlock.scala 519:27]
  wire [5:0] lsqCtrl_io_enq_req_3_bits_pdest; // @[CtrlBlock.scala 519:27]
  wire  lsqCtrl_io_enq_req_3_bits_robIdx_flag; // @[CtrlBlock.scala 519:27]
  wire [4:0] lsqCtrl_io_enq_req_3_bits_robIdx_value; // @[CtrlBlock.scala 519:27]
  wire  lsqCtrl_io_enq_resp_0_lqIdx_flag; // @[CtrlBlock.scala 519:27]
  wire [3:0] lsqCtrl_io_enq_resp_0_lqIdx_value; // @[CtrlBlock.scala 519:27]
  wire  lsqCtrl_io_enq_resp_0_sqIdx_flag; // @[CtrlBlock.scala 519:27]
  wire [3:0] lsqCtrl_io_enq_resp_0_sqIdx_value; // @[CtrlBlock.scala 519:27]
  wire  lsqCtrl_io_enq_resp_1_lqIdx_flag; // @[CtrlBlock.scala 519:27]
  wire [3:0] lsqCtrl_io_enq_resp_1_lqIdx_value; // @[CtrlBlock.scala 519:27]
  wire  lsqCtrl_io_enq_resp_1_sqIdx_flag; // @[CtrlBlock.scala 519:27]
  wire [3:0] lsqCtrl_io_enq_resp_1_sqIdx_value; // @[CtrlBlock.scala 519:27]
  wire  lsqCtrl_io_enq_resp_2_lqIdx_flag; // @[CtrlBlock.scala 519:27]
  wire [3:0] lsqCtrl_io_enq_resp_2_lqIdx_value; // @[CtrlBlock.scala 519:27]
  wire  lsqCtrl_io_enq_resp_2_sqIdx_flag; // @[CtrlBlock.scala 519:27]
  wire [3:0] lsqCtrl_io_enq_resp_2_sqIdx_value; // @[CtrlBlock.scala 519:27]
  wire  lsqCtrl_io_enq_resp_3_lqIdx_flag; // @[CtrlBlock.scala 519:27]
  wire [3:0] lsqCtrl_io_enq_resp_3_lqIdx_value; // @[CtrlBlock.scala 519:27]
  wire  lsqCtrl_io_enq_resp_3_sqIdx_flag; // @[CtrlBlock.scala 519:27]
  wire [3:0] lsqCtrl_io_enq_resp_3_sqIdx_value; // @[CtrlBlock.scala 519:27]
  wire [1:0] lsqCtrl_io_lcommit; // @[CtrlBlock.scala 519:27]
  wire [1:0] lsqCtrl_io_scommit; // @[CtrlBlock.scala 519:27]
  wire [4:0] lsqCtrl_io_lqCancelCnt; // @[CtrlBlock.scala 519:27]
  wire [3:0] lsqCtrl_io_sqCancelCnt; // @[CtrlBlock.scala 519:27]
  wire [1:0] lsqCtrl_io_enqLsq_needAlloc_0; // @[CtrlBlock.scala 519:27]
  wire [1:0] lsqCtrl_io_enqLsq_needAlloc_1; // @[CtrlBlock.scala 519:27]
  wire [1:0] lsqCtrl_io_enqLsq_needAlloc_2; // @[CtrlBlock.scala 519:27]
  wire [1:0] lsqCtrl_io_enqLsq_needAlloc_3; // @[CtrlBlock.scala 519:27]
  wire  lsqCtrl_io_enqLsq_req_0_valid; // @[CtrlBlock.scala 519:27]
  wire  lsqCtrl_io_enqLsq_req_0_bits_cf_trigger_backendEn_0; // @[CtrlBlock.scala 519:27]
  wire  lsqCtrl_io_enqLsq_req_0_bits_cf_trigger_backendEn_1; // @[CtrlBlock.scala 519:27]
  wire [6:0] lsqCtrl_io_enqLsq_req_0_bits_ctrl_fuOpType; // @[CtrlBlock.scala 519:27]
  wire  lsqCtrl_io_enqLsq_req_0_bits_ctrl_rfWen; // @[CtrlBlock.scala 519:27]
  wire  lsqCtrl_io_enqLsq_req_0_bits_ctrl_fpWen; // @[CtrlBlock.scala 519:27]
  wire  lsqCtrl_io_enqLsq_req_0_bits_ctrl_flushPipe; // @[CtrlBlock.scala 519:27]
  wire  lsqCtrl_io_enqLsq_req_0_bits_ctrl_replayInst; // @[CtrlBlock.scala 519:27]
  wire [5:0] lsqCtrl_io_enqLsq_req_0_bits_pdest; // @[CtrlBlock.scala 519:27]
  wire  lsqCtrl_io_enqLsq_req_0_bits_robIdx_flag; // @[CtrlBlock.scala 519:27]
  wire [4:0] lsqCtrl_io_enqLsq_req_0_bits_robIdx_value; // @[CtrlBlock.scala 519:27]
  wire [3:0] lsqCtrl_io_enqLsq_req_0_bits_lqIdx_value; // @[CtrlBlock.scala 519:27]
  wire [3:0] lsqCtrl_io_enqLsq_req_0_bits_sqIdx_value; // @[CtrlBlock.scala 519:27]
  wire  lsqCtrl_io_enqLsq_req_1_valid; // @[CtrlBlock.scala 519:27]
  wire  lsqCtrl_io_enqLsq_req_1_bits_cf_trigger_backendEn_0; // @[CtrlBlock.scala 519:27]
  wire  lsqCtrl_io_enqLsq_req_1_bits_cf_trigger_backendEn_1; // @[CtrlBlock.scala 519:27]
  wire [6:0] lsqCtrl_io_enqLsq_req_1_bits_ctrl_fuOpType; // @[CtrlBlock.scala 519:27]
  wire  lsqCtrl_io_enqLsq_req_1_bits_ctrl_rfWen; // @[CtrlBlock.scala 519:27]
  wire  lsqCtrl_io_enqLsq_req_1_bits_ctrl_fpWen; // @[CtrlBlock.scala 519:27]
  wire  lsqCtrl_io_enqLsq_req_1_bits_ctrl_flushPipe; // @[CtrlBlock.scala 519:27]
  wire  lsqCtrl_io_enqLsq_req_1_bits_ctrl_replayInst; // @[CtrlBlock.scala 519:27]
  wire [5:0] lsqCtrl_io_enqLsq_req_1_bits_pdest; // @[CtrlBlock.scala 519:27]
  wire  lsqCtrl_io_enqLsq_req_1_bits_robIdx_flag; // @[CtrlBlock.scala 519:27]
  wire [4:0] lsqCtrl_io_enqLsq_req_1_bits_robIdx_value; // @[CtrlBlock.scala 519:27]
  wire [3:0] lsqCtrl_io_enqLsq_req_1_bits_lqIdx_value; // @[CtrlBlock.scala 519:27]
  wire [3:0] lsqCtrl_io_enqLsq_req_1_bits_sqIdx_value; // @[CtrlBlock.scala 519:27]
  wire  lsqCtrl_io_enqLsq_req_2_valid; // @[CtrlBlock.scala 519:27]
  wire  lsqCtrl_io_enqLsq_req_2_bits_cf_trigger_backendEn_0; // @[CtrlBlock.scala 519:27]
  wire  lsqCtrl_io_enqLsq_req_2_bits_cf_trigger_backendEn_1; // @[CtrlBlock.scala 519:27]
  wire [6:0] lsqCtrl_io_enqLsq_req_2_bits_ctrl_fuOpType; // @[CtrlBlock.scala 519:27]
  wire  lsqCtrl_io_enqLsq_req_2_bits_ctrl_rfWen; // @[CtrlBlock.scala 519:27]
  wire  lsqCtrl_io_enqLsq_req_2_bits_ctrl_fpWen; // @[CtrlBlock.scala 519:27]
  wire  lsqCtrl_io_enqLsq_req_2_bits_ctrl_flushPipe; // @[CtrlBlock.scala 519:27]
  wire  lsqCtrl_io_enqLsq_req_2_bits_ctrl_replayInst; // @[CtrlBlock.scala 519:27]
  wire [5:0] lsqCtrl_io_enqLsq_req_2_bits_pdest; // @[CtrlBlock.scala 519:27]
  wire  lsqCtrl_io_enqLsq_req_2_bits_robIdx_flag; // @[CtrlBlock.scala 519:27]
  wire [4:0] lsqCtrl_io_enqLsq_req_2_bits_robIdx_value; // @[CtrlBlock.scala 519:27]
  wire [3:0] lsqCtrl_io_enqLsq_req_2_bits_lqIdx_value; // @[CtrlBlock.scala 519:27]
  wire [3:0] lsqCtrl_io_enqLsq_req_2_bits_sqIdx_value; // @[CtrlBlock.scala 519:27]
  wire  lsqCtrl_io_enqLsq_req_3_valid; // @[CtrlBlock.scala 519:27]
  wire  lsqCtrl_io_enqLsq_req_3_bits_cf_trigger_backendEn_0; // @[CtrlBlock.scala 519:27]
  wire  lsqCtrl_io_enqLsq_req_3_bits_cf_trigger_backendEn_1; // @[CtrlBlock.scala 519:27]
  wire [6:0] lsqCtrl_io_enqLsq_req_3_bits_ctrl_fuOpType; // @[CtrlBlock.scala 519:27]
  wire  lsqCtrl_io_enqLsq_req_3_bits_ctrl_rfWen; // @[CtrlBlock.scala 519:27]
  wire  lsqCtrl_io_enqLsq_req_3_bits_ctrl_fpWen; // @[CtrlBlock.scala 519:27]
  wire  lsqCtrl_io_enqLsq_req_3_bits_ctrl_flushPipe; // @[CtrlBlock.scala 519:27]
  wire  lsqCtrl_io_enqLsq_req_3_bits_ctrl_replayInst; // @[CtrlBlock.scala 519:27]
  wire [5:0] lsqCtrl_io_enqLsq_req_3_bits_pdest; // @[CtrlBlock.scala 519:27]
  wire  lsqCtrl_io_enqLsq_req_3_bits_robIdx_flag; // @[CtrlBlock.scala 519:27]
  wire [4:0] lsqCtrl_io_enqLsq_req_3_bits_robIdx_value; // @[CtrlBlock.scala 519:27]
  wire [3:0] lsqCtrl_io_enqLsq_req_3_bits_lqIdx_value; // @[CtrlBlock.scala 519:27]
  wire [3:0] lsqCtrl_io_enqLsq_req_3_bits_sqIdx_value; // @[CtrlBlock.scala 519:27]
  wire  io_cpu_halt_delay_clock; // @[Hold.scala 97:23]
  wire  io_cpu_halt_delay_io_in; // @[Hold.scala 97:23]
  wire  io_cpu_halt_delay_io_out; // @[Hold.scala 97:23]
  wire  pfevent_clock; // @[CtrlBlock.scala 585:23]
  wire  pfevent_reset; // @[CtrlBlock.scala 585:23]
  wire  pfevent_io_distribute_csr_wvalid; // @[CtrlBlock.scala 585:23]
  wire [11:0] pfevent_io_distribute_csr_waddr; // @[CtrlBlock.scala 585:23]
  wire [63:0] pfevent_io_distribute_csr_wdata; // @[CtrlBlock.scala 585:23]
  wire [63:0] pfevent_io_hpmevent_0; // @[CtrlBlock.scala 585:23]
  wire [63:0] pfevent_io_hpmevent_1; // @[CtrlBlock.scala 585:23]
  wire [63:0] pfevent_io_hpmevent_2; // @[CtrlBlock.scala 585:23]
  wire [63:0] pfevent_io_hpmevent_3; // @[CtrlBlock.scala 585:23]
  wire [63:0] pfevent_io_hpmevent_4; // @[CtrlBlock.scala 585:23]
  wire [63:0] pfevent_io_hpmevent_5; // @[CtrlBlock.scala 585:23]
  wire [63:0] pfevent_io_hpmevent_6; // @[CtrlBlock.scala 585:23]
  wire [63:0] pfevent_io_hpmevent_7; // @[CtrlBlock.scala 585:23]
  wire [63:0] pfevent_io_hpmevent_8; // @[CtrlBlock.scala 585:23]
  wire [63:0] pfevent_io_hpmevent_9; // @[CtrlBlock.scala 585:23]
  wire [63:0] pfevent_io_hpmevent_10; // @[CtrlBlock.scala 585:23]
  wire [63:0] pfevent_io_hpmevent_11; // @[CtrlBlock.scala 585:23]
  wire [63:0] pfevent_io_hpmevent_12; // @[CtrlBlock.scala 585:23]
  wire [63:0] pfevent_io_hpmevent_13; // @[CtrlBlock.scala 585:23]
  wire [63:0] pfevent_io_hpmevent_14; // @[CtrlBlock.scala 585:23]
  wire [63:0] pfevent_io_hpmevent_15; // @[CtrlBlock.scala 585:23]
  wire [63:0] pfevent_io_hpmevent_16; // @[CtrlBlock.scala 585:23]
  wire [63:0] pfevent_io_hpmevent_17; // @[CtrlBlock.scala 585:23]
  wire [63:0] pfevent_io_hpmevent_18; // @[CtrlBlock.scala 585:23]
  wire [63:0] pfevent_io_hpmevent_19; // @[CtrlBlock.scala 585:23]
  wire [63:0] pfevent_io_hpmevent_20; // @[CtrlBlock.scala 585:23]
  wire [63:0] pfevent_io_hpmevent_21; // @[CtrlBlock.scala 585:23]
  wire [63:0] pfevent_io_hpmevent_22; // @[CtrlBlock.scala 585:23]
  wire [63:0] pfevent_io_hpmevent_23; // @[CtrlBlock.scala 585:23]
  wire  hpm_clock; // @[PerfCounterUtils.scala 255:21]
  wire [63:0] hpm_io_hpm_event_0; // @[PerfCounterUtils.scala 255:21]
  wire [63:0] hpm_io_hpm_event_1; // @[PerfCounterUtils.scala 255:21]
  wire [63:0] hpm_io_hpm_event_2; // @[PerfCounterUtils.scala 255:21]
  wire [63:0] hpm_io_hpm_event_3; // @[PerfCounterUtils.scala 255:21]
  wire [63:0] hpm_io_hpm_event_4; // @[PerfCounterUtils.scala 255:21]
  wire [63:0] hpm_io_hpm_event_5; // @[PerfCounterUtils.scala 255:21]
  wire [63:0] hpm_io_hpm_event_6; // @[PerfCounterUtils.scala 255:21]
  wire [63:0] hpm_io_hpm_event_7; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_0_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_1_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_2_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_3_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_4_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_5_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_6_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_7_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_8_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_9_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_10_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_11_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_12_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_13_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_14_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_15_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_16_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_17_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_18_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_19_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_20_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_21_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_23_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_24_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_25_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_26_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_27_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_28_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_29_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_30_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_31_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_32_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_33_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_34_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_35_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_36_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_37_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_38_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_39_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_40_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_41_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_42_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_43_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_44_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_45_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_46_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_47_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_48_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_49_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_50_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_51_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_52_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_53_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_54_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_55_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_56_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_57_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_58_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_59_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_60_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_61_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_62_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_63_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_64_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_65_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_66_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_67_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_68_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_69_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_70_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_71_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_72_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_73_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_74_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_75_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_76_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_77_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_78_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_79_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_80_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_81_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_82_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_83_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_84_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_85_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_86_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_87_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_88_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_perf_0_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_perf_1_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_perf_2_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_perf_3_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_perf_4_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_perf_5_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_perf_6_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_perf_7_value; // @[PerfCounterUtils.scala 255:21]
  reg  pcMem_io_wen_0_REG; // @[CtrlBlock.scala 287:33]
  reg [2:0] pcMem_io_waddr_0_REG; // @[CtrlBlock.scala 288:33]
  reg [38:0] pcMem_io_wdata_0_REG_startAddr; // @[CtrlBlock.scala 289:33]
  reg [38:0] pcMem_io_wdata_0_REG_nextLineAddr; // @[CtrlBlock.scala 289:33]
  reg  pcMem_io_wdata_0_REG_isNextMask_0; // @[CtrlBlock.scala 289:33]
  reg  pcMem_io_wdata_0_REG_isNextMask_1; // @[CtrlBlock.scala 289:33]
  reg  pcMem_io_wdata_0_REG_isNextMask_2; // @[CtrlBlock.scala 289:33]
  reg  pcMem_io_wdata_0_REG_isNextMask_3; // @[CtrlBlock.scala 289:33]
  reg  pcMem_io_wdata_0_REG_isNextMask_4; // @[CtrlBlock.scala 289:33]
  reg  pcMem_io_wdata_0_REG_isNextMask_5; // @[CtrlBlock.scala 289:33]
  reg  pcMem_io_wdata_0_REG_isNextMask_6; // @[CtrlBlock.scala 289:33]
  reg  pcMem_io_wdata_0_REG_isNextMask_7; // @[CtrlBlock.scala 289:33]
  reg [2:0] flushPC_REG; // @[CtrlBlock.scala 292:50]
  wire  _GEN_1 = 3'h1 == flushPC_REG ? pcMem_io_rdata_7_isNextMask_1 : pcMem_io_rdata_7_isNextMask_0; // @[NewFtq.scala 91:{42,42}]
  wire  _GEN_2 = 3'h2 == flushPC_REG ? pcMem_io_rdata_7_isNextMask_2 : _GEN_1; // @[NewFtq.scala 91:{42,42}]
  wire  _GEN_3 = 3'h3 == flushPC_REG ? pcMem_io_rdata_7_isNextMask_3 : _GEN_2; // @[NewFtq.scala 91:{42,42}]
  wire  _GEN_4 = 3'h4 == flushPC_REG ? pcMem_io_rdata_7_isNextMask_4 : _GEN_3; // @[NewFtq.scala 91:{42,42}]
  wire  _GEN_5 = 3'h5 == flushPC_REG ? pcMem_io_rdata_7_isNextMask_5 : _GEN_4; // @[NewFtq.scala 91:{42,42}]
  wire  _GEN_6 = 3'h6 == flushPC_REG ? pcMem_io_rdata_7_isNextMask_6 : _GEN_5; // @[NewFtq.scala 91:{42,42}]
  wire  _GEN_7 = 3'h7 == flushPC_REG ? pcMem_io_rdata_7_isNextMask_7 : _GEN_6; // @[NewFtq.scala 91:{42,42}]
  wire [38:0] _flushPC_T_4 = _GEN_7 & pcMem_io_rdata_7_startAddr[4] ? pcMem_io_rdata_7_nextLineAddr :
    pcMem_io_rdata_7_startAddr; // @[NewFtq.scala 91:22]
  wire [3:0] _GEN_1435 = {{1'd0}, flushPC_REG}; // @[NewFtq.scala 92:29]
  wire [3:0] _flushPC_T_8 = pcMem_io_rdata_7_startAddr[4:1] + _GEN_1435; // @[NewFtq.scala 92:29]
  wire [37:0] flushPC_hi = {_flushPC_T_4[38:5],_flushPC_T_8}; // @[Cat.scala 31:58]
  wire [38:0] flushPC = {_flushPC_T_4[38:5],_flushPC_T_8,1'h0}; // @[Cat.scala 31:58]
  reg  flushRedirect_valid_REG; // @[CtrlBlock.scala 295:33]
  reg  flushRedirect_bits_rrobIdx_flag; // @[Reg.scala 16:16]
  reg [4:0] flushRedirect_bits_rrobIdx_value; // @[Reg.scala 16:16]
  reg  flushRedirect_bits_rftqIdx_flag; // @[Reg.scala 16:16]
  reg [2:0] flushRedirect_bits_rftqIdx_value; // @[Reg.scala 16:16]
  reg [2:0] flushRedirect_bits_rftqOffset; // @[Reg.scala 16:16]
  reg  flushRedirect_bits_rlevel; // @[Reg.scala 16:16]
  wire  stage2Redirect_valid = flushRedirect_valid_REG ? flushRedirect_valid_REG : redirectGen_io_stage2Redirect_valid; // @[CtrlBlock.scala 302:27]
  wire  stage2Redirect_bits_robIdx_flag = flushRedirect_valid_REG ? flushRedirect_bits_rrobIdx_flag :
    redirectGen_io_stage2Redirect_bits_robIdx_flag; // @[CtrlBlock.scala 302:27]
  wire [4:0] stage2Redirect_bits_robIdx_value = flushRedirect_valid_REG ? flushRedirect_bits_rrobIdx_value :
    redirectGen_io_stage2Redirect_bits_robIdx_value; // @[CtrlBlock.scala 302:27]
  wire  stage2Redirect_bits_level = flushRedirect_valid_REG ? flushRedirect_bits_rlevel :
    redirectGen_io_stage2Redirect_bits_level; // @[CtrlBlock.scala 302:27]
  reg  redirectForExu_next_valid_REG; // @[BitUtils.scala 28:28]
  reg  redirectForExu_next_bits_rrobIdx_flag; // @[Reg.scala 16:16]
  reg [4:0] redirectForExu_next_bits_rrobIdx_value; // @[Reg.scala 16:16]
  reg  redirectForExu_next_bits_rlevel; // @[Reg.scala 16:16]
  wire  exuRedirect_valid = io_exuRedirect_0_valid & io_exuRedirect_0_bits_redirectValid; // @[CtrlBlock.scala 307:25]
  wire [5:0] _exuRedirect_killedByOlder_flushItself_T_1 = {io_exuRedirect_0_bits_uop_robIdx_flag,
    io_exuRedirect_0_bits_uop_robIdx_value}; // @[CircularQueuePtr.scala 61:50]
  wire [5:0] _exuRedirect_killedByOlder_flushItself_T_2 = {stage2Redirect_bits_robIdx_flag,
    stage2Redirect_bits_robIdx_value}; // @[CircularQueuePtr.scala 61:70]
  wire  _exuRedirect_killedByOlder_flushItself_T_3 = _exuRedirect_killedByOlder_flushItself_T_1 ==
    _exuRedirect_killedByOlder_flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  exuRedirect_killedByOlder_flushItself = stage2Redirect_bits_level & _exuRedirect_killedByOlder_flushItself_T_3; // @[Rob.scala 122:51]
  wire  exuRedirect_killedByOlder_differentFlag = io_exuRedirect_0_bits_uop_robIdx_flag ^
    stage2Redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  exuRedirect_killedByOlder_compare = io_exuRedirect_0_bits_uop_robIdx_value > stage2Redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _exuRedirect_killedByOlder_T = exuRedirect_killedByOlder_differentFlag ^ exuRedirect_killedByOlder_compare; // @[CircularQueuePtr.scala 88:19]
  wire  _exuRedirect_killedByOlder_T_2 = stage2Redirect_valid & (exuRedirect_killedByOlder_flushItself |
    _exuRedirect_killedByOlder_T); // @[Rob.scala 123:20]
  wire [5:0] _exuRedirect_killedByOlder_flushItself_T_6 = {redirectForExu_next_bits_rrobIdx_flag,
    redirectForExu_next_bits_rrobIdx_value}; // @[CircularQueuePtr.scala 61:70]
  wire  _exuRedirect_killedByOlder_flushItself_T_7 = _exuRedirect_killedByOlder_flushItself_T_1 ==
    _exuRedirect_killedByOlder_flushItself_T_6; // @[CircularQueuePtr.scala 61:52]
  wire  exuRedirect_killedByOlder_flushItself_1 = redirectForExu_next_bits_rlevel &
    _exuRedirect_killedByOlder_flushItself_T_7; // @[Rob.scala 122:51]
  wire  exuRedirect_killedByOlder_differentFlag_1 = io_exuRedirect_0_bits_uop_robIdx_flag ^
    redirectForExu_next_bits_rrobIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  exuRedirect_killedByOlder_compare_1 = io_exuRedirect_0_bits_uop_robIdx_value >
    redirectForExu_next_bits_rrobIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _exuRedirect_killedByOlder_T_3 = exuRedirect_killedByOlder_differentFlag_1 ^ exuRedirect_killedByOlder_compare_1
    ; // @[CircularQueuePtr.scala 88:19]
  wire  _exuRedirect_killedByOlder_T_5 = redirectForExu_next_valid_REG & (exuRedirect_killedByOlder_flushItself_1 |
    _exuRedirect_killedByOlder_T_3); // @[Rob.scala 123:20]
  wire [1:0] _exuRedirect_killedByOlder_T_6 = {_exuRedirect_killedByOlder_T_5,_exuRedirect_killedByOlder_T_2}; // @[Rob.scala 126:90]
  wire  exuRedirect_killedByOlder = |_exuRedirect_killedByOlder_T_6; // @[Rob.scala 126:97]
  reg  exuRedirect_delayed_valid_REG; // @[CtrlBlock.scala 310:29]
  reg  exuRedirect_delayed_bits_ruop_cf_pd_isRVC; // @[Reg.scala 16:16]
  reg [1:0] exuRedirect_delayed_bits_ruop_cf_pd_brType; // @[Reg.scala 16:16]
  reg  exuRedirect_delayed_bits_ruop_cf_pd_isCall; // @[Reg.scala 16:16]
  reg  exuRedirect_delayed_bits_ruop_cf_pd_isRet; // @[Reg.scala 16:16]
  reg [19:0] exuRedirect_delayed_bits_ruop_ctrl_imm; // @[Reg.scala 16:16]
  reg  exuRedirect_delayed_bits_rredirect_robIdx_flag; // @[Reg.scala 16:16]
  reg [4:0] exuRedirect_delayed_bits_rredirect_robIdx_value; // @[Reg.scala 16:16]
  reg  exuRedirect_delayed_bits_rredirect_ftqIdx_flag; // @[Reg.scala 16:16]
  reg [2:0] exuRedirect_delayed_bits_rredirect_ftqIdx_value; // @[Reg.scala 16:16]
  reg [2:0] exuRedirect_delayed_bits_rredirect_ftqOffset; // @[Reg.scala 16:16]
  reg [38:0] exuRedirect_delayed_bits_rredirect_cfiUpdate_target; // @[Reg.scala 16:16]
  reg  exuRedirect_delayed_bits_rredirect_cfiUpdate_isMisPred; // @[Reg.scala 16:16]
  wire  exuRedirect_valid_1 = io_exuRedirect_1_valid & io_exuRedirect_1_bits_redirectValid; // @[CtrlBlock.scala 307:25]
  wire [5:0] _exuRedirect_killedByOlder_flushItself_T_9 = {io_exuRedirect_1_bits_uop_robIdx_flag,
    io_exuRedirect_1_bits_uop_robIdx_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _exuRedirect_killedByOlder_flushItself_T_11 = _exuRedirect_killedByOlder_flushItself_T_9 ==
    _exuRedirect_killedByOlder_flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  exuRedirect_killedByOlder_flushItself_2 = stage2Redirect_bits_level &
    _exuRedirect_killedByOlder_flushItself_T_11; // @[Rob.scala 122:51]
  wire  exuRedirect_killedByOlder_differentFlag_2 = io_exuRedirect_1_bits_uop_robIdx_flag ^
    stage2Redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  exuRedirect_killedByOlder_compare_2 = io_exuRedirect_1_bits_uop_robIdx_value > stage2Redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _exuRedirect_killedByOlder_T_7 = exuRedirect_killedByOlder_differentFlag_2 ^ exuRedirect_killedByOlder_compare_2
    ; // @[CircularQueuePtr.scala 88:19]
  wire  _exuRedirect_killedByOlder_T_9 = stage2Redirect_valid & (exuRedirect_killedByOlder_flushItself_2 |
    _exuRedirect_killedByOlder_T_7); // @[Rob.scala 123:20]
  wire  _exuRedirect_killedByOlder_flushItself_T_15 = _exuRedirect_killedByOlder_flushItself_T_9 ==
    _exuRedirect_killedByOlder_flushItself_T_6; // @[CircularQueuePtr.scala 61:52]
  wire  exuRedirect_killedByOlder_flushItself_3 = redirectForExu_next_bits_rlevel &
    _exuRedirect_killedByOlder_flushItself_T_15; // @[Rob.scala 122:51]
  wire  exuRedirect_killedByOlder_differentFlag_3 = io_exuRedirect_1_bits_uop_robIdx_flag ^
    redirectForExu_next_bits_rrobIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  exuRedirect_killedByOlder_compare_3 = io_exuRedirect_1_bits_uop_robIdx_value >
    redirectForExu_next_bits_rrobIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _exuRedirect_killedByOlder_T_10 = exuRedirect_killedByOlder_differentFlag_3 ^
    exuRedirect_killedByOlder_compare_3; // @[CircularQueuePtr.scala 88:19]
  wire  _exuRedirect_killedByOlder_T_12 = redirectForExu_next_valid_REG & (exuRedirect_killedByOlder_flushItself_3 |
    _exuRedirect_killedByOlder_T_10); // @[Rob.scala 123:20]
  wire [1:0] _exuRedirect_killedByOlder_T_13 = {_exuRedirect_killedByOlder_T_12,_exuRedirect_killedByOlder_T_9}; // @[Rob.scala 126:90]
  wire  exuRedirect_killedByOlder_1 = |_exuRedirect_killedByOlder_T_13; // @[Rob.scala 126:97]
  reg  exuRedirect_delayed_valid_REG_1; // @[CtrlBlock.scala 310:29]
  reg  exuRedirect_delayed_bits_r1_uop_cf_pd_isRVC; // @[Reg.scala 16:16]
  reg [1:0] exuRedirect_delayed_bits_r1_uop_cf_pd_brType; // @[Reg.scala 16:16]
  reg  exuRedirect_delayed_bits_r1_uop_cf_pd_isCall; // @[Reg.scala 16:16]
  reg  exuRedirect_delayed_bits_r1_uop_cf_pd_isRet; // @[Reg.scala 16:16]
  reg [19:0] exuRedirect_delayed_bits_r1_uop_ctrl_imm; // @[Reg.scala 16:16]
  reg  exuRedirect_delayed_bits_r1_redirect_robIdx_flag; // @[Reg.scala 16:16]
  reg [4:0] exuRedirect_delayed_bits_r1_redirect_robIdx_value; // @[Reg.scala 16:16]
  reg  exuRedirect_delayed_bits_r1_redirect_ftqIdx_flag; // @[Reg.scala 16:16]
  reg [2:0] exuRedirect_delayed_bits_r1_redirect_ftqIdx_value; // @[Reg.scala 16:16]
  reg [2:0] exuRedirect_delayed_bits_r1_redirect_ftqOffset; // @[Reg.scala 16:16]
  reg  exuRedirect_delayed_bits_r1_redirect_cfiUpdate_taken; // @[Reg.scala 16:16]
  reg  exuRedirect_delayed_bits_r1_redirect_cfiUpdate_isMisPred; // @[Reg.scala 16:16]
  wire  exuRedirect_valid_2 = io_exuRedirect_2_valid & io_exuRedirect_2_bits_redirectValid; // @[CtrlBlock.scala 307:25]
  wire [5:0] _exuRedirect_killedByOlder_flushItself_T_17 = {io_exuRedirect_2_bits_uop_robIdx_flag,
    io_exuRedirect_2_bits_uop_robIdx_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _exuRedirect_killedByOlder_flushItself_T_19 = _exuRedirect_killedByOlder_flushItself_T_17 ==
    _exuRedirect_killedByOlder_flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  exuRedirect_killedByOlder_flushItself_4 = stage2Redirect_bits_level &
    _exuRedirect_killedByOlder_flushItself_T_19; // @[Rob.scala 122:51]
  wire  exuRedirect_killedByOlder_differentFlag_4 = io_exuRedirect_2_bits_uop_robIdx_flag ^
    stage2Redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  exuRedirect_killedByOlder_compare_4 = io_exuRedirect_2_bits_uop_robIdx_value > stage2Redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _exuRedirect_killedByOlder_T_14 = exuRedirect_killedByOlder_differentFlag_4 ^
    exuRedirect_killedByOlder_compare_4; // @[CircularQueuePtr.scala 88:19]
  wire  _exuRedirect_killedByOlder_T_16 = stage2Redirect_valid & (exuRedirect_killedByOlder_flushItself_4 |
    _exuRedirect_killedByOlder_T_14); // @[Rob.scala 123:20]
  wire  _exuRedirect_killedByOlder_flushItself_T_23 = _exuRedirect_killedByOlder_flushItself_T_17 ==
    _exuRedirect_killedByOlder_flushItself_T_6; // @[CircularQueuePtr.scala 61:52]
  wire  exuRedirect_killedByOlder_flushItself_5 = redirectForExu_next_bits_rlevel &
    _exuRedirect_killedByOlder_flushItself_T_23; // @[Rob.scala 122:51]
  wire  exuRedirect_killedByOlder_differentFlag_5 = io_exuRedirect_2_bits_uop_robIdx_flag ^
    redirectForExu_next_bits_rrobIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  exuRedirect_killedByOlder_compare_5 = io_exuRedirect_2_bits_uop_robIdx_value >
    redirectForExu_next_bits_rrobIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _exuRedirect_killedByOlder_T_17 = exuRedirect_killedByOlder_differentFlag_5 ^
    exuRedirect_killedByOlder_compare_5; // @[CircularQueuePtr.scala 88:19]
  wire  _exuRedirect_killedByOlder_T_19 = redirectForExu_next_valid_REG & (exuRedirect_killedByOlder_flushItself_5 |
    _exuRedirect_killedByOlder_T_17); // @[Rob.scala 123:20]
  wire [1:0] _exuRedirect_killedByOlder_T_20 = {_exuRedirect_killedByOlder_T_19,_exuRedirect_killedByOlder_T_16}; // @[Rob.scala 126:90]
  wire  exuRedirect_killedByOlder_2 = |_exuRedirect_killedByOlder_T_20; // @[Rob.scala 126:97]
  reg  exuRedirect_delayed_valid_REG_2; // @[CtrlBlock.scala 310:29]
  reg  exuRedirect_delayed_bits_r2_uop_cf_pd_isRVC; // @[Reg.scala 16:16]
  reg [1:0] exuRedirect_delayed_bits_r2_uop_cf_pd_brType; // @[Reg.scala 16:16]
  reg  exuRedirect_delayed_bits_r2_uop_cf_pd_isCall; // @[Reg.scala 16:16]
  reg  exuRedirect_delayed_bits_r2_uop_cf_pd_isRet; // @[Reg.scala 16:16]
  reg [19:0] exuRedirect_delayed_bits_r2_uop_ctrl_imm; // @[Reg.scala 16:16]
  reg  exuRedirect_delayed_bits_r2_redirect_robIdx_flag; // @[Reg.scala 16:16]
  reg [4:0] exuRedirect_delayed_bits_r2_redirect_robIdx_value; // @[Reg.scala 16:16]
  reg  exuRedirect_delayed_bits_r2_redirect_ftqIdx_flag; // @[Reg.scala 16:16]
  reg [2:0] exuRedirect_delayed_bits_r2_redirect_ftqIdx_value; // @[Reg.scala 16:16]
  reg [2:0] exuRedirect_delayed_bits_r2_redirect_ftqOffset; // @[Reg.scala 16:16]
  reg  exuRedirect_delayed_bits_r2_redirect_cfiUpdate_taken; // @[Reg.scala 16:16]
  reg  exuRedirect_delayed_bits_r2_redirect_cfiUpdate_isMisPred; // @[Reg.scala 16:16]
  wire [5:0] _loadReplay_valid_flushItself_T_1 = {io_memoryViolation_bits_robIdx_flag,
    io_memoryViolation_bits_robIdx_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _loadReplay_valid_flushItself_T_3 = _loadReplay_valid_flushItself_T_1 ==
    _exuRedirect_killedByOlder_flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  loadReplay_valid_flushItself = stage2Redirect_bits_level & _loadReplay_valid_flushItself_T_3; // @[Rob.scala 122:51]
  wire  loadReplay_valid_differentFlag = io_memoryViolation_bits_robIdx_flag ^ stage2Redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  loadReplay_valid_compare = io_memoryViolation_bits_robIdx_value > stage2Redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _loadReplay_valid_T = loadReplay_valid_differentFlag ^ loadReplay_valid_compare; // @[CircularQueuePtr.scala 88:19]
  wire  _loadReplay_valid_T_2 = stage2Redirect_valid & (loadReplay_valid_flushItself | _loadReplay_valid_T); // @[Rob.scala 123:20]
  wire  _loadReplay_valid_flushItself_T_7 = _loadReplay_valid_flushItself_T_1 ==
    _exuRedirect_killedByOlder_flushItself_T_6; // @[CircularQueuePtr.scala 61:52]
  wire  loadReplay_valid_flushItself_1 = redirectForExu_next_bits_rlevel & _loadReplay_valid_flushItself_T_7; // @[Rob.scala 122:51]
  wire  loadReplay_valid_differentFlag_1 = io_memoryViolation_bits_robIdx_flag ^ redirectForExu_next_bits_rrobIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  loadReplay_valid_compare_1 = io_memoryViolation_bits_robIdx_value > redirectForExu_next_bits_rrobIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _loadReplay_valid_T_3 = loadReplay_valid_differentFlag_1 ^ loadReplay_valid_compare_1; // @[CircularQueuePtr.scala 88:19]
  wire  _loadReplay_valid_T_5 = redirectForExu_next_valid_REG & (loadReplay_valid_flushItself_1 | _loadReplay_valid_T_3)
    ; // @[Rob.scala 123:20]
  wire [1:0] _loadReplay_valid_T_6 = {_loadReplay_valid_T_5,_loadReplay_valid_T_2}; // @[Rob.scala 126:90]
  wire  _loadReplay_valid_T_7 = |_loadReplay_valid_T_6; // @[Rob.scala 126:97]
  wire  _loadReplay_valid_T_8 = ~_loadReplay_valid_T_7; // @[CtrlBlock.scala 316:5]
  reg  loadReplay_valid_REG; // @[CtrlBlock.scala 315:30]
  reg  loadReplay_bits_rrobIdx_flag; // @[Reg.scala 16:16]
  reg [4:0] loadReplay_bits_rrobIdx_value; // @[Reg.scala 16:16]
  reg  loadReplay_bits_rftqIdx_flag; // @[Reg.scala 16:16]
  reg [2:0] loadReplay_bits_rftqIdx_value; // @[Reg.scala 16:16]
  reg [2:0] loadReplay_bits_rftqOffset; // @[Reg.scala 16:16]
  reg [2:0] loadReplay_bits_rstFtqIdx_value; // @[Reg.scala 16:16]
  reg [2:0] loadReplay_bits_rstFtqOffset; // @[Reg.scala 16:16]
  reg [2:0] redirectGen_io_redirectPcRead_data_REG; // @[CtrlBlock.scala 321:72]
  wire  _GEN_879 = 3'h1 == redirectGen_io_redirectPcRead_data_REG ? pcMem_io_rdata_2_isNextMask_1 :
    pcMem_io_rdata_2_isNextMask_0; // @[NewFtq.scala 91:{42,42}]
  wire  _GEN_880 = 3'h2 == redirectGen_io_redirectPcRead_data_REG ? pcMem_io_rdata_2_isNextMask_2 : _GEN_879; // @[NewFtq.scala 91:{42,42}]
  wire  _GEN_881 = 3'h3 == redirectGen_io_redirectPcRead_data_REG ? pcMem_io_rdata_2_isNextMask_3 : _GEN_880; // @[NewFtq.scala 91:{42,42}]
  wire  _GEN_882 = 3'h4 == redirectGen_io_redirectPcRead_data_REG ? pcMem_io_rdata_2_isNextMask_4 : _GEN_881; // @[NewFtq.scala 91:{42,42}]
  wire  _GEN_883 = 3'h5 == redirectGen_io_redirectPcRead_data_REG ? pcMem_io_rdata_2_isNextMask_5 : _GEN_882; // @[NewFtq.scala 91:{42,42}]
  wire  _GEN_884 = 3'h6 == redirectGen_io_redirectPcRead_data_REG ? pcMem_io_rdata_2_isNextMask_6 : _GEN_883; // @[NewFtq.scala 91:{42,42}]
  wire  _GEN_885 = 3'h7 == redirectGen_io_redirectPcRead_data_REG ? pcMem_io_rdata_2_isNextMask_7 : _GEN_884; // @[NewFtq.scala 91:{42,42}]
  wire [38:0] _redirectGen_io_redirectPcRead_data_T_4 = _GEN_885 & pcMem_io_rdata_2_startAddr[4] ?
    pcMem_io_rdata_2_nextLineAddr : pcMem_io_rdata_2_startAddr; // @[NewFtq.scala 91:22]
  wire [3:0] _GEN_1436 = {{1'd0}, redirectGen_io_redirectPcRead_data_REG}; // @[NewFtq.scala 92:29]
  wire [3:0] _redirectGen_io_redirectPcRead_data_T_8 = pcMem_io_rdata_2_startAddr[4:1] + _GEN_1436; // @[NewFtq.scala 92:29]
  wire [37:0] redirectGen_io_redirectPcRead_data_hi = {_redirectGen_io_redirectPcRead_data_T_4[38:5],
    _redirectGen_io_redirectPcRead_data_T_8}; // @[Cat.scala 31:58]
  reg [2:0] redirectGen_io_memPredPcRead_data_REG; // @[CtrlBlock.scala 323:71]
  wire  _GEN_887 = 3'h1 == redirectGen_io_memPredPcRead_data_REG ? pcMem_io_rdata_3_isNextMask_1 :
    pcMem_io_rdata_3_isNextMask_0; // @[NewFtq.scala 91:{42,42}]
  wire  _GEN_888 = 3'h2 == redirectGen_io_memPredPcRead_data_REG ? pcMem_io_rdata_3_isNextMask_2 : _GEN_887; // @[NewFtq.scala 91:{42,42}]
  wire  _GEN_889 = 3'h3 == redirectGen_io_memPredPcRead_data_REG ? pcMem_io_rdata_3_isNextMask_3 : _GEN_888; // @[NewFtq.scala 91:{42,42}]
  wire  _GEN_890 = 3'h4 == redirectGen_io_memPredPcRead_data_REG ? pcMem_io_rdata_3_isNextMask_4 : _GEN_889; // @[NewFtq.scala 91:{42,42}]
  wire  _GEN_891 = 3'h5 == redirectGen_io_memPredPcRead_data_REG ? pcMem_io_rdata_3_isNextMask_5 : _GEN_890; // @[NewFtq.scala 91:{42,42}]
  wire  _GEN_892 = 3'h6 == redirectGen_io_memPredPcRead_data_REG ? pcMem_io_rdata_3_isNextMask_6 : _GEN_891; // @[NewFtq.scala 91:{42,42}]
  wire  _GEN_893 = 3'h7 == redirectGen_io_memPredPcRead_data_REG ? pcMem_io_rdata_3_isNextMask_7 : _GEN_892; // @[NewFtq.scala 91:{42,42}]
  wire [38:0] _redirectGen_io_memPredPcRead_data_T_4 = _GEN_893 & pcMem_io_rdata_3_startAddr[4] ?
    pcMem_io_rdata_3_nextLineAddr : pcMem_io_rdata_3_startAddr; // @[NewFtq.scala 91:22]
  wire [3:0] _GEN_1437 = {{1'd0}, redirectGen_io_memPredPcRead_data_REG}; // @[NewFtq.scala 92:29]
  wire [3:0] _redirectGen_io_memPredPcRead_data_T_8 = pcMem_io_rdata_3_startAddr[4:1] + _GEN_1437; // @[NewFtq.scala 92:29]
  wire [37:0] redirectGen_io_memPredPcRead_data_hi = {_redirectGen_io_memPredPcRead_data_T_4[38:5],
    _redirectGen_io_memPredPcRead_data_T_8}; // @[Cat.scala 31:58]
  reg  frontendFlushBits_ftqIdx_flag; // @[Reg.scala 16:16]
  reg [2:0] frontendFlushBits_ftqIdx_value; // @[Reg.scala 16:16]
  reg [2:0] frontendFlushBits_ftqOffset; // @[Reg.scala 16:16]
  reg  frontendFlushBits_level; // @[Reg.scala 16:16]
  wire  is_commit = rob_io_commits_commitValid_0 & rob_io_commits_isCommit & ~rob_io_flushOut_valid; // @[CtrlBlock.scala 337:78]
  reg  io_frontend_toFtq_rob_commits_0_valid_REG; // @[CtrlBlock.scala 338:54]
  reg [2:0] io_frontend_toFtq_rob_commits_0_bits_rcommitType; // @[Reg.scala 16:16]
  reg  io_frontend_toFtq_rob_commits_0_bits_rftqIdx_flag; // @[Reg.scala 16:16]
  reg [2:0] io_frontend_toFtq_rob_commits_0_bits_rftqIdx_value; // @[Reg.scala 16:16]
  reg [2:0] io_frontend_toFtq_rob_commits_0_bits_rftqOffset; // @[Reg.scala 16:16]
  wire  is_commit_1 = rob_io_commits_commitValid_1 & rob_io_commits_isCommit & ~rob_io_flushOut_valid; // @[CtrlBlock.scala 337:78]
  reg  io_frontend_toFtq_rob_commits_1_valid_REG; // @[CtrlBlock.scala 338:54]
  reg [2:0] io_frontend_toFtq_rob_commits_1_bits_rcommitType; // @[Reg.scala 16:16]
  reg  io_frontend_toFtq_rob_commits_1_bits_rftqIdx_flag; // @[Reg.scala 16:16]
  reg [2:0] io_frontend_toFtq_rob_commits_1_bits_rftqIdx_value; // @[Reg.scala 16:16]
  reg [2:0] io_frontend_toFtq_rob_commits_1_bits_rftqOffset; // @[Reg.scala 16:16]
  wire  _io_frontend_toFtq_redirect_bits_T_level = frontendFlushValid_delay_io_out ? frontendFlushBits_level :
    redirectGen_io_stage2Redirect_bits_level; // @[CtrlBlock.scala 342:41]
  wire [38:0] _io_frontend_toFtq_redirect_bits_T_cfiUpdate_target = frontendFlushValid_delay_io_out ? 39'h0 :
    redirectGen_io_stage2Redirect_bits_cfiUpdate_target; // @[CtrlBlock.scala 342:41]
  wire  pc_from_csr = io_robio_toCSR_isXRet | pc_from_csr_delay_io_out; // @[CtrlBlock.scala 350:43]
  wire [38:0] _rob_flush_pc_T_2 = flushPC + 39'h4; // @[CtrlBlock.scala 353:13]
  reg [38:0] rob_flush_pc; // @[Reg.scala 16:16]
  reg [38:0] io_frontend_toFtq_redirect_bits_cfiUpdate_target_REG; // @[CtrlBlock.scala 358:64]
  reg  pendingRedirect; // @[CtrlBlock.scala 362:32]
  reg  REG; // @[CtrlBlock.scala 365:22]
  wire  _GEN_996 = REG ? 1'h0 : pendingRedirect; // @[CtrlBlock.scala 365:58 366:21 362:32]
  reg  decode_io_csrCtrl_REG_fusion_enable; // @[CtrlBlock.scala 403:31]
  reg  decode_io_csrCtrl_REG_wfi_enable; // @[CtrlBlock.scala 403:31]
  reg  decode_io_csrCtrl_REG_svinval_enable; // @[CtrlBlock.scala 403:31]
  reg  decode_io_csrCtrl_REG_singlestep; // @[CtrlBlock.scala 403:31]
  wire  _mdp_foldpc_T = decode_io_out_0_ready & decode_io_out_0_valid; // @[Decoupled.scala 50:35]
  wire  _mdp_foldpc_T_1 = decode_io_out_1_ready & decode_io_out_1_valid; // @[Decoupled.scala 50:35]
  reg  ssit_io_update_REG_valid; // @[CtrlBlock.scala 419:28]
  reg [9:0] ssit_io_update_REG_ldpc; // @[CtrlBlock.scala 419:28]
  reg [9:0] ssit_io_update_REG_stpc; // @[CtrlBlock.scala 419:28]
  reg [4:0] ssit_io_csrCtrl_REG_lvpred_timeout; // @[CtrlBlock.scala 420:29]
  reg  lfst_io_redirect_REG_valid; // @[CtrlBlock.scala 426:30]
  reg  lfst_io_redirect_REG_bits_robIdx_flag; // @[CtrlBlock.scala 426:30]
  reg [4:0] lfst_io_redirect_REG_bits_robIdx_value; // @[CtrlBlock.scala 426:30]
  reg  lfst_io_redirect_REG_bits_level; // @[CtrlBlock.scala 426:30]
  reg  REG_1_0_valid; // @[CtrlBlock.scala 427:32]
  reg  REG_1_0_bits_uop_cf_storeSetHit; // @[CtrlBlock.scala 427:32]
  reg [4:0] REG_1_0_bits_uop_cf_ssid; // @[CtrlBlock.scala 427:32]
  reg [4:0] REG_1_0_bits_uop_robIdx_value; // @[CtrlBlock.scala 427:32]
  reg  REG_1_1_valid; // @[CtrlBlock.scala 427:32]
  reg  REG_1_1_bits_uop_cf_storeSetHit; // @[CtrlBlock.scala 427:32]
  reg [4:0] REG_1_1_bits_uop_cf_ssid; // @[CtrlBlock.scala 427:32]
  reg [4:0] REG_1_1_bits_uop_robIdx_value; // @[CtrlBlock.scala 427:32]
  reg  lfst_io_csrCtrl_REG_lvpred_disable; // @[CtrlBlock.scala 428:29]
  reg  lfst_io_csrCtrl_REG_no_spec_load; // @[CtrlBlock.scala 428:29]
  reg  lfst_io_csrCtrl_REG_storeset_wait_store; // @[CtrlBlock.scala 428:29]
  wire  decodeHasException = io_frontend_cfVec_0_bits_exceptionVec_12 | io_frontend_cfVec_0_bits_exceptionVec_1; // @[CtrlBlock.scala 441:85]
  wire  disableFusion = decode_io_csrCtrl_singlestep | ~decode_io_csrCtrl_fusion_enable; // @[CtrlBlock.scala 442:54]
  wire  _renamePipe_T = stage2Redirect_valid | pendingRedirect; // @[CtrlBlock.scala 451:28]
  reg  renamePipe_valid; // @[PipelineConnect.scala 108:24]
  wire  renamePipe__ready = rename_io_in_0_ready; // @[PipelineConnect.scala 182:21 CtrlBlock.scala 452:22]
  wire  renamePipe_leftFire = decode_io_out_0_valid & renamePipe__ready; // @[PipelineConnect.scala 109:31]
  wire  _GEN_998 = rename_io_in_0_ready ? 1'h0 : renamePipe_valid; // @[PipelineConnect.scala 108:24 110:{25,33}]
  wire  _GEN_999 = renamePipe_leftFire | _GEN_998; // @[PipelineConnect.scala 111:{21,29}]
  reg [9:0] renamePipe_data_cf_foldpc; // @[Reg.scala 16:16]
  reg  renamePipe_data_cf_exceptionVec_1; // @[Reg.scala 16:16]
  reg  renamePipe_data_cf_exceptionVec_2; // @[Reg.scala 16:16]
  reg  renamePipe_data_cf_exceptionVec_12; // @[Reg.scala 16:16]
  reg  renamePipe_data_cf_trigger_frontendHit_0; // @[Reg.scala 16:16]
  reg  renamePipe_data_cf_trigger_frontendHit_1; // @[Reg.scala 16:16]
  reg  renamePipe_data_cf_trigger_frontendHit_2; // @[Reg.scala 16:16]
  reg  renamePipe_data_cf_trigger_frontendHit_3; // @[Reg.scala 16:16]
  reg  renamePipe_data_cf_trigger_backendEn_0; // @[Reg.scala 16:16]
  reg  renamePipe_data_cf_trigger_backendEn_1; // @[Reg.scala 16:16]
  reg  renamePipe_data_cf_pd_isRVC; // @[Reg.scala 16:16]
  reg [1:0] renamePipe_data_cf_pd_brType; // @[Reg.scala 16:16]
  reg  renamePipe_data_cf_pd_isCall; // @[Reg.scala 16:16]
  reg  renamePipe_data_cf_pd_isRet; // @[Reg.scala 16:16]
  reg  renamePipe_data_cf_pred_taken; // @[Reg.scala 16:16]
  reg  renamePipe_data_cf_crossPageIPFFix; // @[Reg.scala 16:16]
  reg  renamePipe_data_cf_ftqPtr_flag; // @[Reg.scala 16:16]
  reg [2:0] renamePipe_data_cf_ftqPtr_value; // @[Reg.scala 16:16]
  reg [2:0] renamePipe_data_cf_ftqOffset; // @[Reg.scala 16:16]
  reg [1:0] renamePipe_data_ctrl_srcType_0; // @[Reg.scala 16:16]
  reg [1:0] renamePipe_data_ctrl_srcType_1; // @[Reg.scala 16:16]
  reg [1:0] renamePipe_data_ctrl_srcType_2; // @[Reg.scala 16:16]
  reg [4:0] renamePipe_data_ctrl_lsrc_0; // @[Reg.scala 16:16]
  reg [4:0] renamePipe_data_ctrl_lsrc_1; // @[Reg.scala 16:16]
  reg [4:0] renamePipe_data_ctrl_ldest; // @[Reg.scala 16:16]
  reg [3:0] renamePipe_data_ctrl_fuType; // @[Reg.scala 16:16]
  reg [6:0] renamePipe_data_ctrl_fuOpType; // @[Reg.scala 16:16]
  reg  renamePipe_data_ctrl_rfWen; // @[Reg.scala 16:16]
  reg  renamePipe_data_ctrl_fpWen; // @[Reg.scala 16:16]
  reg  renamePipe_data_ctrl_isXSTrap; // @[Reg.scala 16:16]
  reg  renamePipe_data_ctrl_noSpecExec; // @[Reg.scala 16:16]
  reg  renamePipe_data_ctrl_blockBackward; // @[Reg.scala 16:16]
  reg  renamePipe_data_ctrl_flushPipe; // @[Reg.scala 16:16]
  reg [3:0] renamePipe_data_ctrl_selImm; // @[Reg.scala 16:16]
  reg [19:0] renamePipe_data_ctrl_imm; // @[Reg.scala 16:16]
  reg  renamePipe_data_ctrl_fpu_isAddSub; // @[Reg.scala 16:16]
  reg  renamePipe_data_ctrl_fpu_typeTagIn; // @[Reg.scala 16:16]
  reg  renamePipe_data_ctrl_fpu_typeTagOut; // @[Reg.scala 16:16]
  reg  renamePipe_data_ctrl_fpu_fromInt; // @[Reg.scala 16:16]
  reg  renamePipe_data_ctrl_fpu_wflags; // @[Reg.scala 16:16]
  reg  renamePipe_data_ctrl_fpu_fpWen; // @[Reg.scala 16:16]
  reg [1:0] renamePipe_data_ctrl_fpu_fmaCmd; // @[Reg.scala 16:16]
  reg  renamePipe_data_ctrl_fpu_div; // @[Reg.scala 16:16]
  reg  renamePipe_data_ctrl_fpu_sqrt; // @[Reg.scala 16:16]
  reg  renamePipe_data_ctrl_fpu_fcvt; // @[Reg.scala 16:16]
  reg [1:0] renamePipe_data_ctrl_fpu_typ; // @[Reg.scala 16:16]
  reg [1:0] renamePipe_data_ctrl_fpu_fmt; // @[Reg.scala 16:16]
  reg  renamePipe_data_ctrl_fpu_ren3; // @[Reg.scala 16:16]
  reg [2:0] renamePipe_data_ctrl_fpu_rm; // @[Reg.scala 16:16]
  reg  renamePipe_data_ctrl_isMove; // @[Reg.scala 16:16]
  wire  _decode_io_fusion_0_T = rename_io_out_0_ready & rename_io_out_0_valid; // @[Decoupled.scala 50:35]
  wire [3:0] _GEN_1085 = fusionDecoder_io_out_0_bits_fuType_valid ? 4'h4 : renamePipe_data_ctrl_fuType; // @[FusionDecoder.scala 475:25 476:17 CtrlBlock.scala 454:26]
  wire [6:0] _GEN_1086 = fusionDecoder_io_out_0_bits_fuOpType_valid ? fusionDecoder_io_out_0_bits_fuOpType_bits :
    renamePipe_data_ctrl_fuOpType; // @[FusionDecoder.scala 478:27 479:19 CtrlBlock.scala 454:26]
  wire [4:0] _GEN_1087 = fusionDecoder_io_out_0_bits_lsrc2_valid ? fusionDecoder_io_out_0_bits_lsrc2_bits :
    renamePipe_data_ctrl_lsrc_1; // @[FusionDecoder.scala 481:24 482:18 CtrlBlock.scala 454:26]
  wire [1:0] _GEN_1088 = fusionDecoder_io_out_0_bits_src2Type_valid ? 2'h0 : renamePipe_data_ctrl_srcType_1; // @[FusionDecoder.scala 484:27 485:21 CtrlBlock.scala 454:26]
  wire  sameFtqPtr = rename_io_in_0_bits_cf_ftqPtr_value == rename_io_in_1_bits_cf_ftqPtr_value; // @[CtrlBlock.scala 469:63]
  wire [2:0] ftqOffsetDiff = rename_io_in_1_bits_cf_ftqOffset - rename_io_in_0_bits_cf_ftqOffset; // @[CtrlBlock.scala 472:40]
  wire  cond1 = sameFtqPtr & ftqOffsetDiff == 3'h1; // @[CtrlBlock.scala 473:32]
  wire  cond2 = sameFtqPtr & ftqOffsetDiff == 3'h2; // @[CtrlBlock.scala 474:32]
  wire  cond3 = ~sameFtqPtr & rename_io_in_1_bits_cf_ftqOffset == 3'h0; // @[CtrlBlock.scala 475:33]
  wire [2:0] _rename_io_in_0_bits_ctrl_commitType_T = cond3 ? 3'h6 : 3'h7; // @[CtrlBlock.scala 477:84]
  wire [2:0] _rename_io_in_0_bits_ctrl_commitType_T_1 = cond2 ? 3'h5 : _rename_io_in_0_bits_ctrl_commitType_T; // @[CtrlBlock.scala 477:68]
  wire [2:0] _rename_io_in_0_bits_ctrl_commitType_T_2 = cond1 ? 3'h4 : _rename_io_in_0_bits_ctrl_commitType_T_1; // @[CtrlBlock.scala 477:52]
  wire  decodeHasException_1 = io_frontend_cfVec_1_bits_exceptionVec_12 | io_frontend_cfVec_1_bits_exceptionVec_1; // @[CtrlBlock.scala 441:85]
  reg  renamePipe_valid_1; // @[PipelineConnect.scala 108:24]
  wire  renamePipe_1_ready = rename_io_in_1_ready; // @[PipelineConnect.scala 182:21 CtrlBlock.scala 452:22]
  wire  renamePipe_leftFire_1 = decode_io_out_1_valid & renamePipe_1_ready; // @[PipelineConnect.scala 109:31]
  wire  _GEN_1094 = rename_io_in_1_ready ? 1'h0 : renamePipe_valid_1; // @[PipelineConnect.scala 108:24 110:{25,33}]
  wire  _GEN_1095 = renamePipe_leftFire_1 | _GEN_1094; // @[PipelineConnect.scala 111:{21,29}]
  reg [9:0] renamePipe_data_1_cf_foldpc; // @[Reg.scala 16:16]
  reg  renamePipe_data_1_cf_exceptionVec_1; // @[Reg.scala 16:16]
  reg  renamePipe_data_1_cf_exceptionVec_2; // @[Reg.scala 16:16]
  reg  renamePipe_data_1_cf_exceptionVec_12; // @[Reg.scala 16:16]
  reg  renamePipe_data_1_cf_trigger_frontendHit_0; // @[Reg.scala 16:16]
  reg  renamePipe_data_1_cf_trigger_frontendHit_1; // @[Reg.scala 16:16]
  reg  renamePipe_data_1_cf_trigger_frontendHit_2; // @[Reg.scala 16:16]
  reg  renamePipe_data_1_cf_trigger_frontendHit_3; // @[Reg.scala 16:16]
  reg  renamePipe_data_1_cf_trigger_backendEn_0; // @[Reg.scala 16:16]
  reg  renamePipe_data_1_cf_trigger_backendEn_1; // @[Reg.scala 16:16]
  reg  renamePipe_data_1_cf_pd_isRVC; // @[Reg.scala 16:16]
  reg [1:0] renamePipe_data_1_cf_pd_brType; // @[Reg.scala 16:16]
  reg  renamePipe_data_1_cf_pd_isCall; // @[Reg.scala 16:16]
  reg  renamePipe_data_1_cf_pd_isRet; // @[Reg.scala 16:16]
  reg  renamePipe_data_1_cf_pred_taken; // @[Reg.scala 16:16]
  reg  renamePipe_data_1_cf_crossPageIPFFix; // @[Reg.scala 16:16]
  reg  renamePipe_data_1_cf_ftqPtr_flag; // @[Reg.scala 16:16]
  reg [2:0] renamePipe_data_1_cf_ftqPtr_value; // @[Reg.scala 16:16]
  reg [2:0] renamePipe_data_1_cf_ftqOffset; // @[Reg.scala 16:16]
  reg [1:0] renamePipe_data_1_ctrl_srcType_0; // @[Reg.scala 16:16]
  reg [1:0] renamePipe_data_1_ctrl_srcType_1; // @[Reg.scala 16:16]
  reg [1:0] renamePipe_data_1_ctrl_srcType_2; // @[Reg.scala 16:16]
  reg [4:0] renamePipe_data_1_ctrl_lsrc_0; // @[Reg.scala 16:16]
  reg [4:0] renamePipe_data_1_ctrl_lsrc_1; // @[Reg.scala 16:16]
  reg [4:0] renamePipe_data_1_ctrl_lsrc_2; // @[Reg.scala 16:16]
  reg [4:0] renamePipe_data_1_ctrl_ldest; // @[Reg.scala 16:16]
  reg [3:0] renamePipe_data_1_ctrl_fuType; // @[Reg.scala 16:16]
  reg [6:0] renamePipe_data_1_ctrl_fuOpType; // @[Reg.scala 16:16]
  reg  renamePipe_data_1_ctrl_rfWen; // @[Reg.scala 16:16]
  reg  renamePipe_data_1_ctrl_fpWen; // @[Reg.scala 16:16]
  reg  renamePipe_data_1_ctrl_isXSTrap; // @[Reg.scala 16:16]
  reg  renamePipe_data_1_ctrl_noSpecExec; // @[Reg.scala 16:16]
  reg  renamePipe_data_1_ctrl_blockBackward; // @[Reg.scala 16:16]
  reg  renamePipe_data_1_ctrl_flushPipe; // @[Reg.scala 16:16]
  reg [3:0] renamePipe_data_1_ctrl_selImm; // @[Reg.scala 16:16]
  reg [19:0] renamePipe_data_1_ctrl_imm; // @[Reg.scala 16:16]
  reg  renamePipe_data_1_ctrl_fpu_isAddSub; // @[Reg.scala 16:16]
  reg  renamePipe_data_1_ctrl_fpu_typeTagIn; // @[Reg.scala 16:16]
  reg  renamePipe_data_1_ctrl_fpu_typeTagOut; // @[Reg.scala 16:16]
  reg  renamePipe_data_1_ctrl_fpu_fromInt; // @[Reg.scala 16:16]
  reg  renamePipe_data_1_ctrl_fpu_wflags; // @[Reg.scala 16:16]
  reg  renamePipe_data_1_ctrl_fpu_fpWen; // @[Reg.scala 16:16]
  reg [1:0] renamePipe_data_1_ctrl_fpu_fmaCmd; // @[Reg.scala 16:16]
  reg  renamePipe_data_1_ctrl_fpu_div; // @[Reg.scala 16:16]
  reg  renamePipe_data_1_ctrl_fpu_sqrt; // @[Reg.scala 16:16]
  reg  renamePipe_data_1_ctrl_fpu_fcvt; // @[Reg.scala 16:16]
  reg [1:0] renamePipe_data_1_ctrl_fpu_typ; // @[Reg.scala 16:16]
  reg [1:0] renamePipe_data_1_ctrl_fpu_fmt; // @[Reg.scala 16:16]
  reg  renamePipe_data_1_ctrl_fpu_ren3; // @[Reg.scala 16:16]
  reg [2:0] renamePipe_data_1_ctrl_fpu_rm; // @[Reg.scala 16:16]
  reg  renamePipe_data_1_ctrl_isMove; // @[Reg.scala 16:16]
  reg  valid; // @[PipelineConnect.scala 108:24]
  wire  leftFire = rename_io_out_0_valid & dispatch_io_fromRename_0_ready; // @[PipelineConnect.scala 109:31]
  wire  _GEN_1181 = dispatch_io_recv_0 ? 1'h0 : valid; // @[PipelineConnect.scala 108:24 110:{25,33}]
  wire  _GEN_1182 = leftFire | _GEN_1181; // @[PipelineConnect.scala 111:{21,29}]
  reg [9:0] data_cf_foldpc; // @[Reg.scala 16:16]
  reg  data_cf_exceptionVec_1; // @[Reg.scala 16:16]
  reg  data_cf_exceptionVec_2; // @[Reg.scala 16:16]
  reg  data_cf_exceptionVec_12; // @[Reg.scala 16:16]
  reg  data_cf_trigger_frontendHit_0; // @[Reg.scala 16:16]
  reg  data_cf_trigger_frontendHit_1; // @[Reg.scala 16:16]
  reg  data_cf_trigger_frontendHit_2; // @[Reg.scala 16:16]
  reg  data_cf_trigger_frontendHit_3; // @[Reg.scala 16:16]
  reg  data_cf_trigger_backendEn_0; // @[Reg.scala 16:16]
  reg  data_cf_trigger_backendEn_1; // @[Reg.scala 16:16]
  reg  data_cf_pd_isRVC; // @[Reg.scala 16:16]
  reg [1:0] data_cf_pd_brType; // @[Reg.scala 16:16]
  reg  data_cf_pd_isCall; // @[Reg.scala 16:16]
  reg  data_cf_pd_isRet; // @[Reg.scala 16:16]
  reg  data_cf_pred_taken; // @[Reg.scala 16:16]
  reg  data_cf_crossPageIPFFix; // @[Reg.scala 16:16]
  reg  data_cf_storeSetHit; // @[Reg.scala 16:16]
  reg  data_cf_loadWaitStrict; // @[Reg.scala 16:16]
  reg [4:0] data_cf_ssid; // @[Reg.scala 16:16]
  reg  data_cf_ftqPtr_flag; // @[Reg.scala 16:16]
  reg [2:0] data_cf_ftqPtr_value; // @[Reg.scala 16:16]
  reg [2:0] data_cf_ftqOffset; // @[Reg.scala 16:16]
  reg [1:0] data_ctrl_srcType_0; // @[Reg.scala 16:16]
  reg [1:0] data_ctrl_srcType_1; // @[Reg.scala 16:16]
  reg [1:0] data_ctrl_srcType_2; // @[Reg.scala 16:16]
  reg [4:0] data_ctrl_ldest; // @[Reg.scala 16:16]
  reg [3:0] data_ctrl_fuType; // @[Reg.scala 16:16]
  reg [6:0] data_ctrl_fuOpType; // @[Reg.scala 16:16]
  reg  data_ctrl_rfWen; // @[Reg.scala 16:16]
  reg  data_ctrl_fpWen; // @[Reg.scala 16:16]
  reg  data_ctrl_isXSTrap; // @[Reg.scala 16:16]
  reg  data_ctrl_noSpecExec; // @[Reg.scala 16:16]
  reg  data_ctrl_blockBackward; // @[Reg.scala 16:16]
  reg  data_ctrl_flushPipe; // @[Reg.scala 16:16]
  reg [3:0] data_ctrl_selImm; // @[Reg.scala 16:16]
  reg [19:0] data_ctrl_imm; // @[Reg.scala 16:16]
  reg [2:0] data_ctrl_commitType; // @[Reg.scala 16:16]
  reg  data_ctrl_fpu_isAddSub; // @[Reg.scala 16:16]
  reg  data_ctrl_fpu_typeTagIn; // @[Reg.scala 16:16]
  reg  data_ctrl_fpu_typeTagOut; // @[Reg.scala 16:16]
  reg  data_ctrl_fpu_fromInt; // @[Reg.scala 16:16]
  reg  data_ctrl_fpu_wflags; // @[Reg.scala 16:16]
  reg  data_ctrl_fpu_fpWen; // @[Reg.scala 16:16]
  reg [1:0] data_ctrl_fpu_fmaCmd; // @[Reg.scala 16:16]
  reg  data_ctrl_fpu_div; // @[Reg.scala 16:16]
  reg  data_ctrl_fpu_sqrt; // @[Reg.scala 16:16]
  reg  data_ctrl_fpu_fcvt; // @[Reg.scala 16:16]
  reg [1:0] data_ctrl_fpu_typ; // @[Reg.scala 16:16]
  reg [1:0] data_ctrl_fpu_fmt; // @[Reg.scala 16:16]
  reg  data_ctrl_fpu_ren3; // @[Reg.scala 16:16]
  reg [2:0] data_ctrl_fpu_rm; // @[Reg.scala 16:16]
  reg  data_ctrl_isMove; // @[Reg.scala 16:16]
  reg [5:0] data_psrc_0; // @[Reg.scala 16:16]
  reg [5:0] data_psrc_1; // @[Reg.scala 16:16]
  reg [5:0] data_psrc_2; // @[Reg.scala 16:16]
  reg [5:0] data_pdest; // @[Reg.scala 16:16]
  reg [5:0] data_old_pdest; // @[Reg.scala 16:16]
  reg  data_robIdx_flag; // @[Reg.scala 16:16]
  reg [4:0] data_robIdx_value; // @[Reg.scala 16:16]
  reg  data_eliminatedMove; // @[Reg.scala 16:16]
  reg  valid_1; // @[PipelineConnect.scala 108:24]
  wire  leftFire_1 = rename_io_out_1_valid & dispatch_io_fromRename_1_ready; // @[PipelineConnect.scala 109:31]
  wire  _GEN_1292 = dispatch_io_recv_1 ? 1'h0 : valid_1; // @[PipelineConnect.scala 108:24 110:{25,33}]
  wire  _GEN_1293 = leftFire_1 | _GEN_1292; // @[PipelineConnect.scala 111:{21,29}]
  reg [9:0] data_1_cf_foldpc; // @[Reg.scala 16:16]
  reg  data_1_cf_exceptionVec_1; // @[Reg.scala 16:16]
  reg  data_1_cf_exceptionVec_2; // @[Reg.scala 16:16]
  reg  data_1_cf_exceptionVec_12; // @[Reg.scala 16:16]
  reg  data_1_cf_trigger_frontendHit_0; // @[Reg.scala 16:16]
  reg  data_1_cf_trigger_frontendHit_1; // @[Reg.scala 16:16]
  reg  data_1_cf_trigger_frontendHit_2; // @[Reg.scala 16:16]
  reg  data_1_cf_trigger_frontendHit_3; // @[Reg.scala 16:16]
  reg  data_1_cf_trigger_backendEn_0; // @[Reg.scala 16:16]
  reg  data_1_cf_trigger_backendEn_1; // @[Reg.scala 16:16]
  reg  data_1_cf_pd_isRVC; // @[Reg.scala 16:16]
  reg [1:0] data_1_cf_pd_brType; // @[Reg.scala 16:16]
  reg  data_1_cf_pd_isCall; // @[Reg.scala 16:16]
  reg  data_1_cf_pd_isRet; // @[Reg.scala 16:16]
  reg  data_1_cf_pred_taken; // @[Reg.scala 16:16]
  reg  data_1_cf_crossPageIPFFix; // @[Reg.scala 16:16]
  reg  data_1_cf_storeSetHit; // @[Reg.scala 16:16]
  reg  data_1_cf_loadWaitStrict; // @[Reg.scala 16:16]
  reg [4:0] data_1_cf_ssid; // @[Reg.scala 16:16]
  reg  data_1_cf_ftqPtr_flag; // @[Reg.scala 16:16]
  reg [2:0] data_1_cf_ftqPtr_value; // @[Reg.scala 16:16]
  reg [2:0] data_1_cf_ftqOffset; // @[Reg.scala 16:16]
  reg [1:0] data_1_ctrl_srcType_0; // @[Reg.scala 16:16]
  reg [1:0] data_1_ctrl_srcType_1; // @[Reg.scala 16:16]
  reg [1:0] data_1_ctrl_srcType_2; // @[Reg.scala 16:16]
  reg [4:0] data_1_ctrl_ldest; // @[Reg.scala 16:16]
  reg [3:0] data_1_ctrl_fuType; // @[Reg.scala 16:16]
  reg [6:0] data_1_ctrl_fuOpType; // @[Reg.scala 16:16]
  reg  data_1_ctrl_rfWen; // @[Reg.scala 16:16]
  reg  data_1_ctrl_fpWen; // @[Reg.scala 16:16]
  reg  data_1_ctrl_isXSTrap; // @[Reg.scala 16:16]
  reg  data_1_ctrl_noSpecExec; // @[Reg.scala 16:16]
  reg  data_1_ctrl_blockBackward; // @[Reg.scala 16:16]
  reg  data_1_ctrl_flushPipe; // @[Reg.scala 16:16]
  reg [3:0] data_1_ctrl_selImm; // @[Reg.scala 16:16]
  reg [19:0] data_1_ctrl_imm; // @[Reg.scala 16:16]
  reg  data_1_ctrl_fpu_isAddSub; // @[Reg.scala 16:16]
  reg  data_1_ctrl_fpu_typeTagIn; // @[Reg.scala 16:16]
  reg  data_1_ctrl_fpu_typeTagOut; // @[Reg.scala 16:16]
  reg  data_1_ctrl_fpu_fromInt; // @[Reg.scala 16:16]
  reg  data_1_ctrl_fpu_wflags; // @[Reg.scala 16:16]
  reg  data_1_ctrl_fpu_fpWen; // @[Reg.scala 16:16]
  reg [1:0] data_1_ctrl_fpu_fmaCmd; // @[Reg.scala 16:16]
  reg  data_1_ctrl_fpu_div; // @[Reg.scala 16:16]
  reg  data_1_ctrl_fpu_sqrt; // @[Reg.scala 16:16]
  reg  data_1_ctrl_fpu_fcvt; // @[Reg.scala 16:16]
  reg [1:0] data_1_ctrl_fpu_typ; // @[Reg.scala 16:16]
  reg [1:0] data_1_ctrl_fpu_fmt; // @[Reg.scala 16:16]
  reg  data_1_ctrl_fpu_ren3; // @[Reg.scala 16:16]
  reg [2:0] data_1_ctrl_fpu_rm; // @[Reg.scala 16:16]
  reg  data_1_ctrl_isMove; // @[Reg.scala 16:16]
  reg [5:0] data_1_psrc_0; // @[Reg.scala 16:16]
  reg [5:0] data_1_psrc_1; // @[Reg.scala 16:16]
  reg [5:0] data_1_psrc_2; // @[Reg.scala 16:16]
  reg [5:0] data_1_pdest; // @[Reg.scala 16:16]
  reg [5:0] data_1_old_pdest; // @[Reg.scala 16:16]
  reg  data_1_robIdx_flag; // @[Reg.scala 16:16]
  reg [4:0] data_1_robIdx_value; // @[Reg.scala 16:16]
  reg  data_1_eliminatedMove; // @[Reg.scala 16:16]
  reg  dispatch_io_singleStep_REG; // @[CtrlBlock.scala 501:36]
  reg [2:0] jumpPcRead0_REG; // @[CtrlBlock.scala 543:52]
  wire  _GEN_1404 = 3'h1 == jumpPcRead0_REG ? pcMem_io_rdata_0_isNextMask_1 : pcMem_io_rdata_0_isNextMask_0; // @[NewFtq.scala 91:{42,42}]
  wire  _GEN_1405 = 3'h2 == jumpPcRead0_REG ? pcMem_io_rdata_0_isNextMask_2 : _GEN_1404; // @[NewFtq.scala 91:{42,42}]
  wire  _GEN_1406 = 3'h3 == jumpPcRead0_REG ? pcMem_io_rdata_0_isNextMask_3 : _GEN_1405; // @[NewFtq.scala 91:{42,42}]
  wire  _GEN_1407 = 3'h4 == jumpPcRead0_REG ? pcMem_io_rdata_0_isNextMask_4 : _GEN_1406; // @[NewFtq.scala 91:{42,42}]
  wire  _GEN_1408 = 3'h5 == jumpPcRead0_REG ? pcMem_io_rdata_0_isNextMask_5 : _GEN_1407; // @[NewFtq.scala 91:{42,42}]
  wire  _GEN_1409 = 3'h6 == jumpPcRead0_REG ? pcMem_io_rdata_0_isNextMask_6 : _GEN_1408; // @[NewFtq.scala 91:{42,42}]
  wire  _GEN_1410 = 3'h7 == jumpPcRead0_REG ? pcMem_io_rdata_0_isNextMask_7 : _GEN_1409; // @[NewFtq.scala 91:{42,42}]
  wire [38:0] _jumpPcRead0_T_4 = _GEN_1410 & pcMem_io_rdata_0_startAddr[4] ? pcMem_io_rdata_0_nextLineAddr :
    pcMem_io_rdata_0_startAddr; // @[NewFtq.scala 91:22]
  wire [3:0] _GEN_1438 = {{1'd0}, jumpPcRead0_REG}; // @[NewFtq.scala 92:29]
  wire [3:0] _jumpPcRead0_T_8 = pcMem_io_rdata_0_startAddr[4:1] + _GEN_1438; // @[NewFtq.scala 92:29]
  wire [37:0] jumpPcRead0_hi = {_jumpPcRead0_T_4[38:5],_jumpPcRead0_T_8}; // @[Cat.scala 31:58]
  wire [3:0] _pcMem_io_raddr_4_new_ptr_T = {io_dispatch_0_bits_cf_ftqPtr_flag,io_dispatch_0_bits_cf_ftqPtr_value}; // @[Cat.scala 31:58]
  wire [3:0] _pcMem_io_raddr_4_new_ptr_T_2 = _pcMem_io_raddr_4_new_ptr_T + 4'h1; // @[CircularQueuePtr.scala 39:46]
  reg  read_from_newest_entry_REG_flag; // @[CtrlBlock.scala 551:39]
  reg [2:0] read_from_newest_entry_REG_value; // @[CtrlBlock.scala 551:39]
  reg  read_from_newest_entry_REG_1_flag; // @[CtrlBlock.scala 551:70]
  reg [2:0] read_from_newest_entry_REG_1_value; // @[CtrlBlock.scala 551:70]
  wire [3:0] _read_from_newest_entry_T = {read_from_newest_entry_REG_flag,read_from_newest_entry_REG_value}; // @[CircularQueuePtr.scala 61:50]
  wire [3:0] _read_from_newest_entry_T_1 = {read_from_newest_entry_REG_1_flag,read_from_newest_entry_REG_1_value}; // @[CircularQueuePtr.scala 61:70]
  wire  read_from_newest_entry = _read_from_newest_entry_T == _read_from_newest_entry_T_1; // @[CircularQueuePtr.scala 61:52]
  reg [38:0] io_jalr_target_REG; // @[CtrlBlock.scala 552:56]
  wire [5:0] _sources_exuOutput_3_valid_flushItself_T_1 = {io_writeback_0_3_bits_uop_robIdx_flag,
    io_writeback_0_3_bits_uop_robIdx_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _sources_exuOutput_3_valid_flushItself_T_3 = _sources_exuOutput_3_valid_flushItself_T_1 ==
    _exuRedirect_killedByOlder_flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  sources_exuOutput_3_valid_flushItself = stage2Redirect_bits_level & _sources_exuOutput_3_valid_flushItself_T_3; // @[Rob.scala 122:51]
  wire  sources_exuOutput_3_valid_differentFlag = io_writeback_0_3_bits_uop_robIdx_flag ^
    stage2Redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  sources_exuOutput_3_valid_compare = io_writeback_0_3_bits_uop_robIdx_value > stage2Redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _sources_exuOutput_3_valid_T = sources_exuOutput_3_valid_differentFlag ^ sources_exuOutput_3_valid_compare; // @[CircularQueuePtr.scala 88:19]
  wire  _sources_exuOutput_3_valid_T_2 = stage2Redirect_valid & (sources_exuOutput_3_valid_flushItself |
    _sources_exuOutput_3_valid_T); // @[Rob.scala 123:20]
  wire  _sources_exuOutput_3_valid_flushItself_T_7 = _sources_exuOutput_3_valid_flushItself_T_1 ==
    _exuRedirect_killedByOlder_flushItself_T_6; // @[CircularQueuePtr.scala 61:52]
  wire  sources_exuOutput_3_valid_flushItself_1 = redirectForExu_next_bits_rlevel &
    _sources_exuOutput_3_valid_flushItself_T_7; // @[Rob.scala 122:51]
  wire  sources_exuOutput_3_valid_differentFlag_1 = io_writeback_0_3_bits_uop_robIdx_flag ^
    redirectForExu_next_bits_rrobIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  sources_exuOutput_3_valid_compare_1 = io_writeback_0_3_bits_uop_robIdx_value >
    redirectForExu_next_bits_rrobIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _sources_exuOutput_3_valid_T_3 = sources_exuOutput_3_valid_differentFlag_1 ^ sources_exuOutput_3_valid_compare_1
    ; // @[CircularQueuePtr.scala 88:19]
  wire  _sources_exuOutput_3_valid_T_5 = redirectForExu_next_valid_REG & (sources_exuOutput_3_valid_flushItself_1 |
    _sources_exuOutput_3_valid_T_3); // @[Rob.scala 123:20]
  wire [1:0] _sources_exuOutput_3_valid_T_6 = {_sources_exuOutput_3_valid_T_5,_sources_exuOutput_3_valid_T_2}; // @[Rob.scala 126:90]
  wire  _sources_exuOutput_3_valid_T_7 = |_sources_exuOutput_3_valid_T_6; // @[Rob.scala 126:97]
  wire [5:0] _sources_exuOutput_4_valid_flushItself_T_1 = {io_writeback_0_4_bits_uop_robIdx_flag,
    io_writeback_0_4_bits_uop_robIdx_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _sources_exuOutput_4_valid_flushItself_T_3 = _sources_exuOutput_4_valid_flushItself_T_1 ==
    _exuRedirect_killedByOlder_flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  sources_exuOutput_4_valid_flushItself = stage2Redirect_bits_level & _sources_exuOutput_4_valid_flushItself_T_3; // @[Rob.scala 122:51]
  wire  sources_exuOutput_4_valid_differentFlag = io_writeback_0_4_bits_uop_robIdx_flag ^
    stage2Redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  sources_exuOutput_4_valid_compare = io_writeback_0_4_bits_uop_robIdx_value > stage2Redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _sources_exuOutput_4_valid_T = sources_exuOutput_4_valid_differentFlag ^ sources_exuOutput_4_valid_compare; // @[CircularQueuePtr.scala 88:19]
  wire  _sources_exuOutput_4_valid_T_2 = stage2Redirect_valid & (sources_exuOutput_4_valid_flushItself |
    _sources_exuOutput_4_valid_T); // @[Rob.scala 123:20]
  wire  _sources_exuOutput_4_valid_flushItself_T_7 = _sources_exuOutput_4_valid_flushItself_T_1 ==
    _exuRedirect_killedByOlder_flushItself_T_6; // @[CircularQueuePtr.scala 61:52]
  wire  sources_exuOutput_4_valid_flushItself_1 = redirectForExu_next_bits_rlevel &
    _sources_exuOutput_4_valid_flushItself_T_7; // @[Rob.scala 122:51]
  wire  sources_exuOutput_4_valid_differentFlag_1 = io_writeback_0_4_bits_uop_robIdx_flag ^
    redirectForExu_next_bits_rrobIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  sources_exuOutput_4_valid_compare_1 = io_writeback_0_4_bits_uop_robIdx_value >
    redirectForExu_next_bits_rrobIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _sources_exuOutput_4_valid_T_3 = sources_exuOutput_4_valid_differentFlag_1 ^ sources_exuOutput_4_valid_compare_1
    ; // @[CircularQueuePtr.scala 88:19]
  wire  _sources_exuOutput_4_valid_T_5 = redirectForExu_next_valid_REG & (sources_exuOutput_4_valid_flushItself_1 |
    _sources_exuOutput_4_valid_T_3); // @[Rob.scala 123:20]
  wire [1:0] _sources_exuOutput_4_valid_T_6 = {_sources_exuOutput_4_valid_T_5,_sources_exuOutput_4_valid_T_2}; // @[Rob.scala 126:90]
  wire  _sources_exuOutput_4_valid_T_7 = |_sources_exuOutput_4_valid_T_6; // @[Rob.scala 126:97]
  wire [5:0] _sources_exuOutput_5_valid_flushItself_T_1 = {io_writeback_0_5_bits_uop_robIdx_flag,
    io_writeback_0_5_bits_uop_robIdx_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _sources_exuOutput_5_valid_flushItself_T_3 = _sources_exuOutput_5_valid_flushItself_T_1 ==
    _exuRedirect_killedByOlder_flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  sources_exuOutput_5_valid_flushItself = stage2Redirect_bits_level & _sources_exuOutput_5_valid_flushItself_T_3; // @[Rob.scala 122:51]
  wire  sources_exuOutput_5_valid_differentFlag = io_writeback_0_5_bits_uop_robIdx_flag ^
    stage2Redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  sources_exuOutput_5_valid_compare = io_writeback_0_5_bits_uop_robIdx_value > stage2Redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _sources_exuOutput_5_valid_T = sources_exuOutput_5_valid_differentFlag ^ sources_exuOutput_5_valid_compare; // @[CircularQueuePtr.scala 88:19]
  wire  _sources_exuOutput_5_valid_T_2 = stage2Redirect_valid & (sources_exuOutput_5_valid_flushItself |
    _sources_exuOutput_5_valid_T); // @[Rob.scala 123:20]
  wire  _sources_exuOutput_5_valid_flushItself_T_7 = _sources_exuOutput_5_valid_flushItself_T_1 ==
    _exuRedirect_killedByOlder_flushItself_T_6; // @[CircularQueuePtr.scala 61:52]
  wire  sources_exuOutput_5_valid_flushItself_1 = redirectForExu_next_bits_rlevel &
    _sources_exuOutput_5_valid_flushItself_T_7; // @[Rob.scala 122:51]
  wire  sources_exuOutput_5_valid_differentFlag_1 = io_writeback_0_5_bits_uop_robIdx_flag ^
    redirectForExu_next_bits_rrobIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  sources_exuOutput_5_valid_compare_1 = io_writeback_0_5_bits_uop_robIdx_value >
    redirectForExu_next_bits_rrobIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _sources_exuOutput_5_valid_T_3 = sources_exuOutput_5_valid_differentFlag_1 ^ sources_exuOutput_5_valid_compare_1
    ; // @[CircularQueuePtr.scala 88:19]
  wire  _sources_exuOutput_5_valid_T_5 = redirectForExu_next_valid_REG & (sources_exuOutput_5_valid_flushItself_1 |
    _sources_exuOutput_5_valid_T_3); // @[Rob.scala 123:20]
  wire [1:0] _sources_exuOutput_5_valid_T_6 = {_sources_exuOutput_5_valid_T_5,_sources_exuOutput_5_valid_T_2}; // @[Rob.scala 126:90]
  wire  _sources_exuOutput_5_valid_T_7 = |_sources_exuOutput_5_valid_T_6; // @[Rob.scala 126:97]
  wire [5:0] _sources_exuOutput_6_valid_flushItself_T_1 = {io_writeback_0_6_bits_uop_robIdx_flag,
    io_writeback_0_6_bits_uop_robIdx_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _sources_exuOutput_6_valid_flushItself_T_3 = _sources_exuOutput_6_valid_flushItself_T_1 ==
    _exuRedirect_killedByOlder_flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  sources_exuOutput_6_valid_flushItself = stage2Redirect_bits_level & _sources_exuOutput_6_valid_flushItself_T_3; // @[Rob.scala 122:51]
  wire  sources_exuOutput_6_valid_differentFlag = io_writeback_0_6_bits_uop_robIdx_flag ^
    stage2Redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  sources_exuOutput_6_valid_compare = io_writeback_0_6_bits_uop_robIdx_value > stage2Redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _sources_exuOutput_6_valid_T = sources_exuOutput_6_valid_differentFlag ^ sources_exuOutput_6_valid_compare; // @[CircularQueuePtr.scala 88:19]
  wire  _sources_exuOutput_6_valid_T_2 = stage2Redirect_valid & (sources_exuOutput_6_valid_flushItself |
    _sources_exuOutput_6_valid_T); // @[Rob.scala 123:20]
  wire  _sources_exuOutput_6_valid_flushItself_T_7 = _sources_exuOutput_6_valid_flushItself_T_1 ==
    _exuRedirect_killedByOlder_flushItself_T_6; // @[CircularQueuePtr.scala 61:52]
  wire  sources_exuOutput_6_valid_flushItself_1 = redirectForExu_next_bits_rlevel &
    _sources_exuOutput_6_valid_flushItself_T_7; // @[Rob.scala 122:51]
  wire  sources_exuOutput_6_valid_differentFlag_1 = io_writeback_0_6_bits_uop_robIdx_flag ^
    redirectForExu_next_bits_rrobIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  sources_exuOutput_6_valid_compare_1 = io_writeback_0_6_bits_uop_robIdx_value >
    redirectForExu_next_bits_rrobIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _sources_exuOutput_6_valid_T_3 = sources_exuOutput_6_valid_differentFlag_1 ^ sources_exuOutput_6_valid_compare_1
    ; // @[CircularQueuePtr.scala 88:19]
  wire  _sources_exuOutput_6_valid_T_5 = redirectForExu_next_valid_REG & (sources_exuOutput_6_valid_flushItself_1 |
    _sources_exuOutput_6_valid_T_3); // @[Rob.scala 123:20]
  wire [1:0] _sources_exuOutput_6_valid_T_6 = {_sources_exuOutput_6_valid_T_5,_sources_exuOutput_6_valid_T_2}; // @[Rob.scala 126:90]
  wire  _sources_exuOutput_6_valid_T_7 = |_sources_exuOutput_6_valid_T_6; // @[Rob.scala 126:97]
  wire [5:0] _sources_exuOutput_7_valid_flushItself_T_1 = {io_writeback_0_7_bits_uop_robIdx_flag,
    io_writeback_0_7_bits_uop_robIdx_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _sources_exuOutput_7_valid_flushItself_T_3 = _sources_exuOutput_7_valid_flushItself_T_1 ==
    _exuRedirect_killedByOlder_flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  sources_exuOutput_7_valid_flushItself = stage2Redirect_bits_level & _sources_exuOutput_7_valid_flushItself_T_3; // @[Rob.scala 122:51]
  wire  sources_exuOutput_7_valid_differentFlag = io_writeback_0_7_bits_uop_robIdx_flag ^
    stage2Redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  sources_exuOutput_7_valid_compare = io_writeback_0_7_bits_uop_robIdx_value > stage2Redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _sources_exuOutput_7_valid_T = sources_exuOutput_7_valid_differentFlag ^ sources_exuOutput_7_valid_compare; // @[CircularQueuePtr.scala 88:19]
  wire  _sources_exuOutput_7_valid_T_2 = stage2Redirect_valid & (sources_exuOutput_7_valid_flushItself |
    _sources_exuOutput_7_valid_T); // @[Rob.scala 123:20]
  wire  _sources_exuOutput_7_valid_flushItself_T_7 = _sources_exuOutput_7_valid_flushItself_T_1 ==
    _exuRedirect_killedByOlder_flushItself_T_6; // @[CircularQueuePtr.scala 61:52]
  wire  sources_exuOutput_7_valid_flushItself_1 = redirectForExu_next_bits_rlevel &
    _sources_exuOutput_7_valid_flushItself_T_7; // @[Rob.scala 122:51]
  wire  sources_exuOutput_7_valid_differentFlag_1 = io_writeback_0_7_bits_uop_robIdx_flag ^
    redirectForExu_next_bits_rrobIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  sources_exuOutput_7_valid_compare_1 = io_writeback_0_7_bits_uop_robIdx_value >
    redirectForExu_next_bits_rrobIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _sources_exuOutput_7_valid_T_3 = sources_exuOutput_7_valid_differentFlag_1 ^ sources_exuOutput_7_valid_compare_1
    ; // @[CircularQueuePtr.scala 88:19]
  wire  _sources_exuOutput_7_valid_T_5 = redirectForExu_next_valid_REG & (sources_exuOutput_7_valid_flushItself_1 |
    _sources_exuOutput_7_valid_T_3); // @[Rob.scala 123:20]
  wire [1:0] _sources_exuOutput_7_valid_T_6 = {_sources_exuOutput_7_valid_T_5,_sources_exuOutput_7_valid_T_2}; // @[Rob.scala 126:90]
  wire  _sources_exuOutput_7_valid_T_7 = |_sources_exuOutput_7_valid_T_6; // @[Rob.scala 126:97]
  wire [5:0] _sources_exuOutput_8_valid_flushItself_T_1 = {io_writeback_0_8_bits_uop_robIdx_flag,
    io_writeback_0_8_bits_uop_robIdx_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _sources_exuOutput_8_valid_flushItself_T_3 = _sources_exuOutput_8_valid_flushItself_T_1 ==
    _exuRedirect_killedByOlder_flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  sources_exuOutput_8_valid_flushItself = stage2Redirect_bits_level & _sources_exuOutput_8_valid_flushItself_T_3; // @[Rob.scala 122:51]
  wire  sources_exuOutput_8_valid_differentFlag = io_writeback_0_8_bits_uop_robIdx_flag ^
    stage2Redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  sources_exuOutput_8_valid_compare = io_writeback_0_8_bits_uop_robIdx_value > stage2Redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _sources_exuOutput_8_valid_T = sources_exuOutput_8_valid_differentFlag ^ sources_exuOutput_8_valid_compare; // @[CircularQueuePtr.scala 88:19]
  wire  _sources_exuOutput_8_valid_T_2 = stage2Redirect_valid & (sources_exuOutput_8_valid_flushItself |
    _sources_exuOutput_8_valid_T); // @[Rob.scala 123:20]
  wire  _sources_exuOutput_8_valid_flushItself_T_7 = _sources_exuOutput_8_valid_flushItself_T_1 ==
    _exuRedirect_killedByOlder_flushItself_T_6; // @[CircularQueuePtr.scala 61:52]
  wire  sources_exuOutput_8_valid_flushItself_1 = redirectForExu_next_bits_rlevel &
    _sources_exuOutput_8_valid_flushItself_T_7; // @[Rob.scala 122:51]
  wire  sources_exuOutput_8_valid_differentFlag_1 = io_writeback_0_8_bits_uop_robIdx_flag ^
    redirectForExu_next_bits_rrobIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  sources_exuOutput_8_valid_compare_1 = io_writeback_0_8_bits_uop_robIdx_value >
    redirectForExu_next_bits_rrobIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _sources_exuOutput_8_valid_T_3 = sources_exuOutput_8_valid_differentFlag_1 ^ sources_exuOutput_8_valid_compare_1
    ; // @[CircularQueuePtr.scala 88:19]
  wire  _sources_exuOutput_8_valid_T_5 = redirectForExu_next_valid_REG & (sources_exuOutput_8_valid_flushItself_1 |
    _sources_exuOutput_8_valid_T_3); // @[Rob.scala 123:20]
  wire [1:0] _sources_exuOutput_8_valid_T_6 = {_sources_exuOutput_8_valid_T_5,_sources_exuOutput_8_valid_T_2}; // @[Rob.scala 126:90]
  wire  _sources_exuOutput_8_valid_T_7 = |_sources_exuOutput_8_valid_T_6; // @[Rob.scala 126:97]
  wire [5:0] _sources_exuOutput_9_valid_flushItself_T_1 = {io_writeback_0_9_bits_uop_robIdx_flag,
    io_writeback_0_9_bits_uop_robIdx_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _sources_exuOutput_9_valid_flushItself_T_3 = _sources_exuOutput_9_valid_flushItself_T_1 ==
    _exuRedirect_killedByOlder_flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  sources_exuOutput_9_valid_flushItself = stage2Redirect_bits_level & _sources_exuOutput_9_valid_flushItself_T_3; // @[Rob.scala 122:51]
  wire  sources_exuOutput_9_valid_differentFlag = io_writeback_0_9_bits_uop_robIdx_flag ^
    stage2Redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  sources_exuOutput_9_valid_compare = io_writeback_0_9_bits_uop_robIdx_value > stage2Redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _sources_exuOutput_9_valid_T = sources_exuOutput_9_valid_differentFlag ^ sources_exuOutput_9_valid_compare; // @[CircularQueuePtr.scala 88:19]
  wire  _sources_exuOutput_9_valid_T_2 = stage2Redirect_valid & (sources_exuOutput_9_valid_flushItself |
    _sources_exuOutput_9_valid_T); // @[Rob.scala 123:20]
  wire  _sources_exuOutput_9_valid_flushItself_T_7 = _sources_exuOutput_9_valid_flushItself_T_1 ==
    _exuRedirect_killedByOlder_flushItself_T_6; // @[CircularQueuePtr.scala 61:52]
  wire  sources_exuOutput_9_valid_flushItself_1 = redirectForExu_next_bits_rlevel &
    _sources_exuOutput_9_valid_flushItself_T_7; // @[Rob.scala 122:51]
  wire  sources_exuOutput_9_valid_differentFlag_1 = io_writeback_0_9_bits_uop_robIdx_flag ^
    redirectForExu_next_bits_rrobIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  sources_exuOutput_9_valid_compare_1 = io_writeback_0_9_bits_uop_robIdx_value >
    redirectForExu_next_bits_rrobIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _sources_exuOutput_9_valid_T_3 = sources_exuOutput_9_valid_differentFlag_1 ^ sources_exuOutput_9_valid_compare_1
    ; // @[CircularQueuePtr.scala 88:19]
  wire  _sources_exuOutput_9_valid_T_5 = redirectForExu_next_valid_REG & (sources_exuOutput_9_valid_flushItself_1 |
    _sources_exuOutput_9_valid_T_3); // @[Rob.scala 123:20]
  wire [1:0] _sources_exuOutput_9_valid_T_6 = {_sources_exuOutput_9_valid_T_5,_sources_exuOutput_9_valid_T_2}; // @[Rob.scala 126:90]
  wire  _sources_exuOutput_9_valid_T_7 = |_sources_exuOutput_9_valid_T_6; // @[Rob.scala 126:97]
  wire [5:0] _sources_exuOutput_0_valid_flushItself_T_9 = {io_writeback_1_0_bits_uop_robIdx_flag,
    io_writeback_1_0_bits_uop_robIdx_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _sources_exuOutput_0_valid_flushItself_T_11 = _sources_exuOutput_0_valid_flushItself_T_9 ==
    _exuRedirect_killedByOlder_flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  sources_exuOutput_0_valid_flushItself_2 = stage2Redirect_bits_level &
    _sources_exuOutput_0_valid_flushItself_T_11; // @[Rob.scala 122:51]
  wire  sources_exuOutput_0_valid_differentFlag_2 = io_writeback_1_0_bits_uop_robIdx_flag ^
    stage2Redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  sources_exuOutput_0_valid_compare_2 = io_writeback_1_0_bits_uop_robIdx_value > stage2Redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _sources_exuOutput_0_valid_T_10 = sources_exuOutput_0_valid_differentFlag_2 ^
    sources_exuOutput_0_valid_compare_2; // @[CircularQueuePtr.scala 88:19]
  wire  _sources_exuOutput_0_valid_T_12 = stage2Redirect_valid & (sources_exuOutput_0_valid_flushItself_2 |
    _sources_exuOutput_0_valid_T_10); // @[Rob.scala 123:20]
  wire  _sources_exuOutput_0_valid_flushItself_T_15 = _sources_exuOutput_0_valid_flushItself_T_9 ==
    _exuRedirect_killedByOlder_flushItself_T_6; // @[CircularQueuePtr.scala 61:52]
  wire  sources_exuOutput_0_valid_flushItself_3 = redirectForExu_next_bits_rlevel &
    _sources_exuOutput_0_valid_flushItself_T_15; // @[Rob.scala 122:51]
  wire  sources_exuOutput_0_valid_differentFlag_3 = io_writeback_1_0_bits_uop_robIdx_flag ^
    redirectForExu_next_bits_rrobIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  sources_exuOutput_0_valid_compare_3 = io_writeback_1_0_bits_uop_robIdx_value >
    redirectForExu_next_bits_rrobIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _sources_exuOutput_0_valid_T_13 = sources_exuOutput_0_valid_differentFlag_3 ^
    sources_exuOutput_0_valid_compare_3; // @[CircularQueuePtr.scala 88:19]
  wire  _sources_exuOutput_0_valid_T_15 = redirectForExu_next_valid_REG & (sources_exuOutput_0_valid_flushItself_3 |
    _sources_exuOutput_0_valid_T_13); // @[Rob.scala 123:20]
  wire [1:0] _sources_exuOutput_0_valid_T_16 = {_sources_exuOutput_0_valid_T_15,_sources_exuOutput_0_valid_T_12}; // @[Rob.scala 126:90]
  wire  _sources_exuOutput_0_valid_T_17 = |_sources_exuOutput_0_valid_T_16; // @[Rob.scala 126:97]
  wire [5:0] _sources_exuOutput_1_valid_flushItself_T_9 = {io_writeback_1_1_bits_uop_robIdx_flag,
    io_writeback_1_1_bits_uop_robIdx_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _sources_exuOutput_1_valid_flushItself_T_11 = _sources_exuOutput_1_valid_flushItself_T_9 ==
    _exuRedirect_killedByOlder_flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  sources_exuOutput_1_valid_flushItself_2 = stage2Redirect_bits_level &
    _sources_exuOutput_1_valid_flushItself_T_11; // @[Rob.scala 122:51]
  wire  sources_exuOutput_1_valid_differentFlag_2 = io_writeback_1_1_bits_uop_robIdx_flag ^
    stage2Redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  sources_exuOutput_1_valid_compare_2 = io_writeback_1_1_bits_uop_robIdx_value > stage2Redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _sources_exuOutput_1_valid_T_10 = sources_exuOutput_1_valid_differentFlag_2 ^
    sources_exuOutput_1_valid_compare_2; // @[CircularQueuePtr.scala 88:19]
  wire  _sources_exuOutput_1_valid_T_12 = stage2Redirect_valid & (sources_exuOutput_1_valid_flushItself_2 |
    _sources_exuOutput_1_valid_T_10); // @[Rob.scala 123:20]
  wire  _sources_exuOutput_1_valid_flushItself_T_15 = _sources_exuOutput_1_valid_flushItself_T_9 ==
    _exuRedirect_killedByOlder_flushItself_T_6; // @[CircularQueuePtr.scala 61:52]
  wire  sources_exuOutput_1_valid_flushItself_3 = redirectForExu_next_bits_rlevel &
    _sources_exuOutput_1_valid_flushItself_T_15; // @[Rob.scala 122:51]
  wire  sources_exuOutput_1_valid_differentFlag_3 = io_writeback_1_1_bits_uop_robIdx_flag ^
    redirectForExu_next_bits_rrobIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  sources_exuOutput_1_valid_compare_3 = io_writeback_1_1_bits_uop_robIdx_value >
    redirectForExu_next_bits_rrobIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _sources_exuOutput_1_valid_T_13 = sources_exuOutput_1_valid_differentFlag_3 ^
    sources_exuOutput_1_valid_compare_3; // @[CircularQueuePtr.scala 88:19]
  wire  _sources_exuOutput_1_valid_T_15 = redirectForExu_next_valid_REG & (sources_exuOutput_1_valid_flushItself_3 |
    _sources_exuOutput_1_valid_T_13); // @[Rob.scala 123:20]
  wire [1:0] _sources_exuOutput_1_valid_T_16 = {_sources_exuOutput_1_valid_T_15,_sources_exuOutput_1_valid_T_12}; // @[Rob.scala 126:90]
  wire  _sources_exuOutput_1_valid_T_17 = |_sources_exuOutput_1_valid_T_16; // @[Rob.scala 126:97]
  wire [5:0] _sources_exuOutput_2_valid_flushItself_T_9 = {io_writeback_1_2_bits_uop_robIdx_flag,
    io_writeback_1_2_bits_uop_robIdx_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _sources_exuOutput_2_valid_flushItself_T_11 = _sources_exuOutput_2_valid_flushItself_T_9 ==
    _exuRedirect_killedByOlder_flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  sources_exuOutput_2_valid_flushItself_2 = stage2Redirect_bits_level &
    _sources_exuOutput_2_valid_flushItself_T_11; // @[Rob.scala 122:51]
  wire  sources_exuOutput_2_valid_differentFlag_2 = io_writeback_1_2_bits_uop_robIdx_flag ^
    stage2Redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  sources_exuOutput_2_valid_compare_2 = io_writeback_1_2_bits_uop_robIdx_value > stage2Redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _sources_exuOutput_2_valid_T_10 = sources_exuOutput_2_valid_differentFlag_2 ^
    sources_exuOutput_2_valid_compare_2; // @[CircularQueuePtr.scala 88:19]
  wire  _sources_exuOutput_2_valid_T_12 = stage2Redirect_valid & (sources_exuOutput_2_valid_flushItself_2 |
    _sources_exuOutput_2_valid_T_10); // @[Rob.scala 123:20]
  wire  _sources_exuOutput_2_valid_flushItself_T_15 = _sources_exuOutput_2_valid_flushItself_T_9 ==
    _exuRedirect_killedByOlder_flushItself_T_6; // @[CircularQueuePtr.scala 61:52]
  wire  sources_exuOutput_2_valid_flushItself_3 = redirectForExu_next_bits_rlevel &
    _sources_exuOutput_2_valid_flushItself_T_15; // @[Rob.scala 122:51]
  wire  sources_exuOutput_2_valid_differentFlag_3 = io_writeback_1_2_bits_uop_robIdx_flag ^
    redirectForExu_next_bits_rrobIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  sources_exuOutput_2_valid_compare_3 = io_writeback_1_2_bits_uop_robIdx_value >
    redirectForExu_next_bits_rrobIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _sources_exuOutput_2_valid_T_13 = sources_exuOutput_2_valid_differentFlag_3 ^
    sources_exuOutput_2_valid_compare_3; // @[CircularQueuePtr.scala 88:19]
  wire  _sources_exuOutput_2_valid_T_15 = redirectForExu_next_valid_REG & (sources_exuOutput_2_valid_flushItself_3 |
    _sources_exuOutput_2_valid_T_13); // @[Rob.scala 123:20]
  wire [1:0] _sources_exuOutput_2_valid_T_16 = {_sources_exuOutput_2_valid_T_15,_sources_exuOutput_2_valid_T_12}; // @[Rob.scala 126:90]
  wire  _sources_exuOutput_2_valid_T_17 = |_sources_exuOutput_2_valid_T_16; // @[Rob.scala 126:97]
  wire [5:0] _sources_exuOutput_3_valid_flushItself_T_9 = {io_writeback_1_3_bits_uop_robIdx_flag,
    io_writeback_1_3_bits_uop_robIdx_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _sources_exuOutput_3_valid_flushItself_T_11 = _sources_exuOutput_3_valid_flushItself_T_9 ==
    _exuRedirect_killedByOlder_flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  sources_exuOutput_3_valid_flushItself_2 = stage2Redirect_bits_level &
    _sources_exuOutput_3_valid_flushItself_T_11; // @[Rob.scala 122:51]
  wire  sources_exuOutput_3_valid_differentFlag_2 = io_writeback_1_3_bits_uop_robIdx_flag ^
    stage2Redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  sources_exuOutput_3_valid_compare_2 = io_writeback_1_3_bits_uop_robIdx_value > stage2Redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _sources_exuOutput_3_valid_T_10 = sources_exuOutput_3_valid_differentFlag_2 ^
    sources_exuOutput_3_valid_compare_2; // @[CircularQueuePtr.scala 88:19]
  wire  _sources_exuOutput_3_valid_T_12 = stage2Redirect_valid & (sources_exuOutput_3_valid_flushItself_2 |
    _sources_exuOutput_3_valid_T_10); // @[Rob.scala 123:20]
  wire  _sources_exuOutput_3_valid_flushItself_T_15 = _sources_exuOutput_3_valid_flushItself_T_9 ==
    _exuRedirect_killedByOlder_flushItself_T_6; // @[CircularQueuePtr.scala 61:52]
  wire  sources_exuOutput_3_valid_flushItself_3 = redirectForExu_next_bits_rlevel &
    _sources_exuOutput_3_valid_flushItself_T_15; // @[Rob.scala 122:51]
  wire  sources_exuOutput_3_valid_differentFlag_3 = io_writeback_1_3_bits_uop_robIdx_flag ^
    redirectForExu_next_bits_rrobIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  sources_exuOutput_3_valid_compare_3 = io_writeback_1_3_bits_uop_robIdx_value >
    redirectForExu_next_bits_rrobIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _sources_exuOutput_3_valid_T_13 = sources_exuOutput_3_valid_differentFlag_3 ^
    sources_exuOutput_3_valid_compare_3; // @[CircularQueuePtr.scala 88:19]
  wire  _sources_exuOutput_3_valid_T_15 = redirectForExu_next_valid_REG & (sources_exuOutput_3_valid_flushItself_3 |
    _sources_exuOutput_3_valid_T_13); // @[Rob.scala 123:20]
  wire [1:0] _sources_exuOutput_3_valid_T_16 = {_sources_exuOutput_3_valid_T_15,_sources_exuOutput_3_valid_T_12}; // @[Rob.scala 126:90]
  wire  _sources_exuOutput_3_valid_T_17 = |_sources_exuOutput_3_valid_T_16; // @[Rob.scala 126:97]
  wire [5:0] _sources_exuOutput_4_valid_flushItself_T_9 = {io_writeback_1_4_bits_uop_robIdx_flag,
    io_writeback_1_4_bits_uop_robIdx_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _sources_exuOutput_4_valid_flushItself_T_11 = _sources_exuOutput_4_valid_flushItself_T_9 ==
    _exuRedirect_killedByOlder_flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  sources_exuOutput_4_valid_flushItself_2 = stage2Redirect_bits_level &
    _sources_exuOutput_4_valid_flushItself_T_11; // @[Rob.scala 122:51]
  wire  sources_exuOutput_4_valid_differentFlag_2 = io_writeback_1_4_bits_uop_robIdx_flag ^
    stage2Redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  sources_exuOutput_4_valid_compare_2 = io_writeback_1_4_bits_uop_robIdx_value > stage2Redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _sources_exuOutput_4_valid_T_10 = sources_exuOutput_4_valid_differentFlag_2 ^
    sources_exuOutput_4_valid_compare_2; // @[CircularQueuePtr.scala 88:19]
  wire  _sources_exuOutput_4_valid_T_12 = stage2Redirect_valid & (sources_exuOutput_4_valid_flushItself_2 |
    _sources_exuOutput_4_valid_T_10); // @[Rob.scala 123:20]
  wire  _sources_exuOutput_4_valid_flushItself_T_15 = _sources_exuOutput_4_valid_flushItself_T_9 ==
    _exuRedirect_killedByOlder_flushItself_T_6; // @[CircularQueuePtr.scala 61:52]
  wire  sources_exuOutput_4_valid_flushItself_3 = redirectForExu_next_bits_rlevel &
    _sources_exuOutput_4_valid_flushItself_T_15; // @[Rob.scala 122:51]
  wire  sources_exuOutput_4_valid_differentFlag_3 = io_writeback_1_4_bits_uop_robIdx_flag ^
    redirectForExu_next_bits_rrobIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  sources_exuOutput_4_valid_compare_3 = io_writeback_1_4_bits_uop_robIdx_value >
    redirectForExu_next_bits_rrobIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _sources_exuOutput_4_valid_T_13 = sources_exuOutput_4_valid_differentFlag_3 ^
    sources_exuOutput_4_valid_compare_3; // @[CircularQueuePtr.scala 88:19]
  wire  _sources_exuOutput_4_valid_T_15 = redirectForExu_next_valid_REG & (sources_exuOutput_4_valid_flushItself_3 |
    _sources_exuOutput_4_valid_T_13); // @[Rob.scala 123:20]
  wire [1:0] _sources_exuOutput_4_valid_T_16 = {_sources_exuOutput_4_valid_T_15,_sources_exuOutput_4_valid_T_12}; // @[Rob.scala 126:90]
  wire  _sources_exuOutput_4_valid_T_17 = |_sources_exuOutput_4_valid_T_16; // @[Rob.scala 126:97]
  wire [5:0] _sources_exuOutput_5_valid_flushItself_T_9 = {io_writeback_1_5_bits_uop_robIdx_flag,
    io_writeback_1_5_bits_uop_robIdx_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _sources_exuOutput_5_valid_flushItself_T_11 = _sources_exuOutput_5_valid_flushItself_T_9 ==
    _exuRedirect_killedByOlder_flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  sources_exuOutput_5_valid_flushItself_2 = stage2Redirect_bits_level &
    _sources_exuOutput_5_valid_flushItself_T_11; // @[Rob.scala 122:51]
  wire  sources_exuOutput_5_valid_differentFlag_2 = io_writeback_1_5_bits_uop_robIdx_flag ^
    stage2Redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  sources_exuOutput_5_valid_compare_2 = io_writeback_1_5_bits_uop_robIdx_value > stage2Redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _sources_exuOutput_5_valid_T_10 = sources_exuOutput_5_valid_differentFlag_2 ^
    sources_exuOutput_5_valid_compare_2; // @[CircularQueuePtr.scala 88:19]
  wire  _sources_exuOutput_5_valid_T_12 = stage2Redirect_valid & (sources_exuOutput_5_valid_flushItself_2 |
    _sources_exuOutput_5_valid_T_10); // @[Rob.scala 123:20]
  wire  _sources_exuOutput_5_valid_flushItself_T_15 = _sources_exuOutput_5_valid_flushItself_T_9 ==
    _exuRedirect_killedByOlder_flushItself_T_6; // @[CircularQueuePtr.scala 61:52]
  wire  sources_exuOutput_5_valid_flushItself_3 = redirectForExu_next_bits_rlevel &
    _sources_exuOutput_5_valid_flushItself_T_15; // @[Rob.scala 122:51]
  wire  sources_exuOutput_5_valid_differentFlag_3 = io_writeback_1_5_bits_uop_robIdx_flag ^
    redirectForExu_next_bits_rrobIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  sources_exuOutput_5_valid_compare_3 = io_writeback_1_5_bits_uop_robIdx_value >
    redirectForExu_next_bits_rrobIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _sources_exuOutput_5_valid_T_13 = sources_exuOutput_5_valid_differentFlag_3 ^
    sources_exuOutput_5_valid_compare_3; // @[CircularQueuePtr.scala 88:19]
  wire  _sources_exuOutput_5_valid_T_15 = redirectForExu_next_valid_REG & (sources_exuOutput_5_valid_flushItself_3 |
    _sources_exuOutput_5_valid_T_13); // @[Rob.scala 123:20]
  wire [1:0] _sources_exuOutput_5_valid_T_16 = {_sources_exuOutput_5_valid_T_15,_sources_exuOutput_5_valid_T_12}; // @[Rob.scala 126:90]
  wire  _sources_exuOutput_5_valid_T_17 = |_sources_exuOutput_5_valid_T_16; // @[Rob.scala 126:97]
  wire [5:0] _sources_exuOutput_6_valid_flushItself_T_9 = {io_writeback_1_6_bits_uop_robIdx_flag,
    io_writeback_1_6_bits_uop_robIdx_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _sources_exuOutput_6_valid_flushItself_T_11 = _sources_exuOutput_6_valid_flushItself_T_9 ==
    _exuRedirect_killedByOlder_flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  sources_exuOutput_6_valid_flushItself_2 = stage2Redirect_bits_level &
    _sources_exuOutput_6_valid_flushItself_T_11; // @[Rob.scala 122:51]
  wire  sources_exuOutput_6_valid_differentFlag_2 = io_writeback_1_6_bits_uop_robIdx_flag ^
    stage2Redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  sources_exuOutput_6_valid_compare_2 = io_writeback_1_6_bits_uop_robIdx_value > stage2Redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _sources_exuOutput_6_valid_T_10 = sources_exuOutput_6_valid_differentFlag_2 ^
    sources_exuOutput_6_valid_compare_2; // @[CircularQueuePtr.scala 88:19]
  wire  _sources_exuOutput_6_valid_T_12 = stage2Redirect_valid & (sources_exuOutput_6_valid_flushItself_2 |
    _sources_exuOutput_6_valid_T_10); // @[Rob.scala 123:20]
  wire  _sources_exuOutput_6_valid_flushItself_T_15 = _sources_exuOutput_6_valid_flushItself_T_9 ==
    _exuRedirect_killedByOlder_flushItself_T_6; // @[CircularQueuePtr.scala 61:52]
  wire  sources_exuOutput_6_valid_flushItself_3 = redirectForExu_next_bits_rlevel &
    _sources_exuOutput_6_valid_flushItself_T_15; // @[Rob.scala 122:51]
  wire  sources_exuOutput_6_valid_differentFlag_3 = io_writeback_1_6_bits_uop_robIdx_flag ^
    redirectForExu_next_bits_rrobIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  sources_exuOutput_6_valid_compare_3 = io_writeback_1_6_bits_uop_robIdx_value >
    redirectForExu_next_bits_rrobIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _sources_exuOutput_6_valid_T_13 = sources_exuOutput_6_valid_differentFlag_3 ^
    sources_exuOutput_6_valid_compare_3; // @[CircularQueuePtr.scala 88:19]
  wire  _sources_exuOutput_6_valid_T_15 = redirectForExu_next_valid_REG & (sources_exuOutput_6_valid_flushItself_3 |
    _sources_exuOutput_6_valid_T_13); // @[Rob.scala 123:20]
  wire [1:0] _sources_exuOutput_6_valid_T_16 = {_sources_exuOutput_6_valid_T_15,_sources_exuOutput_6_valid_T_12}; // @[Rob.scala 126:90]
  wire  _sources_exuOutput_6_valid_T_17 = |_sources_exuOutput_6_valid_T_16; // @[Rob.scala 126:97]
  wire [5:0] _sources_exuOutput_7_valid_flushItself_T_9 = {io_writeback_1_7_bits_uop_robIdx_flag,
    io_writeback_1_7_bits_uop_robIdx_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _sources_exuOutput_7_valid_flushItself_T_11 = _sources_exuOutput_7_valid_flushItself_T_9 ==
    _exuRedirect_killedByOlder_flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  sources_exuOutput_7_valid_flushItself_2 = stage2Redirect_bits_level &
    _sources_exuOutput_7_valid_flushItself_T_11; // @[Rob.scala 122:51]
  wire  sources_exuOutput_7_valid_differentFlag_2 = io_writeback_1_7_bits_uop_robIdx_flag ^
    stage2Redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  sources_exuOutput_7_valid_compare_2 = io_writeback_1_7_bits_uop_robIdx_value > stage2Redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _sources_exuOutput_7_valid_T_10 = sources_exuOutput_7_valid_differentFlag_2 ^
    sources_exuOutput_7_valid_compare_2; // @[CircularQueuePtr.scala 88:19]
  wire  _sources_exuOutput_7_valid_T_12 = stage2Redirect_valid & (sources_exuOutput_7_valid_flushItself_2 |
    _sources_exuOutput_7_valid_T_10); // @[Rob.scala 123:20]
  wire  _sources_exuOutput_7_valid_flushItself_T_15 = _sources_exuOutput_7_valid_flushItself_T_9 ==
    _exuRedirect_killedByOlder_flushItself_T_6; // @[CircularQueuePtr.scala 61:52]
  wire  sources_exuOutput_7_valid_flushItself_3 = redirectForExu_next_bits_rlevel &
    _sources_exuOutput_7_valid_flushItself_T_15; // @[Rob.scala 122:51]
  wire  sources_exuOutput_7_valid_differentFlag_3 = io_writeback_1_7_bits_uop_robIdx_flag ^
    redirectForExu_next_bits_rrobIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  sources_exuOutput_7_valid_compare_3 = io_writeback_1_7_bits_uop_robIdx_value >
    redirectForExu_next_bits_rrobIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _sources_exuOutput_7_valid_T_13 = sources_exuOutput_7_valid_differentFlag_3 ^
    sources_exuOutput_7_valid_compare_3; // @[CircularQueuePtr.scala 88:19]
  wire  _sources_exuOutput_7_valid_T_15 = redirectForExu_next_valid_REG & (sources_exuOutput_7_valid_flushItself_3 |
    _sources_exuOutput_7_valid_T_13); // @[Rob.scala 123:20]
  wire [1:0] _sources_exuOutput_7_valid_T_16 = {_sources_exuOutput_7_valid_T_15,_sources_exuOutput_7_valid_T_12}; // @[Rob.scala 126:90]
  wire  _sources_exuOutput_7_valid_T_17 = |_sources_exuOutput_7_valid_T_16; // @[Rob.scala 126:97]
  wire [5:0] _sources_exuOutput_8_valid_flushItself_T_9 = {io_writeback_1_8_bits_uop_robIdx_flag,
    io_writeback_1_8_bits_uop_robIdx_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _sources_exuOutput_8_valid_flushItself_T_11 = _sources_exuOutput_8_valid_flushItself_T_9 ==
    _exuRedirect_killedByOlder_flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  sources_exuOutput_8_valid_flushItself_2 = stage2Redirect_bits_level &
    _sources_exuOutput_8_valid_flushItself_T_11; // @[Rob.scala 122:51]
  wire  sources_exuOutput_8_valid_differentFlag_2 = io_writeback_1_8_bits_uop_robIdx_flag ^
    stage2Redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  sources_exuOutput_8_valid_compare_2 = io_writeback_1_8_bits_uop_robIdx_value > stage2Redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _sources_exuOutput_8_valid_T_10 = sources_exuOutput_8_valid_differentFlag_2 ^
    sources_exuOutput_8_valid_compare_2; // @[CircularQueuePtr.scala 88:19]
  wire  _sources_exuOutput_8_valid_T_12 = stage2Redirect_valid & (sources_exuOutput_8_valid_flushItself_2 |
    _sources_exuOutput_8_valid_T_10); // @[Rob.scala 123:20]
  wire  _sources_exuOutput_8_valid_flushItself_T_15 = _sources_exuOutput_8_valid_flushItself_T_9 ==
    _exuRedirect_killedByOlder_flushItself_T_6; // @[CircularQueuePtr.scala 61:52]
  wire  sources_exuOutput_8_valid_flushItself_3 = redirectForExu_next_bits_rlevel &
    _sources_exuOutput_8_valid_flushItself_T_15; // @[Rob.scala 122:51]
  wire  sources_exuOutput_8_valid_differentFlag_3 = io_writeback_1_8_bits_uop_robIdx_flag ^
    redirectForExu_next_bits_rrobIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  sources_exuOutput_8_valid_compare_3 = io_writeback_1_8_bits_uop_robIdx_value >
    redirectForExu_next_bits_rrobIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _sources_exuOutput_8_valid_T_13 = sources_exuOutput_8_valid_differentFlag_3 ^
    sources_exuOutput_8_valid_compare_3; // @[CircularQueuePtr.scala 88:19]
  wire  _sources_exuOutput_8_valid_T_15 = redirectForExu_next_valid_REG & (sources_exuOutput_8_valid_flushItself_3 |
    _sources_exuOutput_8_valid_T_13); // @[Rob.scala 123:20]
  wire [1:0] _sources_exuOutput_8_valid_T_16 = {_sources_exuOutput_8_valid_T_15,_sources_exuOutput_8_valid_T_12}; // @[Rob.scala 126:90]
  wire  _sources_exuOutput_8_valid_T_17 = |_sources_exuOutput_8_valid_T_16; // @[Rob.scala 126:97]
  wire [5:0] _sources_exuOutput_9_valid_flushItself_T_9 = {io_writeback_1_9_bits_uop_robIdx_flag,
    io_writeback_1_9_bits_uop_robIdx_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _sources_exuOutput_9_valid_flushItself_T_11 = _sources_exuOutput_9_valid_flushItself_T_9 ==
    _exuRedirect_killedByOlder_flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  sources_exuOutput_9_valid_flushItself_2 = stage2Redirect_bits_level &
    _sources_exuOutput_9_valid_flushItself_T_11; // @[Rob.scala 122:51]
  wire  sources_exuOutput_9_valid_differentFlag_2 = io_writeback_1_9_bits_uop_robIdx_flag ^
    stage2Redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  sources_exuOutput_9_valid_compare_2 = io_writeback_1_9_bits_uop_robIdx_value > stage2Redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _sources_exuOutput_9_valid_T_10 = sources_exuOutput_9_valid_differentFlag_2 ^
    sources_exuOutput_9_valid_compare_2; // @[CircularQueuePtr.scala 88:19]
  wire  _sources_exuOutput_9_valid_T_12 = stage2Redirect_valid & (sources_exuOutput_9_valid_flushItself_2 |
    _sources_exuOutput_9_valid_T_10); // @[Rob.scala 123:20]
  wire  _sources_exuOutput_9_valid_flushItself_T_15 = _sources_exuOutput_9_valid_flushItself_T_9 ==
    _exuRedirect_killedByOlder_flushItself_T_6; // @[CircularQueuePtr.scala 61:52]
  wire  sources_exuOutput_9_valid_flushItself_3 = redirectForExu_next_bits_rlevel &
    _sources_exuOutput_9_valid_flushItself_T_15; // @[Rob.scala 122:51]
  wire  sources_exuOutput_9_valid_differentFlag_3 = io_writeback_1_9_bits_uop_robIdx_flag ^
    redirectForExu_next_bits_rrobIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  sources_exuOutput_9_valid_compare_3 = io_writeback_1_9_bits_uop_robIdx_value >
    redirectForExu_next_bits_rrobIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _sources_exuOutput_9_valid_T_13 = sources_exuOutput_9_valid_differentFlag_3 ^
    sources_exuOutput_9_valid_compare_3; // @[CircularQueuePtr.scala 88:19]
  wire  _sources_exuOutput_9_valid_T_15 = redirectForExu_next_valid_REG & (sources_exuOutput_9_valid_flushItself_3 |
    _sources_exuOutput_9_valid_T_13); // @[Rob.scala 123:20]
  wire [1:0] _sources_exuOutput_9_valid_T_16 = {_sources_exuOutput_9_valid_T_15,_sources_exuOutput_9_valid_T_12}; // @[Rob.scala 126:90]
  wire  _sources_exuOutput_9_valid_T_17 = |_sources_exuOutput_9_valid_T_16; // @[Rob.scala 126:97]
  wire [5:0] _sources_exuOutput_10_valid_flushItself_T_9 = {io_writeback_1_10_bits_uop_robIdx_flag,
    io_writeback_1_10_bits_uop_robIdx_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _sources_exuOutput_10_valid_flushItself_T_11 = _sources_exuOutput_10_valid_flushItself_T_9 ==
    _exuRedirect_killedByOlder_flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  sources_exuOutput_10_valid_flushItself_2 = stage2Redirect_bits_level &
    _sources_exuOutput_10_valid_flushItself_T_11; // @[Rob.scala 122:51]
  wire  sources_exuOutput_10_valid_differentFlag_2 = io_writeback_1_10_bits_uop_robIdx_flag ^
    stage2Redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  sources_exuOutput_10_valid_compare_2 = io_writeback_1_10_bits_uop_robIdx_value >
    stage2Redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _sources_exuOutput_10_valid_T_10 = sources_exuOutput_10_valid_differentFlag_2 ^
    sources_exuOutput_10_valid_compare_2; // @[CircularQueuePtr.scala 88:19]
  wire  _sources_exuOutput_10_valid_T_12 = stage2Redirect_valid & (sources_exuOutput_10_valid_flushItself_2 |
    _sources_exuOutput_10_valid_T_10); // @[Rob.scala 123:20]
  wire  _sources_exuOutput_10_valid_flushItself_T_15 = _sources_exuOutput_10_valid_flushItself_T_9 ==
    _exuRedirect_killedByOlder_flushItself_T_6; // @[CircularQueuePtr.scala 61:52]
  wire  sources_exuOutput_10_valid_flushItself_3 = redirectForExu_next_bits_rlevel &
    _sources_exuOutput_10_valid_flushItself_T_15; // @[Rob.scala 122:51]
  wire  sources_exuOutput_10_valid_differentFlag_3 = io_writeback_1_10_bits_uop_robIdx_flag ^
    redirectForExu_next_bits_rrobIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  sources_exuOutput_10_valid_compare_3 = io_writeback_1_10_bits_uop_robIdx_value >
    redirectForExu_next_bits_rrobIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _sources_exuOutput_10_valid_T_13 = sources_exuOutput_10_valid_differentFlag_3 ^
    sources_exuOutput_10_valid_compare_3; // @[CircularQueuePtr.scala 88:19]
  wire  _sources_exuOutput_10_valid_T_15 = redirectForExu_next_valid_REG & (sources_exuOutput_10_valid_flushItself_3 |
    _sources_exuOutput_10_valid_T_13); // @[Rob.scala 123:20]
  wire [1:0] _sources_exuOutput_10_valid_T_16 = {_sources_exuOutput_10_valid_T_15,_sources_exuOutput_10_valid_T_12}; // @[Rob.scala 126:90]
  wire  _sources_exuOutput_10_valid_T_17 = |_sources_exuOutput_10_valid_T_16; // @[Rob.scala 126:97]
  reg  sources_source_exuOutput_3_valid_REG; // @[CtrlBlock.scala 255:33]
  reg  sources_source_exuOutput_3_bits_REG_uop_cf_exceptionVec_2; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_3_bits_REG_uop_cf_exceptionVec_3; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_3_bits_REG_uop_cf_exceptionVec_8; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_3_bits_REG_uop_cf_exceptionVec_9; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_3_bits_REG_uop_cf_exceptionVec_11; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_3_bits_REG_uop_ctrl_flushPipe; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_3_bits_REG_uop_robIdx_flag; // @[CtrlBlock.scala 256:32]
  reg [4:0] sources_source_exuOutput_3_bits_REG_uop_robIdx_value; // @[CtrlBlock.scala 256:32]
  reg [4:0] sources_source_exuOutput_3_bits_REG_fflags; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_4_valid_REG; // @[CtrlBlock.scala 255:33]
  reg [4:0] sources_source_exuOutput_4_bits_REG_uop_robIdx_value; // @[CtrlBlock.scala 256:32]
  reg [4:0] sources_source_exuOutput_4_bits_REG_fflags; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_5_valid_REG; // @[CtrlBlock.scala 255:33]
  reg [4:0] sources_source_exuOutput_5_bits_REG_uop_robIdx_value; // @[CtrlBlock.scala 256:32]
  reg [4:0] sources_source_exuOutput_5_bits_REG_fflags; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_6_valid_REG; // @[CtrlBlock.scala 255:33]
  reg  sources_source_exuOutput_6_bits_REG_uop_cf_exceptionVec_4; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_6_bits_REG_uop_cf_exceptionVec_5; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_6_bits_REG_uop_cf_exceptionVec_13; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_6_bits_REG_uop_cf_trigger_backendHit_0; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_6_bits_REG_uop_cf_trigger_backendHit_1; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_6_bits_REG_uop_cf_trigger_backendHit_2; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_6_bits_REG_uop_cf_trigger_backendHit_3; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_6_bits_REG_uop_cf_trigger_backendHit_4; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_6_bits_REG_uop_cf_trigger_backendHit_5; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_6_bits_REG_uop_ctrl_flushPipe; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_6_bits_REG_uop_ctrl_replayInst; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_6_bits_REG_uop_robIdx_flag; // @[CtrlBlock.scala 256:32]
  reg [4:0] sources_source_exuOutput_6_bits_REG_uop_robIdx_value; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_7_valid_REG; // @[CtrlBlock.scala 255:33]
  reg  sources_source_exuOutput_7_bits_REG_uop_cf_exceptionVec_4; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_7_bits_REG_uop_cf_exceptionVec_5; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_7_bits_REG_uop_cf_exceptionVec_13; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_7_bits_REG_uop_cf_trigger_backendHit_0; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_7_bits_REG_uop_cf_trigger_backendHit_1; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_7_bits_REG_uop_cf_trigger_backendHit_2; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_7_bits_REG_uop_cf_trigger_backendHit_3; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_7_bits_REG_uop_cf_trigger_backendHit_4; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_7_bits_REG_uop_cf_trigger_backendHit_5; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_7_bits_REG_uop_ctrl_flushPipe; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_7_bits_REG_uop_ctrl_replayInst; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_7_bits_REG_uop_robIdx_flag; // @[CtrlBlock.scala 256:32]
  reg [4:0] sources_source_exuOutput_7_bits_REG_uop_robIdx_value; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_8_valid_REG; // @[CtrlBlock.scala 255:33]
  reg  sources_source_exuOutput_8_bits_REG_uop_cf_exceptionVec_4; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_8_bits_REG_uop_cf_exceptionVec_5; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_8_bits_REG_uop_cf_exceptionVec_6; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_8_bits_REG_uop_cf_exceptionVec_7; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_8_bits_REG_uop_cf_exceptionVec_13; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_8_bits_REG_uop_cf_exceptionVec_15; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_8_bits_REG_uop_cf_trigger_backendHit_0; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_8_bits_REG_uop_cf_trigger_backendHit_1; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_8_bits_REG_uop_cf_trigger_backendHit_2; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_8_bits_REG_uop_cf_trigger_backendHit_3; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_8_bits_REG_uop_cf_trigger_backendHit_4; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_8_bits_REG_uop_cf_trigger_backendHit_5; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_8_bits_REG_uop_robIdx_flag; // @[CtrlBlock.scala 256:32]
  reg [4:0] sources_source_exuOutput_8_bits_REG_uop_robIdx_value; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_9_valid_REG; // @[CtrlBlock.scala 255:33]
  reg  sources_source_exuOutput_9_bits_REG_uop_cf_exceptionVec_6; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_9_bits_REG_uop_cf_exceptionVec_7; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_9_bits_REG_uop_cf_exceptionVec_15; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_9_bits_REG_uop_cf_trigger_backendHit_0; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_9_bits_REG_uop_cf_trigger_backendHit_1; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_9_bits_REG_uop_cf_trigger_backendHit_4; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_9_bits_REG_uop_robIdx_flag; // @[CtrlBlock.scala 256:32]
  reg [4:0] sources_source_exuOutput_9_bits_REG_uop_robIdx_value; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_0_valid_REG_3; // @[CtrlBlock.scala 255:33]
  reg [4:0] sources_source_exuOutput_0_bits_REG_3_uop_robIdx_value; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_0_bits_REG_3_redirectValid; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_0_bits_REG_3_redirect_cfiUpdate_isMisPred; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_1_valid_REG_3; // @[CtrlBlock.scala 255:33]
  reg [4:0] sources_source_exuOutput_1_bits_REG_3_uop_robIdx_value; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_1_bits_REG_3_redirectValid; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_1_bits_REG_3_redirect_cfiUpdate_isMisPred; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_2_valid_REG_3; // @[CtrlBlock.scala 255:33]
  reg  sources_source_exuOutput_2_bits_REG_3_uop_cf_exceptionVec_4; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_2_bits_REG_3_uop_cf_exceptionVec_5; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_2_bits_REG_3_uop_cf_exceptionVec_13; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_2_bits_REG_3_uop_cf_trigger_backendHit_0; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_2_bits_REG_3_uop_cf_trigger_backendHit_1; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_2_bits_REG_3_uop_cf_trigger_backendHit_2; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_2_bits_REG_3_uop_cf_trigger_backendHit_3; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_2_bits_REG_3_uop_cf_trigger_backendHit_4; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_2_bits_REG_3_uop_cf_trigger_backendHit_5; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_2_bits_REG_3_uop_ctrl_flushPipe; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_2_bits_REG_3_uop_ctrl_replayInst; // @[CtrlBlock.scala 256:32]
  reg [4:0] sources_source_exuOutput_2_bits_REG_3_uop_robIdx_value; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_2_bits_REG_3_debug_isMMIO; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_3_valid_REG_3; // @[CtrlBlock.scala 255:33]
  reg  sources_source_exuOutput_3_bits_REG_3_uop_cf_exceptionVec_4; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_3_bits_REG_3_uop_cf_exceptionVec_5; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_3_bits_REG_3_uop_cf_exceptionVec_13; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_3_bits_REG_3_uop_cf_trigger_backendHit_0; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_3_bits_REG_3_uop_cf_trigger_backendHit_1; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_3_bits_REG_3_uop_cf_trigger_backendHit_2; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_3_bits_REG_3_uop_cf_trigger_backendHit_3; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_3_bits_REG_3_uop_cf_trigger_backendHit_4; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_3_bits_REG_3_uop_cf_trigger_backendHit_5; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_3_bits_REG_3_uop_ctrl_flushPipe; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_3_bits_REG_3_uop_ctrl_replayInst; // @[CtrlBlock.scala 256:32]
  reg [4:0] sources_source_exuOutput_3_bits_REG_3_uop_robIdx_value; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_3_bits_REG_3_debug_isMMIO; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_4_valid_REG_3; // @[CtrlBlock.scala 255:33]
  reg  sources_source_exuOutput_4_bits_REG_3_uop_cf_exceptionVec_2; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_4_bits_REG_3_uop_cf_exceptionVec_3; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_4_bits_REG_3_uop_cf_exceptionVec_8; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_4_bits_REG_3_uop_cf_exceptionVec_9; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_4_bits_REG_3_uop_cf_exceptionVec_11; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_4_bits_REG_3_uop_ctrl_flushPipe; // @[CtrlBlock.scala 256:32]
  reg [4:0] sources_source_exuOutput_4_bits_REG_3_uop_robIdx_value; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_4_bits_REG_3_redirectValid; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_4_bits_REG_3_redirect_cfiUpdate_isMisPred; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_4_bits_REG_3_debug_isPerfCnt; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_5_valid_REG_3; // @[CtrlBlock.scala 255:33]
  reg  sources_source_exuOutput_5_bits_REG_3_uop_cf_trigger_backendHit_0; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_5_bits_REG_3_uop_cf_trigger_backendHit_1; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_5_bits_REG_3_uop_cf_trigger_backendHit_2; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_5_bits_REG_3_uop_cf_trigger_backendHit_3; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_5_bits_REG_3_uop_cf_trigger_backendHit_4; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_5_bits_REG_3_uop_cf_trigger_backendHit_5; // @[CtrlBlock.scala 256:32]
  reg [4:0] sources_source_exuOutput_5_bits_REG_3_uop_robIdx_value; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_6_valid_REG_3; // @[CtrlBlock.scala 255:33]
  reg  sources_source_exuOutput_6_bits_REG_3_uop_cf_exceptionVec_2; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_6_bits_REG_3_uop_cf_exceptionVec_3; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_6_bits_REG_3_uop_cf_exceptionVec_8; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_6_bits_REG_3_uop_cf_exceptionVec_9; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_6_bits_REG_3_uop_cf_exceptionVec_11; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_6_bits_REG_3_uop_ctrl_flushPipe; // @[CtrlBlock.scala 256:32]
  reg [4:0] sources_source_exuOutput_6_bits_REG_3_uop_robIdx_value; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_6_bits_REG_3_redirectValid; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_6_bits_REG_3_redirect_cfiUpdate_isMisPred; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_6_bits_REG_3_debug_isPerfCnt; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_7_valid_REG_3; // @[CtrlBlock.scala 255:33]
  reg  sources_source_exuOutput_7_bits_REG_3_uop_cf_exceptionVec_4; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_7_bits_REG_3_uop_cf_exceptionVec_5; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_7_bits_REG_3_uop_cf_exceptionVec_6; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_7_bits_REG_3_uop_cf_exceptionVec_7; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_7_bits_REG_3_uop_cf_exceptionVec_13; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_7_bits_REG_3_uop_cf_exceptionVec_15; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_7_bits_REG_3_uop_cf_trigger_backendHit_0; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_7_bits_REG_3_uop_cf_trigger_backendHit_1; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_7_bits_REG_3_uop_cf_trigger_backendHit_2; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_7_bits_REG_3_uop_cf_trigger_backendHit_3; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_7_bits_REG_3_uop_cf_trigger_backendHit_4; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_7_bits_REG_3_uop_cf_trigger_backendHit_5; // @[CtrlBlock.scala 256:32]
  reg [4:0] sources_source_exuOutput_7_bits_REG_3_uop_robIdx_value; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_7_bits_REG_3_redirectValid; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_7_bits_REG_3_redirect_cfiUpdate_isMisPred; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_7_bits_REG_3_debug_isMMIO; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_7_bits_REG_3_debug_isPerfCnt; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_8_valid_REG_3; // @[CtrlBlock.scala 255:33]
  reg  sources_source_exuOutput_8_bits_REG_3_uop_cf_exceptionVec_4; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_8_bits_REG_3_uop_cf_exceptionVec_5; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_8_bits_REG_3_uop_cf_exceptionVec_6; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_8_bits_REG_3_uop_cf_exceptionVec_7; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_8_bits_REG_3_uop_cf_exceptionVec_13; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_8_bits_REG_3_uop_cf_exceptionVec_15; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_8_bits_REG_3_uop_cf_trigger_backendHit_0; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_8_bits_REG_3_uop_cf_trigger_backendHit_1; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_8_bits_REG_3_uop_cf_trigger_backendHit_2; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_8_bits_REG_3_uop_cf_trigger_backendHit_3; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_8_bits_REG_3_uop_cf_trigger_backendHit_4; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_8_bits_REG_3_uop_cf_trigger_backendHit_5; // @[CtrlBlock.scala 256:32]
  reg [4:0] sources_source_exuOutput_8_bits_REG_3_uop_robIdx_value; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_8_bits_REG_3_redirectValid; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_8_bits_REG_3_redirect_cfiUpdate_isMisPred; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_8_bits_REG_3_debug_isMMIO; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_8_bits_REG_3_debug_isPerfCnt; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_9_valid_REG_3; // @[CtrlBlock.scala 255:33]
  reg [4:0] sources_source_exuOutput_9_bits_REG_3_uop_robIdx_value; // @[CtrlBlock.scala 256:32]
  reg  sources_source_exuOutput_10_valid_REG_3; // @[CtrlBlock.scala 255:33]
  reg [4:0] sources_source_exuOutput_10_bits_REG_3_uop_robIdx_value; // @[CtrlBlock.scala 256:32]
  reg [2:0] io_robio_toCSR_perfinfo_retiredInstr_REG; // @[CtrlBlock.scala 571:50]
  reg  pfevent_io_distribute_csr_REG_wvalid; // @[CtrlBlock.scala 586:39]
  reg [11:0] pfevent_io_distribute_csr_REG_waddr; // @[CtrlBlock.scala 586:39]
  reg [63:0] pfevent_io_distribute_csr_REG_wdata; // @[CtrlBlock.scala 586:39]
  reg [5:0] io_perf_0_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg [5:0] io_perf_0_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  reg [5:0] io_perf_1_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg [5:0] io_perf_1_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  reg [5:0] io_perf_2_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg [5:0] io_perf_2_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  reg [5:0] io_perf_3_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg [5:0] io_perf_3_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  reg [5:0] io_perf_4_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg [5:0] io_perf_4_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  reg [5:0] io_perf_5_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg [5:0] io_perf_5_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  reg [5:0] io_perf_6_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg [5:0] io_perf_6_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  reg [5:0] io_perf_7_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg [5:0] io_perf_7_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  Rob rob ( // @[CtrlBlock.scala 173:23]
    .clock(rob_clock),
    .reset(rob_reset),
    .io_hartId(rob_io_hartId),
    .io_redirect_valid(rob_io_redirect_valid),
    .io_redirect_bits_robIdx_flag(rob_io_redirect_bits_robIdx_flag),
    .io_redirect_bits_robIdx_value(rob_io_redirect_bits_robIdx_value),
    .io_redirect_bits_level(rob_io_redirect_bits_level),
    .io_enq_canAccept(rob_io_enq_canAccept),
    .io_enq_isEmpty(rob_io_enq_isEmpty),
    .io_enq_needAlloc_0(rob_io_enq_needAlloc_0),
    .io_enq_req_0_valid(rob_io_enq_req_0_valid),
    .io_enq_req_0_bits_cf_exceptionVec_1(rob_io_enq_req_0_bits_cf_exceptionVec_1),
    .io_enq_req_0_bits_cf_exceptionVec_2(rob_io_enq_req_0_bits_cf_exceptionVec_2),
    .io_enq_req_0_bits_cf_exceptionVec_12(rob_io_enq_req_0_bits_cf_exceptionVec_12),
    .io_enq_req_0_bits_cf_trigger_frontendHit_0(rob_io_enq_req_0_bits_cf_trigger_frontendHit_0),
    .io_enq_req_0_bits_cf_trigger_frontendHit_1(rob_io_enq_req_0_bits_cf_trigger_frontendHit_1),
    .io_enq_req_0_bits_cf_trigger_frontendHit_2(rob_io_enq_req_0_bits_cf_trigger_frontendHit_2),
    .io_enq_req_0_bits_cf_trigger_frontendHit_3(rob_io_enq_req_0_bits_cf_trigger_frontendHit_3),
    .io_enq_req_0_bits_cf_pd_isRVC(rob_io_enq_req_0_bits_cf_pd_isRVC),
    .io_enq_req_0_bits_cf_crossPageIPFFix(rob_io_enq_req_0_bits_cf_crossPageIPFFix),
    .io_enq_req_0_bits_cf_loadWaitBit(rob_io_enq_req_0_bits_cf_loadWaitBit),
    .io_enq_req_0_bits_cf_ftqPtr_flag(rob_io_enq_req_0_bits_cf_ftqPtr_flag),
    .io_enq_req_0_bits_cf_ftqPtr_value(rob_io_enq_req_0_bits_cf_ftqPtr_value),
    .io_enq_req_0_bits_cf_ftqOffset(rob_io_enq_req_0_bits_cf_ftqOffset),
    .io_enq_req_0_bits_ctrl_ldest(rob_io_enq_req_0_bits_ctrl_ldest),
    .io_enq_req_0_bits_ctrl_fuType(rob_io_enq_req_0_bits_ctrl_fuType),
    .io_enq_req_0_bits_ctrl_fuOpType(rob_io_enq_req_0_bits_ctrl_fuOpType),
    .io_enq_req_0_bits_ctrl_rfWen(rob_io_enq_req_0_bits_ctrl_rfWen),
    .io_enq_req_0_bits_ctrl_fpWen(rob_io_enq_req_0_bits_ctrl_fpWen),
    .io_enq_req_0_bits_ctrl_isXSTrap(rob_io_enq_req_0_bits_ctrl_isXSTrap),
    .io_enq_req_0_bits_ctrl_noSpecExec(rob_io_enq_req_0_bits_ctrl_noSpecExec),
    .io_enq_req_0_bits_ctrl_blockBackward(rob_io_enq_req_0_bits_ctrl_blockBackward),
    .io_enq_req_0_bits_ctrl_flushPipe(rob_io_enq_req_0_bits_ctrl_flushPipe),
    .io_enq_req_0_bits_ctrl_commitType(rob_io_enq_req_0_bits_ctrl_commitType),
    .io_enq_req_0_bits_ctrl_fpu_wflags(rob_io_enq_req_0_bits_ctrl_fpu_wflags),
    .io_enq_req_0_bits_ctrl_isMove(rob_io_enq_req_0_bits_ctrl_isMove),
    .io_enq_req_0_bits_ctrl_singleStep(rob_io_enq_req_0_bits_ctrl_singleStep),
    .io_enq_req_0_bits_pdest(rob_io_enq_req_0_bits_pdest),
    .io_enq_req_0_bits_old_pdest(rob_io_enq_req_0_bits_old_pdest),
    .io_enq_req_0_bits_robIdx_flag(rob_io_enq_req_0_bits_robIdx_flag),
    .io_enq_req_0_bits_robIdx_value(rob_io_enq_req_0_bits_robIdx_value),
    .io_enq_req_0_bits_eliminatedMove(rob_io_enq_req_0_bits_eliminatedMove),
    .io_enq_req_1_valid(rob_io_enq_req_1_valid),
    .io_enq_req_1_bits_cf_exceptionVec_1(rob_io_enq_req_1_bits_cf_exceptionVec_1),
    .io_enq_req_1_bits_cf_exceptionVec_2(rob_io_enq_req_1_bits_cf_exceptionVec_2),
    .io_enq_req_1_bits_cf_exceptionVec_12(rob_io_enq_req_1_bits_cf_exceptionVec_12),
    .io_enq_req_1_bits_cf_trigger_frontendHit_0(rob_io_enq_req_1_bits_cf_trigger_frontendHit_0),
    .io_enq_req_1_bits_cf_trigger_frontendHit_1(rob_io_enq_req_1_bits_cf_trigger_frontendHit_1),
    .io_enq_req_1_bits_cf_trigger_frontendHit_2(rob_io_enq_req_1_bits_cf_trigger_frontendHit_2),
    .io_enq_req_1_bits_cf_trigger_frontendHit_3(rob_io_enq_req_1_bits_cf_trigger_frontendHit_3),
    .io_enq_req_1_bits_cf_pd_isRVC(rob_io_enq_req_1_bits_cf_pd_isRVC),
    .io_enq_req_1_bits_cf_crossPageIPFFix(rob_io_enq_req_1_bits_cf_crossPageIPFFix),
    .io_enq_req_1_bits_cf_loadWaitBit(rob_io_enq_req_1_bits_cf_loadWaitBit),
    .io_enq_req_1_bits_cf_ftqPtr_flag(rob_io_enq_req_1_bits_cf_ftqPtr_flag),
    .io_enq_req_1_bits_cf_ftqPtr_value(rob_io_enq_req_1_bits_cf_ftqPtr_value),
    .io_enq_req_1_bits_cf_ftqOffset(rob_io_enq_req_1_bits_cf_ftqOffset),
    .io_enq_req_1_bits_ctrl_ldest(rob_io_enq_req_1_bits_ctrl_ldest),
    .io_enq_req_1_bits_ctrl_fuType(rob_io_enq_req_1_bits_ctrl_fuType),
    .io_enq_req_1_bits_ctrl_fuOpType(rob_io_enq_req_1_bits_ctrl_fuOpType),
    .io_enq_req_1_bits_ctrl_rfWen(rob_io_enq_req_1_bits_ctrl_rfWen),
    .io_enq_req_1_bits_ctrl_fpWen(rob_io_enq_req_1_bits_ctrl_fpWen),
    .io_enq_req_1_bits_ctrl_isXSTrap(rob_io_enq_req_1_bits_ctrl_isXSTrap),
    .io_enq_req_1_bits_ctrl_noSpecExec(rob_io_enq_req_1_bits_ctrl_noSpecExec),
    .io_enq_req_1_bits_ctrl_blockBackward(rob_io_enq_req_1_bits_ctrl_blockBackward),
    .io_enq_req_1_bits_ctrl_flushPipe(rob_io_enq_req_1_bits_ctrl_flushPipe),
    .io_enq_req_1_bits_ctrl_commitType(rob_io_enq_req_1_bits_ctrl_commitType),
    .io_enq_req_1_bits_ctrl_fpu_wflags(rob_io_enq_req_1_bits_ctrl_fpu_wflags),
    .io_enq_req_1_bits_ctrl_isMove(rob_io_enq_req_1_bits_ctrl_isMove),
    .io_enq_req_1_bits_ctrl_singleStep(rob_io_enq_req_1_bits_ctrl_singleStep),
    .io_enq_req_1_bits_pdest(rob_io_enq_req_1_bits_pdest),
    .io_enq_req_1_bits_old_pdest(rob_io_enq_req_1_bits_old_pdest),
    .io_enq_req_1_bits_robIdx_flag(rob_io_enq_req_1_bits_robIdx_flag),
    .io_enq_req_1_bits_robIdx_value(rob_io_enq_req_1_bits_robIdx_value),
    .io_enq_req_1_bits_eliminatedMove(rob_io_enq_req_1_bits_eliminatedMove),
    .io_flushOut_valid(rob_io_flushOut_valid),
    .io_flushOut_bits_robIdx_flag(rob_io_flushOut_bits_robIdx_flag),
    .io_flushOut_bits_robIdx_value(rob_io_flushOut_bits_robIdx_value),
    .io_flushOut_bits_ftqIdx_flag(rob_io_flushOut_bits_ftqIdx_flag),
    .io_flushOut_bits_ftqIdx_value(rob_io_flushOut_bits_ftqIdx_value),
    .io_flushOut_bits_ftqOffset(rob_io_flushOut_bits_ftqOffset),
    .io_flushOut_bits_level(rob_io_flushOut_bits_level),
    .io_exception_valid(rob_io_exception_valid),
    .io_exception_bits_uop_cf_exceptionVec_0(rob_io_exception_bits_uop_cf_exceptionVec_0),
    .io_exception_bits_uop_cf_exceptionVec_1(rob_io_exception_bits_uop_cf_exceptionVec_1),
    .io_exception_bits_uop_cf_exceptionVec_2(rob_io_exception_bits_uop_cf_exceptionVec_2),
    .io_exception_bits_uop_cf_exceptionVec_3(rob_io_exception_bits_uop_cf_exceptionVec_3),
    .io_exception_bits_uop_cf_exceptionVec_4(rob_io_exception_bits_uop_cf_exceptionVec_4),
    .io_exception_bits_uop_cf_exceptionVec_5(rob_io_exception_bits_uop_cf_exceptionVec_5),
    .io_exception_bits_uop_cf_exceptionVec_6(rob_io_exception_bits_uop_cf_exceptionVec_6),
    .io_exception_bits_uop_cf_exceptionVec_7(rob_io_exception_bits_uop_cf_exceptionVec_7),
    .io_exception_bits_uop_cf_exceptionVec_8(rob_io_exception_bits_uop_cf_exceptionVec_8),
    .io_exception_bits_uop_cf_exceptionVec_9(rob_io_exception_bits_uop_cf_exceptionVec_9),
    .io_exception_bits_uop_cf_exceptionVec_11(rob_io_exception_bits_uop_cf_exceptionVec_11),
    .io_exception_bits_uop_cf_exceptionVec_12(rob_io_exception_bits_uop_cf_exceptionVec_12),
    .io_exception_bits_uop_cf_exceptionVec_13(rob_io_exception_bits_uop_cf_exceptionVec_13),
    .io_exception_bits_uop_cf_exceptionVec_15(rob_io_exception_bits_uop_cf_exceptionVec_15),
    .io_exception_bits_uop_cf_trigger_frontendHit_0(rob_io_exception_bits_uop_cf_trigger_frontendHit_0),
    .io_exception_bits_uop_cf_trigger_frontendHit_1(rob_io_exception_bits_uop_cf_trigger_frontendHit_1),
    .io_exception_bits_uop_cf_trigger_frontendHit_2(rob_io_exception_bits_uop_cf_trigger_frontendHit_2),
    .io_exception_bits_uop_cf_trigger_frontendHit_3(rob_io_exception_bits_uop_cf_trigger_frontendHit_3),
    .io_exception_bits_uop_cf_trigger_backendHit_0(rob_io_exception_bits_uop_cf_trigger_backendHit_0),
    .io_exception_bits_uop_cf_trigger_backendHit_1(rob_io_exception_bits_uop_cf_trigger_backendHit_1),
    .io_exception_bits_uop_cf_trigger_backendHit_2(rob_io_exception_bits_uop_cf_trigger_backendHit_2),
    .io_exception_bits_uop_cf_trigger_backendHit_3(rob_io_exception_bits_uop_cf_trigger_backendHit_3),
    .io_exception_bits_uop_cf_trigger_backendHit_4(rob_io_exception_bits_uop_cf_trigger_backendHit_4),
    .io_exception_bits_uop_cf_trigger_backendHit_5(rob_io_exception_bits_uop_cf_trigger_backendHit_5),
    .io_exception_bits_uop_cf_crossPageIPFFix(rob_io_exception_bits_uop_cf_crossPageIPFFix),
    .io_exception_bits_uop_ctrl_commitType(rob_io_exception_bits_uop_ctrl_commitType),
    .io_exception_bits_uop_ctrl_singleStep(rob_io_exception_bits_uop_ctrl_singleStep),
    .io_exception_bits_isInterrupt(rob_io_exception_bits_isInterrupt),
    .io_writeback_1_0_valid(rob_io_writeback_1_0_valid),
    .io_writeback_1_0_bits_uop_robIdx_value(rob_io_writeback_1_0_bits_uop_robIdx_value),
    .io_writeback_1_0_bits_redirectValid(rob_io_writeback_1_0_bits_redirectValid),
    .io_writeback_1_0_bits_redirect_cfiUpdate_isMisPred(rob_io_writeback_1_0_bits_redirect_cfiUpdate_isMisPred),
    .io_writeback_1_1_valid(rob_io_writeback_1_1_valid),
    .io_writeback_1_1_bits_uop_robIdx_value(rob_io_writeback_1_1_bits_uop_robIdx_value),
    .io_writeback_1_1_bits_redirectValid(rob_io_writeback_1_1_bits_redirectValid),
    .io_writeback_1_1_bits_redirect_cfiUpdate_isMisPred(rob_io_writeback_1_1_bits_redirect_cfiUpdate_isMisPred),
    .io_writeback_1_2_valid(rob_io_writeback_1_2_valid),
    .io_writeback_1_2_bits_uop_cf_exceptionVec_4(rob_io_writeback_1_2_bits_uop_cf_exceptionVec_4),
    .io_writeback_1_2_bits_uop_cf_exceptionVec_5(rob_io_writeback_1_2_bits_uop_cf_exceptionVec_5),
    .io_writeback_1_2_bits_uop_cf_exceptionVec_13(rob_io_writeback_1_2_bits_uop_cf_exceptionVec_13),
    .io_writeback_1_2_bits_uop_cf_trigger_backendHit_0(rob_io_writeback_1_2_bits_uop_cf_trigger_backendHit_0),
    .io_writeback_1_2_bits_uop_cf_trigger_backendHit_1(rob_io_writeback_1_2_bits_uop_cf_trigger_backendHit_1),
    .io_writeback_1_2_bits_uop_cf_trigger_backendHit_2(rob_io_writeback_1_2_bits_uop_cf_trigger_backendHit_2),
    .io_writeback_1_2_bits_uop_cf_trigger_backendHit_3(rob_io_writeback_1_2_bits_uop_cf_trigger_backendHit_3),
    .io_writeback_1_2_bits_uop_cf_trigger_backendHit_4(rob_io_writeback_1_2_bits_uop_cf_trigger_backendHit_4),
    .io_writeback_1_2_bits_uop_cf_trigger_backendHit_5(rob_io_writeback_1_2_bits_uop_cf_trigger_backendHit_5),
    .io_writeback_1_2_bits_uop_ctrl_flushPipe(rob_io_writeback_1_2_bits_uop_ctrl_flushPipe),
    .io_writeback_1_2_bits_uop_ctrl_replayInst(rob_io_writeback_1_2_bits_uop_ctrl_replayInst),
    .io_writeback_1_2_bits_uop_robIdx_value(rob_io_writeback_1_2_bits_uop_robIdx_value),
    .io_writeback_1_2_bits_debug_isMMIO(rob_io_writeback_1_2_bits_debug_isMMIO),
    .io_writeback_1_3_valid(rob_io_writeback_1_3_valid),
    .io_writeback_1_3_bits_uop_cf_exceptionVec_4(rob_io_writeback_1_3_bits_uop_cf_exceptionVec_4),
    .io_writeback_1_3_bits_uop_cf_exceptionVec_5(rob_io_writeback_1_3_bits_uop_cf_exceptionVec_5),
    .io_writeback_1_3_bits_uop_cf_exceptionVec_13(rob_io_writeback_1_3_bits_uop_cf_exceptionVec_13),
    .io_writeback_1_3_bits_uop_cf_trigger_backendHit_0(rob_io_writeback_1_3_bits_uop_cf_trigger_backendHit_0),
    .io_writeback_1_3_bits_uop_cf_trigger_backendHit_1(rob_io_writeback_1_3_bits_uop_cf_trigger_backendHit_1),
    .io_writeback_1_3_bits_uop_cf_trigger_backendHit_2(rob_io_writeback_1_3_bits_uop_cf_trigger_backendHit_2),
    .io_writeback_1_3_bits_uop_cf_trigger_backendHit_3(rob_io_writeback_1_3_bits_uop_cf_trigger_backendHit_3),
    .io_writeback_1_3_bits_uop_cf_trigger_backendHit_4(rob_io_writeback_1_3_bits_uop_cf_trigger_backendHit_4),
    .io_writeback_1_3_bits_uop_cf_trigger_backendHit_5(rob_io_writeback_1_3_bits_uop_cf_trigger_backendHit_5),
    .io_writeback_1_3_bits_uop_ctrl_flushPipe(rob_io_writeback_1_3_bits_uop_ctrl_flushPipe),
    .io_writeback_1_3_bits_uop_ctrl_replayInst(rob_io_writeback_1_3_bits_uop_ctrl_replayInst),
    .io_writeback_1_3_bits_uop_robIdx_value(rob_io_writeback_1_3_bits_uop_robIdx_value),
    .io_writeback_1_3_bits_debug_isMMIO(rob_io_writeback_1_3_bits_debug_isMMIO),
    .io_writeback_1_4_valid(rob_io_writeback_1_4_valid),
    .io_writeback_1_4_bits_uop_cf_exceptionVec_2(rob_io_writeback_1_4_bits_uop_cf_exceptionVec_2),
    .io_writeback_1_4_bits_uop_cf_exceptionVec_3(rob_io_writeback_1_4_bits_uop_cf_exceptionVec_3),
    .io_writeback_1_4_bits_uop_cf_exceptionVec_8(rob_io_writeback_1_4_bits_uop_cf_exceptionVec_8),
    .io_writeback_1_4_bits_uop_cf_exceptionVec_9(rob_io_writeback_1_4_bits_uop_cf_exceptionVec_9),
    .io_writeback_1_4_bits_uop_cf_exceptionVec_11(rob_io_writeback_1_4_bits_uop_cf_exceptionVec_11),
    .io_writeback_1_4_bits_uop_ctrl_flushPipe(rob_io_writeback_1_4_bits_uop_ctrl_flushPipe),
    .io_writeback_1_4_bits_uop_robIdx_value(rob_io_writeback_1_4_bits_uop_robIdx_value),
    .io_writeback_1_4_bits_redirectValid(rob_io_writeback_1_4_bits_redirectValid),
    .io_writeback_1_4_bits_redirect_cfiUpdate_isMisPred(rob_io_writeback_1_4_bits_redirect_cfiUpdate_isMisPred),
    .io_writeback_1_4_bits_debug_isPerfCnt(rob_io_writeback_1_4_bits_debug_isPerfCnt),
    .io_writeback_1_5_valid(rob_io_writeback_1_5_valid),
    .io_writeback_1_5_bits_uop_cf_trigger_backendHit_0(rob_io_writeback_1_5_bits_uop_cf_trigger_backendHit_0),
    .io_writeback_1_5_bits_uop_cf_trigger_backendHit_1(rob_io_writeback_1_5_bits_uop_cf_trigger_backendHit_1),
    .io_writeback_1_5_bits_uop_cf_trigger_backendHit_2(rob_io_writeback_1_5_bits_uop_cf_trigger_backendHit_2),
    .io_writeback_1_5_bits_uop_cf_trigger_backendHit_3(rob_io_writeback_1_5_bits_uop_cf_trigger_backendHit_3),
    .io_writeback_1_5_bits_uop_cf_trigger_backendHit_4(rob_io_writeback_1_5_bits_uop_cf_trigger_backendHit_4),
    .io_writeback_1_5_bits_uop_cf_trigger_backendHit_5(rob_io_writeback_1_5_bits_uop_cf_trigger_backendHit_5),
    .io_writeback_1_5_bits_uop_robIdx_value(rob_io_writeback_1_5_bits_uop_robIdx_value),
    .io_writeback_1_6_valid(rob_io_writeback_1_6_valid),
    .io_writeback_1_6_bits_uop_cf_exceptionVec_2(rob_io_writeback_1_6_bits_uop_cf_exceptionVec_2),
    .io_writeback_1_6_bits_uop_cf_exceptionVec_3(rob_io_writeback_1_6_bits_uop_cf_exceptionVec_3),
    .io_writeback_1_6_bits_uop_cf_exceptionVec_8(rob_io_writeback_1_6_bits_uop_cf_exceptionVec_8),
    .io_writeback_1_6_bits_uop_cf_exceptionVec_9(rob_io_writeback_1_6_bits_uop_cf_exceptionVec_9),
    .io_writeback_1_6_bits_uop_cf_exceptionVec_11(rob_io_writeback_1_6_bits_uop_cf_exceptionVec_11),
    .io_writeback_1_6_bits_uop_ctrl_flushPipe(rob_io_writeback_1_6_bits_uop_ctrl_flushPipe),
    .io_writeback_1_6_bits_uop_robIdx_value(rob_io_writeback_1_6_bits_uop_robIdx_value),
    .io_writeback_1_6_bits_redirectValid(rob_io_writeback_1_6_bits_redirectValid),
    .io_writeback_1_6_bits_redirect_cfiUpdate_isMisPred(rob_io_writeback_1_6_bits_redirect_cfiUpdate_isMisPred),
    .io_writeback_1_6_bits_debug_isPerfCnt(rob_io_writeback_1_6_bits_debug_isPerfCnt),
    .io_writeback_1_7_valid(rob_io_writeback_1_7_valid),
    .io_writeback_1_7_bits_uop_cf_exceptionVec_4(rob_io_writeback_1_7_bits_uop_cf_exceptionVec_4),
    .io_writeback_1_7_bits_uop_cf_exceptionVec_5(rob_io_writeback_1_7_bits_uop_cf_exceptionVec_5),
    .io_writeback_1_7_bits_uop_cf_exceptionVec_6(rob_io_writeback_1_7_bits_uop_cf_exceptionVec_6),
    .io_writeback_1_7_bits_uop_cf_exceptionVec_7(rob_io_writeback_1_7_bits_uop_cf_exceptionVec_7),
    .io_writeback_1_7_bits_uop_cf_exceptionVec_13(rob_io_writeback_1_7_bits_uop_cf_exceptionVec_13),
    .io_writeback_1_7_bits_uop_cf_exceptionVec_15(rob_io_writeback_1_7_bits_uop_cf_exceptionVec_15),
    .io_writeback_1_7_bits_uop_cf_trigger_backendHit_0(rob_io_writeback_1_7_bits_uop_cf_trigger_backendHit_0),
    .io_writeback_1_7_bits_uop_cf_trigger_backendHit_1(rob_io_writeback_1_7_bits_uop_cf_trigger_backendHit_1),
    .io_writeback_1_7_bits_uop_cf_trigger_backendHit_2(rob_io_writeback_1_7_bits_uop_cf_trigger_backendHit_2),
    .io_writeback_1_7_bits_uop_cf_trigger_backendHit_3(rob_io_writeback_1_7_bits_uop_cf_trigger_backendHit_3),
    .io_writeback_1_7_bits_uop_cf_trigger_backendHit_4(rob_io_writeback_1_7_bits_uop_cf_trigger_backendHit_4),
    .io_writeback_1_7_bits_uop_cf_trigger_backendHit_5(rob_io_writeback_1_7_bits_uop_cf_trigger_backendHit_5),
    .io_writeback_1_7_bits_uop_robIdx_value(rob_io_writeback_1_7_bits_uop_robIdx_value),
    .io_writeback_1_7_bits_redirectValid(rob_io_writeback_1_7_bits_redirectValid),
    .io_writeback_1_7_bits_redirect_cfiUpdate_isMisPred(rob_io_writeback_1_7_bits_redirect_cfiUpdate_isMisPred),
    .io_writeback_1_7_bits_debug_isMMIO(rob_io_writeback_1_7_bits_debug_isMMIO),
    .io_writeback_1_7_bits_debug_isPerfCnt(rob_io_writeback_1_7_bits_debug_isPerfCnt),
    .io_writeback_1_8_valid(rob_io_writeback_1_8_valid),
    .io_writeback_1_8_bits_uop_cf_exceptionVec_4(rob_io_writeback_1_8_bits_uop_cf_exceptionVec_4),
    .io_writeback_1_8_bits_uop_cf_exceptionVec_5(rob_io_writeback_1_8_bits_uop_cf_exceptionVec_5),
    .io_writeback_1_8_bits_uop_cf_exceptionVec_6(rob_io_writeback_1_8_bits_uop_cf_exceptionVec_6),
    .io_writeback_1_8_bits_uop_cf_exceptionVec_7(rob_io_writeback_1_8_bits_uop_cf_exceptionVec_7),
    .io_writeback_1_8_bits_uop_cf_exceptionVec_13(rob_io_writeback_1_8_bits_uop_cf_exceptionVec_13),
    .io_writeback_1_8_bits_uop_cf_exceptionVec_15(rob_io_writeback_1_8_bits_uop_cf_exceptionVec_15),
    .io_writeback_1_8_bits_uop_cf_trigger_backendHit_0(rob_io_writeback_1_8_bits_uop_cf_trigger_backendHit_0),
    .io_writeback_1_8_bits_uop_cf_trigger_backendHit_1(rob_io_writeback_1_8_bits_uop_cf_trigger_backendHit_1),
    .io_writeback_1_8_bits_uop_cf_trigger_backendHit_2(rob_io_writeback_1_8_bits_uop_cf_trigger_backendHit_2),
    .io_writeback_1_8_bits_uop_cf_trigger_backendHit_3(rob_io_writeback_1_8_bits_uop_cf_trigger_backendHit_3),
    .io_writeback_1_8_bits_uop_cf_trigger_backendHit_4(rob_io_writeback_1_8_bits_uop_cf_trigger_backendHit_4),
    .io_writeback_1_8_bits_uop_cf_trigger_backendHit_5(rob_io_writeback_1_8_bits_uop_cf_trigger_backendHit_5),
    .io_writeback_1_8_bits_uop_robIdx_value(rob_io_writeback_1_8_bits_uop_robIdx_value),
    .io_writeback_1_8_bits_redirectValid(rob_io_writeback_1_8_bits_redirectValid),
    .io_writeback_1_8_bits_redirect_cfiUpdate_isMisPred(rob_io_writeback_1_8_bits_redirect_cfiUpdate_isMisPred),
    .io_writeback_1_8_bits_debug_isMMIO(rob_io_writeback_1_8_bits_debug_isMMIO),
    .io_writeback_1_8_bits_debug_isPerfCnt(rob_io_writeback_1_8_bits_debug_isPerfCnt),
    .io_writeback_1_9_valid(rob_io_writeback_1_9_valid),
    .io_writeback_1_9_bits_uop_robIdx_value(rob_io_writeback_1_9_bits_uop_robIdx_value),
    .io_writeback_1_10_valid(rob_io_writeback_1_10_valid),
    .io_writeback_1_10_bits_uop_robIdx_value(rob_io_writeback_1_10_bits_uop_robIdx_value),
    .io_writeback_0_3_valid(rob_io_writeback_0_3_valid),
    .io_writeback_0_3_bits_uop_cf_exceptionVec_2(rob_io_writeback_0_3_bits_uop_cf_exceptionVec_2),
    .io_writeback_0_3_bits_uop_cf_exceptionVec_3(rob_io_writeback_0_3_bits_uop_cf_exceptionVec_3),
    .io_writeback_0_3_bits_uop_cf_exceptionVec_8(rob_io_writeback_0_3_bits_uop_cf_exceptionVec_8),
    .io_writeback_0_3_bits_uop_cf_exceptionVec_9(rob_io_writeback_0_3_bits_uop_cf_exceptionVec_9),
    .io_writeback_0_3_bits_uop_cf_exceptionVec_11(rob_io_writeback_0_3_bits_uop_cf_exceptionVec_11),
    .io_writeback_0_3_bits_uop_ctrl_flushPipe(rob_io_writeback_0_3_bits_uop_ctrl_flushPipe),
    .io_writeback_0_3_bits_uop_robIdx_flag(rob_io_writeback_0_3_bits_uop_robIdx_flag),
    .io_writeback_0_3_bits_uop_robIdx_value(rob_io_writeback_0_3_bits_uop_robIdx_value),
    .io_writeback_0_3_bits_fflags(rob_io_writeback_0_3_bits_fflags),
    .io_writeback_0_4_valid(rob_io_writeback_0_4_valid),
    .io_writeback_0_4_bits_uop_robIdx_value(rob_io_writeback_0_4_bits_uop_robIdx_value),
    .io_writeback_0_4_bits_fflags(rob_io_writeback_0_4_bits_fflags),
    .io_writeback_0_5_valid(rob_io_writeback_0_5_valid),
    .io_writeback_0_5_bits_uop_robIdx_value(rob_io_writeback_0_5_bits_uop_robIdx_value),
    .io_writeback_0_5_bits_fflags(rob_io_writeback_0_5_bits_fflags),
    .io_writeback_0_6_valid(rob_io_writeback_0_6_valid),
    .io_writeback_0_6_bits_uop_cf_exceptionVec_4(rob_io_writeback_0_6_bits_uop_cf_exceptionVec_4),
    .io_writeback_0_6_bits_uop_cf_exceptionVec_5(rob_io_writeback_0_6_bits_uop_cf_exceptionVec_5),
    .io_writeback_0_6_bits_uop_cf_exceptionVec_13(rob_io_writeback_0_6_bits_uop_cf_exceptionVec_13),
    .io_writeback_0_6_bits_uop_cf_trigger_backendHit_0(rob_io_writeback_0_6_bits_uop_cf_trigger_backendHit_0),
    .io_writeback_0_6_bits_uop_cf_trigger_backendHit_1(rob_io_writeback_0_6_bits_uop_cf_trigger_backendHit_1),
    .io_writeback_0_6_bits_uop_cf_trigger_backendHit_2(rob_io_writeback_0_6_bits_uop_cf_trigger_backendHit_2),
    .io_writeback_0_6_bits_uop_cf_trigger_backendHit_3(rob_io_writeback_0_6_bits_uop_cf_trigger_backendHit_3),
    .io_writeback_0_6_bits_uop_cf_trigger_backendHit_4(rob_io_writeback_0_6_bits_uop_cf_trigger_backendHit_4),
    .io_writeback_0_6_bits_uop_cf_trigger_backendHit_5(rob_io_writeback_0_6_bits_uop_cf_trigger_backendHit_5),
    .io_writeback_0_6_bits_uop_ctrl_flushPipe(rob_io_writeback_0_6_bits_uop_ctrl_flushPipe),
    .io_writeback_0_6_bits_uop_ctrl_replayInst(rob_io_writeback_0_6_bits_uop_ctrl_replayInst),
    .io_writeback_0_6_bits_uop_robIdx_flag(rob_io_writeback_0_6_bits_uop_robIdx_flag),
    .io_writeback_0_6_bits_uop_robIdx_value(rob_io_writeback_0_6_bits_uop_robIdx_value),
    .io_writeback_0_7_valid(rob_io_writeback_0_7_valid),
    .io_writeback_0_7_bits_uop_cf_exceptionVec_4(rob_io_writeback_0_7_bits_uop_cf_exceptionVec_4),
    .io_writeback_0_7_bits_uop_cf_exceptionVec_5(rob_io_writeback_0_7_bits_uop_cf_exceptionVec_5),
    .io_writeback_0_7_bits_uop_cf_exceptionVec_13(rob_io_writeback_0_7_bits_uop_cf_exceptionVec_13),
    .io_writeback_0_7_bits_uop_cf_trigger_backendHit_0(rob_io_writeback_0_7_bits_uop_cf_trigger_backendHit_0),
    .io_writeback_0_7_bits_uop_cf_trigger_backendHit_1(rob_io_writeback_0_7_bits_uop_cf_trigger_backendHit_1),
    .io_writeback_0_7_bits_uop_cf_trigger_backendHit_2(rob_io_writeback_0_7_bits_uop_cf_trigger_backendHit_2),
    .io_writeback_0_7_bits_uop_cf_trigger_backendHit_3(rob_io_writeback_0_7_bits_uop_cf_trigger_backendHit_3),
    .io_writeback_0_7_bits_uop_cf_trigger_backendHit_4(rob_io_writeback_0_7_bits_uop_cf_trigger_backendHit_4),
    .io_writeback_0_7_bits_uop_cf_trigger_backendHit_5(rob_io_writeback_0_7_bits_uop_cf_trigger_backendHit_5),
    .io_writeback_0_7_bits_uop_ctrl_flushPipe(rob_io_writeback_0_7_bits_uop_ctrl_flushPipe),
    .io_writeback_0_7_bits_uop_ctrl_replayInst(rob_io_writeback_0_7_bits_uop_ctrl_replayInst),
    .io_writeback_0_7_bits_uop_robIdx_flag(rob_io_writeback_0_7_bits_uop_robIdx_flag),
    .io_writeback_0_7_bits_uop_robIdx_value(rob_io_writeback_0_7_bits_uop_robIdx_value),
    .io_writeback_0_8_valid(rob_io_writeback_0_8_valid),
    .io_writeback_0_8_bits_uop_cf_exceptionVec_4(rob_io_writeback_0_8_bits_uop_cf_exceptionVec_4),
    .io_writeback_0_8_bits_uop_cf_exceptionVec_5(rob_io_writeback_0_8_bits_uop_cf_exceptionVec_5),
    .io_writeback_0_8_bits_uop_cf_exceptionVec_6(rob_io_writeback_0_8_bits_uop_cf_exceptionVec_6),
    .io_writeback_0_8_bits_uop_cf_exceptionVec_7(rob_io_writeback_0_8_bits_uop_cf_exceptionVec_7),
    .io_writeback_0_8_bits_uop_cf_exceptionVec_13(rob_io_writeback_0_8_bits_uop_cf_exceptionVec_13),
    .io_writeback_0_8_bits_uop_cf_exceptionVec_15(rob_io_writeback_0_8_bits_uop_cf_exceptionVec_15),
    .io_writeback_0_8_bits_uop_cf_trigger_backendHit_0(rob_io_writeback_0_8_bits_uop_cf_trigger_backendHit_0),
    .io_writeback_0_8_bits_uop_cf_trigger_backendHit_1(rob_io_writeback_0_8_bits_uop_cf_trigger_backendHit_1),
    .io_writeback_0_8_bits_uop_cf_trigger_backendHit_2(rob_io_writeback_0_8_bits_uop_cf_trigger_backendHit_2),
    .io_writeback_0_8_bits_uop_cf_trigger_backendHit_3(rob_io_writeback_0_8_bits_uop_cf_trigger_backendHit_3),
    .io_writeback_0_8_bits_uop_cf_trigger_backendHit_4(rob_io_writeback_0_8_bits_uop_cf_trigger_backendHit_4),
    .io_writeback_0_8_bits_uop_cf_trigger_backendHit_5(rob_io_writeback_0_8_bits_uop_cf_trigger_backendHit_5),
    .io_writeback_0_8_bits_uop_robIdx_flag(rob_io_writeback_0_8_bits_uop_robIdx_flag),
    .io_writeback_0_8_bits_uop_robIdx_value(rob_io_writeback_0_8_bits_uop_robIdx_value),
    .io_writeback_0_9_valid(rob_io_writeback_0_9_valid),
    .io_writeback_0_9_bits_uop_cf_exceptionVec_6(rob_io_writeback_0_9_bits_uop_cf_exceptionVec_6),
    .io_writeback_0_9_bits_uop_cf_exceptionVec_7(rob_io_writeback_0_9_bits_uop_cf_exceptionVec_7),
    .io_writeback_0_9_bits_uop_cf_exceptionVec_15(rob_io_writeback_0_9_bits_uop_cf_exceptionVec_15),
    .io_writeback_0_9_bits_uop_cf_trigger_backendHit_0(rob_io_writeback_0_9_bits_uop_cf_trigger_backendHit_0),
    .io_writeback_0_9_bits_uop_cf_trigger_backendHit_1(rob_io_writeback_0_9_bits_uop_cf_trigger_backendHit_1),
    .io_writeback_0_9_bits_uop_cf_trigger_backendHit_4(rob_io_writeback_0_9_bits_uop_cf_trigger_backendHit_4),
    .io_writeback_0_9_bits_uop_robIdx_flag(rob_io_writeback_0_9_bits_uop_robIdx_flag),
    .io_writeback_0_9_bits_uop_robIdx_value(rob_io_writeback_0_9_bits_uop_robIdx_value),
    .io_commits_isCommit(rob_io_commits_isCommit),
    .io_commits_commitValid_0(rob_io_commits_commitValid_0),
    .io_commits_commitValid_1(rob_io_commits_commitValid_1),
    .io_commits_isWalk(rob_io_commits_isWalk),
    .io_commits_walkValid_0(rob_io_commits_walkValid_0),
    .io_commits_walkValid_1(rob_io_commits_walkValid_1),
    .io_commits_info_0_ldest(rob_io_commits_info_0_ldest),
    .io_commits_info_0_rfWen(rob_io_commits_info_0_rfWen),
    .io_commits_info_0_fpWen(rob_io_commits_info_0_fpWen),
    .io_commits_info_0_wflags(rob_io_commits_info_0_wflags),
    .io_commits_info_0_commitType(rob_io_commits_info_0_commitType),
    .io_commits_info_0_pdest(rob_io_commits_info_0_pdest),
    .io_commits_info_0_old_pdest(rob_io_commits_info_0_old_pdest),
    .io_commits_info_0_ftqIdx_flag(rob_io_commits_info_0_ftqIdx_flag),
    .io_commits_info_0_ftqIdx_value(rob_io_commits_info_0_ftqIdx_value),
    .io_commits_info_0_ftqOffset(rob_io_commits_info_0_ftqOffset),
    .io_commits_info_0_isMove(rob_io_commits_info_0_isMove),
    .io_commits_info_1_ldest(rob_io_commits_info_1_ldest),
    .io_commits_info_1_rfWen(rob_io_commits_info_1_rfWen),
    .io_commits_info_1_fpWen(rob_io_commits_info_1_fpWen),
    .io_commits_info_1_wflags(rob_io_commits_info_1_wflags),
    .io_commits_info_1_commitType(rob_io_commits_info_1_commitType),
    .io_commits_info_1_pdest(rob_io_commits_info_1_pdest),
    .io_commits_info_1_old_pdest(rob_io_commits_info_1_old_pdest),
    .io_commits_info_1_ftqIdx_flag(rob_io_commits_info_1_ftqIdx_flag),
    .io_commits_info_1_ftqIdx_value(rob_io_commits_info_1_ftqIdx_value),
    .io_commits_info_1_ftqOffset(rob_io_commits_info_1_ftqOffset),
    .io_commits_info_1_isMove(rob_io_commits_info_1_isMove),
    .io_lsq_scommit(rob_io_lsq_scommit),
    .io_lsq_pendingld(rob_io_lsq_pendingld),
    .io_lsq_pendingst(rob_io_lsq_pendingst),
    .io_lsq_commit(rob_io_lsq_commit),
    .io_lsq_isMMIO_0(rob_io_lsq_isMMIO_0),
    .io_lsq_isMMIO_1(rob_io_lsq_isMMIO_1),
    .io_lsq_uop_0_robIdx_value(rob_io_lsq_uop_0_robIdx_value),
    .io_lsq_uop_1_robIdx_value(rob_io_lsq_uop_1_robIdx_value),
    .io_csr_intrBitSet(rob_io_csr_intrBitSet),
    .io_csr_wfiEvent(rob_io_csr_wfiEvent),
    .io_csr_fflags_valid(rob_io_csr_fflags_valid),
    .io_csr_fflags_bits(rob_io_csr_fflags_bits),
    .io_csr_dirty_fs(rob_io_csr_dirty_fs),
    .io_csr_perfinfo_retiredInstr(rob_io_csr_perfinfo_retiredInstr),
    .io_cpu_halt(rob_io_cpu_halt),
    .io_wfi_enable(rob_io_wfi_enable),
    .io_perf_0_value(rob_io_perf_0_value),
    .io_perf_1_value(rob_io_perf_1_value),
    .io_perf_2_value(rob_io_perf_2_value),
    .io_perf_3_value(rob_io_perf_3_value),
    .io_perf_4_value(rob_io_perf_4_value),
    .io_perf_5_value(rob_io_perf_5_value),
    .io_perf_6_value(rob_io_perf_6_value),
    .io_perf_7_value(rob_io_perf_7_value),
    .io_perf_8_value(rob_io_perf_8_value),
    .io_perf_9_value(rob_io_perf_9_value),
    .io_perf_10_value(rob_io_perf_10_value),
    .io_perf_11_value(rob_io_perf_11_value),
    .io_perf_12_value(rob_io_perf_12_value),
    .io_perf_13_value(rob_io_perf_13_value),
    .io_perf_14_value(rob_io_perf_14_value),
    .io_perf_15_value(rob_io_perf_15_value),
    .io_perf_16_value(rob_io_perf_16_value),
    .io_perf_17_value(rob_io_perf_17_value)
  );
  Dispatch2Rs_3 dispatch2 ( // @[CtrlBlock.scala 181:51]
    .io_in_0_ready(dispatch2_io_in_0_ready),
    .io_in_1_ready(dispatch2_io_in_1_ready),
    .io_in_1_bits_ctrl_fuType(dispatch2_io_in_1_bits_ctrl_fuType),
    .io_out_0_ready(dispatch2_io_out_0_ready),
    .io_out_1_ready(dispatch2_io_out_1_ready)
  );
  Dispatch2Rs_1 dispatch2_1 ( // @[CtrlBlock.scala 181:51]
    .clock(dispatch2_1_clock),
    .reset(dispatch2_1_reset),
    .io_redirect_valid(dispatch2_1_io_redirect_valid),
    .io_redirect_bits_robIdx_flag(dispatch2_1_io_redirect_bits_robIdx_flag),
    .io_redirect_bits_robIdx_value(dispatch2_1_io_redirect_bits_robIdx_value),
    .io_redirect_bits_level(dispatch2_1_io_redirect_bits_level),
    .io_in_0_ready(dispatch2_1_io_in_0_ready),
    .io_in_0_valid(dispatch2_1_io_in_0_valid),
    .io_in_0_bits_cf_foldpc(dispatch2_1_io_in_0_bits_cf_foldpc),
    .io_in_0_bits_cf_trigger_backendEn_0(dispatch2_1_io_in_0_bits_cf_trigger_backendEn_0),
    .io_in_0_bits_cf_trigger_backendEn_1(dispatch2_1_io_in_0_bits_cf_trigger_backendEn_1),
    .io_in_0_bits_cf_pd_isRVC(dispatch2_1_io_in_0_bits_cf_pd_isRVC),
    .io_in_0_bits_cf_pd_brType(dispatch2_1_io_in_0_bits_cf_pd_brType),
    .io_in_0_bits_cf_pd_isCall(dispatch2_1_io_in_0_bits_cf_pd_isCall),
    .io_in_0_bits_cf_pd_isRet(dispatch2_1_io_in_0_bits_cf_pd_isRet),
    .io_in_0_bits_cf_pred_taken(dispatch2_1_io_in_0_bits_cf_pred_taken),
    .io_in_0_bits_cf_storeSetHit(dispatch2_1_io_in_0_bits_cf_storeSetHit),
    .io_in_0_bits_cf_waitForRobIdx_flag(dispatch2_1_io_in_0_bits_cf_waitForRobIdx_flag),
    .io_in_0_bits_cf_waitForRobIdx_value(dispatch2_1_io_in_0_bits_cf_waitForRobIdx_value),
    .io_in_0_bits_cf_loadWaitBit(dispatch2_1_io_in_0_bits_cf_loadWaitBit),
    .io_in_0_bits_cf_loadWaitStrict(dispatch2_1_io_in_0_bits_cf_loadWaitStrict),
    .io_in_0_bits_cf_ssid(dispatch2_1_io_in_0_bits_cf_ssid),
    .io_in_0_bits_cf_ftqPtr_flag(dispatch2_1_io_in_0_bits_cf_ftqPtr_flag),
    .io_in_0_bits_cf_ftqPtr_value(dispatch2_1_io_in_0_bits_cf_ftqPtr_value),
    .io_in_0_bits_cf_ftqOffset(dispatch2_1_io_in_0_bits_cf_ftqOffset),
    .io_in_0_bits_ctrl_srcType_0(dispatch2_1_io_in_0_bits_ctrl_srcType_0),
    .io_in_0_bits_ctrl_srcType_1(dispatch2_1_io_in_0_bits_ctrl_srcType_1),
    .io_in_0_bits_ctrl_fuType(dispatch2_1_io_in_0_bits_ctrl_fuType),
    .io_in_0_bits_ctrl_fuOpType(dispatch2_1_io_in_0_bits_ctrl_fuOpType),
    .io_in_0_bits_ctrl_rfWen(dispatch2_1_io_in_0_bits_ctrl_rfWen),
    .io_in_0_bits_ctrl_fpWen(dispatch2_1_io_in_0_bits_ctrl_fpWen),
    .io_in_0_bits_ctrl_flushPipe(dispatch2_1_io_in_0_bits_ctrl_flushPipe),
    .io_in_0_bits_ctrl_imm(dispatch2_1_io_in_0_bits_ctrl_imm),
    .io_in_0_bits_ctrl_replayInst(dispatch2_1_io_in_0_bits_ctrl_replayInst),
    .io_in_0_bits_psrc_0(dispatch2_1_io_in_0_bits_psrc_0),
    .io_in_0_bits_psrc_1(dispatch2_1_io_in_0_bits_psrc_1),
    .io_in_0_bits_pdest(dispatch2_1_io_in_0_bits_pdest),
    .io_in_0_bits_robIdx_flag(dispatch2_1_io_in_0_bits_robIdx_flag),
    .io_in_0_bits_robIdx_value(dispatch2_1_io_in_0_bits_robIdx_value),
    .io_in_1_ready(dispatch2_1_io_in_1_ready),
    .io_in_1_valid(dispatch2_1_io_in_1_valid),
    .io_in_1_bits_cf_foldpc(dispatch2_1_io_in_1_bits_cf_foldpc),
    .io_in_1_bits_cf_trigger_backendEn_0(dispatch2_1_io_in_1_bits_cf_trigger_backendEn_0),
    .io_in_1_bits_cf_trigger_backendEn_1(dispatch2_1_io_in_1_bits_cf_trigger_backendEn_1),
    .io_in_1_bits_cf_pd_isRVC(dispatch2_1_io_in_1_bits_cf_pd_isRVC),
    .io_in_1_bits_cf_pd_brType(dispatch2_1_io_in_1_bits_cf_pd_brType),
    .io_in_1_bits_cf_pd_isCall(dispatch2_1_io_in_1_bits_cf_pd_isCall),
    .io_in_1_bits_cf_pd_isRet(dispatch2_1_io_in_1_bits_cf_pd_isRet),
    .io_in_1_bits_cf_pred_taken(dispatch2_1_io_in_1_bits_cf_pred_taken),
    .io_in_1_bits_cf_storeSetHit(dispatch2_1_io_in_1_bits_cf_storeSetHit),
    .io_in_1_bits_cf_waitForRobIdx_flag(dispatch2_1_io_in_1_bits_cf_waitForRobIdx_flag),
    .io_in_1_bits_cf_waitForRobIdx_value(dispatch2_1_io_in_1_bits_cf_waitForRobIdx_value),
    .io_in_1_bits_cf_loadWaitBit(dispatch2_1_io_in_1_bits_cf_loadWaitBit),
    .io_in_1_bits_cf_loadWaitStrict(dispatch2_1_io_in_1_bits_cf_loadWaitStrict),
    .io_in_1_bits_cf_ssid(dispatch2_1_io_in_1_bits_cf_ssid),
    .io_in_1_bits_cf_ftqPtr_flag(dispatch2_1_io_in_1_bits_cf_ftqPtr_flag),
    .io_in_1_bits_cf_ftqPtr_value(dispatch2_1_io_in_1_bits_cf_ftqPtr_value),
    .io_in_1_bits_cf_ftqOffset(dispatch2_1_io_in_1_bits_cf_ftqOffset),
    .io_in_1_bits_ctrl_srcType_0(dispatch2_1_io_in_1_bits_ctrl_srcType_0),
    .io_in_1_bits_ctrl_srcType_1(dispatch2_1_io_in_1_bits_ctrl_srcType_1),
    .io_in_1_bits_ctrl_fuType(dispatch2_1_io_in_1_bits_ctrl_fuType),
    .io_in_1_bits_ctrl_fuOpType(dispatch2_1_io_in_1_bits_ctrl_fuOpType),
    .io_in_1_bits_ctrl_rfWen(dispatch2_1_io_in_1_bits_ctrl_rfWen),
    .io_in_1_bits_ctrl_fpWen(dispatch2_1_io_in_1_bits_ctrl_fpWen),
    .io_in_1_bits_ctrl_flushPipe(dispatch2_1_io_in_1_bits_ctrl_flushPipe),
    .io_in_1_bits_ctrl_imm(dispatch2_1_io_in_1_bits_ctrl_imm),
    .io_in_1_bits_ctrl_replayInst(dispatch2_1_io_in_1_bits_ctrl_replayInst),
    .io_in_1_bits_psrc_0(dispatch2_1_io_in_1_bits_psrc_0),
    .io_in_1_bits_psrc_1(dispatch2_1_io_in_1_bits_psrc_1),
    .io_in_1_bits_pdest(dispatch2_1_io_in_1_bits_pdest),
    .io_in_1_bits_robIdx_flag(dispatch2_1_io_in_1_bits_robIdx_flag),
    .io_in_1_bits_robIdx_value(dispatch2_1_io_in_1_bits_robIdx_value),
    .io_in_2_ready(dispatch2_1_io_in_2_ready),
    .io_in_2_valid(dispatch2_1_io_in_2_valid),
    .io_in_2_bits_cf_foldpc(dispatch2_1_io_in_2_bits_cf_foldpc),
    .io_in_2_bits_cf_trigger_backendEn_0(dispatch2_1_io_in_2_bits_cf_trigger_backendEn_0),
    .io_in_2_bits_cf_trigger_backendEn_1(dispatch2_1_io_in_2_bits_cf_trigger_backendEn_1),
    .io_in_2_bits_cf_pd_isRVC(dispatch2_1_io_in_2_bits_cf_pd_isRVC),
    .io_in_2_bits_cf_pd_brType(dispatch2_1_io_in_2_bits_cf_pd_brType),
    .io_in_2_bits_cf_pd_isCall(dispatch2_1_io_in_2_bits_cf_pd_isCall),
    .io_in_2_bits_cf_pd_isRet(dispatch2_1_io_in_2_bits_cf_pd_isRet),
    .io_in_2_bits_cf_pred_taken(dispatch2_1_io_in_2_bits_cf_pred_taken),
    .io_in_2_bits_cf_storeSetHit(dispatch2_1_io_in_2_bits_cf_storeSetHit),
    .io_in_2_bits_cf_waitForRobIdx_flag(dispatch2_1_io_in_2_bits_cf_waitForRobIdx_flag),
    .io_in_2_bits_cf_waitForRobIdx_value(dispatch2_1_io_in_2_bits_cf_waitForRobIdx_value),
    .io_in_2_bits_cf_loadWaitBit(dispatch2_1_io_in_2_bits_cf_loadWaitBit),
    .io_in_2_bits_cf_loadWaitStrict(dispatch2_1_io_in_2_bits_cf_loadWaitStrict),
    .io_in_2_bits_cf_ssid(dispatch2_1_io_in_2_bits_cf_ssid),
    .io_in_2_bits_cf_ftqPtr_flag(dispatch2_1_io_in_2_bits_cf_ftqPtr_flag),
    .io_in_2_bits_cf_ftqPtr_value(dispatch2_1_io_in_2_bits_cf_ftqPtr_value),
    .io_in_2_bits_cf_ftqOffset(dispatch2_1_io_in_2_bits_cf_ftqOffset),
    .io_in_2_bits_ctrl_srcType_0(dispatch2_1_io_in_2_bits_ctrl_srcType_0),
    .io_in_2_bits_ctrl_srcType_1(dispatch2_1_io_in_2_bits_ctrl_srcType_1),
    .io_in_2_bits_ctrl_fuType(dispatch2_1_io_in_2_bits_ctrl_fuType),
    .io_in_2_bits_ctrl_fuOpType(dispatch2_1_io_in_2_bits_ctrl_fuOpType),
    .io_in_2_bits_ctrl_rfWen(dispatch2_1_io_in_2_bits_ctrl_rfWen),
    .io_in_2_bits_ctrl_fpWen(dispatch2_1_io_in_2_bits_ctrl_fpWen),
    .io_in_2_bits_ctrl_flushPipe(dispatch2_1_io_in_2_bits_ctrl_flushPipe),
    .io_in_2_bits_ctrl_imm(dispatch2_1_io_in_2_bits_ctrl_imm),
    .io_in_2_bits_ctrl_replayInst(dispatch2_1_io_in_2_bits_ctrl_replayInst),
    .io_in_2_bits_psrc_0(dispatch2_1_io_in_2_bits_psrc_0),
    .io_in_2_bits_psrc_1(dispatch2_1_io_in_2_bits_psrc_1),
    .io_in_2_bits_pdest(dispatch2_1_io_in_2_bits_pdest),
    .io_in_2_bits_robIdx_flag(dispatch2_1_io_in_2_bits_robIdx_flag),
    .io_in_2_bits_robIdx_value(dispatch2_1_io_in_2_bits_robIdx_value),
    .io_in_3_ready(dispatch2_1_io_in_3_ready),
    .io_in_3_valid(dispatch2_1_io_in_3_valid),
    .io_in_3_bits_cf_foldpc(dispatch2_1_io_in_3_bits_cf_foldpc),
    .io_in_3_bits_cf_trigger_backendEn_0(dispatch2_1_io_in_3_bits_cf_trigger_backendEn_0),
    .io_in_3_bits_cf_trigger_backendEn_1(dispatch2_1_io_in_3_bits_cf_trigger_backendEn_1),
    .io_in_3_bits_cf_pd_isRVC(dispatch2_1_io_in_3_bits_cf_pd_isRVC),
    .io_in_3_bits_cf_pd_brType(dispatch2_1_io_in_3_bits_cf_pd_brType),
    .io_in_3_bits_cf_pd_isCall(dispatch2_1_io_in_3_bits_cf_pd_isCall),
    .io_in_3_bits_cf_pd_isRet(dispatch2_1_io_in_3_bits_cf_pd_isRet),
    .io_in_3_bits_cf_pred_taken(dispatch2_1_io_in_3_bits_cf_pred_taken),
    .io_in_3_bits_cf_storeSetHit(dispatch2_1_io_in_3_bits_cf_storeSetHit),
    .io_in_3_bits_cf_waitForRobIdx_flag(dispatch2_1_io_in_3_bits_cf_waitForRobIdx_flag),
    .io_in_3_bits_cf_waitForRobIdx_value(dispatch2_1_io_in_3_bits_cf_waitForRobIdx_value),
    .io_in_3_bits_cf_loadWaitBit(dispatch2_1_io_in_3_bits_cf_loadWaitBit),
    .io_in_3_bits_cf_loadWaitStrict(dispatch2_1_io_in_3_bits_cf_loadWaitStrict),
    .io_in_3_bits_cf_ssid(dispatch2_1_io_in_3_bits_cf_ssid),
    .io_in_3_bits_cf_ftqPtr_flag(dispatch2_1_io_in_3_bits_cf_ftqPtr_flag),
    .io_in_3_bits_cf_ftqPtr_value(dispatch2_1_io_in_3_bits_cf_ftqPtr_value),
    .io_in_3_bits_cf_ftqOffset(dispatch2_1_io_in_3_bits_cf_ftqOffset),
    .io_in_3_bits_ctrl_srcType_0(dispatch2_1_io_in_3_bits_ctrl_srcType_0),
    .io_in_3_bits_ctrl_srcType_1(dispatch2_1_io_in_3_bits_ctrl_srcType_1),
    .io_in_3_bits_ctrl_fuType(dispatch2_1_io_in_3_bits_ctrl_fuType),
    .io_in_3_bits_ctrl_fuOpType(dispatch2_1_io_in_3_bits_ctrl_fuOpType),
    .io_in_3_bits_ctrl_rfWen(dispatch2_1_io_in_3_bits_ctrl_rfWen),
    .io_in_3_bits_ctrl_fpWen(dispatch2_1_io_in_3_bits_ctrl_fpWen),
    .io_in_3_bits_ctrl_flushPipe(dispatch2_1_io_in_3_bits_ctrl_flushPipe),
    .io_in_3_bits_ctrl_imm(dispatch2_1_io_in_3_bits_ctrl_imm),
    .io_in_3_bits_ctrl_replayInst(dispatch2_1_io_in_3_bits_ctrl_replayInst),
    .io_in_3_bits_psrc_0(dispatch2_1_io_in_3_bits_psrc_0),
    .io_in_3_bits_psrc_1(dispatch2_1_io_in_3_bits_psrc_1),
    .io_in_3_bits_pdest(dispatch2_1_io_in_3_bits_pdest),
    .io_in_3_bits_robIdx_flag(dispatch2_1_io_in_3_bits_robIdx_flag),
    .io_in_3_bits_robIdx_value(dispatch2_1_io_in_3_bits_robIdx_value),
    .io_readIntState_0_req(dispatch2_1_io_readIntState_0_req),
    .io_readIntState_0_resp(dispatch2_1_io_readIntState_0_resp),
    .io_readIntState_1_req(dispatch2_1_io_readIntState_1_req),
    .io_readIntState_1_resp(dispatch2_1_io_readIntState_1_resp),
    .io_readIntState_2_req(dispatch2_1_io_readIntState_2_req),
    .io_readIntState_2_resp(dispatch2_1_io_readIntState_2_resp),
    .io_readIntState_3_req(dispatch2_1_io_readIntState_3_req),
    .io_readIntState_3_resp(dispatch2_1_io_readIntState_3_resp),
    .io_readIntState_4_req(dispatch2_1_io_readIntState_4_req),
    .io_readIntState_4_resp(dispatch2_1_io_readIntState_4_resp),
    .io_readIntState_5_req(dispatch2_1_io_readIntState_5_req),
    .io_readIntState_5_resp(dispatch2_1_io_readIntState_5_resp),
    .io_readFpState_0_req(dispatch2_1_io_readFpState_0_req),
    .io_readFpState_0_resp(dispatch2_1_io_readFpState_0_resp),
    .io_readFpState_1_req(dispatch2_1_io_readFpState_1_req),
    .io_readFpState_1_resp(dispatch2_1_io_readFpState_1_resp),
    .io_out_0_ready(dispatch2_1_io_out_0_ready),
    .io_out_0_valid(dispatch2_1_io_out_0_valid),
    .io_out_0_bits_cf_foldpc(dispatch2_1_io_out_0_bits_cf_foldpc),
    .io_out_0_bits_cf_trigger_backendEn_0(dispatch2_1_io_out_0_bits_cf_trigger_backendEn_0),
    .io_out_0_bits_cf_trigger_backendEn_1(dispatch2_1_io_out_0_bits_cf_trigger_backendEn_1),
    .io_out_0_bits_cf_pd_isRVC(dispatch2_1_io_out_0_bits_cf_pd_isRVC),
    .io_out_0_bits_cf_pd_brType(dispatch2_1_io_out_0_bits_cf_pd_brType),
    .io_out_0_bits_cf_pd_isCall(dispatch2_1_io_out_0_bits_cf_pd_isCall),
    .io_out_0_bits_cf_pd_isRet(dispatch2_1_io_out_0_bits_cf_pd_isRet),
    .io_out_0_bits_cf_pred_taken(dispatch2_1_io_out_0_bits_cf_pred_taken),
    .io_out_0_bits_cf_storeSetHit(dispatch2_1_io_out_0_bits_cf_storeSetHit),
    .io_out_0_bits_cf_waitForRobIdx_flag(dispatch2_1_io_out_0_bits_cf_waitForRobIdx_flag),
    .io_out_0_bits_cf_waitForRobIdx_value(dispatch2_1_io_out_0_bits_cf_waitForRobIdx_value),
    .io_out_0_bits_cf_loadWaitBit(dispatch2_1_io_out_0_bits_cf_loadWaitBit),
    .io_out_0_bits_cf_loadWaitStrict(dispatch2_1_io_out_0_bits_cf_loadWaitStrict),
    .io_out_0_bits_cf_ssid(dispatch2_1_io_out_0_bits_cf_ssid),
    .io_out_0_bits_cf_ftqPtr_flag(dispatch2_1_io_out_0_bits_cf_ftqPtr_flag),
    .io_out_0_bits_cf_ftqPtr_value(dispatch2_1_io_out_0_bits_cf_ftqPtr_value),
    .io_out_0_bits_cf_ftqOffset(dispatch2_1_io_out_0_bits_cf_ftqOffset),
    .io_out_0_bits_ctrl_srcType_0(dispatch2_1_io_out_0_bits_ctrl_srcType_0),
    .io_out_0_bits_ctrl_fuType(dispatch2_1_io_out_0_bits_ctrl_fuType),
    .io_out_0_bits_ctrl_fuOpType(dispatch2_1_io_out_0_bits_ctrl_fuOpType),
    .io_out_0_bits_ctrl_rfWen(dispatch2_1_io_out_0_bits_ctrl_rfWen),
    .io_out_0_bits_ctrl_fpWen(dispatch2_1_io_out_0_bits_ctrl_fpWen),
    .io_out_0_bits_ctrl_imm(dispatch2_1_io_out_0_bits_ctrl_imm),
    .io_out_0_bits_srcState_0(dispatch2_1_io_out_0_bits_srcState_0),
    .io_out_0_bits_psrc_0(dispatch2_1_io_out_0_bits_psrc_0),
    .io_out_0_bits_psrc_1(dispatch2_1_io_out_0_bits_psrc_1),
    .io_out_0_bits_pdest(dispatch2_1_io_out_0_bits_pdest),
    .io_out_0_bits_robIdx_flag(dispatch2_1_io_out_0_bits_robIdx_flag),
    .io_out_0_bits_robIdx_value(dispatch2_1_io_out_0_bits_robIdx_value),
    .io_out_0_bits_lqIdx_flag(dispatch2_1_io_out_0_bits_lqIdx_flag),
    .io_out_0_bits_lqIdx_value(dispatch2_1_io_out_0_bits_lqIdx_value),
    .io_out_0_bits_sqIdx_flag(dispatch2_1_io_out_0_bits_sqIdx_flag),
    .io_out_0_bits_sqIdx_value(dispatch2_1_io_out_0_bits_sqIdx_value),
    .io_out_1_ready(dispatch2_1_io_out_1_ready),
    .io_out_1_valid(dispatch2_1_io_out_1_valid),
    .io_out_1_bits_cf_foldpc(dispatch2_1_io_out_1_bits_cf_foldpc),
    .io_out_1_bits_cf_trigger_backendEn_0(dispatch2_1_io_out_1_bits_cf_trigger_backendEn_0),
    .io_out_1_bits_cf_trigger_backendEn_1(dispatch2_1_io_out_1_bits_cf_trigger_backendEn_1),
    .io_out_1_bits_cf_pd_isRVC(dispatch2_1_io_out_1_bits_cf_pd_isRVC),
    .io_out_1_bits_cf_pd_brType(dispatch2_1_io_out_1_bits_cf_pd_brType),
    .io_out_1_bits_cf_pd_isCall(dispatch2_1_io_out_1_bits_cf_pd_isCall),
    .io_out_1_bits_cf_pd_isRet(dispatch2_1_io_out_1_bits_cf_pd_isRet),
    .io_out_1_bits_cf_pred_taken(dispatch2_1_io_out_1_bits_cf_pred_taken),
    .io_out_1_bits_cf_storeSetHit(dispatch2_1_io_out_1_bits_cf_storeSetHit),
    .io_out_1_bits_cf_waitForRobIdx_flag(dispatch2_1_io_out_1_bits_cf_waitForRobIdx_flag),
    .io_out_1_bits_cf_waitForRobIdx_value(dispatch2_1_io_out_1_bits_cf_waitForRobIdx_value),
    .io_out_1_bits_cf_loadWaitBit(dispatch2_1_io_out_1_bits_cf_loadWaitBit),
    .io_out_1_bits_cf_loadWaitStrict(dispatch2_1_io_out_1_bits_cf_loadWaitStrict),
    .io_out_1_bits_cf_ssid(dispatch2_1_io_out_1_bits_cf_ssid),
    .io_out_1_bits_cf_ftqPtr_flag(dispatch2_1_io_out_1_bits_cf_ftqPtr_flag),
    .io_out_1_bits_cf_ftqPtr_value(dispatch2_1_io_out_1_bits_cf_ftqPtr_value),
    .io_out_1_bits_cf_ftqOffset(dispatch2_1_io_out_1_bits_cf_ftqOffset),
    .io_out_1_bits_ctrl_srcType_0(dispatch2_1_io_out_1_bits_ctrl_srcType_0),
    .io_out_1_bits_ctrl_fuType(dispatch2_1_io_out_1_bits_ctrl_fuType),
    .io_out_1_bits_ctrl_fuOpType(dispatch2_1_io_out_1_bits_ctrl_fuOpType),
    .io_out_1_bits_ctrl_rfWen(dispatch2_1_io_out_1_bits_ctrl_rfWen),
    .io_out_1_bits_ctrl_fpWen(dispatch2_1_io_out_1_bits_ctrl_fpWen),
    .io_out_1_bits_ctrl_imm(dispatch2_1_io_out_1_bits_ctrl_imm),
    .io_out_1_bits_srcState_0(dispatch2_1_io_out_1_bits_srcState_0),
    .io_out_1_bits_psrc_0(dispatch2_1_io_out_1_bits_psrc_0),
    .io_out_1_bits_psrc_1(dispatch2_1_io_out_1_bits_psrc_1),
    .io_out_1_bits_pdest(dispatch2_1_io_out_1_bits_pdest),
    .io_out_1_bits_robIdx_flag(dispatch2_1_io_out_1_bits_robIdx_flag),
    .io_out_1_bits_robIdx_value(dispatch2_1_io_out_1_bits_robIdx_value),
    .io_out_1_bits_lqIdx_flag(dispatch2_1_io_out_1_bits_lqIdx_flag),
    .io_out_1_bits_lqIdx_value(dispatch2_1_io_out_1_bits_lqIdx_value),
    .io_out_1_bits_sqIdx_flag(dispatch2_1_io_out_1_bits_sqIdx_flag),
    .io_out_1_bits_sqIdx_value(dispatch2_1_io_out_1_bits_sqIdx_value),
    .io_out_2_ready(dispatch2_1_io_out_2_ready),
    .io_out_2_valid(dispatch2_1_io_out_2_valid),
    .io_out_2_bits_cf_foldpc(dispatch2_1_io_out_2_bits_cf_foldpc),
    .io_out_2_bits_cf_trigger_backendEn_0(dispatch2_1_io_out_2_bits_cf_trigger_backendEn_0),
    .io_out_2_bits_cf_trigger_backendEn_1(dispatch2_1_io_out_2_bits_cf_trigger_backendEn_1),
    .io_out_2_bits_cf_pd_isRVC(dispatch2_1_io_out_2_bits_cf_pd_isRVC),
    .io_out_2_bits_cf_pd_brType(dispatch2_1_io_out_2_bits_cf_pd_brType),
    .io_out_2_bits_cf_pd_isCall(dispatch2_1_io_out_2_bits_cf_pd_isCall),
    .io_out_2_bits_cf_pd_isRet(dispatch2_1_io_out_2_bits_cf_pd_isRet),
    .io_out_2_bits_cf_pred_taken(dispatch2_1_io_out_2_bits_cf_pred_taken),
    .io_out_2_bits_cf_storeSetHit(dispatch2_1_io_out_2_bits_cf_storeSetHit),
    .io_out_2_bits_cf_waitForRobIdx_flag(dispatch2_1_io_out_2_bits_cf_waitForRobIdx_flag),
    .io_out_2_bits_cf_waitForRobIdx_value(dispatch2_1_io_out_2_bits_cf_waitForRobIdx_value),
    .io_out_2_bits_cf_loadWaitBit(dispatch2_1_io_out_2_bits_cf_loadWaitBit),
    .io_out_2_bits_cf_loadWaitStrict(dispatch2_1_io_out_2_bits_cf_loadWaitStrict),
    .io_out_2_bits_cf_ssid(dispatch2_1_io_out_2_bits_cf_ssid),
    .io_out_2_bits_cf_ftqPtr_flag(dispatch2_1_io_out_2_bits_cf_ftqPtr_flag),
    .io_out_2_bits_cf_ftqPtr_value(dispatch2_1_io_out_2_bits_cf_ftqPtr_value),
    .io_out_2_bits_cf_ftqOffset(dispatch2_1_io_out_2_bits_cf_ftqOffset),
    .io_out_2_bits_ctrl_srcType_0(dispatch2_1_io_out_2_bits_ctrl_srcType_0),
    .io_out_2_bits_ctrl_fuType(dispatch2_1_io_out_2_bits_ctrl_fuType),
    .io_out_2_bits_ctrl_fuOpType(dispatch2_1_io_out_2_bits_ctrl_fuOpType),
    .io_out_2_bits_ctrl_rfWen(dispatch2_1_io_out_2_bits_ctrl_rfWen),
    .io_out_2_bits_ctrl_fpWen(dispatch2_1_io_out_2_bits_ctrl_fpWen),
    .io_out_2_bits_ctrl_imm(dispatch2_1_io_out_2_bits_ctrl_imm),
    .io_out_2_bits_srcState_0(dispatch2_1_io_out_2_bits_srcState_0),
    .io_out_2_bits_psrc_0(dispatch2_1_io_out_2_bits_psrc_0),
    .io_out_2_bits_pdest(dispatch2_1_io_out_2_bits_pdest),
    .io_out_2_bits_robIdx_flag(dispatch2_1_io_out_2_bits_robIdx_flag),
    .io_out_2_bits_robIdx_value(dispatch2_1_io_out_2_bits_robIdx_value),
    .io_out_2_bits_lqIdx_flag(dispatch2_1_io_out_2_bits_lqIdx_flag),
    .io_out_2_bits_lqIdx_value(dispatch2_1_io_out_2_bits_lqIdx_value),
    .io_out_2_bits_sqIdx_flag(dispatch2_1_io_out_2_bits_sqIdx_flag),
    .io_out_2_bits_sqIdx_value(dispatch2_1_io_out_2_bits_sqIdx_value),
    .io_out_3_ready(dispatch2_1_io_out_3_ready),
    .io_out_3_valid(dispatch2_1_io_out_3_valid),
    .io_out_3_bits_cf_foldpc(dispatch2_1_io_out_3_bits_cf_foldpc),
    .io_out_3_bits_cf_trigger_backendEn_0(dispatch2_1_io_out_3_bits_cf_trigger_backendEn_0),
    .io_out_3_bits_cf_trigger_backendEn_1(dispatch2_1_io_out_3_bits_cf_trigger_backendEn_1),
    .io_out_3_bits_cf_pd_isRVC(dispatch2_1_io_out_3_bits_cf_pd_isRVC),
    .io_out_3_bits_cf_pd_brType(dispatch2_1_io_out_3_bits_cf_pd_brType),
    .io_out_3_bits_cf_pd_isCall(dispatch2_1_io_out_3_bits_cf_pd_isCall),
    .io_out_3_bits_cf_pd_isRet(dispatch2_1_io_out_3_bits_cf_pd_isRet),
    .io_out_3_bits_cf_pred_taken(dispatch2_1_io_out_3_bits_cf_pred_taken),
    .io_out_3_bits_cf_storeSetHit(dispatch2_1_io_out_3_bits_cf_storeSetHit),
    .io_out_3_bits_cf_waitForRobIdx_flag(dispatch2_1_io_out_3_bits_cf_waitForRobIdx_flag),
    .io_out_3_bits_cf_waitForRobIdx_value(dispatch2_1_io_out_3_bits_cf_waitForRobIdx_value),
    .io_out_3_bits_cf_loadWaitBit(dispatch2_1_io_out_3_bits_cf_loadWaitBit),
    .io_out_3_bits_cf_loadWaitStrict(dispatch2_1_io_out_3_bits_cf_loadWaitStrict),
    .io_out_3_bits_cf_ssid(dispatch2_1_io_out_3_bits_cf_ssid),
    .io_out_3_bits_cf_ftqPtr_flag(dispatch2_1_io_out_3_bits_cf_ftqPtr_flag),
    .io_out_3_bits_cf_ftqPtr_value(dispatch2_1_io_out_3_bits_cf_ftqPtr_value),
    .io_out_3_bits_cf_ftqOffset(dispatch2_1_io_out_3_bits_cf_ftqOffset),
    .io_out_3_bits_ctrl_srcType_0(dispatch2_1_io_out_3_bits_ctrl_srcType_0),
    .io_out_3_bits_ctrl_fuType(dispatch2_1_io_out_3_bits_ctrl_fuType),
    .io_out_3_bits_ctrl_fuOpType(dispatch2_1_io_out_3_bits_ctrl_fuOpType),
    .io_out_3_bits_ctrl_rfWen(dispatch2_1_io_out_3_bits_ctrl_rfWen),
    .io_out_3_bits_ctrl_fpWen(dispatch2_1_io_out_3_bits_ctrl_fpWen),
    .io_out_3_bits_ctrl_imm(dispatch2_1_io_out_3_bits_ctrl_imm),
    .io_out_3_bits_srcState_0(dispatch2_1_io_out_3_bits_srcState_0),
    .io_out_3_bits_psrc_0(dispatch2_1_io_out_3_bits_psrc_0),
    .io_out_3_bits_pdest(dispatch2_1_io_out_3_bits_pdest),
    .io_out_3_bits_robIdx_flag(dispatch2_1_io_out_3_bits_robIdx_flag),
    .io_out_3_bits_robIdx_value(dispatch2_1_io_out_3_bits_robIdx_value),
    .io_out_3_bits_lqIdx_flag(dispatch2_1_io_out_3_bits_lqIdx_flag),
    .io_out_3_bits_lqIdx_value(dispatch2_1_io_out_3_bits_lqIdx_value),
    .io_out_3_bits_sqIdx_flag(dispatch2_1_io_out_3_bits_sqIdx_flag),
    .io_out_3_bits_sqIdx_value(dispatch2_1_io_out_3_bits_sqIdx_value),
    .io_out_4_ready(dispatch2_1_io_out_4_ready),
    .io_out_4_valid(dispatch2_1_io_out_4_valid),
    .io_out_4_bits_cf_foldpc(dispatch2_1_io_out_4_bits_cf_foldpc),
    .io_out_4_bits_cf_trigger_backendEn_0(dispatch2_1_io_out_4_bits_cf_trigger_backendEn_0),
    .io_out_4_bits_cf_trigger_backendEn_1(dispatch2_1_io_out_4_bits_cf_trigger_backendEn_1),
    .io_out_4_bits_cf_pd_isRVC(dispatch2_1_io_out_4_bits_cf_pd_isRVC),
    .io_out_4_bits_cf_pd_brType(dispatch2_1_io_out_4_bits_cf_pd_brType),
    .io_out_4_bits_cf_pd_isCall(dispatch2_1_io_out_4_bits_cf_pd_isCall),
    .io_out_4_bits_cf_pd_isRet(dispatch2_1_io_out_4_bits_cf_pd_isRet),
    .io_out_4_bits_cf_pred_taken(dispatch2_1_io_out_4_bits_cf_pred_taken),
    .io_out_4_bits_cf_storeSetHit(dispatch2_1_io_out_4_bits_cf_storeSetHit),
    .io_out_4_bits_cf_waitForRobIdx_flag(dispatch2_1_io_out_4_bits_cf_waitForRobIdx_flag),
    .io_out_4_bits_cf_waitForRobIdx_value(dispatch2_1_io_out_4_bits_cf_waitForRobIdx_value),
    .io_out_4_bits_cf_loadWaitBit(dispatch2_1_io_out_4_bits_cf_loadWaitBit),
    .io_out_4_bits_cf_loadWaitStrict(dispatch2_1_io_out_4_bits_cf_loadWaitStrict),
    .io_out_4_bits_cf_ssid(dispatch2_1_io_out_4_bits_cf_ssid),
    .io_out_4_bits_cf_ftqPtr_flag(dispatch2_1_io_out_4_bits_cf_ftqPtr_flag),
    .io_out_4_bits_cf_ftqPtr_value(dispatch2_1_io_out_4_bits_cf_ftqPtr_value),
    .io_out_4_bits_cf_ftqOffset(dispatch2_1_io_out_4_bits_cf_ftqOffset),
    .io_out_4_bits_ctrl_srcType_0(dispatch2_1_io_out_4_bits_ctrl_srcType_0),
    .io_out_4_bits_ctrl_fuType(dispatch2_1_io_out_4_bits_ctrl_fuType),
    .io_out_4_bits_ctrl_fuOpType(dispatch2_1_io_out_4_bits_ctrl_fuOpType),
    .io_out_4_bits_ctrl_rfWen(dispatch2_1_io_out_4_bits_ctrl_rfWen),
    .io_out_4_bits_ctrl_fpWen(dispatch2_1_io_out_4_bits_ctrl_fpWen),
    .io_out_4_bits_ctrl_imm(dispatch2_1_io_out_4_bits_ctrl_imm),
    .io_out_4_bits_srcState_0(dispatch2_1_io_out_4_bits_srcState_0),
    .io_out_4_bits_psrc_0(dispatch2_1_io_out_4_bits_psrc_0),
    .io_out_4_bits_pdest(dispatch2_1_io_out_4_bits_pdest),
    .io_out_4_bits_robIdx_flag(dispatch2_1_io_out_4_bits_robIdx_flag),
    .io_out_4_bits_robIdx_value(dispatch2_1_io_out_4_bits_robIdx_value),
    .io_out_4_bits_lqIdx_flag(dispatch2_1_io_out_4_bits_lqIdx_flag),
    .io_out_4_bits_lqIdx_value(dispatch2_1_io_out_4_bits_lqIdx_value),
    .io_out_4_bits_sqIdx_flag(dispatch2_1_io_out_4_bits_sqIdx_flag),
    .io_out_4_bits_sqIdx_value(dispatch2_1_io_out_4_bits_sqIdx_value),
    .io_out_5_ready(dispatch2_1_io_out_5_ready),
    .io_out_5_valid(dispatch2_1_io_out_5_valid),
    .io_out_5_bits_cf_foldpc(dispatch2_1_io_out_5_bits_cf_foldpc),
    .io_out_5_bits_cf_trigger_backendEn_0(dispatch2_1_io_out_5_bits_cf_trigger_backendEn_0),
    .io_out_5_bits_cf_trigger_backendEn_1(dispatch2_1_io_out_5_bits_cf_trigger_backendEn_1),
    .io_out_5_bits_cf_pd_isRVC(dispatch2_1_io_out_5_bits_cf_pd_isRVC),
    .io_out_5_bits_cf_pd_brType(dispatch2_1_io_out_5_bits_cf_pd_brType),
    .io_out_5_bits_cf_pd_isCall(dispatch2_1_io_out_5_bits_cf_pd_isCall),
    .io_out_5_bits_cf_pd_isRet(dispatch2_1_io_out_5_bits_cf_pd_isRet),
    .io_out_5_bits_cf_pred_taken(dispatch2_1_io_out_5_bits_cf_pred_taken),
    .io_out_5_bits_cf_storeSetHit(dispatch2_1_io_out_5_bits_cf_storeSetHit),
    .io_out_5_bits_cf_waitForRobIdx_flag(dispatch2_1_io_out_5_bits_cf_waitForRobIdx_flag),
    .io_out_5_bits_cf_waitForRobIdx_value(dispatch2_1_io_out_5_bits_cf_waitForRobIdx_value),
    .io_out_5_bits_cf_loadWaitBit(dispatch2_1_io_out_5_bits_cf_loadWaitBit),
    .io_out_5_bits_cf_loadWaitStrict(dispatch2_1_io_out_5_bits_cf_loadWaitStrict),
    .io_out_5_bits_cf_ssid(dispatch2_1_io_out_5_bits_cf_ssid),
    .io_out_5_bits_cf_ftqPtr_flag(dispatch2_1_io_out_5_bits_cf_ftqPtr_flag),
    .io_out_5_bits_cf_ftqPtr_value(dispatch2_1_io_out_5_bits_cf_ftqPtr_value),
    .io_out_5_bits_cf_ftqOffset(dispatch2_1_io_out_5_bits_cf_ftqOffset),
    .io_out_5_bits_ctrl_srcType_0(dispatch2_1_io_out_5_bits_ctrl_srcType_0),
    .io_out_5_bits_ctrl_fuType(dispatch2_1_io_out_5_bits_ctrl_fuType),
    .io_out_5_bits_ctrl_fuOpType(dispatch2_1_io_out_5_bits_ctrl_fuOpType),
    .io_out_5_bits_ctrl_rfWen(dispatch2_1_io_out_5_bits_ctrl_rfWen),
    .io_out_5_bits_ctrl_fpWen(dispatch2_1_io_out_5_bits_ctrl_fpWen),
    .io_out_5_bits_ctrl_imm(dispatch2_1_io_out_5_bits_ctrl_imm),
    .io_out_5_bits_srcState_0(dispatch2_1_io_out_5_bits_srcState_0),
    .io_out_5_bits_psrc_0(dispatch2_1_io_out_5_bits_psrc_0),
    .io_out_5_bits_pdest(dispatch2_1_io_out_5_bits_pdest),
    .io_out_5_bits_robIdx_flag(dispatch2_1_io_out_5_bits_robIdx_flag),
    .io_out_5_bits_robIdx_value(dispatch2_1_io_out_5_bits_robIdx_value),
    .io_out_5_bits_lqIdx_flag(dispatch2_1_io_out_5_bits_lqIdx_flag),
    .io_out_5_bits_lqIdx_value(dispatch2_1_io_out_5_bits_lqIdx_value),
    .io_out_5_bits_sqIdx_flag(dispatch2_1_io_out_5_bits_sqIdx_flag),
    .io_out_5_bits_sqIdx_value(dispatch2_1_io_out_5_bits_sqIdx_value),
    .io_enqLsq_canAccept(dispatch2_1_io_enqLsq_canAccept),
    .io_enqLsq_needAlloc_0(dispatch2_1_io_enqLsq_needAlloc_0),
    .io_enqLsq_needAlloc_1(dispatch2_1_io_enqLsq_needAlloc_1),
    .io_enqLsq_needAlloc_2(dispatch2_1_io_enqLsq_needAlloc_2),
    .io_enqLsq_needAlloc_3(dispatch2_1_io_enqLsq_needAlloc_3),
    .io_enqLsq_req_0_valid(dispatch2_1_io_enqLsq_req_0_valid),
    .io_enqLsq_req_0_bits_cf_trigger_backendEn_0(dispatch2_1_io_enqLsq_req_0_bits_cf_trigger_backendEn_0),
    .io_enqLsq_req_0_bits_cf_trigger_backendEn_1(dispatch2_1_io_enqLsq_req_0_bits_cf_trigger_backendEn_1),
    .io_enqLsq_req_0_bits_ctrl_fuOpType(dispatch2_1_io_enqLsq_req_0_bits_ctrl_fuOpType),
    .io_enqLsq_req_0_bits_ctrl_rfWen(dispatch2_1_io_enqLsq_req_0_bits_ctrl_rfWen),
    .io_enqLsq_req_0_bits_ctrl_fpWen(dispatch2_1_io_enqLsq_req_0_bits_ctrl_fpWen),
    .io_enqLsq_req_0_bits_ctrl_flushPipe(dispatch2_1_io_enqLsq_req_0_bits_ctrl_flushPipe),
    .io_enqLsq_req_0_bits_ctrl_replayInst(dispatch2_1_io_enqLsq_req_0_bits_ctrl_replayInst),
    .io_enqLsq_req_0_bits_pdest(dispatch2_1_io_enqLsq_req_0_bits_pdest),
    .io_enqLsq_req_0_bits_robIdx_flag(dispatch2_1_io_enqLsq_req_0_bits_robIdx_flag),
    .io_enqLsq_req_0_bits_robIdx_value(dispatch2_1_io_enqLsq_req_0_bits_robIdx_value),
    .io_enqLsq_req_1_valid(dispatch2_1_io_enqLsq_req_1_valid),
    .io_enqLsq_req_1_bits_cf_trigger_backendEn_0(dispatch2_1_io_enqLsq_req_1_bits_cf_trigger_backendEn_0),
    .io_enqLsq_req_1_bits_cf_trigger_backendEn_1(dispatch2_1_io_enqLsq_req_1_bits_cf_trigger_backendEn_1),
    .io_enqLsq_req_1_bits_ctrl_fuOpType(dispatch2_1_io_enqLsq_req_1_bits_ctrl_fuOpType),
    .io_enqLsq_req_1_bits_ctrl_rfWen(dispatch2_1_io_enqLsq_req_1_bits_ctrl_rfWen),
    .io_enqLsq_req_1_bits_ctrl_fpWen(dispatch2_1_io_enqLsq_req_1_bits_ctrl_fpWen),
    .io_enqLsq_req_1_bits_ctrl_flushPipe(dispatch2_1_io_enqLsq_req_1_bits_ctrl_flushPipe),
    .io_enqLsq_req_1_bits_ctrl_replayInst(dispatch2_1_io_enqLsq_req_1_bits_ctrl_replayInst),
    .io_enqLsq_req_1_bits_pdest(dispatch2_1_io_enqLsq_req_1_bits_pdest),
    .io_enqLsq_req_1_bits_robIdx_flag(dispatch2_1_io_enqLsq_req_1_bits_robIdx_flag),
    .io_enqLsq_req_1_bits_robIdx_value(dispatch2_1_io_enqLsq_req_1_bits_robIdx_value),
    .io_enqLsq_req_2_valid(dispatch2_1_io_enqLsq_req_2_valid),
    .io_enqLsq_req_2_bits_cf_trigger_backendEn_0(dispatch2_1_io_enqLsq_req_2_bits_cf_trigger_backendEn_0),
    .io_enqLsq_req_2_bits_cf_trigger_backendEn_1(dispatch2_1_io_enqLsq_req_2_bits_cf_trigger_backendEn_1),
    .io_enqLsq_req_2_bits_ctrl_fuOpType(dispatch2_1_io_enqLsq_req_2_bits_ctrl_fuOpType),
    .io_enqLsq_req_2_bits_ctrl_rfWen(dispatch2_1_io_enqLsq_req_2_bits_ctrl_rfWen),
    .io_enqLsq_req_2_bits_ctrl_fpWen(dispatch2_1_io_enqLsq_req_2_bits_ctrl_fpWen),
    .io_enqLsq_req_2_bits_ctrl_flushPipe(dispatch2_1_io_enqLsq_req_2_bits_ctrl_flushPipe),
    .io_enqLsq_req_2_bits_ctrl_replayInst(dispatch2_1_io_enqLsq_req_2_bits_ctrl_replayInst),
    .io_enqLsq_req_2_bits_pdest(dispatch2_1_io_enqLsq_req_2_bits_pdest),
    .io_enqLsq_req_2_bits_robIdx_flag(dispatch2_1_io_enqLsq_req_2_bits_robIdx_flag),
    .io_enqLsq_req_2_bits_robIdx_value(dispatch2_1_io_enqLsq_req_2_bits_robIdx_value),
    .io_enqLsq_req_3_valid(dispatch2_1_io_enqLsq_req_3_valid),
    .io_enqLsq_req_3_bits_cf_trigger_backendEn_0(dispatch2_1_io_enqLsq_req_3_bits_cf_trigger_backendEn_0),
    .io_enqLsq_req_3_bits_cf_trigger_backendEn_1(dispatch2_1_io_enqLsq_req_3_bits_cf_trigger_backendEn_1),
    .io_enqLsq_req_3_bits_ctrl_fuOpType(dispatch2_1_io_enqLsq_req_3_bits_ctrl_fuOpType),
    .io_enqLsq_req_3_bits_ctrl_rfWen(dispatch2_1_io_enqLsq_req_3_bits_ctrl_rfWen),
    .io_enqLsq_req_3_bits_ctrl_fpWen(dispatch2_1_io_enqLsq_req_3_bits_ctrl_fpWen),
    .io_enqLsq_req_3_bits_ctrl_flushPipe(dispatch2_1_io_enqLsq_req_3_bits_ctrl_flushPipe),
    .io_enqLsq_req_3_bits_ctrl_replayInst(dispatch2_1_io_enqLsq_req_3_bits_ctrl_replayInst),
    .io_enqLsq_req_3_bits_pdest(dispatch2_1_io_enqLsq_req_3_bits_pdest),
    .io_enqLsq_req_3_bits_robIdx_flag(dispatch2_1_io_enqLsq_req_3_bits_robIdx_flag),
    .io_enqLsq_req_3_bits_robIdx_value(dispatch2_1_io_enqLsq_req_3_bits_robIdx_value),
    .io_enqLsq_resp_0_lqIdx_flag(dispatch2_1_io_enqLsq_resp_0_lqIdx_flag),
    .io_enqLsq_resp_0_lqIdx_value(dispatch2_1_io_enqLsq_resp_0_lqIdx_value),
    .io_enqLsq_resp_0_sqIdx_flag(dispatch2_1_io_enqLsq_resp_0_sqIdx_flag),
    .io_enqLsq_resp_0_sqIdx_value(dispatch2_1_io_enqLsq_resp_0_sqIdx_value),
    .io_enqLsq_resp_1_lqIdx_flag(dispatch2_1_io_enqLsq_resp_1_lqIdx_flag),
    .io_enqLsq_resp_1_lqIdx_value(dispatch2_1_io_enqLsq_resp_1_lqIdx_value),
    .io_enqLsq_resp_1_sqIdx_flag(dispatch2_1_io_enqLsq_resp_1_sqIdx_flag),
    .io_enqLsq_resp_1_sqIdx_value(dispatch2_1_io_enqLsq_resp_1_sqIdx_value),
    .io_enqLsq_resp_2_lqIdx_flag(dispatch2_1_io_enqLsq_resp_2_lqIdx_flag),
    .io_enqLsq_resp_2_lqIdx_value(dispatch2_1_io_enqLsq_resp_2_lqIdx_value),
    .io_enqLsq_resp_2_sqIdx_flag(dispatch2_1_io_enqLsq_resp_2_sqIdx_flag),
    .io_enqLsq_resp_2_sqIdx_value(dispatch2_1_io_enqLsq_resp_2_sqIdx_value),
    .io_enqLsq_resp_3_lqIdx_flag(dispatch2_1_io_enqLsq_resp_3_lqIdx_flag),
    .io_enqLsq_resp_3_lqIdx_value(dispatch2_1_io_enqLsq_resp_3_lqIdx_value),
    .io_enqLsq_resp_3_sqIdx_flag(dispatch2_1_io_enqLsq_resp_3_sqIdx_flag),
    .io_enqLsq_resp_3_sqIdx_value(dispatch2_1_io_enqLsq_resp_3_sqIdx_value)
  );
  Dispatch2Rs_5 dispatch2_2 ( // @[CtrlBlock.scala 181:51]
    .io_in_0_ready(dispatch2_2_io_in_0_ready),
    .io_out_0_ready(dispatch2_2_io_out_0_ready)
  );
  DecodeStage decode ( // @[CtrlBlock.scala 263:22]
    .clock(decode_clock),
    .io_in_0_ready(decode_io_in_0_ready),
    .io_in_0_valid(decode_io_in_0_valid),
    .io_in_0_bits_instr(decode_io_in_0_bits_instr),
    .io_in_0_bits_foldpc(decode_io_in_0_bits_foldpc),
    .io_in_0_bits_exceptionVec_1(decode_io_in_0_bits_exceptionVec_1),
    .io_in_0_bits_exceptionVec_12(decode_io_in_0_bits_exceptionVec_12),
    .io_in_0_bits_trigger_frontendHit_0(decode_io_in_0_bits_trigger_frontendHit_0),
    .io_in_0_bits_trigger_frontendHit_1(decode_io_in_0_bits_trigger_frontendHit_1),
    .io_in_0_bits_trigger_frontendHit_2(decode_io_in_0_bits_trigger_frontendHit_2),
    .io_in_0_bits_trigger_frontendHit_3(decode_io_in_0_bits_trigger_frontendHit_3),
    .io_in_0_bits_trigger_backendEn_0(decode_io_in_0_bits_trigger_backendEn_0),
    .io_in_0_bits_trigger_backendEn_1(decode_io_in_0_bits_trigger_backendEn_1),
    .io_in_0_bits_pd_isRVC(decode_io_in_0_bits_pd_isRVC),
    .io_in_0_bits_pd_brType(decode_io_in_0_bits_pd_brType),
    .io_in_0_bits_pd_isCall(decode_io_in_0_bits_pd_isCall),
    .io_in_0_bits_pd_isRet(decode_io_in_0_bits_pd_isRet),
    .io_in_0_bits_pred_taken(decode_io_in_0_bits_pred_taken),
    .io_in_0_bits_crossPageIPFFix(decode_io_in_0_bits_crossPageIPFFix),
    .io_in_0_bits_ftqPtr_flag(decode_io_in_0_bits_ftqPtr_flag),
    .io_in_0_bits_ftqPtr_value(decode_io_in_0_bits_ftqPtr_value),
    .io_in_0_bits_ftqOffset(decode_io_in_0_bits_ftqOffset),
    .io_in_1_ready(decode_io_in_1_ready),
    .io_in_1_valid(decode_io_in_1_valid),
    .io_in_1_bits_instr(decode_io_in_1_bits_instr),
    .io_in_1_bits_foldpc(decode_io_in_1_bits_foldpc),
    .io_in_1_bits_exceptionVec_1(decode_io_in_1_bits_exceptionVec_1),
    .io_in_1_bits_exceptionVec_12(decode_io_in_1_bits_exceptionVec_12),
    .io_in_1_bits_trigger_frontendHit_0(decode_io_in_1_bits_trigger_frontendHit_0),
    .io_in_1_bits_trigger_frontendHit_1(decode_io_in_1_bits_trigger_frontendHit_1),
    .io_in_1_bits_trigger_frontendHit_2(decode_io_in_1_bits_trigger_frontendHit_2),
    .io_in_1_bits_trigger_frontendHit_3(decode_io_in_1_bits_trigger_frontendHit_3),
    .io_in_1_bits_trigger_backendEn_0(decode_io_in_1_bits_trigger_backendEn_0),
    .io_in_1_bits_trigger_backendEn_1(decode_io_in_1_bits_trigger_backendEn_1),
    .io_in_1_bits_pd_isRVC(decode_io_in_1_bits_pd_isRVC),
    .io_in_1_bits_pd_brType(decode_io_in_1_bits_pd_brType),
    .io_in_1_bits_pd_isCall(decode_io_in_1_bits_pd_isCall),
    .io_in_1_bits_pd_isRet(decode_io_in_1_bits_pd_isRet),
    .io_in_1_bits_pred_taken(decode_io_in_1_bits_pred_taken),
    .io_in_1_bits_crossPageIPFFix(decode_io_in_1_bits_crossPageIPFFix),
    .io_in_1_bits_ftqPtr_flag(decode_io_in_1_bits_ftqPtr_flag),
    .io_in_1_bits_ftqPtr_value(decode_io_in_1_bits_ftqPtr_value),
    .io_in_1_bits_ftqOffset(decode_io_in_1_bits_ftqOffset),
    .io_out_0_ready(decode_io_out_0_ready),
    .io_out_0_valid(decode_io_out_0_valid),
    .io_out_0_bits_cf_foldpc(decode_io_out_0_bits_cf_foldpc),
    .io_out_0_bits_cf_exceptionVec_1(decode_io_out_0_bits_cf_exceptionVec_1),
    .io_out_0_bits_cf_exceptionVec_2(decode_io_out_0_bits_cf_exceptionVec_2),
    .io_out_0_bits_cf_exceptionVec_12(decode_io_out_0_bits_cf_exceptionVec_12),
    .io_out_0_bits_cf_trigger_frontendHit_0(decode_io_out_0_bits_cf_trigger_frontendHit_0),
    .io_out_0_bits_cf_trigger_frontendHit_1(decode_io_out_0_bits_cf_trigger_frontendHit_1),
    .io_out_0_bits_cf_trigger_frontendHit_2(decode_io_out_0_bits_cf_trigger_frontendHit_2),
    .io_out_0_bits_cf_trigger_frontendHit_3(decode_io_out_0_bits_cf_trigger_frontendHit_3),
    .io_out_0_bits_cf_trigger_backendEn_0(decode_io_out_0_bits_cf_trigger_backendEn_0),
    .io_out_0_bits_cf_trigger_backendEn_1(decode_io_out_0_bits_cf_trigger_backendEn_1),
    .io_out_0_bits_cf_pd_isRVC(decode_io_out_0_bits_cf_pd_isRVC),
    .io_out_0_bits_cf_pd_brType(decode_io_out_0_bits_cf_pd_brType),
    .io_out_0_bits_cf_pd_isCall(decode_io_out_0_bits_cf_pd_isCall),
    .io_out_0_bits_cf_pd_isRet(decode_io_out_0_bits_cf_pd_isRet),
    .io_out_0_bits_cf_pred_taken(decode_io_out_0_bits_cf_pred_taken),
    .io_out_0_bits_cf_crossPageIPFFix(decode_io_out_0_bits_cf_crossPageIPFFix),
    .io_out_0_bits_cf_ftqPtr_flag(decode_io_out_0_bits_cf_ftqPtr_flag),
    .io_out_0_bits_cf_ftqPtr_value(decode_io_out_0_bits_cf_ftqPtr_value),
    .io_out_0_bits_cf_ftqOffset(decode_io_out_0_bits_cf_ftqOffset),
    .io_out_0_bits_ctrl_srcType_0(decode_io_out_0_bits_ctrl_srcType_0),
    .io_out_0_bits_ctrl_srcType_1(decode_io_out_0_bits_ctrl_srcType_1),
    .io_out_0_bits_ctrl_srcType_2(decode_io_out_0_bits_ctrl_srcType_2),
    .io_out_0_bits_ctrl_lsrc_0(decode_io_out_0_bits_ctrl_lsrc_0),
    .io_out_0_bits_ctrl_lsrc_1(decode_io_out_0_bits_ctrl_lsrc_1),
    .io_out_0_bits_ctrl_ldest(decode_io_out_0_bits_ctrl_ldest),
    .io_out_0_bits_ctrl_fuType(decode_io_out_0_bits_ctrl_fuType),
    .io_out_0_bits_ctrl_fuOpType(decode_io_out_0_bits_ctrl_fuOpType),
    .io_out_0_bits_ctrl_rfWen(decode_io_out_0_bits_ctrl_rfWen),
    .io_out_0_bits_ctrl_fpWen(decode_io_out_0_bits_ctrl_fpWen),
    .io_out_0_bits_ctrl_isXSTrap(decode_io_out_0_bits_ctrl_isXSTrap),
    .io_out_0_bits_ctrl_noSpecExec(decode_io_out_0_bits_ctrl_noSpecExec),
    .io_out_0_bits_ctrl_blockBackward(decode_io_out_0_bits_ctrl_blockBackward),
    .io_out_0_bits_ctrl_flushPipe(decode_io_out_0_bits_ctrl_flushPipe),
    .io_out_0_bits_ctrl_selImm(decode_io_out_0_bits_ctrl_selImm),
    .io_out_0_bits_ctrl_imm(decode_io_out_0_bits_ctrl_imm),
    .io_out_0_bits_ctrl_fpu_isAddSub(decode_io_out_0_bits_ctrl_fpu_isAddSub),
    .io_out_0_bits_ctrl_fpu_typeTagIn(decode_io_out_0_bits_ctrl_fpu_typeTagIn),
    .io_out_0_bits_ctrl_fpu_typeTagOut(decode_io_out_0_bits_ctrl_fpu_typeTagOut),
    .io_out_0_bits_ctrl_fpu_fromInt(decode_io_out_0_bits_ctrl_fpu_fromInt),
    .io_out_0_bits_ctrl_fpu_wflags(decode_io_out_0_bits_ctrl_fpu_wflags),
    .io_out_0_bits_ctrl_fpu_fpWen(decode_io_out_0_bits_ctrl_fpu_fpWen),
    .io_out_0_bits_ctrl_fpu_fmaCmd(decode_io_out_0_bits_ctrl_fpu_fmaCmd),
    .io_out_0_bits_ctrl_fpu_div(decode_io_out_0_bits_ctrl_fpu_div),
    .io_out_0_bits_ctrl_fpu_sqrt(decode_io_out_0_bits_ctrl_fpu_sqrt),
    .io_out_0_bits_ctrl_fpu_fcvt(decode_io_out_0_bits_ctrl_fpu_fcvt),
    .io_out_0_bits_ctrl_fpu_typ(decode_io_out_0_bits_ctrl_fpu_typ),
    .io_out_0_bits_ctrl_fpu_fmt(decode_io_out_0_bits_ctrl_fpu_fmt),
    .io_out_0_bits_ctrl_fpu_ren3(decode_io_out_0_bits_ctrl_fpu_ren3),
    .io_out_0_bits_ctrl_fpu_rm(decode_io_out_0_bits_ctrl_fpu_rm),
    .io_out_0_bits_ctrl_isMove(decode_io_out_0_bits_ctrl_isMove),
    .io_out_1_ready(decode_io_out_1_ready),
    .io_out_1_valid(decode_io_out_1_valid),
    .io_out_1_bits_cf_foldpc(decode_io_out_1_bits_cf_foldpc),
    .io_out_1_bits_cf_exceptionVec_1(decode_io_out_1_bits_cf_exceptionVec_1),
    .io_out_1_bits_cf_exceptionVec_2(decode_io_out_1_bits_cf_exceptionVec_2),
    .io_out_1_bits_cf_exceptionVec_12(decode_io_out_1_bits_cf_exceptionVec_12),
    .io_out_1_bits_cf_trigger_frontendHit_0(decode_io_out_1_bits_cf_trigger_frontendHit_0),
    .io_out_1_bits_cf_trigger_frontendHit_1(decode_io_out_1_bits_cf_trigger_frontendHit_1),
    .io_out_1_bits_cf_trigger_frontendHit_2(decode_io_out_1_bits_cf_trigger_frontendHit_2),
    .io_out_1_bits_cf_trigger_frontendHit_3(decode_io_out_1_bits_cf_trigger_frontendHit_3),
    .io_out_1_bits_cf_trigger_backendEn_0(decode_io_out_1_bits_cf_trigger_backendEn_0),
    .io_out_1_bits_cf_trigger_backendEn_1(decode_io_out_1_bits_cf_trigger_backendEn_1),
    .io_out_1_bits_cf_pd_isRVC(decode_io_out_1_bits_cf_pd_isRVC),
    .io_out_1_bits_cf_pd_brType(decode_io_out_1_bits_cf_pd_brType),
    .io_out_1_bits_cf_pd_isCall(decode_io_out_1_bits_cf_pd_isCall),
    .io_out_1_bits_cf_pd_isRet(decode_io_out_1_bits_cf_pd_isRet),
    .io_out_1_bits_cf_pred_taken(decode_io_out_1_bits_cf_pred_taken),
    .io_out_1_bits_cf_crossPageIPFFix(decode_io_out_1_bits_cf_crossPageIPFFix),
    .io_out_1_bits_cf_ftqPtr_flag(decode_io_out_1_bits_cf_ftqPtr_flag),
    .io_out_1_bits_cf_ftqPtr_value(decode_io_out_1_bits_cf_ftqPtr_value),
    .io_out_1_bits_cf_ftqOffset(decode_io_out_1_bits_cf_ftqOffset),
    .io_out_1_bits_ctrl_srcType_0(decode_io_out_1_bits_ctrl_srcType_0),
    .io_out_1_bits_ctrl_srcType_1(decode_io_out_1_bits_ctrl_srcType_1),
    .io_out_1_bits_ctrl_srcType_2(decode_io_out_1_bits_ctrl_srcType_2),
    .io_out_1_bits_ctrl_lsrc_0(decode_io_out_1_bits_ctrl_lsrc_0),
    .io_out_1_bits_ctrl_lsrc_1(decode_io_out_1_bits_ctrl_lsrc_1),
    .io_out_1_bits_ctrl_lsrc_2(decode_io_out_1_bits_ctrl_lsrc_2),
    .io_out_1_bits_ctrl_ldest(decode_io_out_1_bits_ctrl_ldest),
    .io_out_1_bits_ctrl_fuType(decode_io_out_1_bits_ctrl_fuType),
    .io_out_1_bits_ctrl_fuOpType(decode_io_out_1_bits_ctrl_fuOpType),
    .io_out_1_bits_ctrl_rfWen(decode_io_out_1_bits_ctrl_rfWen),
    .io_out_1_bits_ctrl_fpWen(decode_io_out_1_bits_ctrl_fpWen),
    .io_out_1_bits_ctrl_isXSTrap(decode_io_out_1_bits_ctrl_isXSTrap),
    .io_out_1_bits_ctrl_noSpecExec(decode_io_out_1_bits_ctrl_noSpecExec),
    .io_out_1_bits_ctrl_blockBackward(decode_io_out_1_bits_ctrl_blockBackward),
    .io_out_1_bits_ctrl_flushPipe(decode_io_out_1_bits_ctrl_flushPipe),
    .io_out_1_bits_ctrl_selImm(decode_io_out_1_bits_ctrl_selImm),
    .io_out_1_bits_ctrl_imm(decode_io_out_1_bits_ctrl_imm),
    .io_out_1_bits_ctrl_fpu_isAddSub(decode_io_out_1_bits_ctrl_fpu_isAddSub),
    .io_out_1_bits_ctrl_fpu_typeTagIn(decode_io_out_1_bits_ctrl_fpu_typeTagIn),
    .io_out_1_bits_ctrl_fpu_typeTagOut(decode_io_out_1_bits_ctrl_fpu_typeTagOut),
    .io_out_1_bits_ctrl_fpu_fromInt(decode_io_out_1_bits_ctrl_fpu_fromInt),
    .io_out_1_bits_ctrl_fpu_wflags(decode_io_out_1_bits_ctrl_fpu_wflags),
    .io_out_1_bits_ctrl_fpu_fpWen(decode_io_out_1_bits_ctrl_fpu_fpWen),
    .io_out_1_bits_ctrl_fpu_fmaCmd(decode_io_out_1_bits_ctrl_fpu_fmaCmd),
    .io_out_1_bits_ctrl_fpu_div(decode_io_out_1_bits_ctrl_fpu_div),
    .io_out_1_bits_ctrl_fpu_sqrt(decode_io_out_1_bits_ctrl_fpu_sqrt),
    .io_out_1_bits_ctrl_fpu_fcvt(decode_io_out_1_bits_ctrl_fpu_fcvt),
    .io_out_1_bits_ctrl_fpu_typ(decode_io_out_1_bits_ctrl_fpu_typ),
    .io_out_1_bits_ctrl_fpu_fmt(decode_io_out_1_bits_ctrl_fpu_fmt),
    .io_out_1_bits_ctrl_fpu_ren3(decode_io_out_1_bits_ctrl_fpu_ren3),
    .io_out_1_bits_ctrl_fpu_rm(decode_io_out_1_bits_ctrl_fpu_rm),
    .io_out_1_bits_ctrl_isMove(decode_io_out_1_bits_ctrl_isMove),
    .io_intRat_0_0_hold(decode_io_intRat_0_0_hold),
    .io_intRat_0_0_addr(decode_io_intRat_0_0_addr),
    .io_intRat_0_1_hold(decode_io_intRat_0_1_hold),
    .io_intRat_0_1_addr(decode_io_intRat_0_1_addr),
    .io_intRat_0_2_hold(decode_io_intRat_0_2_hold),
    .io_intRat_0_2_addr(decode_io_intRat_0_2_addr),
    .io_intRat_1_0_hold(decode_io_intRat_1_0_hold),
    .io_intRat_1_0_addr(decode_io_intRat_1_0_addr),
    .io_intRat_1_1_hold(decode_io_intRat_1_1_hold),
    .io_intRat_1_1_addr(decode_io_intRat_1_1_addr),
    .io_intRat_1_2_hold(decode_io_intRat_1_2_hold),
    .io_intRat_1_2_addr(decode_io_intRat_1_2_addr),
    .io_fpRat_0_0_hold(decode_io_fpRat_0_0_hold),
    .io_fpRat_0_0_addr(decode_io_fpRat_0_0_addr),
    .io_fpRat_0_1_hold(decode_io_fpRat_0_1_hold),
    .io_fpRat_0_1_addr(decode_io_fpRat_0_1_addr),
    .io_fpRat_0_2_hold(decode_io_fpRat_0_2_hold),
    .io_fpRat_0_2_addr(decode_io_fpRat_0_2_addr),
    .io_fpRat_0_3_hold(decode_io_fpRat_0_3_hold),
    .io_fpRat_0_3_addr(decode_io_fpRat_0_3_addr),
    .io_fpRat_1_0_hold(decode_io_fpRat_1_0_hold),
    .io_fpRat_1_0_addr(decode_io_fpRat_1_0_addr),
    .io_fpRat_1_1_hold(decode_io_fpRat_1_1_hold),
    .io_fpRat_1_1_addr(decode_io_fpRat_1_1_addr),
    .io_fpRat_1_2_hold(decode_io_fpRat_1_2_hold),
    .io_fpRat_1_2_addr(decode_io_fpRat_1_2_addr),
    .io_fpRat_1_3_hold(decode_io_fpRat_1_3_hold),
    .io_fpRat_1_3_addr(decode_io_fpRat_1_3_addr),
    .io_csrCtrl_fusion_enable(decode_io_csrCtrl_fusion_enable),
    .io_csrCtrl_wfi_enable(decode_io_csrCtrl_wfi_enable),
    .io_csrCtrl_svinval_enable(decode_io_csrCtrl_svinval_enable),
    .io_csrCtrl_singlestep(decode_io_csrCtrl_singlestep),
    .io_fusion_0(decode_io_fusion_0),
    .io_perf_0_value(decode_io_perf_0_value),
    .io_perf_1_value(decode_io_perf_1_value),
    .io_perf_2_value(decode_io_perf_2_value),
    .io_perf_3_value(decode_io_perf_3_value)
  );
  FusionDecoder fusionDecoder ( // @[CtrlBlock.scala 264:29]
    .clock(fusionDecoder_clock),
    .reset(fusionDecoder_reset),
    .io_in_0_valid(fusionDecoder_io_in_0_valid),
    .io_in_0_bits(fusionDecoder_io_in_0_bits),
    .io_in_1_valid(fusionDecoder_io_in_1_valid),
    .io_in_1_bits(fusionDecoder_io_in_1_bits),
    .io_inReady_0(fusionDecoder_io_inReady_0),
    .io_dec_0_fuOpType(fusionDecoder_io_dec_0_fuOpType),
    .io_out_0_valid(fusionDecoder_io_out_0_valid),
    .io_out_0_bits_fuType_valid(fusionDecoder_io_out_0_bits_fuType_valid),
    .io_out_0_bits_fuOpType_valid(fusionDecoder_io_out_0_bits_fuOpType_valid),
    .io_out_0_bits_fuOpType_bits(fusionDecoder_io_out_0_bits_fuOpType_bits),
    .io_out_0_bits_lsrc2_valid(fusionDecoder_io_out_0_bits_lsrc2_valid),
    .io_out_0_bits_lsrc2_bits(fusionDecoder_io_out_0_bits_lsrc2_bits),
    .io_out_0_bits_src2Type_valid(fusionDecoder_io_out_0_bits_src2Type_valid),
    .io_info_0_rs2FromRs1(fusionDecoder_io_info_0_rs2FromRs1),
    .io_info_0_rs2FromRs2(fusionDecoder_io_info_0_rs2FromRs2),
    .io_info_0_rs2FromZero(fusionDecoder_io_info_0_rs2FromZero),
    .io_clear_0(fusionDecoder_io_clear_0),
    .io_clear_1(fusionDecoder_io_clear_1)
  );
  RenameTableWrapper rat ( // @[CtrlBlock.scala 265:19]
    .clock(rat_clock),
    .reset(rat_reset),
    .io_redirect(rat_io_redirect),
    .io_robCommits_isCommit(rat_io_robCommits_isCommit),
    .io_robCommits_commitValid_0(rat_io_robCommits_commitValid_0),
    .io_robCommits_commitValid_1(rat_io_robCommits_commitValid_1),
    .io_robCommits_isWalk(rat_io_robCommits_isWalk),
    .io_robCommits_walkValid_0(rat_io_robCommits_walkValid_0),
    .io_robCommits_walkValid_1(rat_io_robCommits_walkValid_1),
    .io_robCommits_info_0_ldest(rat_io_robCommits_info_0_ldest),
    .io_robCommits_info_0_rfWen(rat_io_robCommits_info_0_rfWen),
    .io_robCommits_info_0_fpWen(rat_io_robCommits_info_0_fpWen),
    .io_robCommits_info_0_pdest(rat_io_robCommits_info_0_pdest),
    .io_robCommits_info_1_ldest(rat_io_robCommits_info_1_ldest),
    .io_robCommits_info_1_rfWen(rat_io_robCommits_info_1_rfWen),
    .io_robCommits_info_1_fpWen(rat_io_robCommits_info_1_fpWen),
    .io_robCommits_info_1_pdest(rat_io_robCommits_info_1_pdest),
    .io_intReadPorts_0_0_hold(rat_io_intReadPorts_0_0_hold),
    .io_intReadPorts_0_0_addr(rat_io_intReadPorts_0_0_addr),
    .io_intReadPorts_0_0_data(rat_io_intReadPorts_0_0_data),
    .io_intReadPorts_0_1_hold(rat_io_intReadPorts_0_1_hold),
    .io_intReadPorts_0_1_addr(rat_io_intReadPorts_0_1_addr),
    .io_intReadPorts_0_1_data(rat_io_intReadPorts_0_1_data),
    .io_intReadPorts_0_2_hold(rat_io_intReadPorts_0_2_hold),
    .io_intReadPorts_0_2_addr(rat_io_intReadPorts_0_2_addr),
    .io_intReadPorts_0_2_data(rat_io_intReadPorts_0_2_data),
    .io_intReadPorts_1_0_hold(rat_io_intReadPorts_1_0_hold),
    .io_intReadPorts_1_0_addr(rat_io_intReadPorts_1_0_addr),
    .io_intReadPorts_1_0_data(rat_io_intReadPorts_1_0_data),
    .io_intReadPorts_1_1_hold(rat_io_intReadPorts_1_1_hold),
    .io_intReadPorts_1_1_addr(rat_io_intReadPorts_1_1_addr),
    .io_intReadPorts_1_1_data(rat_io_intReadPorts_1_1_data),
    .io_intReadPorts_1_2_hold(rat_io_intReadPorts_1_2_hold),
    .io_intReadPorts_1_2_addr(rat_io_intReadPorts_1_2_addr),
    .io_intReadPorts_1_2_data(rat_io_intReadPorts_1_2_data),
    .io_intRenamePorts_0_wen(rat_io_intRenamePorts_0_wen),
    .io_intRenamePorts_0_addr(rat_io_intRenamePorts_0_addr),
    .io_intRenamePorts_0_data(rat_io_intRenamePorts_0_data),
    .io_intRenamePorts_1_wen(rat_io_intRenamePorts_1_wen),
    .io_intRenamePorts_1_addr(rat_io_intRenamePorts_1_addr),
    .io_intRenamePorts_1_data(rat_io_intRenamePorts_1_data),
    .io_fpReadPorts_0_0_hold(rat_io_fpReadPorts_0_0_hold),
    .io_fpReadPorts_0_0_addr(rat_io_fpReadPorts_0_0_addr),
    .io_fpReadPorts_0_0_data(rat_io_fpReadPorts_0_0_data),
    .io_fpReadPorts_0_1_hold(rat_io_fpReadPorts_0_1_hold),
    .io_fpReadPorts_0_1_addr(rat_io_fpReadPorts_0_1_addr),
    .io_fpReadPorts_0_1_data(rat_io_fpReadPorts_0_1_data),
    .io_fpReadPorts_0_2_hold(rat_io_fpReadPorts_0_2_hold),
    .io_fpReadPorts_0_2_addr(rat_io_fpReadPorts_0_2_addr),
    .io_fpReadPorts_0_2_data(rat_io_fpReadPorts_0_2_data),
    .io_fpReadPorts_0_3_hold(rat_io_fpReadPorts_0_3_hold),
    .io_fpReadPorts_0_3_addr(rat_io_fpReadPorts_0_3_addr),
    .io_fpReadPorts_0_3_data(rat_io_fpReadPorts_0_3_data),
    .io_fpReadPorts_1_0_hold(rat_io_fpReadPorts_1_0_hold),
    .io_fpReadPorts_1_0_addr(rat_io_fpReadPorts_1_0_addr),
    .io_fpReadPorts_1_0_data(rat_io_fpReadPorts_1_0_data),
    .io_fpReadPorts_1_1_hold(rat_io_fpReadPorts_1_1_hold),
    .io_fpReadPorts_1_1_addr(rat_io_fpReadPorts_1_1_addr),
    .io_fpReadPorts_1_1_data(rat_io_fpReadPorts_1_1_data),
    .io_fpReadPorts_1_2_hold(rat_io_fpReadPorts_1_2_hold),
    .io_fpReadPorts_1_2_addr(rat_io_fpReadPorts_1_2_addr),
    .io_fpReadPorts_1_2_data(rat_io_fpReadPorts_1_2_data),
    .io_fpReadPorts_1_3_hold(rat_io_fpReadPorts_1_3_hold),
    .io_fpReadPorts_1_3_addr(rat_io_fpReadPorts_1_3_addr),
    .io_fpReadPorts_1_3_data(rat_io_fpReadPorts_1_3_data),
    .io_fpRenamePorts_0_wen(rat_io_fpRenamePorts_0_wen),
    .io_fpRenamePorts_0_addr(rat_io_fpRenamePorts_0_addr),
    .io_fpRenamePorts_0_data(rat_io_fpRenamePorts_0_data),
    .io_fpRenamePorts_1_wen(rat_io_fpRenamePorts_1_wen),
    .io_fpRenamePorts_1_addr(rat_io_fpRenamePorts_1_addr),
    .io_fpRenamePorts_1_data(rat_io_fpRenamePorts_1_data),
    .io_debug_int_rat_0(rat_io_debug_int_rat_0),
    .io_debug_int_rat_1(rat_io_debug_int_rat_1),
    .io_debug_int_rat_2(rat_io_debug_int_rat_2),
    .io_debug_int_rat_3(rat_io_debug_int_rat_3),
    .io_debug_int_rat_4(rat_io_debug_int_rat_4),
    .io_debug_int_rat_5(rat_io_debug_int_rat_5),
    .io_debug_int_rat_6(rat_io_debug_int_rat_6),
    .io_debug_int_rat_7(rat_io_debug_int_rat_7),
    .io_debug_int_rat_8(rat_io_debug_int_rat_8),
    .io_debug_int_rat_9(rat_io_debug_int_rat_9),
    .io_debug_int_rat_10(rat_io_debug_int_rat_10),
    .io_debug_int_rat_11(rat_io_debug_int_rat_11),
    .io_debug_int_rat_12(rat_io_debug_int_rat_12),
    .io_debug_int_rat_13(rat_io_debug_int_rat_13),
    .io_debug_int_rat_14(rat_io_debug_int_rat_14),
    .io_debug_int_rat_15(rat_io_debug_int_rat_15),
    .io_debug_int_rat_16(rat_io_debug_int_rat_16),
    .io_debug_int_rat_17(rat_io_debug_int_rat_17),
    .io_debug_int_rat_18(rat_io_debug_int_rat_18),
    .io_debug_int_rat_19(rat_io_debug_int_rat_19),
    .io_debug_int_rat_20(rat_io_debug_int_rat_20),
    .io_debug_int_rat_21(rat_io_debug_int_rat_21),
    .io_debug_int_rat_22(rat_io_debug_int_rat_22),
    .io_debug_int_rat_23(rat_io_debug_int_rat_23),
    .io_debug_int_rat_24(rat_io_debug_int_rat_24),
    .io_debug_int_rat_25(rat_io_debug_int_rat_25),
    .io_debug_int_rat_26(rat_io_debug_int_rat_26),
    .io_debug_int_rat_27(rat_io_debug_int_rat_27),
    .io_debug_int_rat_28(rat_io_debug_int_rat_28),
    .io_debug_int_rat_29(rat_io_debug_int_rat_29),
    .io_debug_int_rat_30(rat_io_debug_int_rat_30),
    .io_debug_int_rat_31(rat_io_debug_int_rat_31),
    .io_debug_fp_rat_0(rat_io_debug_fp_rat_0),
    .io_debug_fp_rat_1(rat_io_debug_fp_rat_1),
    .io_debug_fp_rat_2(rat_io_debug_fp_rat_2),
    .io_debug_fp_rat_3(rat_io_debug_fp_rat_3),
    .io_debug_fp_rat_4(rat_io_debug_fp_rat_4),
    .io_debug_fp_rat_5(rat_io_debug_fp_rat_5),
    .io_debug_fp_rat_6(rat_io_debug_fp_rat_6),
    .io_debug_fp_rat_7(rat_io_debug_fp_rat_7),
    .io_debug_fp_rat_8(rat_io_debug_fp_rat_8),
    .io_debug_fp_rat_9(rat_io_debug_fp_rat_9),
    .io_debug_fp_rat_10(rat_io_debug_fp_rat_10),
    .io_debug_fp_rat_11(rat_io_debug_fp_rat_11),
    .io_debug_fp_rat_12(rat_io_debug_fp_rat_12),
    .io_debug_fp_rat_13(rat_io_debug_fp_rat_13),
    .io_debug_fp_rat_14(rat_io_debug_fp_rat_14),
    .io_debug_fp_rat_15(rat_io_debug_fp_rat_15),
    .io_debug_fp_rat_16(rat_io_debug_fp_rat_16),
    .io_debug_fp_rat_17(rat_io_debug_fp_rat_17),
    .io_debug_fp_rat_18(rat_io_debug_fp_rat_18),
    .io_debug_fp_rat_19(rat_io_debug_fp_rat_19),
    .io_debug_fp_rat_20(rat_io_debug_fp_rat_20),
    .io_debug_fp_rat_21(rat_io_debug_fp_rat_21),
    .io_debug_fp_rat_22(rat_io_debug_fp_rat_22),
    .io_debug_fp_rat_23(rat_io_debug_fp_rat_23),
    .io_debug_fp_rat_24(rat_io_debug_fp_rat_24),
    .io_debug_fp_rat_25(rat_io_debug_fp_rat_25),
    .io_debug_fp_rat_26(rat_io_debug_fp_rat_26),
    .io_debug_fp_rat_27(rat_io_debug_fp_rat_27),
    .io_debug_fp_rat_28(rat_io_debug_fp_rat_28),
    .io_debug_fp_rat_29(rat_io_debug_fp_rat_29),
    .io_debug_fp_rat_30(rat_io_debug_fp_rat_30),
    .io_debug_fp_rat_31(rat_io_debug_fp_rat_31)
  );
  SSIT ssit ( // @[CtrlBlock.scala 266:20]
    .clock(ssit_clock),
    .reset(ssit_reset),
    .io_raddr_0(ssit_io_raddr_0),
    .io_raddr_1(ssit_io_raddr_1),
    .io_rdata_0_valid(ssit_io_rdata_0_valid),
    .io_rdata_0_ssid(ssit_io_rdata_0_ssid),
    .io_rdata_0_strict(ssit_io_rdata_0_strict),
    .io_rdata_1_valid(ssit_io_rdata_1_valid),
    .io_rdata_1_ssid(ssit_io_rdata_1_ssid),
    .io_rdata_1_strict(ssit_io_rdata_1_strict),
    .io_update_valid(ssit_io_update_valid),
    .io_update_ldpc(ssit_io_update_ldpc),
    .io_update_stpc(ssit_io_update_stpc),
    .io_csrCtrl_lvpred_timeout(ssit_io_csrCtrl_lvpred_timeout)
  );
  Rename rename ( // @[CtrlBlock.scala 268:22]
    .clock(rename_clock),
    .reset(rename_reset),
    .io_redirect_valid(rename_io_redirect_valid),
    .io_redirect_bits_robIdx_flag(rename_io_redirect_bits_robIdx_flag),
    .io_redirect_bits_robIdx_value(rename_io_redirect_bits_robIdx_value),
    .io_redirect_bits_level(rename_io_redirect_bits_level),
    .io_robCommits_isCommit(rename_io_robCommits_isCommit),
    .io_robCommits_commitValid_0(rename_io_robCommits_commitValid_0),
    .io_robCommits_commitValid_1(rename_io_robCommits_commitValid_1),
    .io_robCommits_isWalk(rename_io_robCommits_isWalk),
    .io_robCommits_walkValid_0(rename_io_robCommits_walkValid_0),
    .io_robCommits_walkValid_1(rename_io_robCommits_walkValid_1),
    .io_robCommits_info_0_ldest(rename_io_robCommits_info_0_ldest),
    .io_robCommits_info_0_rfWen(rename_io_robCommits_info_0_rfWen),
    .io_robCommits_info_0_fpWen(rename_io_robCommits_info_0_fpWen),
    .io_robCommits_info_0_pdest(rename_io_robCommits_info_0_pdest),
    .io_robCommits_info_0_old_pdest(rename_io_robCommits_info_0_old_pdest),
    .io_robCommits_info_0_isMove(rename_io_robCommits_info_0_isMove),
    .io_robCommits_info_1_ldest(rename_io_robCommits_info_1_ldest),
    .io_robCommits_info_1_rfWen(rename_io_robCommits_info_1_rfWen),
    .io_robCommits_info_1_fpWen(rename_io_robCommits_info_1_fpWen),
    .io_robCommits_info_1_pdest(rename_io_robCommits_info_1_pdest),
    .io_robCommits_info_1_old_pdest(rename_io_robCommits_info_1_old_pdest),
    .io_robCommits_info_1_isMove(rename_io_robCommits_info_1_isMove),
    .io_in_0_ready(rename_io_in_0_ready),
    .io_in_0_valid(rename_io_in_0_valid),
    .io_in_0_bits_cf_foldpc(rename_io_in_0_bits_cf_foldpc),
    .io_in_0_bits_cf_exceptionVec_1(rename_io_in_0_bits_cf_exceptionVec_1),
    .io_in_0_bits_cf_exceptionVec_2(rename_io_in_0_bits_cf_exceptionVec_2),
    .io_in_0_bits_cf_exceptionVec_12(rename_io_in_0_bits_cf_exceptionVec_12),
    .io_in_0_bits_cf_trigger_frontendHit_0(rename_io_in_0_bits_cf_trigger_frontendHit_0),
    .io_in_0_bits_cf_trigger_frontendHit_1(rename_io_in_0_bits_cf_trigger_frontendHit_1),
    .io_in_0_bits_cf_trigger_frontendHit_2(rename_io_in_0_bits_cf_trigger_frontendHit_2),
    .io_in_0_bits_cf_trigger_frontendHit_3(rename_io_in_0_bits_cf_trigger_frontendHit_3),
    .io_in_0_bits_cf_trigger_backendEn_0(rename_io_in_0_bits_cf_trigger_backendEn_0),
    .io_in_0_bits_cf_trigger_backendEn_1(rename_io_in_0_bits_cf_trigger_backendEn_1),
    .io_in_0_bits_cf_pd_isRVC(rename_io_in_0_bits_cf_pd_isRVC),
    .io_in_0_bits_cf_pd_brType(rename_io_in_0_bits_cf_pd_brType),
    .io_in_0_bits_cf_pd_isCall(rename_io_in_0_bits_cf_pd_isCall),
    .io_in_0_bits_cf_pd_isRet(rename_io_in_0_bits_cf_pd_isRet),
    .io_in_0_bits_cf_pred_taken(rename_io_in_0_bits_cf_pred_taken),
    .io_in_0_bits_cf_crossPageIPFFix(rename_io_in_0_bits_cf_crossPageIPFFix),
    .io_in_0_bits_cf_ftqPtr_flag(rename_io_in_0_bits_cf_ftqPtr_flag),
    .io_in_0_bits_cf_ftqPtr_value(rename_io_in_0_bits_cf_ftqPtr_value),
    .io_in_0_bits_cf_ftqOffset(rename_io_in_0_bits_cf_ftqOffset),
    .io_in_0_bits_ctrl_srcType_0(rename_io_in_0_bits_ctrl_srcType_0),
    .io_in_0_bits_ctrl_srcType_1(rename_io_in_0_bits_ctrl_srcType_1),
    .io_in_0_bits_ctrl_srcType_2(rename_io_in_0_bits_ctrl_srcType_2),
    .io_in_0_bits_ctrl_lsrc_0(rename_io_in_0_bits_ctrl_lsrc_0),
    .io_in_0_bits_ctrl_lsrc_1(rename_io_in_0_bits_ctrl_lsrc_1),
    .io_in_0_bits_ctrl_ldest(rename_io_in_0_bits_ctrl_ldest),
    .io_in_0_bits_ctrl_fuType(rename_io_in_0_bits_ctrl_fuType),
    .io_in_0_bits_ctrl_fuOpType(rename_io_in_0_bits_ctrl_fuOpType),
    .io_in_0_bits_ctrl_rfWen(rename_io_in_0_bits_ctrl_rfWen),
    .io_in_0_bits_ctrl_fpWen(rename_io_in_0_bits_ctrl_fpWen),
    .io_in_0_bits_ctrl_isXSTrap(rename_io_in_0_bits_ctrl_isXSTrap),
    .io_in_0_bits_ctrl_noSpecExec(rename_io_in_0_bits_ctrl_noSpecExec),
    .io_in_0_bits_ctrl_blockBackward(rename_io_in_0_bits_ctrl_blockBackward),
    .io_in_0_bits_ctrl_flushPipe(rename_io_in_0_bits_ctrl_flushPipe),
    .io_in_0_bits_ctrl_selImm(rename_io_in_0_bits_ctrl_selImm),
    .io_in_0_bits_ctrl_imm(rename_io_in_0_bits_ctrl_imm),
    .io_in_0_bits_ctrl_commitType(rename_io_in_0_bits_ctrl_commitType),
    .io_in_0_bits_ctrl_fpu_isAddSub(rename_io_in_0_bits_ctrl_fpu_isAddSub),
    .io_in_0_bits_ctrl_fpu_typeTagIn(rename_io_in_0_bits_ctrl_fpu_typeTagIn),
    .io_in_0_bits_ctrl_fpu_typeTagOut(rename_io_in_0_bits_ctrl_fpu_typeTagOut),
    .io_in_0_bits_ctrl_fpu_fromInt(rename_io_in_0_bits_ctrl_fpu_fromInt),
    .io_in_0_bits_ctrl_fpu_wflags(rename_io_in_0_bits_ctrl_fpu_wflags),
    .io_in_0_bits_ctrl_fpu_fpWen(rename_io_in_0_bits_ctrl_fpu_fpWen),
    .io_in_0_bits_ctrl_fpu_fmaCmd(rename_io_in_0_bits_ctrl_fpu_fmaCmd),
    .io_in_0_bits_ctrl_fpu_div(rename_io_in_0_bits_ctrl_fpu_div),
    .io_in_0_bits_ctrl_fpu_sqrt(rename_io_in_0_bits_ctrl_fpu_sqrt),
    .io_in_0_bits_ctrl_fpu_fcvt(rename_io_in_0_bits_ctrl_fpu_fcvt),
    .io_in_0_bits_ctrl_fpu_typ(rename_io_in_0_bits_ctrl_fpu_typ),
    .io_in_0_bits_ctrl_fpu_fmt(rename_io_in_0_bits_ctrl_fpu_fmt),
    .io_in_0_bits_ctrl_fpu_ren3(rename_io_in_0_bits_ctrl_fpu_ren3),
    .io_in_0_bits_ctrl_fpu_rm(rename_io_in_0_bits_ctrl_fpu_rm),
    .io_in_0_bits_ctrl_isMove(rename_io_in_0_bits_ctrl_isMove),
    .io_in_1_ready(rename_io_in_1_ready),
    .io_in_1_valid(rename_io_in_1_valid),
    .io_in_1_bits_cf_foldpc(rename_io_in_1_bits_cf_foldpc),
    .io_in_1_bits_cf_exceptionVec_1(rename_io_in_1_bits_cf_exceptionVec_1),
    .io_in_1_bits_cf_exceptionVec_2(rename_io_in_1_bits_cf_exceptionVec_2),
    .io_in_1_bits_cf_exceptionVec_12(rename_io_in_1_bits_cf_exceptionVec_12),
    .io_in_1_bits_cf_trigger_frontendHit_0(rename_io_in_1_bits_cf_trigger_frontendHit_0),
    .io_in_1_bits_cf_trigger_frontendHit_1(rename_io_in_1_bits_cf_trigger_frontendHit_1),
    .io_in_1_bits_cf_trigger_frontendHit_2(rename_io_in_1_bits_cf_trigger_frontendHit_2),
    .io_in_1_bits_cf_trigger_frontendHit_3(rename_io_in_1_bits_cf_trigger_frontendHit_3),
    .io_in_1_bits_cf_trigger_backendEn_0(rename_io_in_1_bits_cf_trigger_backendEn_0),
    .io_in_1_bits_cf_trigger_backendEn_1(rename_io_in_1_bits_cf_trigger_backendEn_1),
    .io_in_1_bits_cf_pd_isRVC(rename_io_in_1_bits_cf_pd_isRVC),
    .io_in_1_bits_cf_pd_brType(rename_io_in_1_bits_cf_pd_brType),
    .io_in_1_bits_cf_pd_isCall(rename_io_in_1_bits_cf_pd_isCall),
    .io_in_1_bits_cf_pd_isRet(rename_io_in_1_bits_cf_pd_isRet),
    .io_in_1_bits_cf_pred_taken(rename_io_in_1_bits_cf_pred_taken),
    .io_in_1_bits_cf_crossPageIPFFix(rename_io_in_1_bits_cf_crossPageIPFFix),
    .io_in_1_bits_cf_ftqPtr_flag(rename_io_in_1_bits_cf_ftqPtr_flag),
    .io_in_1_bits_cf_ftqPtr_value(rename_io_in_1_bits_cf_ftqPtr_value),
    .io_in_1_bits_cf_ftqOffset(rename_io_in_1_bits_cf_ftqOffset),
    .io_in_1_bits_ctrl_srcType_0(rename_io_in_1_bits_ctrl_srcType_0),
    .io_in_1_bits_ctrl_srcType_1(rename_io_in_1_bits_ctrl_srcType_1),
    .io_in_1_bits_ctrl_srcType_2(rename_io_in_1_bits_ctrl_srcType_2),
    .io_in_1_bits_ctrl_lsrc_0(rename_io_in_1_bits_ctrl_lsrc_0),
    .io_in_1_bits_ctrl_lsrc_1(rename_io_in_1_bits_ctrl_lsrc_1),
    .io_in_1_bits_ctrl_lsrc_2(rename_io_in_1_bits_ctrl_lsrc_2),
    .io_in_1_bits_ctrl_ldest(rename_io_in_1_bits_ctrl_ldest),
    .io_in_1_bits_ctrl_fuType(rename_io_in_1_bits_ctrl_fuType),
    .io_in_1_bits_ctrl_fuOpType(rename_io_in_1_bits_ctrl_fuOpType),
    .io_in_1_bits_ctrl_rfWen(rename_io_in_1_bits_ctrl_rfWen),
    .io_in_1_bits_ctrl_fpWen(rename_io_in_1_bits_ctrl_fpWen),
    .io_in_1_bits_ctrl_isXSTrap(rename_io_in_1_bits_ctrl_isXSTrap),
    .io_in_1_bits_ctrl_noSpecExec(rename_io_in_1_bits_ctrl_noSpecExec),
    .io_in_1_bits_ctrl_blockBackward(rename_io_in_1_bits_ctrl_blockBackward),
    .io_in_1_bits_ctrl_flushPipe(rename_io_in_1_bits_ctrl_flushPipe),
    .io_in_1_bits_ctrl_selImm(rename_io_in_1_bits_ctrl_selImm),
    .io_in_1_bits_ctrl_imm(rename_io_in_1_bits_ctrl_imm),
    .io_in_1_bits_ctrl_fpu_isAddSub(rename_io_in_1_bits_ctrl_fpu_isAddSub),
    .io_in_1_bits_ctrl_fpu_typeTagIn(rename_io_in_1_bits_ctrl_fpu_typeTagIn),
    .io_in_1_bits_ctrl_fpu_typeTagOut(rename_io_in_1_bits_ctrl_fpu_typeTagOut),
    .io_in_1_bits_ctrl_fpu_fromInt(rename_io_in_1_bits_ctrl_fpu_fromInt),
    .io_in_1_bits_ctrl_fpu_wflags(rename_io_in_1_bits_ctrl_fpu_wflags),
    .io_in_1_bits_ctrl_fpu_fpWen(rename_io_in_1_bits_ctrl_fpu_fpWen),
    .io_in_1_bits_ctrl_fpu_fmaCmd(rename_io_in_1_bits_ctrl_fpu_fmaCmd),
    .io_in_1_bits_ctrl_fpu_div(rename_io_in_1_bits_ctrl_fpu_div),
    .io_in_1_bits_ctrl_fpu_sqrt(rename_io_in_1_bits_ctrl_fpu_sqrt),
    .io_in_1_bits_ctrl_fpu_fcvt(rename_io_in_1_bits_ctrl_fpu_fcvt),
    .io_in_1_bits_ctrl_fpu_typ(rename_io_in_1_bits_ctrl_fpu_typ),
    .io_in_1_bits_ctrl_fpu_fmt(rename_io_in_1_bits_ctrl_fpu_fmt),
    .io_in_1_bits_ctrl_fpu_ren3(rename_io_in_1_bits_ctrl_fpu_ren3),
    .io_in_1_bits_ctrl_fpu_rm(rename_io_in_1_bits_ctrl_fpu_rm),
    .io_in_1_bits_ctrl_isMove(rename_io_in_1_bits_ctrl_isMove),
    .io_fusionInfo_0_rs2FromRs1(rename_io_fusionInfo_0_rs2FromRs1),
    .io_fusionInfo_0_rs2FromRs2(rename_io_fusionInfo_0_rs2FromRs2),
    .io_fusionInfo_0_rs2FromZero(rename_io_fusionInfo_0_rs2FromZero),
    .io_ssit_0_valid(rename_io_ssit_0_valid),
    .io_ssit_0_ssid(rename_io_ssit_0_ssid),
    .io_ssit_0_strict(rename_io_ssit_0_strict),
    .io_ssit_1_valid(rename_io_ssit_1_valid),
    .io_ssit_1_ssid(rename_io_ssit_1_ssid),
    .io_ssit_1_strict(rename_io_ssit_1_strict),
    .io_intReadPorts_0_0(rename_io_intReadPorts_0_0),
    .io_intReadPorts_0_1(rename_io_intReadPorts_0_1),
    .io_intReadPorts_0_2(rename_io_intReadPorts_0_2),
    .io_intReadPorts_1_0(rename_io_intReadPorts_1_0),
    .io_intReadPorts_1_1(rename_io_intReadPorts_1_1),
    .io_intReadPorts_1_2(rename_io_intReadPorts_1_2),
    .io_fpReadPorts_0_0(rename_io_fpReadPorts_0_0),
    .io_fpReadPorts_0_1(rename_io_fpReadPorts_0_1),
    .io_fpReadPorts_0_2(rename_io_fpReadPorts_0_2),
    .io_fpReadPorts_0_3(rename_io_fpReadPorts_0_3),
    .io_fpReadPorts_1_0(rename_io_fpReadPorts_1_0),
    .io_fpReadPorts_1_1(rename_io_fpReadPorts_1_1),
    .io_fpReadPorts_1_2(rename_io_fpReadPorts_1_2),
    .io_fpReadPorts_1_3(rename_io_fpReadPorts_1_3),
    .io_intRenamePorts_0_wen(rename_io_intRenamePorts_0_wen),
    .io_intRenamePorts_0_addr(rename_io_intRenamePorts_0_addr),
    .io_intRenamePorts_0_data(rename_io_intRenamePorts_0_data),
    .io_intRenamePorts_1_wen(rename_io_intRenamePorts_1_wen),
    .io_intRenamePorts_1_addr(rename_io_intRenamePorts_1_addr),
    .io_intRenamePorts_1_data(rename_io_intRenamePorts_1_data),
    .io_fpRenamePorts_0_wen(rename_io_fpRenamePorts_0_wen),
    .io_fpRenamePorts_0_addr(rename_io_fpRenamePorts_0_addr),
    .io_fpRenamePorts_0_data(rename_io_fpRenamePorts_0_data),
    .io_fpRenamePorts_1_wen(rename_io_fpRenamePorts_1_wen),
    .io_fpRenamePorts_1_addr(rename_io_fpRenamePorts_1_addr),
    .io_fpRenamePorts_1_data(rename_io_fpRenamePorts_1_data),
    .io_out_0_ready(rename_io_out_0_ready),
    .io_out_0_valid(rename_io_out_0_valid),
    .io_out_0_bits_cf_foldpc(rename_io_out_0_bits_cf_foldpc),
    .io_out_0_bits_cf_exceptionVec_1(rename_io_out_0_bits_cf_exceptionVec_1),
    .io_out_0_bits_cf_exceptionVec_2(rename_io_out_0_bits_cf_exceptionVec_2),
    .io_out_0_bits_cf_exceptionVec_12(rename_io_out_0_bits_cf_exceptionVec_12),
    .io_out_0_bits_cf_trigger_frontendHit_0(rename_io_out_0_bits_cf_trigger_frontendHit_0),
    .io_out_0_bits_cf_trigger_frontendHit_1(rename_io_out_0_bits_cf_trigger_frontendHit_1),
    .io_out_0_bits_cf_trigger_frontendHit_2(rename_io_out_0_bits_cf_trigger_frontendHit_2),
    .io_out_0_bits_cf_trigger_frontendHit_3(rename_io_out_0_bits_cf_trigger_frontendHit_3),
    .io_out_0_bits_cf_trigger_backendEn_0(rename_io_out_0_bits_cf_trigger_backendEn_0),
    .io_out_0_bits_cf_trigger_backendEn_1(rename_io_out_0_bits_cf_trigger_backendEn_1),
    .io_out_0_bits_cf_pd_isRVC(rename_io_out_0_bits_cf_pd_isRVC),
    .io_out_0_bits_cf_pd_brType(rename_io_out_0_bits_cf_pd_brType),
    .io_out_0_bits_cf_pd_isCall(rename_io_out_0_bits_cf_pd_isCall),
    .io_out_0_bits_cf_pd_isRet(rename_io_out_0_bits_cf_pd_isRet),
    .io_out_0_bits_cf_pred_taken(rename_io_out_0_bits_cf_pred_taken),
    .io_out_0_bits_cf_crossPageIPFFix(rename_io_out_0_bits_cf_crossPageIPFFix),
    .io_out_0_bits_cf_storeSetHit(rename_io_out_0_bits_cf_storeSetHit),
    .io_out_0_bits_cf_loadWaitStrict(rename_io_out_0_bits_cf_loadWaitStrict),
    .io_out_0_bits_cf_ssid(rename_io_out_0_bits_cf_ssid),
    .io_out_0_bits_cf_ftqPtr_flag(rename_io_out_0_bits_cf_ftqPtr_flag),
    .io_out_0_bits_cf_ftqPtr_value(rename_io_out_0_bits_cf_ftqPtr_value),
    .io_out_0_bits_cf_ftqOffset(rename_io_out_0_bits_cf_ftqOffset),
    .io_out_0_bits_ctrl_srcType_0(rename_io_out_0_bits_ctrl_srcType_0),
    .io_out_0_bits_ctrl_srcType_1(rename_io_out_0_bits_ctrl_srcType_1),
    .io_out_0_bits_ctrl_srcType_2(rename_io_out_0_bits_ctrl_srcType_2),
    .io_out_0_bits_ctrl_ldest(rename_io_out_0_bits_ctrl_ldest),
    .io_out_0_bits_ctrl_fuType(rename_io_out_0_bits_ctrl_fuType),
    .io_out_0_bits_ctrl_fuOpType(rename_io_out_0_bits_ctrl_fuOpType),
    .io_out_0_bits_ctrl_rfWen(rename_io_out_0_bits_ctrl_rfWen),
    .io_out_0_bits_ctrl_fpWen(rename_io_out_0_bits_ctrl_fpWen),
    .io_out_0_bits_ctrl_isXSTrap(rename_io_out_0_bits_ctrl_isXSTrap),
    .io_out_0_bits_ctrl_noSpecExec(rename_io_out_0_bits_ctrl_noSpecExec),
    .io_out_0_bits_ctrl_blockBackward(rename_io_out_0_bits_ctrl_blockBackward),
    .io_out_0_bits_ctrl_flushPipe(rename_io_out_0_bits_ctrl_flushPipe),
    .io_out_0_bits_ctrl_selImm(rename_io_out_0_bits_ctrl_selImm),
    .io_out_0_bits_ctrl_imm(rename_io_out_0_bits_ctrl_imm),
    .io_out_0_bits_ctrl_commitType(rename_io_out_0_bits_ctrl_commitType),
    .io_out_0_bits_ctrl_fpu_isAddSub(rename_io_out_0_bits_ctrl_fpu_isAddSub),
    .io_out_0_bits_ctrl_fpu_typeTagIn(rename_io_out_0_bits_ctrl_fpu_typeTagIn),
    .io_out_0_bits_ctrl_fpu_typeTagOut(rename_io_out_0_bits_ctrl_fpu_typeTagOut),
    .io_out_0_bits_ctrl_fpu_fromInt(rename_io_out_0_bits_ctrl_fpu_fromInt),
    .io_out_0_bits_ctrl_fpu_wflags(rename_io_out_0_bits_ctrl_fpu_wflags),
    .io_out_0_bits_ctrl_fpu_fpWen(rename_io_out_0_bits_ctrl_fpu_fpWen),
    .io_out_0_bits_ctrl_fpu_fmaCmd(rename_io_out_0_bits_ctrl_fpu_fmaCmd),
    .io_out_0_bits_ctrl_fpu_div(rename_io_out_0_bits_ctrl_fpu_div),
    .io_out_0_bits_ctrl_fpu_sqrt(rename_io_out_0_bits_ctrl_fpu_sqrt),
    .io_out_0_bits_ctrl_fpu_fcvt(rename_io_out_0_bits_ctrl_fpu_fcvt),
    .io_out_0_bits_ctrl_fpu_typ(rename_io_out_0_bits_ctrl_fpu_typ),
    .io_out_0_bits_ctrl_fpu_fmt(rename_io_out_0_bits_ctrl_fpu_fmt),
    .io_out_0_bits_ctrl_fpu_ren3(rename_io_out_0_bits_ctrl_fpu_ren3),
    .io_out_0_bits_ctrl_fpu_rm(rename_io_out_0_bits_ctrl_fpu_rm),
    .io_out_0_bits_ctrl_isMove(rename_io_out_0_bits_ctrl_isMove),
    .io_out_0_bits_psrc_0(rename_io_out_0_bits_psrc_0),
    .io_out_0_bits_psrc_1(rename_io_out_0_bits_psrc_1),
    .io_out_0_bits_psrc_2(rename_io_out_0_bits_psrc_2),
    .io_out_0_bits_pdest(rename_io_out_0_bits_pdest),
    .io_out_0_bits_old_pdest(rename_io_out_0_bits_old_pdest),
    .io_out_0_bits_robIdx_flag(rename_io_out_0_bits_robIdx_flag),
    .io_out_0_bits_robIdx_value(rename_io_out_0_bits_robIdx_value),
    .io_out_0_bits_eliminatedMove(rename_io_out_0_bits_eliminatedMove),
    .io_out_1_valid(rename_io_out_1_valid),
    .io_out_1_bits_cf_foldpc(rename_io_out_1_bits_cf_foldpc),
    .io_out_1_bits_cf_exceptionVec_1(rename_io_out_1_bits_cf_exceptionVec_1),
    .io_out_1_bits_cf_exceptionVec_2(rename_io_out_1_bits_cf_exceptionVec_2),
    .io_out_1_bits_cf_exceptionVec_12(rename_io_out_1_bits_cf_exceptionVec_12),
    .io_out_1_bits_cf_trigger_frontendHit_0(rename_io_out_1_bits_cf_trigger_frontendHit_0),
    .io_out_1_bits_cf_trigger_frontendHit_1(rename_io_out_1_bits_cf_trigger_frontendHit_1),
    .io_out_1_bits_cf_trigger_frontendHit_2(rename_io_out_1_bits_cf_trigger_frontendHit_2),
    .io_out_1_bits_cf_trigger_frontendHit_3(rename_io_out_1_bits_cf_trigger_frontendHit_3),
    .io_out_1_bits_cf_trigger_backendEn_0(rename_io_out_1_bits_cf_trigger_backendEn_0),
    .io_out_1_bits_cf_trigger_backendEn_1(rename_io_out_1_bits_cf_trigger_backendEn_1),
    .io_out_1_bits_cf_pd_isRVC(rename_io_out_1_bits_cf_pd_isRVC),
    .io_out_1_bits_cf_pd_brType(rename_io_out_1_bits_cf_pd_brType),
    .io_out_1_bits_cf_pd_isCall(rename_io_out_1_bits_cf_pd_isCall),
    .io_out_1_bits_cf_pd_isRet(rename_io_out_1_bits_cf_pd_isRet),
    .io_out_1_bits_cf_pred_taken(rename_io_out_1_bits_cf_pred_taken),
    .io_out_1_bits_cf_crossPageIPFFix(rename_io_out_1_bits_cf_crossPageIPFFix),
    .io_out_1_bits_cf_storeSetHit(rename_io_out_1_bits_cf_storeSetHit),
    .io_out_1_bits_cf_loadWaitStrict(rename_io_out_1_bits_cf_loadWaitStrict),
    .io_out_1_bits_cf_ssid(rename_io_out_1_bits_cf_ssid),
    .io_out_1_bits_cf_ftqPtr_flag(rename_io_out_1_bits_cf_ftqPtr_flag),
    .io_out_1_bits_cf_ftqPtr_value(rename_io_out_1_bits_cf_ftqPtr_value),
    .io_out_1_bits_cf_ftqOffset(rename_io_out_1_bits_cf_ftqOffset),
    .io_out_1_bits_ctrl_srcType_0(rename_io_out_1_bits_ctrl_srcType_0),
    .io_out_1_bits_ctrl_srcType_1(rename_io_out_1_bits_ctrl_srcType_1),
    .io_out_1_bits_ctrl_srcType_2(rename_io_out_1_bits_ctrl_srcType_2),
    .io_out_1_bits_ctrl_ldest(rename_io_out_1_bits_ctrl_ldest),
    .io_out_1_bits_ctrl_fuType(rename_io_out_1_bits_ctrl_fuType),
    .io_out_1_bits_ctrl_fuOpType(rename_io_out_1_bits_ctrl_fuOpType),
    .io_out_1_bits_ctrl_rfWen(rename_io_out_1_bits_ctrl_rfWen),
    .io_out_1_bits_ctrl_fpWen(rename_io_out_1_bits_ctrl_fpWen),
    .io_out_1_bits_ctrl_isXSTrap(rename_io_out_1_bits_ctrl_isXSTrap),
    .io_out_1_bits_ctrl_noSpecExec(rename_io_out_1_bits_ctrl_noSpecExec),
    .io_out_1_bits_ctrl_blockBackward(rename_io_out_1_bits_ctrl_blockBackward),
    .io_out_1_bits_ctrl_flushPipe(rename_io_out_1_bits_ctrl_flushPipe),
    .io_out_1_bits_ctrl_selImm(rename_io_out_1_bits_ctrl_selImm),
    .io_out_1_bits_ctrl_imm(rename_io_out_1_bits_ctrl_imm),
    .io_out_1_bits_ctrl_fpu_isAddSub(rename_io_out_1_bits_ctrl_fpu_isAddSub),
    .io_out_1_bits_ctrl_fpu_typeTagIn(rename_io_out_1_bits_ctrl_fpu_typeTagIn),
    .io_out_1_bits_ctrl_fpu_typeTagOut(rename_io_out_1_bits_ctrl_fpu_typeTagOut),
    .io_out_1_bits_ctrl_fpu_fromInt(rename_io_out_1_bits_ctrl_fpu_fromInt),
    .io_out_1_bits_ctrl_fpu_wflags(rename_io_out_1_bits_ctrl_fpu_wflags),
    .io_out_1_bits_ctrl_fpu_fpWen(rename_io_out_1_bits_ctrl_fpu_fpWen),
    .io_out_1_bits_ctrl_fpu_fmaCmd(rename_io_out_1_bits_ctrl_fpu_fmaCmd),
    .io_out_1_bits_ctrl_fpu_div(rename_io_out_1_bits_ctrl_fpu_div),
    .io_out_1_bits_ctrl_fpu_sqrt(rename_io_out_1_bits_ctrl_fpu_sqrt),
    .io_out_1_bits_ctrl_fpu_fcvt(rename_io_out_1_bits_ctrl_fpu_fcvt),
    .io_out_1_bits_ctrl_fpu_typ(rename_io_out_1_bits_ctrl_fpu_typ),
    .io_out_1_bits_ctrl_fpu_fmt(rename_io_out_1_bits_ctrl_fpu_fmt),
    .io_out_1_bits_ctrl_fpu_ren3(rename_io_out_1_bits_ctrl_fpu_ren3),
    .io_out_1_bits_ctrl_fpu_rm(rename_io_out_1_bits_ctrl_fpu_rm),
    .io_out_1_bits_ctrl_isMove(rename_io_out_1_bits_ctrl_isMove),
    .io_out_1_bits_psrc_0(rename_io_out_1_bits_psrc_0),
    .io_out_1_bits_psrc_1(rename_io_out_1_bits_psrc_1),
    .io_out_1_bits_psrc_2(rename_io_out_1_bits_psrc_2),
    .io_out_1_bits_pdest(rename_io_out_1_bits_pdest),
    .io_out_1_bits_old_pdest(rename_io_out_1_bits_old_pdest),
    .io_out_1_bits_robIdx_flag(rename_io_out_1_bits_robIdx_flag),
    .io_out_1_bits_robIdx_value(rename_io_out_1_bits_robIdx_value),
    .io_out_1_bits_eliminatedMove(rename_io_out_1_bits_eliminatedMove),
    .io_perf_0_value(rename_io_perf_0_value),
    .io_perf_1_value(rename_io_perf_1_value),
    .io_perf_2_value(rename_io_perf_2_value),
    .io_perf_3_value(rename_io_perf_3_value),
    .io_perf_4_value(rename_io_perf_4_value),
    .io_perf_5_value(rename_io_perf_5_value),
    .io_perf_6_value(rename_io_perf_6_value),
    .io_perf_7_value(rename_io_perf_7_value),
    .io_perf_8_value(rename_io_perf_8_value),
    .io_perf_9_value(rename_io_perf_9_value),
    .io_perf_10_value(rename_io_perf_10_value),
    .io_perf_11_value(rename_io_perf_11_value),
    .io_perf_12_value(rename_io_perf_12_value),
    .io_perf_13_value(rename_io_perf_13_value)
  );
  Dispatch dispatch ( // @[CtrlBlock.scala 269:24]
    .clock(dispatch_clock),
    .reset(dispatch_reset),
    .io_fromRename_0_ready(dispatch_io_fromRename_0_ready),
    .io_fromRename_0_valid(dispatch_io_fromRename_0_valid),
    .io_fromRename_0_bits_cf_foldpc(dispatch_io_fromRename_0_bits_cf_foldpc),
    .io_fromRename_0_bits_cf_exceptionVec_1(dispatch_io_fromRename_0_bits_cf_exceptionVec_1),
    .io_fromRename_0_bits_cf_exceptionVec_2(dispatch_io_fromRename_0_bits_cf_exceptionVec_2),
    .io_fromRename_0_bits_cf_exceptionVec_12(dispatch_io_fromRename_0_bits_cf_exceptionVec_12),
    .io_fromRename_0_bits_cf_trigger_frontendHit_0(dispatch_io_fromRename_0_bits_cf_trigger_frontendHit_0),
    .io_fromRename_0_bits_cf_trigger_frontendHit_1(dispatch_io_fromRename_0_bits_cf_trigger_frontendHit_1),
    .io_fromRename_0_bits_cf_trigger_frontendHit_2(dispatch_io_fromRename_0_bits_cf_trigger_frontendHit_2),
    .io_fromRename_0_bits_cf_trigger_frontendHit_3(dispatch_io_fromRename_0_bits_cf_trigger_frontendHit_3),
    .io_fromRename_0_bits_cf_trigger_backendEn_0(dispatch_io_fromRename_0_bits_cf_trigger_backendEn_0),
    .io_fromRename_0_bits_cf_trigger_backendEn_1(dispatch_io_fromRename_0_bits_cf_trigger_backendEn_1),
    .io_fromRename_0_bits_cf_pd_isRVC(dispatch_io_fromRename_0_bits_cf_pd_isRVC),
    .io_fromRename_0_bits_cf_pd_brType(dispatch_io_fromRename_0_bits_cf_pd_brType),
    .io_fromRename_0_bits_cf_pd_isCall(dispatch_io_fromRename_0_bits_cf_pd_isCall),
    .io_fromRename_0_bits_cf_pd_isRet(dispatch_io_fromRename_0_bits_cf_pd_isRet),
    .io_fromRename_0_bits_cf_pred_taken(dispatch_io_fromRename_0_bits_cf_pred_taken),
    .io_fromRename_0_bits_cf_crossPageIPFFix(dispatch_io_fromRename_0_bits_cf_crossPageIPFFix),
    .io_fromRename_0_bits_cf_storeSetHit(dispatch_io_fromRename_0_bits_cf_storeSetHit),
    .io_fromRename_0_bits_cf_loadWaitStrict(dispatch_io_fromRename_0_bits_cf_loadWaitStrict),
    .io_fromRename_0_bits_cf_ssid(dispatch_io_fromRename_0_bits_cf_ssid),
    .io_fromRename_0_bits_cf_ftqPtr_flag(dispatch_io_fromRename_0_bits_cf_ftqPtr_flag),
    .io_fromRename_0_bits_cf_ftqPtr_value(dispatch_io_fromRename_0_bits_cf_ftqPtr_value),
    .io_fromRename_0_bits_cf_ftqOffset(dispatch_io_fromRename_0_bits_cf_ftqOffset),
    .io_fromRename_0_bits_ctrl_srcType_0(dispatch_io_fromRename_0_bits_ctrl_srcType_0),
    .io_fromRename_0_bits_ctrl_srcType_1(dispatch_io_fromRename_0_bits_ctrl_srcType_1),
    .io_fromRename_0_bits_ctrl_srcType_2(dispatch_io_fromRename_0_bits_ctrl_srcType_2),
    .io_fromRename_0_bits_ctrl_ldest(dispatch_io_fromRename_0_bits_ctrl_ldest),
    .io_fromRename_0_bits_ctrl_fuType(dispatch_io_fromRename_0_bits_ctrl_fuType),
    .io_fromRename_0_bits_ctrl_fuOpType(dispatch_io_fromRename_0_bits_ctrl_fuOpType),
    .io_fromRename_0_bits_ctrl_rfWen(dispatch_io_fromRename_0_bits_ctrl_rfWen),
    .io_fromRename_0_bits_ctrl_fpWen(dispatch_io_fromRename_0_bits_ctrl_fpWen),
    .io_fromRename_0_bits_ctrl_isXSTrap(dispatch_io_fromRename_0_bits_ctrl_isXSTrap),
    .io_fromRename_0_bits_ctrl_noSpecExec(dispatch_io_fromRename_0_bits_ctrl_noSpecExec),
    .io_fromRename_0_bits_ctrl_blockBackward(dispatch_io_fromRename_0_bits_ctrl_blockBackward),
    .io_fromRename_0_bits_ctrl_flushPipe(dispatch_io_fromRename_0_bits_ctrl_flushPipe),
    .io_fromRename_0_bits_ctrl_selImm(dispatch_io_fromRename_0_bits_ctrl_selImm),
    .io_fromRename_0_bits_ctrl_imm(dispatch_io_fromRename_0_bits_ctrl_imm),
    .io_fromRename_0_bits_ctrl_commitType(dispatch_io_fromRename_0_bits_ctrl_commitType),
    .io_fromRename_0_bits_ctrl_fpu_isAddSub(dispatch_io_fromRename_0_bits_ctrl_fpu_isAddSub),
    .io_fromRename_0_bits_ctrl_fpu_typeTagIn(dispatch_io_fromRename_0_bits_ctrl_fpu_typeTagIn),
    .io_fromRename_0_bits_ctrl_fpu_typeTagOut(dispatch_io_fromRename_0_bits_ctrl_fpu_typeTagOut),
    .io_fromRename_0_bits_ctrl_fpu_fromInt(dispatch_io_fromRename_0_bits_ctrl_fpu_fromInt),
    .io_fromRename_0_bits_ctrl_fpu_wflags(dispatch_io_fromRename_0_bits_ctrl_fpu_wflags),
    .io_fromRename_0_bits_ctrl_fpu_fpWen(dispatch_io_fromRename_0_bits_ctrl_fpu_fpWen),
    .io_fromRename_0_bits_ctrl_fpu_fmaCmd(dispatch_io_fromRename_0_bits_ctrl_fpu_fmaCmd),
    .io_fromRename_0_bits_ctrl_fpu_div(dispatch_io_fromRename_0_bits_ctrl_fpu_div),
    .io_fromRename_0_bits_ctrl_fpu_sqrt(dispatch_io_fromRename_0_bits_ctrl_fpu_sqrt),
    .io_fromRename_0_bits_ctrl_fpu_fcvt(dispatch_io_fromRename_0_bits_ctrl_fpu_fcvt),
    .io_fromRename_0_bits_ctrl_fpu_typ(dispatch_io_fromRename_0_bits_ctrl_fpu_typ),
    .io_fromRename_0_bits_ctrl_fpu_fmt(dispatch_io_fromRename_0_bits_ctrl_fpu_fmt),
    .io_fromRename_0_bits_ctrl_fpu_ren3(dispatch_io_fromRename_0_bits_ctrl_fpu_ren3),
    .io_fromRename_0_bits_ctrl_fpu_rm(dispatch_io_fromRename_0_bits_ctrl_fpu_rm),
    .io_fromRename_0_bits_ctrl_isMove(dispatch_io_fromRename_0_bits_ctrl_isMove),
    .io_fromRename_0_bits_psrc_0(dispatch_io_fromRename_0_bits_psrc_0),
    .io_fromRename_0_bits_psrc_1(dispatch_io_fromRename_0_bits_psrc_1),
    .io_fromRename_0_bits_psrc_2(dispatch_io_fromRename_0_bits_psrc_2),
    .io_fromRename_0_bits_pdest(dispatch_io_fromRename_0_bits_pdest),
    .io_fromRename_0_bits_old_pdest(dispatch_io_fromRename_0_bits_old_pdest),
    .io_fromRename_0_bits_robIdx_flag(dispatch_io_fromRename_0_bits_robIdx_flag),
    .io_fromRename_0_bits_robIdx_value(dispatch_io_fromRename_0_bits_robIdx_value),
    .io_fromRename_0_bits_eliminatedMove(dispatch_io_fromRename_0_bits_eliminatedMove),
    .io_fromRename_1_ready(dispatch_io_fromRename_1_ready),
    .io_fromRename_1_valid(dispatch_io_fromRename_1_valid),
    .io_fromRename_1_bits_cf_foldpc(dispatch_io_fromRename_1_bits_cf_foldpc),
    .io_fromRename_1_bits_cf_exceptionVec_1(dispatch_io_fromRename_1_bits_cf_exceptionVec_1),
    .io_fromRename_1_bits_cf_exceptionVec_2(dispatch_io_fromRename_1_bits_cf_exceptionVec_2),
    .io_fromRename_1_bits_cf_exceptionVec_12(dispatch_io_fromRename_1_bits_cf_exceptionVec_12),
    .io_fromRename_1_bits_cf_trigger_frontendHit_0(dispatch_io_fromRename_1_bits_cf_trigger_frontendHit_0),
    .io_fromRename_1_bits_cf_trigger_frontendHit_1(dispatch_io_fromRename_1_bits_cf_trigger_frontendHit_1),
    .io_fromRename_1_bits_cf_trigger_frontendHit_2(dispatch_io_fromRename_1_bits_cf_trigger_frontendHit_2),
    .io_fromRename_1_bits_cf_trigger_frontendHit_3(dispatch_io_fromRename_1_bits_cf_trigger_frontendHit_3),
    .io_fromRename_1_bits_cf_trigger_backendEn_0(dispatch_io_fromRename_1_bits_cf_trigger_backendEn_0),
    .io_fromRename_1_bits_cf_trigger_backendEn_1(dispatch_io_fromRename_1_bits_cf_trigger_backendEn_1),
    .io_fromRename_1_bits_cf_pd_isRVC(dispatch_io_fromRename_1_bits_cf_pd_isRVC),
    .io_fromRename_1_bits_cf_pd_brType(dispatch_io_fromRename_1_bits_cf_pd_brType),
    .io_fromRename_1_bits_cf_pd_isCall(dispatch_io_fromRename_1_bits_cf_pd_isCall),
    .io_fromRename_1_bits_cf_pd_isRet(dispatch_io_fromRename_1_bits_cf_pd_isRet),
    .io_fromRename_1_bits_cf_pred_taken(dispatch_io_fromRename_1_bits_cf_pred_taken),
    .io_fromRename_1_bits_cf_crossPageIPFFix(dispatch_io_fromRename_1_bits_cf_crossPageIPFFix),
    .io_fromRename_1_bits_cf_storeSetHit(dispatch_io_fromRename_1_bits_cf_storeSetHit),
    .io_fromRename_1_bits_cf_loadWaitStrict(dispatch_io_fromRename_1_bits_cf_loadWaitStrict),
    .io_fromRename_1_bits_cf_ssid(dispatch_io_fromRename_1_bits_cf_ssid),
    .io_fromRename_1_bits_cf_ftqPtr_flag(dispatch_io_fromRename_1_bits_cf_ftqPtr_flag),
    .io_fromRename_1_bits_cf_ftqPtr_value(dispatch_io_fromRename_1_bits_cf_ftqPtr_value),
    .io_fromRename_1_bits_cf_ftqOffset(dispatch_io_fromRename_1_bits_cf_ftqOffset),
    .io_fromRename_1_bits_ctrl_srcType_0(dispatch_io_fromRename_1_bits_ctrl_srcType_0),
    .io_fromRename_1_bits_ctrl_srcType_1(dispatch_io_fromRename_1_bits_ctrl_srcType_1),
    .io_fromRename_1_bits_ctrl_srcType_2(dispatch_io_fromRename_1_bits_ctrl_srcType_2),
    .io_fromRename_1_bits_ctrl_ldest(dispatch_io_fromRename_1_bits_ctrl_ldest),
    .io_fromRename_1_bits_ctrl_fuType(dispatch_io_fromRename_1_bits_ctrl_fuType),
    .io_fromRename_1_bits_ctrl_fuOpType(dispatch_io_fromRename_1_bits_ctrl_fuOpType),
    .io_fromRename_1_bits_ctrl_rfWen(dispatch_io_fromRename_1_bits_ctrl_rfWen),
    .io_fromRename_1_bits_ctrl_fpWen(dispatch_io_fromRename_1_bits_ctrl_fpWen),
    .io_fromRename_1_bits_ctrl_isXSTrap(dispatch_io_fromRename_1_bits_ctrl_isXSTrap),
    .io_fromRename_1_bits_ctrl_noSpecExec(dispatch_io_fromRename_1_bits_ctrl_noSpecExec),
    .io_fromRename_1_bits_ctrl_blockBackward(dispatch_io_fromRename_1_bits_ctrl_blockBackward),
    .io_fromRename_1_bits_ctrl_flushPipe(dispatch_io_fromRename_1_bits_ctrl_flushPipe),
    .io_fromRename_1_bits_ctrl_selImm(dispatch_io_fromRename_1_bits_ctrl_selImm),
    .io_fromRename_1_bits_ctrl_imm(dispatch_io_fromRename_1_bits_ctrl_imm),
    .io_fromRename_1_bits_ctrl_fpu_isAddSub(dispatch_io_fromRename_1_bits_ctrl_fpu_isAddSub),
    .io_fromRename_1_bits_ctrl_fpu_typeTagIn(dispatch_io_fromRename_1_bits_ctrl_fpu_typeTagIn),
    .io_fromRename_1_bits_ctrl_fpu_typeTagOut(dispatch_io_fromRename_1_bits_ctrl_fpu_typeTagOut),
    .io_fromRename_1_bits_ctrl_fpu_fromInt(dispatch_io_fromRename_1_bits_ctrl_fpu_fromInt),
    .io_fromRename_1_bits_ctrl_fpu_wflags(dispatch_io_fromRename_1_bits_ctrl_fpu_wflags),
    .io_fromRename_1_bits_ctrl_fpu_fpWen(dispatch_io_fromRename_1_bits_ctrl_fpu_fpWen),
    .io_fromRename_1_bits_ctrl_fpu_fmaCmd(dispatch_io_fromRename_1_bits_ctrl_fpu_fmaCmd),
    .io_fromRename_1_bits_ctrl_fpu_div(dispatch_io_fromRename_1_bits_ctrl_fpu_div),
    .io_fromRename_1_bits_ctrl_fpu_sqrt(dispatch_io_fromRename_1_bits_ctrl_fpu_sqrt),
    .io_fromRename_1_bits_ctrl_fpu_fcvt(dispatch_io_fromRename_1_bits_ctrl_fpu_fcvt),
    .io_fromRename_1_bits_ctrl_fpu_typ(dispatch_io_fromRename_1_bits_ctrl_fpu_typ),
    .io_fromRename_1_bits_ctrl_fpu_fmt(dispatch_io_fromRename_1_bits_ctrl_fpu_fmt),
    .io_fromRename_1_bits_ctrl_fpu_ren3(dispatch_io_fromRename_1_bits_ctrl_fpu_ren3),
    .io_fromRename_1_bits_ctrl_fpu_rm(dispatch_io_fromRename_1_bits_ctrl_fpu_rm),
    .io_fromRename_1_bits_ctrl_isMove(dispatch_io_fromRename_1_bits_ctrl_isMove),
    .io_fromRename_1_bits_psrc_0(dispatch_io_fromRename_1_bits_psrc_0),
    .io_fromRename_1_bits_psrc_1(dispatch_io_fromRename_1_bits_psrc_1),
    .io_fromRename_1_bits_psrc_2(dispatch_io_fromRename_1_bits_psrc_2),
    .io_fromRename_1_bits_pdest(dispatch_io_fromRename_1_bits_pdest),
    .io_fromRename_1_bits_old_pdest(dispatch_io_fromRename_1_bits_old_pdest),
    .io_fromRename_1_bits_robIdx_flag(dispatch_io_fromRename_1_bits_robIdx_flag),
    .io_fromRename_1_bits_robIdx_value(dispatch_io_fromRename_1_bits_robIdx_value),
    .io_fromRename_1_bits_eliminatedMove(dispatch_io_fromRename_1_bits_eliminatedMove),
    .io_recv_0(dispatch_io_recv_0),
    .io_recv_1(dispatch_io_recv_1),
    .io_enqRob_canAccept(dispatch_io_enqRob_canAccept),
    .io_enqRob_isEmpty(dispatch_io_enqRob_isEmpty),
    .io_enqRob_needAlloc_0(dispatch_io_enqRob_needAlloc_0),
    .io_enqRob_req_0_valid(dispatch_io_enqRob_req_0_valid),
    .io_enqRob_req_0_bits_cf_exceptionVec_1(dispatch_io_enqRob_req_0_bits_cf_exceptionVec_1),
    .io_enqRob_req_0_bits_cf_exceptionVec_2(dispatch_io_enqRob_req_0_bits_cf_exceptionVec_2),
    .io_enqRob_req_0_bits_cf_exceptionVec_12(dispatch_io_enqRob_req_0_bits_cf_exceptionVec_12),
    .io_enqRob_req_0_bits_cf_trigger_frontendHit_0(dispatch_io_enqRob_req_0_bits_cf_trigger_frontendHit_0),
    .io_enqRob_req_0_bits_cf_trigger_frontendHit_1(dispatch_io_enqRob_req_0_bits_cf_trigger_frontendHit_1),
    .io_enqRob_req_0_bits_cf_trigger_frontendHit_2(dispatch_io_enqRob_req_0_bits_cf_trigger_frontendHit_2),
    .io_enqRob_req_0_bits_cf_trigger_frontendHit_3(dispatch_io_enqRob_req_0_bits_cf_trigger_frontendHit_3),
    .io_enqRob_req_0_bits_cf_pd_isRVC(dispatch_io_enqRob_req_0_bits_cf_pd_isRVC),
    .io_enqRob_req_0_bits_cf_crossPageIPFFix(dispatch_io_enqRob_req_0_bits_cf_crossPageIPFFix),
    .io_enqRob_req_0_bits_cf_loadWaitBit(dispatch_io_enqRob_req_0_bits_cf_loadWaitBit),
    .io_enqRob_req_0_bits_cf_ftqPtr_flag(dispatch_io_enqRob_req_0_bits_cf_ftqPtr_flag),
    .io_enqRob_req_0_bits_cf_ftqPtr_value(dispatch_io_enqRob_req_0_bits_cf_ftqPtr_value),
    .io_enqRob_req_0_bits_cf_ftqOffset(dispatch_io_enqRob_req_0_bits_cf_ftqOffset),
    .io_enqRob_req_0_bits_ctrl_ldest(dispatch_io_enqRob_req_0_bits_ctrl_ldest),
    .io_enqRob_req_0_bits_ctrl_fuType(dispatch_io_enqRob_req_0_bits_ctrl_fuType),
    .io_enqRob_req_0_bits_ctrl_fuOpType(dispatch_io_enqRob_req_0_bits_ctrl_fuOpType),
    .io_enqRob_req_0_bits_ctrl_rfWen(dispatch_io_enqRob_req_0_bits_ctrl_rfWen),
    .io_enqRob_req_0_bits_ctrl_fpWen(dispatch_io_enqRob_req_0_bits_ctrl_fpWen),
    .io_enqRob_req_0_bits_ctrl_isXSTrap(dispatch_io_enqRob_req_0_bits_ctrl_isXSTrap),
    .io_enqRob_req_0_bits_ctrl_noSpecExec(dispatch_io_enqRob_req_0_bits_ctrl_noSpecExec),
    .io_enqRob_req_0_bits_ctrl_blockBackward(dispatch_io_enqRob_req_0_bits_ctrl_blockBackward),
    .io_enqRob_req_0_bits_ctrl_flushPipe(dispatch_io_enqRob_req_0_bits_ctrl_flushPipe),
    .io_enqRob_req_0_bits_ctrl_commitType(dispatch_io_enqRob_req_0_bits_ctrl_commitType),
    .io_enqRob_req_0_bits_ctrl_fpu_wflags(dispatch_io_enqRob_req_0_bits_ctrl_fpu_wflags),
    .io_enqRob_req_0_bits_ctrl_isMove(dispatch_io_enqRob_req_0_bits_ctrl_isMove),
    .io_enqRob_req_0_bits_ctrl_singleStep(dispatch_io_enqRob_req_0_bits_ctrl_singleStep),
    .io_enqRob_req_0_bits_pdest(dispatch_io_enqRob_req_0_bits_pdest),
    .io_enqRob_req_0_bits_old_pdest(dispatch_io_enqRob_req_0_bits_old_pdest),
    .io_enqRob_req_0_bits_robIdx_flag(dispatch_io_enqRob_req_0_bits_robIdx_flag),
    .io_enqRob_req_0_bits_robIdx_value(dispatch_io_enqRob_req_0_bits_robIdx_value),
    .io_enqRob_req_0_bits_eliminatedMove(dispatch_io_enqRob_req_0_bits_eliminatedMove),
    .io_enqRob_req_1_valid(dispatch_io_enqRob_req_1_valid),
    .io_enqRob_req_1_bits_cf_exceptionVec_1(dispatch_io_enqRob_req_1_bits_cf_exceptionVec_1),
    .io_enqRob_req_1_bits_cf_exceptionVec_2(dispatch_io_enqRob_req_1_bits_cf_exceptionVec_2),
    .io_enqRob_req_1_bits_cf_exceptionVec_12(dispatch_io_enqRob_req_1_bits_cf_exceptionVec_12),
    .io_enqRob_req_1_bits_cf_trigger_frontendHit_0(dispatch_io_enqRob_req_1_bits_cf_trigger_frontendHit_0),
    .io_enqRob_req_1_bits_cf_trigger_frontendHit_1(dispatch_io_enqRob_req_1_bits_cf_trigger_frontendHit_1),
    .io_enqRob_req_1_bits_cf_trigger_frontendHit_2(dispatch_io_enqRob_req_1_bits_cf_trigger_frontendHit_2),
    .io_enqRob_req_1_bits_cf_trigger_frontendHit_3(dispatch_io_enqRob_req_1_bits_cf_trigger_frontendHit_3),
    .io_enqRob_req_1_bits_cf_pd_isRVC(dispatch_io_enqRob_req_1_bits_cf_pd_isRVC),
    .io_enqRob_req_1_bits_cf_crossPageIPFFix(dispatch_io_enqRob_req_1_bits_cf_crossPageIPFFix),
    .io_enqRob_req_1_bits_cf_loadWaitBit(dispatch_io_enqRob_req_1_bits_cf_loadWaitBit),
    .io_enqRob_req_1_bits_cf_ftqPtr_flag(dispatch_io_enqRob_req_1_bits_cf_ftqPtr_flag),
    .io_enqRob_req_1_bits_cf_ftqPtr_value(dispatch_io_enqRob_req_1_bits_cf_ftqPtr_value),
    .io_enqRob_req_1_bits_cf_ftqOffset(dispatch_io_enqRob_req_1_bits_cf_ftqOffset),
    .io_enqRob_req_1_bits_ctrl_ldest(dispatch_io_enqRob_req_1_bits_ctrl_ldest),
    .io_enqRob_req_1_bits_ctrl_fuType(dispatch_io_enqRob_req_1_bits_ctrl_fuType),
    .io_enqRob_req_1_bits_ctrl_fuOpType(dispatch_io_enqRob_req_1_bits_ctrl_fuOpType),
    .io_enqRob_req_1_bits_ctrl_rfWen(dispatch_io_enqRob_req_1_bits_ctrl_rfWen),
    .io_enqRob_req_1_bits_ctrl_fpWen(dispatch_io_enqRob_req_1_bits_ctrl_fpWen),
    .io_enqRob_req_1_bits_ctrl_isXSTrap(dispatch_io_enqRob_req_1_bits_ctrl_isXSTrap),
    .io_enqRob_req_1_bits_ctrl_noSpecExec(dispatch_io_enqRob_req_1_bits_ctrl_noSpecExec),
    .io_enqRob_req_1_bits_ctrl_blockBackward(dispatch_io_enqRob_req_1_bits_ctrl_blockBackward),
    .io_enqRob_req_1_bits_ctrl_flushPipe(dispatch_io_enqRob_req_1_bits_ctrl_flushPipe),
    .io_enqRob_req_1_bits_ctrl_commitType(dispatch_io_enqRob_req_1_bits_ctrl_commitType),
    .io_enqRob_req_1_bits_ctrl_fpu_wflags(dispatch_io_enqRob_req_1_bits_ctrl_fpu_wflags),
    .io_enqRob_req_1_bits_ctrl_isMove(dispatch_io_enqRob_req_1_bits_ctrl_isMove),
    .io_enqRob_req_1_bits_ctrl_singleStep(dispatch_io_enqRob_req_1_bits_ctrl_singleStep),
    .io_enqRob_req_1_bits_pdest(dispatch_io_enqRob_req_1_bits_pdest),
    .io_enqRob_req_1_bits_old_pdest(dispatch_io_enqRob_req_1_bits_old_pdest),
    .io_enqRob_req_1_bits_robIdx_flag(dispatch_io_enqRob_req_1_bits_robIdx_flag),
    .io_enqRob_req_1_bits_robIdx_value(dispatch_io_enqRob_req_1_bits_robIdx_value),
    .io_enqRob_req_1_bits_eliminatedMove(dispatch_io_enqRob_req_1_bits_eliminatedMove),
    .io_allocPregs_0_isInt(dispatch_io_allocPregs_0_isInt),
    .io_allocPregs_0_isFp(dispatch_io_allocPregs_0_isFp),
    .io_allocPregs_0_preg(dispatch_io_allocPregs_0_preg),
    .io_allocPregs_1_isInt(dispatch_io_allocPregs_1_isInt),
    .io_allocPregs_1_isFp(dispatch_io_allocPregs_1_isFp),
    .io_allocPregs_1_preg(dispatch_io_allocPregs_1_preg),
    .io_toIntDq_canAccept(dispatch_io_toIntDq_canAccept),
    .io_toIntDq_needAlloc_0(dispatch_io_toIntDq_needAlloc_0),
    .io_toIntDq_needAlloc_1(dispatch_io_toIntDq_needAlloc_1),
    .io_toIntDq_req_0_valid(dispatch_io_toIntDq_req_0_valid),
    .io_toIntDq_req_0_bits_cf_foldpc(dispatch_io_toIntDq_req_0_bits_cf_foldpc),
    .io_toIntDq_req_0_bits_cf_trigger_backendEn_0(dispatch_io_toIntDq_req_0_bits_cf_trigger_backendEn_0),
    .io_toIntDq_req_0_bits_cf_trigger_backendEn_1(dispatch_io_toIntDq_req_0_bits_cf_trigger_backendEn_1),
    .io_toIntDq_req_0_bits_cf_pd_isRVC(dispatch_io_toIntDq_req_0_bits_cf_pd_isRVC),
    .io_toIntDq_req_0_bits_cf_pd_brType(dispatch_io_toIntDq_req_0_bits_cf_pd_brType),
    .io_toIntDq_req_0_bits_cf_pd_isCall(dispatch_io_toIntDq_req_0_bits_cf_pd_isCall),
    .io_toIntDq_req_0_bits_cf_pd_isRet(dispatch_io_toIntDq_req_0_bits_cf_pd_isRet),
    .io_toIntDq_req_0_bits_cf_pred_taken(dispatch_io_toIntDq_req_0_bits_cf_pred_taken),
    .io_toIntDq_req_0_bits_cf_storeSetHit(dispatch_io_toIntDq_req_0_bits_cf_storeSetHit),
    .io_toIntDq_req_0_bits_cf_waitForRobIdx_flag(dispatch_io_toIntDq_req_0_bits_cf_waitForRobIdx_flag),
    .io_toIntDq_req_0_bits_cf_waitForRobIdx_value(dispatch_io_toIntDq_req_0_bits_cf_waitForRobIdx_value),
    .io_toIntDq_req_0_bits_cf_loadWaitBit(dispatch_io_toIntDq_req_0_bits_cf_loadWaitBit),
    .io_toIntDq_req_0_bits_cf_loadWaitStrict(dispatch_io_toIntDq_req_0_bits_cf_loadWaitStrict),
    .io_toIntDq_req_0_bits_cf_ssid(dispatch_io_toIntDq_req_0_bits_cf_ssid),
    .io_toIntDq_req_0_bits_cf_ftqPtr_flag(dispatch_io_toIntDq_req_0_bits_cf_ftqPtr_flag),
    .io_toIntDq_req_0_bits_cf_ftqPtr_value(dispatch_io_toIntDq_req_0_bits_cf_ftqPtr_value),
    .io_toIntDq_req_0_bits_cf_ftqOffset(dispatch_io_toIntDq_req_0_bits_cf_ftqOffset),
    .io_toIntDq_req_0_bits_ctrl_srcType_0(dispatch_io_toIntDq_req_0_bits_ctrl_srcType_0),
    .io_toIntDq_req_0_bits_ctrl_srcType_1(dispatch_io_toIntDq_req_0_bits_ctrl_srcType_1),
    .io_toIntDq_req_0_bits_ctrl_srcType_2(dispatch_io_toIntDq_req_0_bits_ctrl_srcType_2),
    .io_toIntDq_req_0_bits_ctrl_fuType(dispatch_io_toIntDq_req_0_bits_ctrl_fuType),
    .io_toIntDq_req_0_bits_ctrl_fuOpType(dispatch_io_toIntDq_req_0_bits_ctrl_fuOpType),
    .io_toIntDq_req_0_bits_ctrl_rfWen(dispatch_io_toIntDq_req_0_bits_ctrl_rfWen),
    .io_toIntDq_req_0_bits_ctrl_fpWen(dispatch_io_toIntDq_req_0_bits_ctrl_fpWen),
    .io_toIntDq_req_0_bits_ctrl_flushPipe(dispatch_io_toIntDq_req_0_bits_ctrl_flushPipe),
    .io_toIntDq_req_0_bits_ctrl_selImm(dispatch_io_toIntDq_req_0_bits_ctrl_selImm),
    .io_toIntDq_req_0_bits_ctrl_imm(dispatch_io_toIntDq_req_0_bits_ctrl_imm),
    .io_toIntDq_req_0_bits_ctrl_fpu_isAddSub(dispatch_io_toIntDq_req_0_bits_ctrl_fpu_isAddSub),
    .io_toIntDq_req_0_bits_ctrl_fpu_typeTagIn(dispatch_io_toIntDq_req_0_bits_ctrl_fpu_typeTagIn),
    .io_toIntDq_req_0_bits_ctrl_fpu_typeTagOut(dispatch_io_toIntDq_req_0_bits_ctrl_fpu_typeTagOut),
    .io_toIntDq_req_0_bits_ctrl_fpu_fromInt(dispatch_io_toIntDq_req_0_bits_ctrl_fpu_fromInt),
    .io_toIntDq_req_0_bits_ctrl_fpu_wflags(dispatch_io_toIntDq_req_0_bits_ctrl_fpu_wflags),
    .io_toIntDq_req_0_bits_ctrl_fpu_fpWen(dispatch_io_toIntDq_req_0_bits_ctrl_fpu_fpWen),
    .io_toIntDq_req_0_bits_ctrl_fpu_fmaCmd(dispatch_io_toIntDq_req_0_bits_ctrl_fpu_fmaCmd),
    .io_toIntDq_req_0_bits_ctrl_fpu_div(dispatch_io_toIntDq_req_0_bits_ctrl_fpu_div),
    .io_toIntDq_req_0_bits_ctrl_fpu_sqrt(dispatch_io_toIntDq_req_0_bits_ctrl_fpu_sqrt),
    .io_toIntDq_req_0_bits_ctrl_fpu_fcvt(dispatch_io_toIntDq_req_0_bits_ctrl_fpu_fcvt),
    .io_toIntDq_req_0_bits_ctrl_fpu_typ(dispatch_io_toIntDq_req_0_bits_ctrl_fpu_typ),
    .io_toIntDq_req_0_bits_ctrl_fpu_fmt(dispatch_io_toIntDq_req_0_bits_ctrl_fpu_fmt),
    .io_toIntDq_req_0_bits_ctrl_fpu_ren3(dispatch_io_toIntDq_req_0_bits_ctrl_fpu_ren3),
    .io_toIntDq_req_0_bits_ctrl_fpu_rm(dispatch_io_toIntDq_req_0_bits_ctrl_fpu_rm),
    .io_toIntDq_req_0_bits_psrc_0(dispatch_io_toIntDq_req_0_bits_psrc_0),
    .io_toIntDq_req_0_bits_psrc_1(dispatch_io_toIntDq_req_0_bits_psrc_1),
    .io_toIntDq_req_0_bits_psrc_2(dispatch_io_toIntDq_req_0_bits_psrc_2),
    .io_toIntDq_req_0_bits_pdest(dispatch_io_toIntDq_req_0_bits_pdest),
    .io_toIntDq_req_0_bits_robIdx_flag(dispatch_io_toIntDq_req_0_bits_robIdx_flag),
    .io_toIntDq_req_0_bits_robIdx_value(dispatch_io_toIntDq_req_0_bits_robIdx_value),
    .io_toIntDq_req_1_valid(dispatch_io_toIntDq_req_1_valid),
    .io_toIntDq_req_1_bits_cf_foldpc(dispatch_io_toIntDq_req_1_bits_cf_foldpc),
    .io_toIntDq_req_1_bits_cf_trigger_backendEn_0(dispatch_io_toIntDq_req_1_bits_cf_trigger_backendEn_0),
    .io_toIntDq_req_1_bits_cf_trigger_backendEn_1(dispatch_io_toIntDq_req_1_bits_cf_trigger_backendEn_1),
    .io_toIntDq_req_1_bits_cf_pd_isRVC(dispatch_io_toIntDq_req_1_bits_cf_pd_isRVC),
    .io_toIntDq_req_1_bits_cf_pd_brType(dispatch_io_toIntDq_req_1_bits_cf_pd_brType),
    .io_toIntDq_req_1_bits_cf_pd_isCall(dispatch_io_toIntDq_req_1_bits_cf_pd_isCall),
    .io_toIntDq_req_1_bits_cf_pd_isRet(dispatch_io_toIntDq_req_1_bits_cf_pd_isRet),
    .io_toIntDq_req_1_bits_cf_pred_taken(dispatch_io_toIntDq_req_1_bits_cf_pred_taken),
    .io_toIntDq_req_1_bits_cf_storeSetHit(dispatch_io_toIntDq_req_1_bits_cf_storeSetHit),
    .io_toIntDq_req_1_bits_cf_waitForRobIdx_flag(dispatch_io_toIntDq_req_1_bits_cf_waitForRobIdx_flag),
    .io_toIntDq_req_1_bits_cf_waitForRobIdx_value(dispatch_io_toIntDq_req_1_bits_cf_waitForRobIdx_value),
    .io_toIntDq_req_1_bits_cf_loadWaitBit(dispatch_io_toIntDq_req_1_bits_cf_loadWaitBit),
    .io_toIntDq_req_1_bits_cf_loadWaitStrict(dispatch_io_toIntDq_req_1_bits_cf_loadWaitStrict),
    .io_toIntDq_req_1_bits_cf_ssid(dispatch_io_toIntDq_req_1_bits_cf_ssid),
    .io_toIntDq_req_1_bits_cf_ftqPtr_flag(dispatch_io_toIntDq_req_1_bits_cf_ftqPtr_flag),
    .io_toIntDq_req_1_bits_cf_ftqPtr_value(dispatch_io_toIntDq_req_1_bits_cf_ftqPtr_value),
    .io_toIntDq_req_1_bits_cf_ftqOffset(dispatch_io_toIntDq_req_1_bits_cf_ftqOffset),
    .io_toIntDq_req_1_bits_ctrl_srcType_0(dispatch_io_toIntDq_req_1_bits_ctrl_srcType_0),
    .io_toIntDq_req_1_bits_ctrl_srcType_1(dispatch_io_toIntDq_req_1_bits_ctrl_srcType_1),
    .io_toIntDq_req_1_bits_ctrl_srcType_2(dispatch_io_toIntDq_req_1_bits_ctrl_srcType_2),
    .io_toIntDq_req_1_bits_ctrl_fuType(dispatch_io_toIntDq_req_1_bits_ctrl_fuType),
    .io_toIntDq_req_1_bits_ctrl_fuOpType(dispatch_io_toIntDq_req_1_bits_ctrl_fuOpType),
    .io_toIntDq_req_1_bits_ctrl_rfWen(dispatch_io_toIntDq_req_1_bits_ctrl_rfWen),
    .io_toIntDq_req_1_bits_ctrl_fpWen(dispatch_io_toIntDq_req_1_bits_ctrl_fpWen),
    .io_toIntDq_req_1_bits_ctrl_flushPipe(dispatch_io_toIntDq_req_1_bits_ctrl_flushPipe),
    .io_toIntDq_req_1_bits_ctrl_selImm(dispatch_io_toIntDq_req_1_bits_ctrl_selImm),
    .io_toIntDq_req_1_bits_ctrl_imm(dispatch_io_toIntDq_req_1_bits_ctrl_imm),
    .io_toIntDq_req_1_bits_ctrl_fpu_isAddSub(dispatch_io_toIntDq_req_1_bits_ctrl_fpu_isAddSub),
    .io_toIntDq_req_1_bits_ctrl_fpu_typeTagIn(dispatch_io_toIntDq_req_1_bits_ctrl_fpu_typeTagIn),
    .io_toIntDq_req_1_bits_ctrl_fpu_typeTagOut(dispatch_io_toIntDq_req_1_bits_ctrl_fpu_typeTagOut),
    .io_toIntDq_req_1_bits_ctrl_fpu_fromInt(dispatch_io_toIntDq_req_1_bits_ctrl_fpu_fromInt),
    .io_toIntDq_req_1_bits_ctrl_fpu_wflags(dispatch_io_toIntDq_req_1_bits_ctrl_fpu_wflags),
    .io_toIntDq_req_1_bits_ctrl_fpu_fpWen(dispatch_io_toIntDq_req_1_bits_ctrl_fpu_fpWen),
    .io_toIntDq_req_1_bits_ctrl_fpu_fmaCmd(dispatch_io_toIntDq_req_1_bits_ctrl_fpu_fmaCmd),
    .io_toIntDq_req_1_bits_ctrl_fpu_div(dispatch_io_toIntDq_req_1_bits_ctrl_fpu_div),
    .io_toIntDq_req_1_bits_ctrl_fpu_sqrt(dispatch_io_toIntDq_req_1_bits_ctrl_fpu_sqrt),
    .io_toIntDq_req_1_bits_ctrl_fpu_fcvt(dispatch_io_toIntDq_req_1_bits_ctrl_fpu_fcvt),
    .io_toIntDq_req_1_bits_ctrl_fpu_typ(dispatch_io_toIntDq_req_1_bits_ctrl_fpu_typ),
    .io_toIntDq_req_1_bits_ctrl_fpu_fmt(dispatch_io_toIntDq_req_1_bits_ctrl_fpu_fmt),
    .io_toIntDq_req_1_bits_ctrl_fpu_ren3(dispatch_io_toIntDq_req_1_bits_ctrl_fpu_ren3),
    .io_toIntDq_req_1_bits_ctrl_fpu_rm(dispatch_io_toIntDq_req_1_bits_ctrl_fpu_rm),
    .io_toIntDq_req_1_bits_psrc_0(dispatch_io_toIntDq_req_1_bits_psrc_0),
    .io_toIntDq_req_1_bits_psrc_1(dispatch_io_toIntDq_req_1_bits_psrc_1),
    .io_toIntDq_req_1_bits_psrc_2(dispatch_io_toIntDq_req_1_bits_psrc_2),
    .io_toIntDq_req_1_bits_pdest(dispatch_io_toIntDq_req_1_bits_pdest),
    .io_toIntDq_req_1_bits_robIdx_flag(dispatch_io_toIntDq_req_1_bits_robIdx_flag),
    .io_toIntDq_req_1_bits_robIdx_value(dispatch_io_toIntDq_req_1_bits_robIdx_value),
    .io_toFpDq_canAccept(dispatch_io_toFpDq_canAccept),
    .io_toFpDq_needAlloc_0(dispatch_io_toFpDq_needAlloc_0),
    .io_toFpDq_needAlloc_1(dispatch_io_toFpDq_needAlloc_1),
    .io_toFpDq_req_0_valid(dispatch_io_toFpDq_req_0_valid),
    .io_toFpDq_req_0_bits_cf_foldpc(dispatch_io_toFpDq_req_0_bits_cf_foldpc),
    .io_toFpDq_req_0_bits_cf_trigger_backendEn_0(dispatch_io_toFpDq_req_0_bits_cf_trigger_backendEn_0),
    .io_toFpDq_req_0_bits_cf_trigger_backendEn_1(dispatch_io_toFpDq_req_0_bits_cf_trigger_backendEn_1),
    .io_toFpDq_req_0_bits_cf_pd_isRVC(dispatch_io_toFpDq_req_0_bits_cf_pd_isRVC),
    .io_toFpDq_req_0_bits_cf_pd_brType(dispatch_io_toFpDq_req_0_bits_cf_pd_brType),
    .io_toFpDq_req_0_bits_cf_pd_isCall(dispatch_io_toFpDq_req_0_bits_cf_pd_isCall),
    .io_toFpDq_req_0_bits_cf_pd_isRet(dispatch_io_toFpDq_req_0_bits_cf_pd_isRet),
    .io_toFpDq_req_0_bits_cf_pred_taken(dispatch_io_toFpDq_req_0_bits_cf_pred_taken),
    .io_toFpDq_req_0_bits_cf_storeSetHit(dispatch_io_toFpDq_req_0_bits_cf_storeSetHit),
    .io_toFpDq_req_0_bits_cf_waitForRobIdx_flag(dispatch_io_toFpDq_req_0_bits_cf_waitForRobIdx_flag),
    .io_toFpDq_req_0_bits_cf_waitForRobIdx_value(dispatch_io_toFpDq_req_0_bits_cf_waitForRobIdx_value),
    .io_toFpDq_req_0_bits_cf_loadWaitBit(dispatch_io_toFpDq_req_0_bits_cf_loadWaitBit),
    .io_toFpDq_req_0_bits_cf_loadWaitStrict(dispatch_io_toFpDq_req_0_bits_cf_loadWaitStrict),
    .io_toFpDq_req_0_bits_cf_ssid(dispatch_io_toFpDq_req_0_bits_cf_ssid),
    .io_toFpDq_req_0_bits_cf_ftqPtr_flag(dispatch_io_toFpDq_req_0_bits_cf_ftqPtr_flag),
    .io_toFpDq_req_0_bits_cf_ftqPtr_value(dispatch_io_toFpDq_req_0_bits_cf_ftqPtr_value),
    .io_toFpDq_req_0_bits_cf_ftqOffset(dispatch_io_toFpDq_req_0_bits_cf_ftqOffset),
    .io_toFpDq_req_0_bits_ctrl_srcType_0(dispatch_io_toFpDq_req_0_bits_ctrl_srcType_0),
    .io_toFpDq_req_0_bits_ctrl_srcType_1(dispatch_io_toFpDq_req_0_bits_ctrl_srcType_1),
    .io_toFpDq_req_0_bits_ctrl_srcType_2(dispatch_io_toFpDq_req_0_bits_ctrl_srcType_2),
    .io_toFpDq_req_0_bits_ctrl_fuType(dispatch_io_toFpDq_req_0_bits_ctrl_fuType),
    .io_toFpDq_req_0_bits_ctrl_fuOpType(dispatch_io_toFpDq_req_0_bits_ctrl_fuOpType),
    .io_toFpDq_req_0_bits_ctrl_rfWen(dispatch_io_toFpDq_req_0_bits_ctrl_rfWen),
    .io_toFpDq_req_0_bits_ctrl_fpWen(dispatch_io_toFpDq_req_0_bits_ctrl_fpWen),
    .io_toFpDq_req_0_bits_ctrl_flushPipe(dispatch_io_toFpDq_req_0_bits_ctrl_flushPipe),
    .io_toFpDq_req_0_bits_ctrl_selImm(dispatch_io_toFpDq_req_0_bits_ctrl_selImm),
    .io_toFpDq_req_0_bits_ctrl_imm(dispatch_io_toFpDq_req_0_bits_ctrl_imm),
    .io_toFpDq_req_0_bits_ctrl_fpu_isAddSub(dispatch_io_toFpDq_req_0_bits_ctrl_fpu_isAddSub),
    .io_toFpDq_req_0_bits_ctrl_fpu_typeTagIn(dispatch_io_toFpDq_req_0_bits_ctrl_fpu_typeTagIn),
    .io_toFpDq_req_0_bits_ctrl_fpu_typeTagOut(dispatch_io_toFpDq_req_0_bits_ctrl_fpu_typeTagOut),
    .io_toFpDq_req_0_bits_ctrl_fpu_fromInt(dispatch_io_toFpDq_req_0_bits_ctrl_fpu_fromInt),
    .io_toFpDq_req_0_bits_ctrl_fpu_wflags(dispatch_io_toFpDq_req_0_bits_ctrl_fpu_wflags),
    .io_toFpDq_req_0_bits_ctrl_fpu_fpWen(dispatch_io_toFpDq_req_0_bits_ctrl_fpu_fpWen),
    .io_toFpDq_req_0_bits_ctrl_fpu_fmaCmd(dispatch_io_toFpDq_req_0_bits_ctrl_fpu_fmaCmd),
    .io_toFpDq_req_0_bits_ctrl_fpu_div(dispatch_io_toFpDq_req_0_bits_ctrl_fpu_div),
    .io_toFpDq_req_0_bits_ctrl_fpu_sqrt(dispatch_io_toFpDq_req_0_bits_ctrl_fpu_sqrt),
    .io_toFpDq_req_0_bits_ctrl_fpu_fcvt(dispatch_io_toFpDq_req_0_bits_ctrl_fpu_fcvt),
    .io_toFpDq_req_0_bits_ctrl_fpu_typ(dispatch_io_toFpDq_req_0_bits_ctrl_fpu_typ),
    .io_toFpDq_req_0_bits_ctrl_fpu_fmt(dispatch_io_toFpDq_req_0_bits_ctrl_fpu_fmt),
    .io_toFpDq_req_0_bits_ctrl_fpu_ren3(dispatch_io_toFpDq_req_0_bits_ctrl_fpu_ren3),
    .io_toFpDq_req_0_bits_ctrl_fpu_rm(dispatch_io_toFpDq_req_0_bits_ctrl_fpu_rm),
    .io_toFpDq_req_0_bits_psrc_0(dispatch_io_toFpDq_req_0_bits_psrc_0),
    .io_toFpDq_req_0_bits_psrc_1(dispatch_io_toFpDq_req_0_bits_psrc_1),
    .io_toFpDq_req_0_bits_psrc_2(dispatch_io_toFpDq_req_0_bits_psrc_2),
    .io_toFpDq_req_0_bits_pdest(dispatch_io_toFpDq_req_0_bits_pdest),
    .io_toFpDq_req_0_bits_robIdx_flag(dispatch_io_toFpDq_req_0_bits_robIdx_flag),
    .io_toFpDq_req_0_bits_robIdx_value(dispatch_io_toFpDq_req_0_bits_robIdx_value),
    .io_toFpDq_req_1_valid(dispatch_io_toFpDq_req_1_valid),
    .io_toFpDq_req_1_bits_cf_foldpc(dispatch_io_toFpDq_req_1_bits_cf_foldpc),
    .io_toFpDq_req_1_bits_cf_trigger_backendEn_0(dispatch_io_toFpDq_req_1_bits_cf_trigger_backendEn_0),
    .io_toFpDq_req_1_bits_cf_trigger_backendEn_1(dispatch_io_toFpDq_req_1_bits_cf_trigger_backendEn_1),
    .io_toFpDq_req_1_bits_cf_pd_isRVC(dispatch_io_toFpDq_req_1_bits_cf_pd_isRVC),
    .io_toFpDq_req_1_bits_cf_pd_brType(dispatch_io_toFpDq_req_1_bits_cf_pd_brType),
    .io_toFpDq_req_1_bits_cf_pd_isCall(dispatch_io_toFpDq_req_1_bits_cf_pd_isCall),
    .io_toFpDq_req_1_bits_cf_pd_isRet(dispatch_io_toFpDq_req_1_bits_cf_pd_isRet),
    .io_toFpDq_req_1_bits_cf_pred_taken(dispatch_io_toFpDq_req_1_bits_cf_pred_taken),
    .io_toFpDq_req_1_bits_cf_storeSetHit(dispatch_io_toFpDq_req_1_bits_cf_storeSetHit),
    .io_toFpDq_req_1_bits_cf_waitForRobIdx_flag(dispatch_io_toFpDq_req_1_bits_cf_waitForRobIdx_flag),
    .io_toFpDq_req_1_bits_cf_waitForRobIdx_value(dispatch_io_toFpDq_req_1_bits_cf_waitForRobIdx_value),
    .io_toFpDq_req_1_bits_cf_loadWaitBit(dispatch_io_toFpDq_req_1_bits_cf_loadWaitBit),
    .io_toFpDq_req_1_bits_cf_loadWaitStrict(dispatch_io_toFpDq_req_1_bits_cf_loadWaitStrict),
    .io_toFpDq_req_1_bits_cf_ssid(dispatch_io_toFpDq_req_1_bits_cf_ssid),
    .io_toFpDq_req_1_bits_cf_ftqPtr_flag(dispatch_io_toFpDq_req_1_bits_cf_ftqPtr_flag),
    .io_toFpDq_req_1_bits_cf_ftqPtr_value(dispatch_io_toFpDq_req_1_bits_cf_ftqPtr_value),
    .io_toFpDq_req_1_bits_cf_ftqOffset(dispatch_io_toFpDq_req_1_bits_cf_ftqOffset),
    .io_toFpDq_req_1_bits_ctrl_srcType_0(dispatch_io_toFpDq_req_1_bits_ctrl_srcType_0),
    .io_toFpDq_req_1_bits_ctrl_srcType_1(dispatch_io_toFpDq_req_1_bits_ctrl_srcType_1),
    .io_toFpDq_req_1_bits_ctrl_srcType_2(dispatch_io_toFpDq_req_1_bits_ctrl_srcType_2),
    .io_toFpDq_req_1_bits_ctrl_fuType(dispatch_io_toFpDq_req_1_bits_ctrl_fuType),
    .io_toFpDq_req_1_bits_ctrl_fuOpType(dispatch_io_toFpDq_req_1_bits_ctrl_fuOpType),
    .io_toFpDq_req_1_bits_ctrl_rfWen(dispatch_io_toFpDq_req_1_bits_ctrl_rfWen),
    .io_toFpDq_req_1_bits_ctrl_fpWen(dispatch_io_toFpDq_req_1_bits_ctrl_fpWen),
    .io_toFpDq_req_1_bits_ctrl_flushPipe(dispatch_io_toFpDq_req_1_bits_ctrl_flushPipe),
    .io_toFpDq_req_1_bits_ctrl_selImm(dispatch_io_toFpDq_req_1_bits_ctrl_selImm),
    .io_toFpDq_req_1_bits_ctrl_imm(dispatch_io_toFpDq_req_1_bits_ctrl_imm),
    .io_toFpDq_req_1_bits_ctrl_fpu_isAddSub(dispatch_io_toFpDq_req_1_bits_ctrl_fpu_isAddSub),
    .io_toFpDq_req_1_bits_ctrl_fpu_typeTagIn(dispatch_io_toFpDq_req_1_bits_ctrl_fpu_typeTagIn),
    .io_toFpDq_req_1_bits_ctrl_fpu_typeTagOut(dispatch_io_toFpDq_req_1_bits_ctrl_fpu_typeTagOut),
    .io_toFpDq_req_1_bits_ctrl_fpu_fromInt(dispatch_io_toFpDq_req_1_bits_ctrl_fpu_fromInt),
    .io_toFpDq_req_1_bits_ctrl_fpu_wflags(dispatch_io_toFpDq_req_1_bits_ctrl_fpu_wflags),
    .io_toFpDq_req_1_bits_ctrl_fpu_fpWen(dispatch_io_toFpDq_req_1_bits_ctrl_fpu_fpWen),
    .io_toFpDq_req_1_bits_ctrl_fpu_fmaCmd(dispatch_io_toFpDq_req_1_bits_ctrl_fpu_fmaCmd),
    .io_toFpDq_req_1_bits_ctrl_fpu_div(dispatch_io_toFpDq_req_1_bits_ctrl_fpu_div),
    .io_toFpDq_req_1_bits_ctrl_fpu_sqrt(dispatch_io_toFpDq_req_1_bits_ctrl_fpu_sqrt),
    .io_toFpDq_req_1_bits_ctrl_fpu_fcvt(dispatch_io_toFpDq_req_1_bits_ctrl_fpu_fcvt),
    .io_toFpDq_req_1_bits_ctrl_fpu_typ(dispatch_io_toFpDq_req_1_bits_ctrl_fpu_typ),
    .io_toFpDq_req_1_bits_ctrl_fpu_fmt(dispatch_io_toFpDq_req_1_bits_ctrl_fpu_fmt),
    .io_toFpDq_req_1_bits_ctrl_fpu_ren3(dispatch_io_toFpDq_req_1_bits_ctrl_fpu_ren3),
    .io_toFpDq_req_1_bits_ctrl_fpu_rm(dispatch_io_toFpDq_req_1_bits_ctrl_fpu_rm),
    .io_toFpDq_req_1_bits_psrc_0(dispatch_io_toFpDq_req_1_bits_psrc_0),
    .io_toFpDq_req_1_bits_psrc_1(dispatch_io_toFpDq_req_1_bits_psrc_1),
    .io_toFpDq_req_1_bits_psrc_2(dispatch_io_toFpDq_req_1_bits_psrc_2),
    .io_toFpDq_req_1_bits_pdest(dispatch_io_toFpDq_req_1_bits_pdest),
    .io_toFpDq_req_1_bits_robIdx_flag(dispatch_io_toFpDq_req_1_bits_robIdx_flag),
    .io_toFpDq_req_1_bits_robIdx_value(dispatch_io_toFpDq_req_1_bits_robIdx_value),
    .io_toLsDq_canAccept(dispatch_io_toLsDq_canAccept),
    .io_toLsDq_needAlloc_0(dispatch_io_toLsDq_needAlloc_0),
    .io_toLsDq_needAlloc_1(dispatch_io_toLsDq_needAlloc_1),
    .io_toLsDq_req_0_valid(dispatch_io_toLsDq_req_0_valid),
    .io_toLsDq_req_0_bits_cf_foldpc(dispatch_io_toLsDq_req_0_bits_cf_foldpc),
    .io_toLsDq_req_0_bits_cf_trigger_backendEn_0(dispatch_io_toLsDq_req_0_bits_cf_trigger_backendEn_0),
    .io_toLsDq_req_0_bits_cf_trigger_backendEn_1(dispatch_io_toLsDq_req_0_bits_cf_trigger_backendEn_1),
    .io_toLsDq_req_0_bits_cf_pd_isRVC(dispatch_io_toLsDq_req_0_bits_cf_pd_isRVC),
    .io_toLsDq_req_0_bits_cf_pd_brType(dispatch_io_toLsDq_req_0_bits_cf_pd_brType),
    .io_toLsDq_req_0_bits_cf_pd_isCall(dispatch_io_toLsDq_req_0_bits_cf_pd_isCall),
    .io_toLsDq_req_0_bits_cf_pd_isRet(dispatch_io_toLsDq_req_0_bits_cf_pd_isRet),
    .io_toLsDq_req_0_bits_cf_pred_taken(dispatch_io_toLsDq_req_0_bits_cf_pred_taken),
    .io_toLsDq_req_0_bits_cf_storeSetHit(dispatch_io_toLsDq_req_0_bits_cf_storeSetHit),
    .io_toLsDq_req_0_bits_cf_waitForRobIdx_flag(dispatch_io_toLsDq_req_0_bits_cf_waitForRobIdx_flag),
    .io_toLsDq_req_0_bits_cf_waitForRobIdx_value(dispatch_io_toLsDq_req_0_bits_cf_waitForRobIdx_value),
    .io_toLsDq_req_0_bits_cf_loadWaitBit(dispatch_io_toLsDq_req_0_bits_cf_loadWaitBit),
    .io_toLsDq_req_0_bits_cf_loadWaitStrict(dispatch_io_toLsDq_req_0_bits_cf_loadWaitStrict),
    .io_toLsDq_req_0_bits_cf_ssid(dispatch_io_toLsDq_req_0_bits_cf_ssid),
    .io_toLsDq_req_0_bits_cf_ftqPtr_flag(dispatch_io_toLsDq_req_0_bits_cf_ftqPtr_flag),
    .io_toLsDq_req_0_bits_cf_ftqPtr_value(dispatch_io_toLsDq_req_0_bits_cf_ftqPtr_value),
    .io_toLsDq_req_0_bits_cf_ftqOffset(dispatch_io_toLsDq_req_0_bits_cf_ftqOffset),
    .io_toLsDq_req_0_bits_ctrl_srcType_0(dispatch_io_toLsDq_req_0_bits_ctrl_srcType_0),
    .io_toLsDq_req_0_bits_ctrl_srcType_1(dispatch_io_toLsDq_req_0_bits_ctrl_srcType_1),
    .io_toLsDq_req_0_bits_ctrl_srcType_2(dispatch_io_toLsDq_req_0_bits_ctrl_srcType_2),
    .io_toLsDq_req_0_bits_ctrl_fuType(dispatch_io_toLsDq_req_0_bits_ctrl_fuType),
    .io_toLsDq_req_0_bits_ctrl_fuOpType(dispatch_io_toLsDq_req_0_bits_ctrl_fuOpType),
    .io_toLsDq_req_0_bits_ctrl_rfWen(dispatch_io_toLsDq_req_0_bits_ctrl_rfWen),
    .io_toLsDq_req_0_bits_ctrl_fpWen(dispatch_io_toLsDq_req_0_bits_ctrl_fpWen),
    .io_toLsDq_req_0_bits_ctrl_flushPipe(dispatch_io_toLsDq_req_0_bits_ctrl_flushPipe),
    .io_toLsDq_req_0_bits_ctrl_selImm(dispatch_io_toLsDq_req_0_bits_ctrl_selImm),
    .io_toLsDq_req_0_bits_ctrl_imm(dispatch_io_toLsDq_req_0_bits_ctrl_imm),
    .io_toLsDq_req_0_bits_ctrl_fpu_isAddSub(dispatch_io_toLsDq_req_0_bits_ctrl_fpu_isAddSub),
    .io_toLsDq_req_0_bits_ctrl_fpu_typeTagIn(dispatch_io_toLsDq_req_0_bits_ctrl_fpu_typeTagIn),
    .io_toLsDq_req_0_bits_ctrl_fpu_typeTagOut(dispatch_io_toLsDq_req_0_bits_ctrl_fpu_typeTagOut),
    .io_toLsDq_req_0_bits_ctrl_fpu_fromInt(dispatch_io_toLsDq_req_0_bits_ctrl_fpu_fromInt),
    .io_toLsDq_req_0_bits_ctrl_fpu_wflags(dispatch_io_toLsDq_req_0_bits_ctrl_fpu_wflags),
    .io_toLsDq_req_0_bits_ctrl_fpu_fpWen(dispatch_io_toLsDq_req_0_bits_ctrl_fpu_fpWen),
    .io_toLsDq_req_0_bits_ctrl_fpu_fmaCmd(dispatch_io_toLsDq_req_0_bits_ctrl_fpu_fmaCmd),
    .io_toLsDq_req_0_bits_ctrl_fpu_div(dispatch_io_toLsDq_req_0_bits_ctrl_fpu_div),
    .io_toLsDq_req_0_bits_ctrl_fpu_sqrt(dispatch_io_toLsDq_req_0_bits_ctrl_fpu_sqrt),
    .io_toLsDq_req_0_bits_ctrl_fpu_fcvt(dispatch_io_toLsDq_req_0_bits_ctrl_fpu_fcvt),
    .io_toLsDq_req_0_bits_ctrl_fpu_typ(dispatch_io_toLsDq_req_0_bits_ctrl_fpu_typ),
    .io_toLsDq_req_0_bits_ctrl_fpu_fmt(dispatch_io_toLsDq_req_0_bits_ctrl_fpu_fmt),
    .io_toLsDq_req_0_bits_ctrl_fpu_ren3(dispatch_io_toLsDq_req_0_bits_ctrl_fpu_ren3),
    .io_toLsDq_req_0_bits_ctrl_fpu_rm(dispatch_io_toLsDq_req_0_bits_ctrl_fpu_rm),
    .io_toLsDq_req_0_bits_psrc_0(dispatch_io_toLsDq_req_0_bits_psrc_0),
    .io_toLsDq_req_0_bits_psrc_1(dispatch_io_toLsDq_req_0_bits_psrc_1),
    .io_toLsDq_req_0_bits_psrc_2(dispatch_io_toLsDq_req_0_bits_psrc_2),
    .io_toLsDq_req_0_bits_pdest(dispatch_io_toLsDq_req_0_bits_pdest),
    .io_toLsDq_req_0_bits_robIdx_flag(dispatch_io_toLsDq_req_0_bits_robIdx_flag),
    .io_toLsDq_req_0_bits_robIdx_value(dispatch_io_toLsDq_req_0_bits_robIdx_value),
    .io_toLsDq_req_1_valid(dispatch_io_toLsDq_req_1_valid),
    .io_toLsDq_req_1_bits_cf_foldpc(dispatch_io_toLsDq_req_1_bits_cf_foldpc),
    .io_toLsDq_req_1_bits_cf_trigger_backendEn_0(dispatch_io_toLsDq_req_1_bits_cf_trigger_backendEn_0),
    .io_toLsDq_req_1_bits_cf_trigger_backendEn_1(dispatch_io_toLsDq_req_1_bits_cf_trigger_backendEn_1),
    .io_toLsDq_req_1_bits_cf_pd_isRVC(dispatch_io_toLsDq_req_1_bits_cf_pd_isRVC),
    .io_toLsDq_req_1_bits_cf_pd_brType(dispatch_io_toLsDq_req_1_bits_cf_pd_brType),
    .io_toLsDq_req_1_bits_cf_pd_isCall(dispatch_io_toLsDq_req_1_bits_cf_pd_isCall),
    .io_toLsDq_req_1_bits_cf_pd_isRet(dispatch_io_toLsDq_req_1_bits_cf_pd_isRet),
    .io_toLsDq_req_1_bits_cf_pred_taken(dispatch_io_toLsDq_req_1_bits_cf_pred_taken),
    .io_toLsDq_req_1_bits_cf_storeSetHit(dispatch_io_toLsDq_req_1_bits_cf_storeSetHit),
    .io_toLsDq_req_1_bits_cf_waitForRobIdx_flag(dispatch_io_toLsDq_req_1_bits_cf_waitForRobIdx_flag),
    .io_toLsDq_req_1_bits_cf_waitForRobIdx_value(dispatch_io_toLsDq_req_1_bits_cf_waitForRobIdx_value),
    .io_toLsDq_req_1_bits_cf_loadWaitBit(dispatch_io_toLsDq_req_1_bits_cf_loadWaitBit),
    .io_toLsDq_req_1_bits_cf_loadWaitStrict(dispatch_io_toLsDq_req_1_bits_cf_loadWaitStrict),
    .io_toLsDq_req_1_bits_cf_ssid(dispatch_io_toLsDq_req_1_bits_cf_ssid),
    .io_toLsDq_req_1_bits_cf_ftqPtr_flag(dispatch_io_toLsDq_req_1_bits_cf_ftqPtr_flag),
    .io_toLsDq_req_1_bits_cf_ftqPtr_value(dispatch_io_toLsDq_req_1_bits_cf_ftqPtr_value),
    .io_toLsDq_req_1_bits_cf_ftqOffset(dispatch_io_toLsDq_req_1_bits_cf_ftqOffset),
    .io_toLsDq_req_1_bits_ctrl_srcType_0(dispatch_io_toLsDq_req_1_bits_ctrl_srcType_0),
    .io_toLsDq_req_1_bits_ctrl_srcType_1(dispatch_io_toLsDq_req_1_bits_ctrl_srcType_1),
    .io_toLsDq_req_1_bits_ctrl_srcType_2(dispatch_io_toLsDq_req_1_bits_ctrl_srcType_2),
    .io_toLsDq_req_1_bits_ctrl_fuType(dispatch_io_toLsDq_req_1_bits_ctrl_fuType),
    .io_toLsDq_req_1_bits_ctrl_fuOpType(dispatch_io_toLsDq_req_1_bits_ctrl_fuOpType),
    .io_toLsDq_req_1_bits_ctrl_rfWen(dispatch_io_toLsDq_req_1_bits_ctrl_rfWen),
    .io_toLsDq_req_1_bits_ctrl_fpWen(dispatch_io_toLsDq_req_1_bits_ctrl_fpWen),
    .io_toLsDq_req_1_bits_ctrl_flushPipe(dispatch_io_toLsDq_req_1_bits_ctrl_flushPipe),
    .io_toLsDq_req_1_bits_ctrl_selImm(dispatch_io_toLsDq_req_1_bits_ctrl_selImm),
    .io_toLsDq_req_1_bits_ctrl_imm(dispatch_io_toLsDq_req_1_bits_ctrl_imm),
    .io_toLsDq_req_1_bits_ctrl_fpu_isAddSub(dispatch_io_toLsDq_req_1_bits_ctrl_fpu_isAddSub),
    .io_toLsDq_req_1_bits_ctrl_fpu_typeTagIn(dispatch_io_toLsDq_req_1_bits_ctrl_fpu_typeTagIn),
    .io_toLsDq_req_1_bits_ctrl_fpu_typeTagOut(dispatch_io_toLsDq_req_1_bits_ctrl_fpu_typeTagOut),
    .io_toLsDq_req_1_bits_ctrl_fpu_fromInt(dispatch_io_toLsDq_req_1_bits_ctrl_fpu_fromInt),
    .io_toLsDq_req_1_bits_ctrl_fpu_wflags(dispatch_io_toLsDq_req_1_bits_ctrl_fpu_wflags),
    .io_toLsDq_req_1_bits_ctrl_fpu_fpWen(dispatch_io_toLsDq_req_1_bits_ctrl_fpu_fpWen),
    .io_toLsDq_req_1_bits_ctrl_fpu_fmaCmd(dispatch_io_toLsDq_req_1_bits_ctrl_fpu_fmaCmd),
    .io_toLsDq_req_1_bits_ctrl_fpu_div(dispatch_io_toLsDq_req_1_bits_ctrl_fpu_div),
    .io_toLsDq_req_1_bits_ctrl_fpu_sqrt(dispatch_io_toLsDq_req_1_bits_ctrl_fpu_sqrt),
    .io_toLsDq_req_1_bits_ctrl_fpu_fcvt(dispatch_io_toLsDq_req_1_bits_ctrl_fpu_fcvt),
    .io_toLsDq_req_1_bits_ctrl_fpu_typ(dispatch_io_toLsDq_req_1_bits_ctrl_fpu_typ),
    .io_toLsDq_req_1_bits_ctrl_fpu_fmt(dispatch_io_toLsDq_req_1_bits_ctrl_fpu_fmt),
    .io_toLsDq_req_1_bits_ctrl_fpu_ren3(dispatch_io_toLsDq_req_1_bits_ctrl_fpu_ren3),
    .io_toLsDq_req_1_bits_ctrl_fpu_rm(dispatch_io_toLsDq_req_1_bits_ctrl_fpu_rm),
    .io_toLsDq_req_1_bits_psrc_0(dispatch_io_toLsDq_req_1_bits_psrc_0),
    .io_toLsDq_req_1_bits_psrc_1(dispatch_io_toLsDq_req_1_bits_psrc_1),
    .io_toLsDq_req_1_bits_psrc_2(dispatch_io_toLsDq_req_1_bits_psrc_2),
    .io_toLsDq_req_1_bits_pdest(dispatch_io_toLsDq_req_1_bits_pdest),
    .io_toLsDq_req_1_bits_robIdx_flag(dispatch_io_toLsDq_req_1_bits_robIdx_flag),
    .io_toLsDq_req_1_bits_robIdx_value(dispatch_io_toLsDq_req_1_bits_robIdx_value),
    .io_redirect_valid(dispatch_io_redirect_valid),
    .io_singleStep(dispatch_io_singleStep),
    .io_lfst_req_0_valid(dispatch_io_lfst_req_0_valid),
    .io_lfst_req_0_bits_isstore(dispatch_io_lfst_req_0_bits_isstore),
    .io_lfst_req_0_bits_ssid(dispatch_io_lfst_req_0_bits_ssid),
    .io_lfst_req_0_bits_robIdx_flag(dispatch_io_lfst_req_0_bits_robIdx_flag),
    .io_lfst_req_0_bits_robIdx_value(dispatch_io_lfst_req_0_bits_robIdx_value),
    .io_lfst_req_1_valid(dispatch_io_lfst_req_1_valid),
    .io_lfst_req_1_bits_isstore(dispatch_io_lfst_req_1_bits_isstore),
    .io_lfst_req_1_bits_ssid(dispatch_io_lfst_req_1_bits_ssid),
    .io_lfst_req_1_bits_robIdx_flag(dispatch_io_lfst_req_1_bits_robIdx_flag),
    .io_lfst_req_1_bits_robIdx_value(dispatch_io_lfst_req_1_bits_robIdx_value),
    .io_lfst_resp_0_bits_shouldWait(dispatch_io_lfst_resp_0_bits_shouldWait),
    .io_lfst_resp_0_bits_robIdx_flag(dispatch_io_lfst_resp_0_bits_robIdx_flag),
    .io_lfst_resp_0_bits_robIdx_value(dispatch_io_lfst_resp_0_bits_robIdx_value),
    .io_lfst_resp_1_bits_shouldWait(dispatch_io_lfst_resp_1_bits_shouldWait),
    .io_lfst_resp_1_bits_robIdx_flag(dispatch_io_lfst_resp_1_bits_robIdx_flag),
    .io_lfst_resp_1_bits_robIdx_value(dispatch_io_lfst_resp_1_bits_robIdx_value),
    .io_perf_0_value(dispatch_io_perf_0_value),
    .io_perf_1_value(dispatch_io_perf_1_value),
    .io_perf_2_value(dispatch_io_perf_2_value),
    .io_perf_3_value(dispatch_io_perf_3_value),
    .io_perf_5_value(dispatch_io_perf_5_value),
    .io_perf_6_value(dispatch_io_perf_6_value),
    .io_perf_7_value(dispatch_io_perf_7_value),
    .io_perf_8_value(dispatch_io_perf_8_value)
  );
  DispatchQueue intDq ( // @[CtrlBlock.scala 270:21]
    .clock(intDq_clock),
    .reset(intDq_reset),
    .io_enq_canAccept(intDq_io_enq_canAccept),
    .io_enq_needAlloc_0(intDq_io_enq_needAlloc_0),
    .io_enq_needAlloc_1(intDq_io_enq_needAlloc_1),
    .io_enq_req_0_valid(intDq_io_enq_req_0_valid),
    .io_enq_req_0_bits_cf_foldpc(intDq_io_enq_req_0_bits_cf_foldpc),
    .io_enq_req_0_bits_cf_trigger_backendEn_0(intDq_io_enq_req_0_bits_cf_trigger_backendEn_0),
    .io_enq_req_0_bits_cf_trigger_backendEn_1(intDq_io_enq_req_0_bits_cf_trigger_backendEn_1),
    .io_enq_req_0_bits_cf_pd_isRVC(intDq_io_enq_req_0_bits_cf_pd_isRVC),
    .io_enq_req_0_bits_cf_pd_brType(intDq_io_enq_req_0_bits_cf_pd_brType),
    .io_enq_req_0_bits_cf_pd_isCall(intDq_io_enq_req_0_bits_cf_pd_isCall),
    .io_enq_req_0_bits_cf_pd_isRet(intDq_io_enq_req_0_bits_cf_pd_isRet),
    .io_enq_req_0_bits_cf_pred_taken(intDq_io_enq_req_0_bits_cf_pred_taken),
    .io_enq_req_0_bits_cf_storeSetHit(intDq_io_enq_req_0_bits_cf_storeSetHit),
    .io_enq_req_0_bits_cf_waitForRobIdx_flag(intDq_io_enq_req_0_bits_cf_waitForRobIdx_flag),
    .io_enq_req_0_bits_cf_waitForRobIdx_value(intDq_io_enq_req_0_bits_cf_waitForRobIdx_value),
    .io_enq_req_0_bits_cf_loadWaitBit(intDq_io_enq_req_0_bits_cf_loadWaitBit),
    .io_enq_req_0_bits_cf_loadWaitStrict(intDq_io_enq_req_0_bits_cf_loadWaitStrict),
    .io_enq_req_0_bits_cf_ssid(intDq_io_enq_req_0_bits_cf_ssid),
    .io_enq_req_0_bits_cf_ftqPtr_flag(intDq_io_enq_req_0_bits_cf_ftqPtr_flag),
    .io_enq_req_0_bits_cf_ftqPtr_value(intDq_io_enq_req_0_bits_cf_ftqPtr_value),
    .io_enq_req_0_bits_cf_ftqOffset(intDq_io_enq_req_0_bits_cf_ftqOffset),
    .io_enq_req_0_bits_ctrl_srcType_0(intDq_io_enq_req_0_bits_ctrl_srcType_0),
    .io_enq_req_0_bits_ctrl_srcType_1(intDq_io_enq_req_0_bits_ctrl_srcType_1),
    .io_enq_req_0_bits_ctrl_srcType_2(intDq_io_enq_req_0_bits_ctrl_srcType_2),
    .io_enq_req_0_bits_ctrl_fuType(intDq_io_enq_req_0_bits_ctrl_fuType),
    .io_enq_req_0_bits_ctrl_fuOpType(intDq_io_enq_req_0_bits_ctrl_fuOpType),
    .io_enq_req_0_bits_ctrl_rfWen(intDq_io_enq_req_0_bits_ctrl_rfWen),
    .io_enq_req_0_bits_ctrl_fpWen(intDq_io_enq_req_0_bits_ctrl_fpWen),
    .io_enq_req_0_bits_ctrl_flushPipe(intDq_io_enq_req_0_bits_ctrl_flushPipe),
    .io_enq_req_0_bits_ctrl_selImm(intDq_io_enq_req_0_bits_ctrl_selImm),
    .io_enq_req_0_bits_ctrl_imm(intDq_io_enq_req_0_bits_ctrl_imm),
    .io_enq_req_0_bits_ctrl_fpu_isAddSub(intDq_io_enq_req_0_bits_ctrl_fpu_isAddSub),
    .io_enq_req_0_bits_ctrl_fpu_typeTagIn(intDq_io_enq_req_0_bits_ctrl_fpu_typeTagIn),
    .io_enq_req_0_bits_ctrl_fpu_typeTagOut(intDq_io_enq_req_0_bits_ctrl_fpu_typeTagOut),
    .io_enq_req_0_bits_ctrl_fpu_fromInt(intDq_io_enq_req_0_bits_ctrl_fpu_fromInt),
    .io_enq_req_0_bits_ctrl_fpu_wflags(intDq_io_enq_req_0_bits_ctrl_fpu_wflags),
    .io_enq_req_0_bits_ctrl_fpu_fpWen(intDq_io_enq_req_0_bits_ctrl_fpu_fpWen),
    .io_enq_req_0_bits_ctrl_fpu_fmaCmd(intDq_io_enq_req_0_bits_ctrl_fpu_fmaCmd),
    .io_enq_req_0_bits_ctrl_fpu_div(intDq_io_enq_req_0_bits_ctrl_fpu_div),
    .io_enq_req_0_bits_ctrl_fpu_sqrt(intDq_io_enq_req_0_bits_ctrl_fpu_sqrt),
    .io_enq_req_0_bits_ctrl_fpu_fcvt(intDq_io_enq_req_0_bits_ctrl_fpu_fcvt),
    .io_enq_req_0_bits_ctrl_fpu_typ(intDq_io_enq_req_0_bits_ctrl_fpu_typ),
    .io_enq_req_0_bits_ctrl_fpu_fmt(intDq_io_enq_req_0_bits_ctrl_fpu_fmt),
    .io_enq_req_0_bits_ctrl_fpu_ren3(intDq_io_enq_req_0_bits_ctrl_fpu_ren3),
    .io_enq_req_0_bits_ctrl_fpu_rm(intDq_io_enq_req_0_bits_ctrl_fpu_rm),
    .io_enq_req_0_bits_psrc_0(intDq_io_enq_req_0_bits_psrc_0),
    .io_enq_req_0_bits_psrc_1(intDq_io_enq_req_0_bits_psrc_1),
    .io_enq_req_0_bits_psrc_2(intDq_io_enq_req_0_bits_psrc_2),
    .io_enq_req_0_bits_pdest(intDq_io_enq_req_0_bits_pdest),
    .io_enq_req_0_bits_robIdx_flag(intDq_io_enq_req_0_bits_robIdx_flag),
    .io_enq_req_0_bits_robIdx_value(intDq_io_enq_req_0_bits_robIdx_value),
    .io_enq_req_1_valid(intDq_io_enq_req_1_valid),
    .io_enq_req_1_bits_cf_foldpc(intDq_io_enq_req_1_bits_cf_foldpc),
    .io_enq_req_1_bits_cf_trigger_backendEn_0(intDq_io_enq_req_1_bits_cf_trigger_backendEn_0),
    .io_enq_req_1_bits_cf_trigger_backendEn_1(intDq_io_enq_req_1_bits_cf_trigger_backendEn_1),
    .io_enq_req_1_bits_cf_pd_isRVC(intDq_io_enq_req_1_bits_cf_pd_isRVC),
    .io_enq_req_1_bits_cf_pd_brType(intDq_io_enq_req_1_bits_cf_pd_brType),
    .io_enq_req_1_bits_cf_pd_isCall(intDq_io_enq_req_1_bits_cf_pd_isCall),
    .io_enq_req_1_bits_cf_pd_isRet(intDq_io_enq_req_1_bits_cf_pd_isRet),
    .io_enq_req_1_bits_cf_pred_taken(intDq_io_enq_req_1_bits_cf_pred_taken),
    .io_enq_req_1_bits_cf_storeSetHit(intDq_io_enq_req_1_bits_cf_storeSetHit),
    .io_enq_req_1_bits_cf_waitForRobIdx_flag(intDq_io_enq_req_1_bits_cf_waitForRobIdx_flag),
    .io_enq_req_1_bits_cf_waitForRobIdx_value(intDq_io_enq_req_1_bits_cf_waitForRobIdx_value),
    .io_enq_req_1_bits_cf_loadWaitBit(intDq_io_enq_req_1_bits_cf_loadWaitBit),
    .io_enq_req_1_bits_cf_loadWaitStrict(intDq_io_enq_req_1_bits_cf_loadWaitStrict),
    .io_enq_req_1_bits_cf_ssid(intDq_io_enq_req_1_bits_cf_ssid),
    .io_enq_req_1_bits_cf_ftqPtr_flag(intDq_io_enq_req_1_bits_cf_ftqPtr_flag),
    .io_enq_req_1_bits_cf_ftqPtr_value(intDq_io_enq_req_1_bits_cf_ftqPtr_value),
    .io_enq_req_1_bits_cf_ftqOffset(intDq_io_enq_req_1_bits_cf_ftqOffset),
    .io_enq_req_1_bits_ctrl_srcType_0(intDq_io_enq_req_1_bits_ctrl_srcType_0),
    .io_enq_req_1_bits_ctrl_srcType_1(intDq_io_enq_req_1_bits_ctrl_srcType_1),
    .io_enq_req_1_bits_ctrl_srcType_2(intDq_io_enq_req_1_bits_ctrl_srcType_2),
    .io_enq_req_1_bits_ctrl_fuType(intDq_io_enq_req_1_bits_ctrl_fuType),
    .io_enq_req_1_bits_ctrl_fuOpType(intDq_io_enq_req_1_bits_ctrl_fuOpType),
    .io_enq_req_1_bits_ctrl_rfWen(intDq_io_enq_req_1_bits_ctrl_rfWen),
    .io_enq_req_1_bits_ctrl_fpWen(intDq_io_enq_req_1_bits_ctrl_fpWen),
    .io_enq_req_1_bits_ctrl_flushPipe(intDq_io_enq_req_1_bits_ctrl_flushPipe),
    .io_enq_req_1_bits_ctrl_selImm(intDq_io_enq_req_1_bits_ctrl_selImm),
    .io_enq_req_1_bits_ctrl_imm(intDq_io_enq_req_1_bits_ctrl_imm),
    .io_enq_req_1_bits_ctrl_fpu_isAddSub(intDq_io_enq_req_1_bits_ctrl_fpu_isAddSub),
    .io_enq_req_1_bits_ctrl_fpu_typeTagIn(intDq_io_enq_req_1_bits_ctrl_fpu_typeTagIn),
    .io_enq_req_1_bits_ctrl_fpu_typeTagOut(intDq_io_enq_req_1_bits_ctrl_fpu_typeTagOut),
    .io_enq_req_1_bits_ctrl_fpu_fromInt(intDq_io_enq_req_1_bits_ctrl_fpu_fromInt),
    .io_enq_req_1_bits_ctrl_fpu_wflags(intDq_io_enq_req_1_bits_ctrl_fpu_wflags),
    .io_enq_req_1_bits_ctrl_fpu_fpWen(intDq_io_enq_req_1_bits_ctrl_fpu_fpWen),
    .io_enq_req_1_bits_ctrl_fpu_fmaCmd(intDq_io_enq_req_1_bits_ctrl_fpu_fmaCmd),
    .io_enq_req_1_bits_ctrl_fpu_div(intDq_io_enq_req_1_bits_ctrl_fpu_div),
    .io_enq_req_1_bits_ctrl_fpu_sqrt(intDq_io_enq_req_1_bits_ctrl_fpu_sqrt),
    .io_enq_req_1_bits_ctrl_fpu_fcvt(intDq_io_enq_req_1_bits_ctrl_fpu_fcvt),
    .io_enq_req_1_bits_ctrl_fpu_typ(intDq_io_enq_req_1_bits_ctrl_fpu_typ),
    .io_enq_req_1_bits_ctrl_fpu_fmt(intDq_io_enq_req_1_bits_ctrl_fpu_fmt),
    .io_enq_req_1_bits_ctrl_fpu_ren3(intDq_io_enq_req_1_bits_ctrl_fpu_ren3),
    .io_enq_req_1_bits_ctrl_fpu_rm(intDq_io_enq_req_1_bits_ctrl_fpu_rm),
    .io_enq_req_1_bits_psrc_0(intDq_io_enq_req_1_bits_psrc_0),
    .io_enq_req_1_bits_psrc_1(intDq_io_enq_req_1_bits_psrc_1),
    .io_enq_req_1_bits_psrc_2(intDq_io_enq_req_1_bits_psrc_2),
    .io_enq_req_1_bits_pdest(intDq_io_enq_req_1_bits_pdest),
    .io_enq_req_1_bits_robIdx_flag(intDq_io_enq_req_1_bits_robIdx_flag),
    .io_enq_req_1_bits_robIdx_value(intDq_io_enq_req_1_bits_robIdx_value),
    .io_deq_0_ready(intDq_io_deq_0_ready),
    .io_deq_0_valid(intDq_io_deq_0_valid),
    .io_deq_0_bits_cf_foldpc(intDq_io_deq_0_bits_cf_foldpc),
    .io_deq_0_bits_cf_trigger_backendEn_0(intDq_io_deq_0_bits_cf_trigger_backendEn_0),
    .io_deq_0_bits_cf_trigger_backendEn_1(intDq_io_deq_0_bits_cf_trigger_backendEn_1),
    .io_deq_0_bits_cf_pd_isRVC(intDq_io_deq_0_bits_cf_pd_isRVC),
    .io_deq_0_bits_cf_pd_brType(intDq_io_deq_0_bits_cf_pd_brType),
    .io_deq_0_bits_cf_pd_isCall(intDq_io_deq_0_bits_cf_pd_isCall),
    .io_deq_0_bits_cf_pd_isRet(intDq_io_deq_0_bits_cf_pd_isRet),
    .io_deq_0_bits_cf_pred_taken(intDq_io_deq_0_bits_cf_pred_taken),
    .io_deq_0_bits_cf_storeSetHit(intDq_io_deq_0_bits_cf_storeSetHit),
    .io_deq_0_bits_cf_waitForRobIdx_flag(intDq_io_deq_0_bits_cf_waitForRobIdx_flag),
    .io_deq_0_bits_cf_waitForRobIdx_value(intDq_io_deq_0_bits_cf_waitForRobIdx_value),
    .io_deq_0_bits_cf_loadWaitBit(intDq_io_deq_0_bits_cf_loadWaitBit),
    .io_deq_0_bits_cf_loadWaitStrict(intDq_io_deq_0_bits_cf_loadWaitStrict),
    .io_deq_0_bits_cf_ssid(intDq_io_deq_0_bits_cf_ssid),
    .io_deq_0_bits_cf_ftqPtr_flag(intDq_io_deq_0_bits_cf_ftqPtr_flag),
    .io_deq_0_bits_cf_ftqPtr_value(intDq_io_deq_0_bits_cf_ftqPtr_value),
    .io_deq_0_bits_cf_ftqOffset(intDq_io_deq_0_bits_cf_ftqOffset),
    .io_deq_0_bits_ctrl_srcType_0(intDq_io_deq_0_bits_ctrl_srcType_0),
    .io_deq_0_bits_ctrl_srcType_1(intDq_io_deq_0_bits_ctrl_srcType_1),
    .io_deq_0_bits_ctrl_srcType_2(intDq_io_deq_0_bits_ctrl_srcType_2),
    .io_deq_0_bits_ctrl_fuType(intDq_io_deq_0_bits_ctrl_fuType),
    .io_deq_0_bits_ctrl_fuOpType(intDq_io_deq_0_bits_ctrl_fuOpType),
    .io_deq_0_bits_ctrl_rfWen(intDq_io_deq_0_bits_ctrl_rfWen),
    .io_deq_0_bits_ctrl_fpWen(intDq_io_deq_0_bits_ctrl_fpWen),
    .io_deq_0_bits_ctrl_flushPipe(intDq_io_deq_0_bits_ctrl_flushPipe),
    .io_deq_0_bits_ctrl_selImm(intDq_io_deq_0_bits_ctrl_selImm),
    .io_deq_0_bits_ctrl_imm(intDq_io_deq_0_bits_ctrl_imm),
    .io_deq_0_bits_ctrl_fpu_isAddSub(intDq_io_deq_0_bits_ctrl_fpu_isAddSub),
    .io_deq_0_bits_ctrl_fpu_typeTagIn(intDq_io_deq_0_bits_ctrl_fpu_typeTagIn),
    .io_deq_0_bits_ctrl_fpu_typeTagOut(intDq_io_deq_0_bits_ctrl_fpu_typeTagOut),
    .io_deq_0_bits_ctrl_fpu_fromInt(intDq_io_deq_0_bits_ctrl_fpu_fromInt),
    .io_deq_0_bits_ctrl_fpu_wflags(intDq_io_deq_0_bits_ctrl_fpu_wflags),
    .io_deq_0_bits_ctrl_fpu_fpWen(intDq_io_deq_0_bits_ctrl_fpu_fpWen),
    .io_deq_0_bits_ctrl_fpu_fmaCmd(intDq_io_deq_0_bits_ctrl_fpu_fmaCmd),
    .io_deq_0_bits_ctrl_fpu_div(intDq_io_deq_0_bits_ctrl_fpu_div),
    .io_deq_0_bits_ctrl_fpu_sqrt(intDq_io_deq_0_bits_ctrl_fpu_sqrt),
    .io_deq_0_bits_ctrl_fpu_fcvt(intDq_io_deq_0_bits_ctrl_fpu_fcvt),
    .io_deq_0_bits_ctrl_fpu_typ(intDq_io_deq_0_bits_ctrl_fpu_typ),
    .io_deq_0_bits_ctrl_fpu_fmt(intDq_io_deq_0_bits_ctrl_fpu_fmt),
    .io_deq_0_bits_ctrl_fpu_ren3(intDq_io_deq_0_bits_ctrl_fpu_ren3),
    .io_deq_0_bits_ctrl_fpu_rm(intDq_io_deq_0_bits_ctrl_fpu_rm),
    .io_deq_0_bits_ctrl_replayInst(intDq_io_deq_0_bits_ctrl_replayInst),
    .io_deq_0_bits_psrc_0(intDq_io_deq_0_bits_psrc_0),
    .io_deq_0_bits_psrc_1(intDq_io_deq_0_bits_psrc_1),
    .io_deq_0_bits_psrc_2(intDq_io_deq_0_bits_psrc_2),
    .io_deq_0_bits_pdest(intDq_io_deq_0_bits_pdest),
    .io_deq_0_bits_robIdx_flag(intDq_io_deq_0_bits_robIdx_flag),
    .io_deq_0_bits_robIdx_value(intDq_io_deq_0_bits_robIdx_value),
    .io_deq_0_bits_lqIdx_flag(intDq_io_deq_0_bits_lqIdx_flag),
    .io_deq_0_bits_lqIdx_value(intDq_io_deq_0_bits_lqIdx_value),
    .io_deq_0_bits_sqIdx_flag(intDq_io_deq_0_bits_sqIdx_flag),
    .io_deq_0_bits_sqIdx_value(intDq_io_deq_0_bits_sqIdx_value),
    .io_deq_1_ready(intDq_io_deq_1_ready),
    .io_deq_1_valid(intDq_io_deq_1_valid),
    .io_deq_1_bits_cf_foldpc(intDq_io_deq_1_bits_cf_foldpc),
    .io_deq_1_bits_cf_trigger_backendEn_0(intDq_io_deq_1_bits_cf_trigger_backendEn_0),
    .io_deq_1_bits_cf_trigger_backendEn_1(intDq_io_deq_1_bits_cf_trigger_backendEn_1),
    .io_deq_1_bits_cf_pd_isRVC(intDq_io_deq_1_bits_cf_pd_isRVC),
    .io_deq_1_bits_cf_pd_brType(intDq_io_deq_1_bits_cf_pd_brType),
    .io_deq_1_bits_cf_pd_isCall(intDq_io_deq_1_bits_cf_pd_isCall),
    .io_deq_1_bits_cf_pd_isRet(intDq_io_deq_1_bits_cf_pd_isRet),
    .io_deq_1_bits_cf_pred_taken(intDq_io_deq_1_bits_cf_pred_taken),
    .io_deq_1_bits_cf_storeSetHit(intDq_io_deq_1_bits_cf_storeSetHit),
    .io_deq_1_bits_cf_waitForRobIdx_flag(intDq_io_deq_1_bits_cf_waitForRobIdx_flag),
    .io_deq_1_bits_cf_waitForRobIdx_value(intDq_io_deq_1_bits_cf_waitForRobIdx_value),
    .io_deq_1_bits_cf_loadWaitBit(intDq_io_deq_1_bits_cf_loadWaitBit),
    .io_deq_1_bits_cf_loadWaitStrict(intDq_io_deq_1_bits_cf_loadWaitStrict),
    .io_deq_1_bits_cf_ssid(intDq_io_deq_1_bits_cf_ssid),
    .io_deq_1_bits_cf_ftqPtr_flag(intDq_io_deq_1_bits_cf_ftqPtr_flag),
    .io_deq_1_bits_cf_ftqPtr_value(intDq_io_deq_1_bits_cf_ftqPtr_value),
    .io_deq_1_bits_cf_ftqOffset(intDq_io_deq_1_bits_cf_ftqOffset),
    .io_deq_1_bits_ctrl_srcType_0(intDq_io_deq_1_bits_ctrl_srcType_0),
    .io_deq_1_bits_ctrl_srcType_1(intDq_io_deq_1_bits_ctrl_srcType_1),
    .io_deq_1_bits_ctrl_fuType(intDq_io_deq_1_bits_ctrl_fuType),
    .io_deq_1_bits_ctrl_fuOpType(intDq_io_deq_1_bits_ctrl_fuOpType),
    .io_deq_1_bits_ctrl_rfWen(intDq_io_deq_1_bits_ctrl_rfWen),
    .io_deq_1_bits_ctrl_fpWen(intDq_io_deq_1_bits_ctrl_fpWen),
    .io_deq_1_bits_ctrl_flushPipe(intDq_io_deq_1_bits_ctrl_flushPipe),
    .io_deq_1_bits_ctrl_selImm(intDq_io_deq_1_bits_ctrl_selImm),
    .io_deq_1_bits_ctrl_imm(intDq_io_deq_1_bits_ctrl_imm),
    .io_deq_1_bits_ctrl_replayInst(intDq_io_deq_1_bits_ctrl_replayInst),
    .io_deq_1_bits_psrc_0(intDq_io_deq_1_bits_psrc_0),
    .io_deq_1_bits_psrc_1(intDq_io_deq_1_bits_psrc_1),
    .io_deq_1_bits_pdest(intDq_io_deq_1_bits_pdest),
    .io_deq_1_bits_robIdx_flag(intDq_io_deq_1_bits_robIdx_flag),
    .io_deq_1_bits_robIdx_value(intDq_io_deq_1_bits_robIdx_value),
    .io_deq_1_bits_lqIdx_flag(intDq_io_deq_1_bits_lqIdx_flag),
    .io_deq_1_bits_lqIdx_value(intDq_io_deq_1_bits_lqIdx_value),
    .io_deq_1_bits_sqIdx_flag(intDq_io_deq_1_bits_sqIdx_flag),
    .io_deq_1_bits_sqIdx_value(intDq_io_deq_1_bits_sqIdx_value),
    .io_deq_2_ready(intDq_io_deq_2_ready),
    .io_deq_2_valid(intDq_io_deq_2_valid),
    .io_deq_2_bits_cf_foldpc(intDq_io_deq_2_bits_cf_foldpc),
    .io_deq_2_bits_cf_trigger_backendEn_0(intDq_io_deq_2_bits_cf_trigger_backendEn_0),
    .io_deq_2_bits_cf_trigger_backendEn_1(intDq_io_deq_2_bits_cf_trigger_backendEn_1),
    .io_deq_2_bits_cf_pd_isRVC(intDq_io_deq_2_bits_cf_pd_isRVC),
    .io_deq_2_bits_cf_pd_brType(intDq_io_deq_2_bits_cf_pd_brType),
    .io_deq_2_bits_cf_pd_isCall(intDq_io_deq_2_bits_cf_pd_isCall),
    .io_deq_2_bits_cf_pd_isRet(intDq_io_deq_2_bits_cf_pd_isRet),
    .io_deq_2_bits_cf_pred_taken(intDq_io_deq_2_bits_cf_pred_taken),
    .io_deq_2_bits_cf_storeSetHit(intDq_io_deq_2_bits_cf_storeSetHit),
    .io_deq_2_bits_cf_waitForRobIdx_flag(intDq_io_deq_2_bits_cf_waitForRobIdx_flag),
    .io_deq_2_bits_cf_waitForRobIdx_value(intDq_io_deq_2_bits_cf_waitForRobIdx_value),
    .io_deq_2_bits_cf_loadWaitBit(intDq_io_deq_2_bits_cf_loadWaitBit),
    .io_deq_2_bits_cf_loadWaitStrict(intDq_io_deq_2_bits_cf_loadWaitStrict),
    .io_deq_2_bits_cf_ssid(intDq_io_deq_2_bits_cf_ssid),
    .io_deq_2_bits_cf_ftqPtr_flag(intDq_io_deq_2_bits_cf_ftqPtr_flag),
    .io_deq_2_bits_cf_ftqPtr_value(intDq_io_deq_2_bits_cf_ftqPtr_value),
    .io_deq_2_bits_cf_ftqOffset(intDq_io_deq_2_bits_cf_ftqOffset),
    .io_deq_2_bits_ctrl_srcType_0(intDq_io_deq_2_bits_ctrl_srcType_0),
    .io_deq_2_bits_ctrl_srcType_1(intDq_io_deq_2_bits_ctrl_srcType_1),
    .io_deq_2_bits_ctrl_fuType(intDq_io_deq_2_bits_ctrl_fuType),
    .io_deq_2_bits_ctrl_fuOpType(intDq_io_deq_2_bits_ctrl_fuOpType),
    .io_deq_2_bits_ctrl_rfWen(intDq_io_deq_2_bits_ctrl_rfWen),
    .io_deq_2_bits_ctrl_fpWen(intDq_io_deq_2_bits_ctrl_fpWen),
    .io_deq_2_bits_ctrl_flushPipe(intDq_io_deq_2_bits_ctrl_flushPipe),
    .io_deq_2_bits_ctrl_imm(intDq_io_deq_2_bits_ctrl_imm),
    .io_deq_2_bits_ctrl_replayInst(intDq_io_deq_2_bits_ctrl_replayInst),
    .io_deq_2_bits_psrc_0(intDq_io_deq_2_bits_psrc_0),
    .io_deq_2_bits_psrc_1(intDq_io_deq_2_bits_psrc_1),
    .io_deq_2_bits_pdest(intDq_io_deq_2_bits_pdest),
    .io_deq_2_bits_robIdx_flag(intDq_io_deq_2_bits_robIdx_flag),
    .io_deq_2_bits_robIdx_value(intDq_io_deq_2_bits_robIdx_value),
    .io_deq_3_ready(intDq_io_deq_3_ready),
    .io_deq_3_valid(intDq_io_deq_3_valid),
    .io_deq_3_bits_cf_foldpc(intDq_io_deq_3_bits_cf_foldpc),
    .io_deq_3_bits_cf_trigger_backendEn_0(intDq_io_deq_3_bits_cf_trigger_backendEn_0),
    .io_deq_3_bits_cf_trigger_backendEn_1(intDq_io_deq_3_bits_cf_trigger_backendEn_1),
    .io_deq_3_bits_cf_pd_isRVC(intDq_io_deq_3_bits_cf_pd_isRVC),
    .io_deq_3_bits_cf_pd_brType(intDq_io_deq_3_bits_cf_pd_brType),
    .io_deq_3_bits_cf_pd_isCall(intDq_io_deq_3_bits_cf_pd_isCall),
    .io_deq_3_bits_cf_pd_isRet(intDq_io_deq_3_bits_cf_pd_isRet),
    .io_deq_3_bits_cf_pred_taken(intDq_io_deq_3_bits_cf_pred_taken),
    .io_deq_3_bits_cf_storeSetHit(intDq_io_deq_3_bits_cf_storeSetHit),
    .io_deq_3_bits_cf_waitForRobIdx_flag(intDq_io_deq_3_bits_cf_waitForRobIdx_flag),
    .io_deq_3_bits_cf_waitForRobIdx_value(intDq_io_deq_3_bits_cf_waitForRobIdx_value),
    .io_deq_3_bits_cf_loadWaitBit(intDq_io_deq_3_bits_cf_loadWaitBit),
    .io_deq_3_bits_cf_loadWaitStrict(intDq_io_deq_3_bits_cf_loadWaitStrict),
    .io_deq_3_bits_cf_ssid(intDq_io_deq_3_bits_cf_ssid),
    .io_deq_3_bits_cf_ftqPtr_flag(intDq_io_deq_3_bits_cf_ftqPtr_flag),
    .io_deq_3_bits_cf_ftqPtr_value(intDq_io_deq_3_bits_cf_ftqPtr_value),
    .io_deq_3_bits_cf_ftqOffset(intDq_io_deq_3_bits_cf_ftqOffset),
    .io_deq_3_bits_ctrl_srcType_0(intDq_io_deq_3_bits_ctrl_srcType_0),
    .io_deq_3_bits_ctrl_srcType_1(intDq_io_deq_3_bits_ctrl_srcType_1),
    .io_deq_3_bits_ctrl_fuType(intDq_io_deq_3_bits_ctrl_fuType),
    .io_deq_3_bits_ctrl_fuOpType(intDq_io_deq_3_bits_ctrl_fuOpType),
    .io_deq_3_bits_ctrl_rfWen(intDq_io_deq_3_bits_ctrl_rfWen),
    .io_deq_3_bits_ctrl_fpWen(intDq_io_deq_3_bits_ctrl_fpWen),
    .io_deq_3_bits_ctrl_flushPipe(intDq_io_deq_3_bits_ctrl_flushPipe),
    .io_deq_3_bits_ctrl_imm(intDq_io_deq_3_bits_ctrl_imm),
    .io_deq_3_bits_ctrl_replayInst(intDq_io_deq_3_bits_ctrl_replayInst),
    .io_deq_3_bits_psrc_0(intDq_io_deq_3_bits_psrc_0),
    .io_deq_3_bits_psrc_1(intDq_io_deq_3_bits_psrc_1),
    .io_deq_3_bits_pdest(intDq_io_deq_3_bits_pdest),
    .io_deq_3_bits_robIdx_flag(intDq_io_deq_3_bits_robIdx_flag),
    .io_deq_3_bits_robIdx_value(intDq_io_deq_3_bits_robIdx_value),
    .io_redirect_valid(intDq_io_redirect_valid),
    .io_redirect_bits_robIdx_flag(intDq_io_redirect_bits_robIdx_flag),
    .io_redirect_bits_robIdx_value(intDq_io_redirect_bits_robIdx_value),
    .io_redirect_bits_level(intDq_io_redirect_bits_level),
    .io_deqNext_0_cf_ftqPtr_value(intDq_io_deqNext_0_cf_ftqPtr_value),
    .io_deqNext_0_cf_ftqOffset(intDq_io_deqNext_0_cf_ftqOffset),
    .io_deqNext_0_ctrl_srcType_0(intDq_io_deqNext_0_ctrl_srcType_0),
    .io_deqNext_0_ctrl_srcType_1(intDq_io_deqNext_0_ctrl_srcType_1),
    .io_deqNext_0_ctrl_srcType_2(intDq_io_deqNext_0_ctrl_srcType_2),
    .io_deqNext_0_ctrl_fuType(intDq_io_deqNext_0_ctrl_fuType),
    .io_deqNext_0_ctrl_fuOpType(intDq_io_deqNext_0_ctrl_fuOpType),
    .io_deqNext_0_ctrl_rfWen(intDq_io_deqNext_0_ctrl_rfWen),
    .io_deqNext_0_ctrl_fpWen(intDq_io_deqNext_0_ctrl_fpWen),
    .io_deqNext_0_ctrl_flushPipe(intDq_io_deqNext_0_ctrl_flushPipe),
    .io_deqNext_0_ctrl_selImm(intDq_io_deqNext_0_ctrl_selImm),
    .io_deqNext_0_ctrl_imm(intDq_io_deqNext_0_ctrl_imm),
    .io_deqNext_0_ctrl_replayInst(intDq_io_deqNext_0_ctrl_replayInst),
    .io_deqNext_0_psrc_0(intDq_io_deqNext_0_psrc_0),
    .io_deqNext_0_psrc_1(intDq_io_deqNext_0_psrc_1),
    .io_deqNext_0_psrc_2(intDq_io_deqNext_0_psrc_2),
    .io_deqNext_0_pdest(intDq_io_deqNext_0_pdest),
    .io_deqNext_0_robIdx_flag(intDq_io_deqNext_0_robIdx_flag),
    .io_deqNext_0_robIdx_value(intDq_io_deqNext_0_robIdx_value),
    .io_deqNext_0_lqIdx_flag(intDq_io_deqNext_0_lqIdx_flag),
    .io_deqNext_0_lqIdx_value(intDq_io_deqNext_0_lqIdx_value),
    .io_deqNext_0_sqIdx_flag(intDq_io_deqNext_0_sqIdx_flag),
    .io_deqNext_0_sqIdx_value(intDq_io_deqNext_0_sqIdx_value),
    .io_deqNext_1_cf_ftqPtr_value(intDq_io_deqNext_1_cf_ftqPtr_value),
    .io_deqNext_1_cf_ftqOffset(intDq_io_deqNext_1_cf_ftqOffset),
    .io_deqNext_1_ctrl_srcType_0(intDq_io_deqNext_1_ctrl_srcType_0),
    .io_deqNext_1_ctrl_srcType_1(intDq_io_deqNext_1_ctrl_srcType_1),
    .io_deqNext_1_ctrl_srcType_2(intDq_io_deqNext_1_ctrl_srcType_2),
    .io_deqNext_1_ctrl_fuType(intDq_io_deqNext_1_ctrl_fuType),
    .io_deqNext_1_ctrl_fuOpType(intDq_io_deqNext_1_ctrl_fuOpType),
    .io_deqNext_1_ctrl_rfWen(intDq_io_deqNext_1_ctrl_rfWen),
    .io_deqNext_1_ctrl_fpWen(intDq_io_deqNext_1_ctrl_fpWen),
    .io_deqNext_1_ctrl_flushPipe(intDq_io_deqNext_1_ctrl_flushPipe),
    .io_deqNext_1_ctrl_selImm(intDq_io_deqNext_1_ctrl_selImm),
    .io_deqNext_1_ctrl_imm(intDq_io_deqNext_1_ctrl_imm),
    .io_deqNext_1_ctrl_replayInst(intDq_io_deqNext_1_ctrl_replayInst),
    .io_deqNext_1_psrc_0(intDq_io_deqNext_1_psrc_0),
    .io_deqNext_1_psrc_1(intDq_io_deqNext_1_psrc_1),
    .io_deqNext_1_psrc_2(intDq_io_deqNext_1_psrc_2),
    .io_deqNext_1_pdest(intDq_io_deqNext_1_pdest),
    .io_deqNext_1_robIdx_flag(intDq_io_deqNext_1_robIdx_flag),
    .io_deqNext_1_robIdx_value(intDq_io_deqNext_1_robIdx_value),
    .io_deqNext_1_lqIdx_flag(intDq_io_deqNext_1_lqIdx_flag),
    .io_deqNext_1_lqIdx_value(intDq_io_deqNext_1_lqIdx_value),
    .io_deqNext_1_sqIdx_flag(intDq_io_deqNext_1_sqIdx_flag),
    .io_deqNext_1_sqIdx_value(intDq_io_deqNext_1_sqIdx_value),
    .io_deqNext_2_cf_ftqPtr_value(intDq_io_deqNext_2_cf_ftqPtr_value),
    .io_deqNext_2_cf_ftqOffset(intDq_io_deqNext_2_cf_ftqOffset),
    .io_deqNext_2_ctrl_srcType_0(intDq_io_deqNext_2_ctrl_srcType_0),
    .io_deqNext_2_ctrl_srcType_1(intDq_io_deqNext_2_ctrl_srcType_1),
    .io_deqNext_2_ctrl_srcType_2(intDq_io_deqNext_2_ctrl_srcType_2),
    .io_deqNext_2_ctrl_fuType(intDq_io_deqNext_2_ctrl_fuType),
    .io_deqNext_2_ctrl_fuOpType(intDq_io_deqNext_2_ctrl_fuOpType),
    .io_deqNext_2_ctrl_rfWen(intDq_io_deqNext_2_ctrl_rfWen),
    .io_deqNext_2_ctrl_fpWen(intDq_io_deqNext_2_ctrl_fpWen),
    .io_deqNext_2_ctrl_flushPipe(intDq_io_deqNext_2_ctrl_flushPipe),
    .io_deqNext_2_ctrl_selImm(intDq_io_deqNext_2_ctrl_selImm),
    .io_deqNext_2_ctrl_imm(intDq_io_deqNext_2_ctrl_imm),
    .io_deqNext_2_ctrl_replayInst(intDq_io_deqNext_2_ctrl_replayInst),
    .io_deqNext_2_psrc_0(intDq_io_deqNext_2_psrc_0),
    .io_deqNext_2_psrc_1(intDq_io_deqNext_2_psrc_1),
    .io_deqNext_2_psrc_2(intDq_io_deqNext_2_psrc_2),
    .io_deqNext_2_pdest(intDq_io_deqNext_2_pdest),
    .io_deqNext_2_robIdx_flag(intDq_io_deqNext_2_robIdx_flag),
    .io_deqNext_2_robIdx_value(intDq_io_deqNext_2_robIdx_value),
    .io_deqNext_2_lqIdx_flag(intDq_io_deqNext_2_lqIdx_flag),
    .io_deqNext_2_lqIdx_value(intDq_io_deqNext_2_lqIdx_value),
    .io_deqNext_2_sqIdx_flag(intDq_io_deqNext_2_sqIdx_flag),
    .io_deqNext_2_sqIdx_value(intDq_io_deqNext_2_sqIdx_value),
    .io_deqNext_3_cf_ftqPtr_value(intDq_io_deqNext_3_cf_ftqPtr_value),
    .io_deqNext_3_cf_ftqOffset(intDq_io_deqNext_3_cf_ftqOffset),
    .io_deqNext_3_ctrl_srcType_0(intDq_io_deqNext_3_ctrl_srcType_0),
    .io_deqNext_3_ctrl_srcType_1(intDq_io_deqNext_3_ctrl_srcType_1),
    .io_deqNext_3_ctrl_srcType_2(intDq_io_deqNext_3_ctrl_srcType_2),
    .io_deqNext_3_ctrl_fuType(intDq_io_deqNext_3_ctrl_fuType),
    .io_deqNext_3_ctrl_fuOpType(intDq_io_deqNext_3_ctrl_fuOpType),
    .io_deqNext_3_ctrl_rfWen(intDq_io_deqNext_3_ctrl_rfWen),
    .io_deqNext_3_ctrl_fpWen(intDq_io_deqNext_3_ctrl_fpWen),
    .io_deqNext_3_ctrl_flushPipe(intDq_io_deqNext_3_ctrl_flushPipe),
    .io_deqNext_3_ctrl_selImm(intDq_io_deqNext_3_ctrl_selImm),
    .io_deqNext_3_ctrl_imm(intDq_io_deqNext_3_ctrl_imm),
    .io_deqNext_3_ctrl_replayInst(intDq_io_deqNext_3_ctrl_replayInst),
    .io_deqNext_3_psrc_0(intDq_io_deqNext_3_psrc_0),
    .io_deqNext_3_psrc_1(intDq_io_deqNext_3_psrc_1),
    .io_deqNext_3_psrc_2(intDq_io_deqNext_3_psrc_2),
    .io_deqNext_3_pdest(intDq_io_deqNext_3_pdest),
    .io_deqNext_3_robIdx_flag(intDq_io_deqNext_3_robIdx_flag),
    .io_deqNext_3_robIdx_value(intDq_io_deqNext_3_robIdx_value),
    .io_deqNext_3_lqIdx_flag(intDq_io_deqNext_3_lqIdx_flag),
    .io_deqNext_3_lqIdx_value(intDq_io_deqNext_3_lqIdx_value),
    .io_deqNext_3_sqIdx_flag(intDq_io_deqNext_3_sqIdx_flag),
    .io_deqNext_3_sqIdx_value(intDq_io_deqNext_3_sqIdx_value),
    .io_perf_0_value(intDq_io_perf_0_value),
    .io_perf_1_value(intDq_io_perf_1_value),
    .io_perf_2_value(intDq_io_perf_2_value),
    .io_perf_3_value(intDq_io_perf_3_value),
    .io_perf_4_value(intDq_io_perf_4_value),
    .io_perf_5_value(intDq_io_perf_5_value),
    .io_perf_6_value(intDq_io_perf_6_value),
    .io_perf_7_value(intDq_io_perf_7_value)
  );
  DispatchQueue fpDq ( // @[CtrlBlock.scala 271:20]
    .clock(fpDq_clock),
    .reset(fpDq_reset),
    .io_enq_canAccept(fpDq_io_enq_canAccept),
    .io_enq_needAlloc_0(fpDq_io_enq_needAlloc_0),
    .io_enq_needAlloc_1(fpDq_io_enq_needAlloc_1),
    .io_enq_req_0_valid(fpDq_io_enq_req_0_valid),
    .io_enq_req_0_bits_cf_foldpc(fpDq_io_enq_req_0_bits_cf_foldpc),
    .io_enq_req_0_bits_cf_trigger_backendEn_0(fpDq_io_enq_req_0_bits_cf_trigger_backendEn_0),
    .io_enq_req_0_bits_cf_trigger_backendEn_1(fpDq_io_enq_req_0_bits_cf_trigger_backendEn_1),
    .io_enq_req_0_bits_cf_pd_isRVC(fpDq_io_enq_req_0_bits_cf_pd_isRVC),
    .io_enq_req_0_bits_cf_pd_brType(fpDq_io_enq_req_0_bits_cf_pd_brType),
    .io_enq_req_0_bits_cf_pd_isCall(fpDq_io_enq_req_0_bits_cf_pd_isCall),
    .io_enq_req_0_bits_cf_pd_isRet(fpDq_io_enq_req_0_bits_cf_pd_isRet),
    .io_enq_req_0_bits_cf_pred_taken(fpDq_io_enq_req_0_bits_cf_pred_taken),
    .io_enq_req_0_bits_cf_storeSetHit(fpDq_io_enq_req_0_bits_cf_storeSetHit),
    .io_enq_req_0_bits_cf_waitForRobIdx_flag(fpDq_io_enq_req_0_bits_cf_waitForRobIdx_flag),
    .io_enq_req_0_bits_cf_waitForRobIdx_value(fpDq_io_enq_req_0_bits_cf_waitForRobIdx_value),
    .io_enq_req_0_bits_cf_loadWaitBit(fpDq_io_enq_req_0_bits_cf_loadWaitBit),
    .io_enq_req_0_bits_cf_loadWaitStrict(fpDq_io_enq_req_0_bits_cf_loadWaitStrict),
    .io_enq_req_0_bits_cf_ssid(fpDq_io_enq_req_0_bits_cf_ssid),
    .io_enq_req_0_bits_cf_ftqPtr_flag(fpDq_io_enq_req_0_bits_cf_ftqPtr_flag),
    .io_enq_req_0_bits_cf_ftqPtr_value(fpDq_io_enq_req_0_bits_cf_ftqPtr_value),
    .io_enq_req_0_bits_cf_ftqOffset(fpDq_io_enq_req_0_bits_cf_ftqOffset),
    .io_enq_req_0_bits_ctrl_srcType_0(fpDq_io_enq_req_0_bits_ctrl_srcType_0),
    .io_enq_req_0_bits_ctrl_srcType_1(fpDq_io_enq_req_0_bits_ctrl_srcType_1),
    .io_enq_req_0_bits_ctrl_srcType_2(fpDq_io_enq_req_0_bits_ctrl_srcType_2),
    .io_enq_req_0_bits_ctrl_fuType(fpDq_io_enq_req_0_bits_ctrl_fuType),
    .io_enq_req_0_bits_ctrl_fuOpType(fpDq_io_enq_req_0_bits_ctrl_fuOpType),
    .io_enq_req_0_bits_ctrl_rfWen(fpDq_io_enq_req_0_bits_ctrl_rfWen),
    .io_enq_req_0_bits_ctrl_fpWen(fpDq_io_enq_req_0_bits_ctrl_fpWen),
    .io_enq_req_0_bits_ctrl_flushPipe(fpDq_io_enq_req_0_bits_ctrl_flushPipe),
    .io_enq_req_0_bits_ctrl_selImm(fpDq_io_enq_req_0_bits_ctrl_selImm),
    .io_enq_req_0_bits_ctrl_imm(fpDq_io_enq_req_0_bits_ctrl_imm),
    .io_enq_req_0_bits_ctrl_fpu_isAddSub(fpDq_io_enq_req_0_bits_ctrl_fpu_isAddSub),
    .io_enq_req_0_bits_ctrl_fpu_typeTagIn(fpDq_io_enq_req_0_bits_ctrl_fpu_typeTagIn),
    .io_enq_req_0_bits_ctrl_fpu_typeTagOut(fpDq_io_enq_req_0_bits_ctrl_fpu_typeTagOut),
    .io_enq_req_0_bits_ctrl_fpu_fromInt(fpDq_io_enq_req_0_bits_ctrl_fpu_fromInt),
    .io_enq_req_0_bits_ctrl_fpu_wflags(fpDq_io_enq_req_0_bits_ctrl_fpu_wflags),
    .io_enq_req_0_bits_ctrl_fpu_fpWen(fpDq_io_enq_req_0_bits_ctrl_fpu_fpWen),
    .io_enq_req_0_bits_ctrl_fpu_fmaCmd(fpDq_io_enq_req_0_bits_ctrl_fpu_fmaCmd),
    .io_enq_req_0_bits_ctrl_fpu_div(fpDq_io_enq_req_0_bits_ctrl_fpu_div),
    .io_enq_req_0_bits_ctrl_fpu_sqrt(fpDq_io_enq_req_0_bits_ctrl_fpu_sqrt),
    .io_enq_req_0_bits_ctrl_fpu_fcvt(fpDq_io_enq_req_0_bits_ctrl_fpu_fcvt),
    .io_enq_req_0_bits_ctrl_fpu_typ(fpDq_io_enq_req_0_bits_ctrl_fpu_typ),
    .io_enq_req_0_bits_ctrl_fpu_fmt(fpDq_io_enq_req_0_bits_ctrl_fpu_fmt),
    .io_enq_req_0_bits_ctrl_fpu_ren3(fpDq_io_enq_req_0_bits_ctrl_fpu_ren3),
    .io_enq_req_0_bits_ctrl_fpu_rm(fpDq_io_enq_req_0_bits_ctrl_fpu_rm),
    .io_enq_req_0_bits_psrc_0(fpDq_io_enq_req_0_bits_psrc_0),
    .io_enq_req_0_bits_psrc_1(fpDq_io_enq_req_0_bits_psrc_1),
    .io_enq_req_0_bits_psrc_2(fpDq_io_enq_req_0_bits_psrc_2),
    .io_enq_req_0_bits_pdest(fpDq_io_enq_req_0_bits_pdest),
    .io_enq_req_0_bits_robIdx_flag(fpDq_io_enq_req_0_bits_robIdx_flag),
    .io_enq_req_0_bits_robIdx_value(fpDq_io_enq_req_0_bits_robIdx_value),
    .io_enq_req_1_valid(fpDq_io_enq_req_1_valid),
    .io_enq_req_1_bits_cf_foldpc(fpDq_io_enq_req_1_bits_cf_foldpc),
    .io_enq_req_1_bits_cf_trigger_backendEn_0(fpDq_io_enq_req_1_bits_cf_trigger_backendEn_0),
    .io_enq_req_1_bits_cf_trigger_backendEn_1(fpDq_io_enq_req_1_bits_cf_trigger_backendEn_1),
    .io_enq_req_1_bits_cf_pd_isRVC(fpDq_io_enq_req_1_bits_cf_pd_isRVC),
    .io_enq_req_1_bits_cf_pd_brType(fpDq_io_enq_req_1_bits_cf_pd_brType),
    .io_enq_req_1_bits_cf_pd_isCall(fpDq_io_enq_req_1_bits_cf_pd_isCall),
    .io_enq_req_1_bits_cf_pd_isRet(fpDq_io_enq_req_1_bits_cf_pd_isRet),
    .io_enq_req_1_bits_cf_pred_taken(fpDq_io_enq_req_1_bits_cf_pred_taken),
    .io_enq_req_1_bits_cf_storeSetHit(fpDq_io_enq_req_1_bits_cf_storeSetHit),
    .io_enq_req_1_bits_cf_waitForRobIdx_flag(fpDq_io_enq_req_1_bits_cf_waitForRobIdx_flag),
    .io_enq_req_1_bits_cf_waitForRobIdx_value(fpDq_io_enq_req_1_bits_cf_waitForRobIdx_value),
    .io_enq_req_1_bits_cf_loadWaitBit(fpDq_io_enq_req_1_bits_cf_loadWaitBit),
    .io_enq_req_1_bits_cf_loadWaitStrict(fpDq_io_enq_req_1_bits_cf_loadWaitStrict),
    .io_enq_req_1_bits_cf_ssid(fpDq_io_enq_req_1_bits_cf_ssid),
    .io_enq_req_1_bits_cf_ftqPtr_flag(fpDq_io_enq_req_1_bits_cf_ftqPtr_flag),
    .io_enq_req_1_bits_cf_ftqPtr_value(fpDq_io_enq_req_1_bits_cf_ftqPtr_value),
    .io_enq_req_1_bits_cf_ftqOffset(fpDq_io_enq_req_1_bits_cf_ftqOffset),
    .io_enq_req_1_bits_ctrl_srcType_0(fpDq_io_enq_req_1_bits_ctrl_srcType_0),
    .io_enq_req_1_bits_ctrl_srcType_1(fpDq_io_enq_req_1_bits_ctrl_srcType_1),
    .io_enq_req_1_bits_ctrl_srcType_2(fpDq_io_enq_req_1_bits_ctrl_srcType_2),
    .io_enq_req_1_bits_ctrl_fuType(fpDq_io_enq_req_1_bits_ctrl_fuType),
    .io_enq_req_1_bits_ctrl_fuOpType(fpDq_io_enq_req_1_bits_ctrl_fuOpType),
    .io_enq_req_1_bits_ctrl_rfWen(fpDq_io_enq_req_1_bits_ctrl_rfWen),
    .io_enq_req_1_bits_ctrl_fpWen(fpDq_io_enq_req_1_bits_ctrl_fpWen),
    .io_enq_req_1_bits_ctrl_flushPipe(fpDq_io_enq_req_1_bits_ctrl_flushPipe),
    .io_enq_req_1_bits_ctrl_selImm(fpDq_io_enq_req_1_bits_ctrl_selImm),
    .io_enq_req_1_bits_ctrl_imm(fpDq_io_enq_req_1_bits_ctrl_imm),
    .io_enq_req_1_bits_ctrl_fpu_isAddSub(fpDq_io_enq_req_1_bits_ctrl_fpu_isAddSub),
    .io_enq_req_1_bits_ctrl_fpu_typeTagIn(fpDq_io_enq_req_1_bits_ctrl_fpu_typeTagIn),
    .io_enq_req_1_bits_ctrl_fpu_typeTagOut(fpDq_io_enq_req_1_bits_ctrl_fpu_typeTagOut),
    .io_enq_req_1_bits_ctrl_fpu_fromInt(fpDq_io_enq_req_1_bits_ctrl_fpu_fromInt),
    .io_enq_req_1_bits_ctrl_fpu_wflags(fpDq_io_enq_req_1_bits_ctrl_fpu_wflags),
    .io_enq_req_1_bits_ctrl_fpu_fpWen(fpDq_io_enq_req_1_bits_ctrl_fpu_fpWen),
    .io_enq_req_1_bits_ctrl_fpu_fmaCmd(fpDq_io_enq_req_1_bits_ctrl_fpu_fmaCmd),
    .io_enq_req_1_bits_ctrl_fpu_div(fpDq_io_enq_req_1_bits_ctrl_fpu_div),
    .io_enq_req_1_bits_ctrl_fpu_sqrt(fpDq_io_enq_req_1_bits_ctrl_fpu_sqrt),
    .io_enq_req_1_bits_ctrl_fpu_fcvt(fpDq_io_enq_req_1_bits_ctrl_fpu_fcvt),
    .io_enq_req_1_bits_ctrl_fpu_typ(fpDq_io_enq_req_1_bits_ctrl_fpu_typ),
    .io_enq_req_1_bits_ctrl_fpu_fmt(fpDq_io_enq_req_1_bits_ctrl_fpu_fmt),
    .io_enq_req_1_bits_ctrl_fpu_ren3(fpDq_io_enq_req_1_bits_ctrl_fpu_ren3),
    .io_enq_req_1_bits_ctrl_fpu_rm(fpDq_io_enq_req_1_bits_ctrl_fpu_rm),
    .io_enq_req_1_bits_psrc_0(fpDq_io_enq_req_1_bits_psrc_0),
    .io_enq_req_1_bits_psrc_1(fpDq_io_enq_req_1_bits_psrc_1),
    .io_enq_req_1_bits_psrc_2(fpDq_io_enq_req_1_bits_psrc_2),
    .io_enq_req_1_bits_pdest(fpDq_io_enq_req_1_bits_pdest),
    .io_enq_req_1_bits_robIdx_flag(fpDq_io_enq_req_1_bits_robIdx_flag),
    .io_enq_req_1_bits_robIdx_value(fpDq_io_enq_req_1_bits_robIdx_value),
    .io_deq_0_ready(fpDq_io_deq_0_ready),
    .io_deq_0_valid(fpDq_io_deq_0_valid),
    .io_deq_0_bits_cf_foldpc(fpDq_io_deq_0_bits_cf_foldpc),
    .io_deq_0_bits_cf_trigger_backendEn_0(fpDq_io_deq_0_bits_cf_trigger_backendEn_0),
    .io_deq_0_bits_cf_trigger_backendEn_1(fpDq_io_deq_0_bits_cf_trigger_backendEn_1),
    .io_deq_0_bits_cf_pd_isRVC(fpDq_io_deq_0_bits_cf_pd_isRVC),
    .io_deq_0_bits_cf_pd_brType(fpDq_io_deq_0_bits_cf_pd_brType),
    .io_deq_0_bits_cf_pd_isCall(fpDq_io_deq_0_bits_cf_pd_isCall),
    .io_deq_0_bits_cf_pd_isRet(fpDq_io_deq_0_bits_cf_pd_isRet),
    .io_deq_0_bits_cf_pred_taken(fpDq_io_deq_0_bits_cf_pred_taken),
    .io_deq_0_bits_cf_storeSetHit(fpDq_io_deq_0_bits_cf_storeSetHit),
    .io_deq_0_bits_cf_waitForRobIdx_flag(fpDq_io_deq_0_bits_cf_waitForRobIdx_flag),
    .io_deq_0_bits_cf_waitForRobIdx_value(fpDq_io_deq_0_bits_cf_waitForRobIdx_value),
    .io_deq_0_bits_cf_loadWaitBit(fpDq_io_deq_0_bits_cf_loadWaitBit),
    .io_deq_0_bits_cf_loadWaitStrict(fpDq_io_deq_0_bits_cf_loadWaitStrict),
    .io_deq_0_bits_cf_ssid(fpDq_io_deq_0_bits_cf_ssid),
    .io_deq_0_bits_cf_ftqPtr_flag(fpDq_io_deq_0_bits_cf_ftqPtr_flag),
    .io_deq_0_bits_cf_ftqPtr_value(fpDq_io_deq_0_bits_cf_ftqPtr_value),
    .io_deq_0_bits_cf_ftqOffset(fpDq_io_deq_0_bits_cf_ftqOffset),
    .io_deq_0_bits_ctrl_srcType_0(fpDq_io_deq_0_bits_ctrl_srcType_0),
    .io_deq_0_bits_ctrl_srcType_1(fpDq_io_deq_0_bits_ctrl_srcType_1),
    .io_deq_0_bits_ctrl_srcType_2(fpDq_io_deq_0_bits_ctrl_srcType_2),
    .io_deq_0_bits_ctrl_fuType(fpDq_io_deq_0_bits_ctrl_fuType),
    .io_deq_0_bits_ctrl_fuOpType(fpDq_io_deq_0_bits_ctrl_fuOpType),
    .io_deq_0_bits_ctrl_rfWen(fpDq_io_deq_0_bits_ctrl_rfWen),
    .io_deq_0_bits_ctrl_fpWen(fpDq_io_deq_0_bits_ctrl_fpWen),
    .io_deq_0_bits_ctrl_flushPipe(fpDq_io_deq_0_bits_ctrl_flushPipe),
    .io_deq_0_bits_ctrl_selImm(fpDq_io_deq_0_bits_ctrl_selImm),
    .io_deq_0_bits_ctrl_imm(fpDq_io_deq_0_bits_ctrl_imm),
    .io_deq_0_bits_ctrl_fpu_isAddSub(fpDq_io_deq_0_bits_ctrl_fpu_isAddSub),
    .io_deq_0_bits_ctrl_fpu_typeTagIn(fpDq_io_deq_0_bits_ctrl_fpu_typeTagIn),
    .io_deq_0_bits_ctrl_fpu_typeTagOut(fpDq_io_deq_0_bits_ctrl_fpu_typeTagOut),
    .io_deq_0_bits_ctrl_fpu_fromInt(fpDq_io_deq_0_bits_ctrl_fpu_fromInt),
    .io_deq_0_bits_ctrl_fpu_wflags(fpDq_io_deq_0_bits_ctrl_fpu_wflags),
    .io_deq_0_bits_ctrl_fpu_fpWen(fpDq_io_deq_0_bits_ctrl_fpu_fpWen),
    .io_deq_0_bits_ctrl_fpu_fmaCmd(fpDq_io_deq_0_bits_ctrl_fpu_fmaCmd),
    .io_deq_0_bits_ctrl_fpu_div(fpDq_io_deq_0_bits_ctrl_fpu_div),
    .io_deq_0_bits_ctrl_fpu_sqrt(fpDq_io_deq_0_bits_ctrl_fpu_sqrt),
    .io_deq_0_bits_ctrl_fpu_fcvt(fpDq_io_deq_0_bits_ctrl_fpu_fcvt),
    .io_deq_0_bits_ctrl_fpu_typ(fpDq_io_deq_0_bits_ctrl_fpu_typ),
    .io_deq_0_bits_ctrl_fpu_fmt(fpDq_io_deq_0_bits_ctrl_fpu_fmt),
    .io_deq_0_bits_ctrl_fpu_ren3(fpDq_io_deq_0_bits_ctrl_fpu_ren3),
    .io_deq_0_bits_ctrl_fpu_rm(fpDq_io_deq_0_bits_ctrl_fpu_rm),
    .io_deq_0_bits_ctrl_replayInst(fpDq_io_deq_0_bits_ctrl_replayInst),
    .io_deq_0_bits_psrc_0(fpDq_io_deq_0_bits_psrc_0),
    .io_deq_0_bits_psrc_1(fpDq_io_deq_0_bits_psrc_1),
    .io_deq_0_bits_psrc_2(fpDq_io_deq_0_bits_psrc_2),
    .io_deq_0_bits_pdest(fpDq_io_deq_0_bits_pdest),
    .io_deq_0_bits_robIdx_flag(fpDq_io_deq_0_bits_robIdx_flag),
    .io_deq_0_bits_robIdx_value(fpDq_io_deq_0_bits_robIdx_value),
    .io_deq_0_bits_lqIdx_flag(fpDq_io_deq_0_bits_lqIdx_flag),
    .io_deq_0_bits_lqIdx_value(fpDq_io_deq_0_bits_lqIdx_value),
    .io_deq_0_bits_sqIdx_flag(fpDq_io_deq_0_bits_sqIdx_flag),
    .io_deq_0_bits_sqIdx_value(fpDq_io_deq_0_bits_sqIdx_value),
    .io_deq_1_ready(fpDq_io_deq_1_ready),
    .io_deq_1_valid(fpDq_io_deq_1_valid),
    .io_deq_1_bits_cf_foldpc(fpDq_io_deq_1_bits_cf_foldpc),
    .io_deq_1_bits_cf_trigger_backendEn_0(fpDq_io_deq_1_bits_cf_trigger_backendEn_0),
    .io_deq_1_bits_cf_trigger_backendEn_1(fpDq_io_deq_1_bits_cf_trigger_backendEn_1),
    .io_deq_1_bits_cf_pd_isRVC(fpDq_io_deq_1_bits_cf_pd_isRVC),
    .io_deq_1_bits_cf_pd_brType(fpDq_io_deq_1_bits_cf_pd_brType),
    .io_deq_1_bits_cf_pd_isCall(fpDq_io_deq_1_bits_cf_pd_isCall),
    .io_deq_1_bits_cf_pd_isRet(fpDq_io_deq_1_bits_cf_pd_isRet),
    .io_deq_1_bits_cf_pred_taken(fpDq_io_deq_1_bits_cf_pred_taken),
    .io_deq_1_bits_cf_storeSetHit(fpDq_io_deq_1_bits_cf_storeSetHit),
    .io_deq_1_bits_cf_waitForRobIdx_flag(fpDq_io_deq_1_bits_cf_waitForRobIdx_flag),
    .io_deq_1_bits_cf_waitForRobIdx_value(fpDq_io_deq_1_bits_cf_waitForRobIdx_value),
    .io_deq_1_bits_cf_loadWaitBit(fpDq_io_deq_1_bits_cf_loadWaitBit),
    .io_deq_1_bits_cf_loadWaitStrict(fpDq_io_deq_1_bits_cf_loadWaitStrict),
    .io_deq_1_bits_cf_ssid(fpDq_io_deq_1_bits_cf_ssid),
    .io_deq_1_bits_cf_ftqPtr_flag(fpDq_io_deq_1_bits_cf_ftqPtr_flag),
    .io_deq_1_bits_cf_ftqPtr_value(fpDq_io_deq_1_bits_cf_ftqPtr_value),
    .io_deq_1_bits_cf_ftqOffset(fpDq_io_deq_1_bits_cf_ftqOffset),
    .io_deq_1_bits_ctrl_srcType_0(fpDq_io_deq_1_bits_ctrl_srcType_0),
    .io_deq_1_bits_ctrl_srcType_1(fpDq_io_deq_1_bits_ctrl_srcType_1),
    .io_deq_1_bits_ctrl_fuType(fpDq_io_deq_1_bits_ctrl_fuType),
    .io_deq_1_bits_ctrl_fuOpType(fpDq_io_deq_1_bits_ctrl_fuOpType),
    .io_deq_1_bits_ctrl_rfWen(fpDq_io_deq_1_bits_ctrl_rfWen),
    .io_deq_1_bits_ctrl_fpWen(fpDq_io_deq_1_bits_ctrl_fpWen),
    .io_deq_1_bits_ctrl_flushPipe(fpDq_io_deq_1_bits_ctrl_flushPipe),
    .io_deq_1_bits_ctrl_selImm(fpDq_io_deq_1_bits_ctrl_selImm),
    .io_deq_1_bits_ctrl_imm(fpDq_io_deq_1_bits_ctrl_imm),
    .io_deq_1_bits_ctrl_replayInst(fpDq_io_deq_1_bits_ctrl_replayInst),
    .io_deq_1_bits_psrc_0(fpDq_io_deq_1_bits_psrc_0),
    .io_deq_1_bits_psrc_1(fpDq_io_deq_1_bits_psrc_1),
    .io_deq_1_bits_pdest(fpDq_io_deq_1_bits_pdest),
    .io_deq_1_bits_robIdx_flag(fpDq_io_deq_1_bits_robIdx_flag),
    .io_deq_1_bits_robIdx_value(fpDq_io_deq_1_bits_robIdx_value),
    .io_deq_1_bits_lqIdx_flag(fpDq_io_deq_1_bits_lqIdx_flag),
    .io_deq_1_bits_lqIdx_value(fpDq_io_deq_1_bits_lqIdx_value),
    .io_deq_1_bits_sqIdx_flag(fpDq_io_deq_1_bits_sqIdx_flag),
    .io_deq_1_bits_sqIdx_value(fpDq_io_deq_1_bits_sqIdx_value),
    .io_deq_2_ready(fpDq_io_deq_2_ready),
    .io_deq_2_valid(fpDq_io_deq_2_valid),
    .io_deq_2_bits_cf_foldpc(fpDq_io_deq_2_bits_cf_foldpc),
    .io_deq_2_bits_cf_trigger_backendEn_0(fpDq_io_deq_2_bits_cf_trigger_backendEn_0),
    .io_deq_2_bits_cf_trigger_backendEn_1(fpDq_io_deq_2_bits_cf_trigger_backendEn_1),
    .io_deq_2_bits_cf_pd_isRVC(fpDq_io_deq_2_bits_cf_pd_isRVC),
    .io_deq_2_bits_cf_pd_brType(fpDq_io_deq_2_bits_cf_pd_brType),
    .io_deq_2_bits_cf_pd_isCall(fpDq_io_deq_2_bits_cf_pd_isCall),
    .io_deq_2_bits_cf_pd_isRet(fpDq_io_deq_2_bits_cf_pd_isRet),
    .io_deq_2_bits_cf_pred_taken(fpDq_io_deq_2_bits_cf_pred_taken),
    .io_deq_2_bits_cf_storeSetHit(fpDq_io_deq_2_bits_cf_storeSetHit),
    .io_deq_2_bits_cf_waitForRobIdx_flag(fpDq_io_deq_2_bits_cf_waitForRobIdx_flag),
    .io_deq_2_bits_cf_waitForRobIdx_value(fpDq_io_deq_2_bits_cf_waitForRobIdx_value),
    .io_deq_2_bits_cf_loadWaitBit(fpDq_io_deq_2_bits_cf_loadWaitBit),
    .io_deq_2_bits_cf_loadWaitStrict(fpDq_io_deq_2_bits_cf_loadWaitStrict),
    .io_deq_2_bits_cf_ssid(fpDq_io_deq_2_bits_cf_ssid),
    .io_deq_2_bits_cf_ftqPtr_flag(fpDq_io_deq_2_bits_cf_ftqPtr_flag),
    .io_deq_2_bits_cf_ftqPtr_value(fpDq_io_deq_2_bits_cf_ftqPtr_value),
    .io_deq_2_bits_cf_ftqOffset(fpDq_io_deq_2_bits_cf_ftqOffset),
    .io_deq_2_bits_ctrl_srcType_0(fpDq_io_deq_2_bits_ctrl_srcType_0),
    .io_deq_2_bits_ctrl_srcType_1(fpDq_io_deq_2_bits_ctrl_srcType_1),
    .io_deq_2_bits_ctrl_fuType(fpDq_io_deq_2_bits_ctrl_fuType),
    .io_deq_2_bits_ctrl_fuOpType(fpDq_io_deq_2_bits_ctrl_fuOpType),
    .io_deq_2_bits_ctrl_rfWen(fpDq_io_deq_2_bits_ctrl_rfWen),
    .io_deq_2_bits_ctrl_fpWen(fpDq_io_deq_2_bits_ctrl_fpWen),
    .io_deq_2_bits_ctrl_flushPipe(fpDq_io_deq_2_bits_ctrl_flushPipe),
    .io_deq_2_bits_ctrl_imm(fpDq_io_deq_2_bits_ctrl_imm),
    .io_deq_2_bits_ctrl_replayInst(fpDq_io_deq_2_bits_ctrl_replayInst),
    .io_deq_2_bits_psrc_0(fpDq_io_deq_2_bits_psrc_0),
    .io_deq_2_bits_psrc_1(fpDq_io_deq_2_bits_psrc_1),
    .io_deq_2_bits_pdest(fpDq_io_deq_2_bits_pdest),
    .io_deq_2_bits_robIdx_flag(fpDq_io_deq_2_bits_robIdx_flag),
    .io_deq_2_bits_robIdx_value(fpDq_io_deq_2_bits_robIdx_value),
    .io_deq_3_ready(fpDq_io_deq_3_ready),
    .io_deq_3_valid(fpDq_io_deq_3_valid),
    .io_deq_3_bits_cf_foldpc(fpDq_io_deq_3_bits_cf_foldpc),
    .io_deq_3_bits_cf_trigger_backendEn_0(fpDq_io_deq_3_bits_cf_trigger_backendEn_0),
    .io_deq_3_bits_cf_trigger_backendEn_1(fpDq_io_deq_3_bits_cf_trigger_backendEn_1),
    .io_deq_3_bits_cf_pd_isRVC(fpDq_io_deq_3_bits_cf_pd_isRVC),
    .io_deq_3_bits_cf_pd_brType(fpDq_io_deq_3_bits_cf_pd_brType),
    .io_deq_3_bits_cf_pd_isCall(fpDq_io_deq_3_bits_cf_pd_isCall),
    .io_deq_3_bits_cf_pd_isRet(fpDq_io_deq_3_bits_cf_pd_isRet),
    .io_deq_3_bits_cf_pred_taken(fpDq_io_deq_3_bits_cf_pred_taken),
    .io_deq_3_bits_cf_storeSetHit(fpDq_io_deq_3_bits_cf_storeSetHit),
    .io_deq_3_bits_cf_waitForRobIdx_flag(fpDq_io_deq_3_bits_cf_waitForRobIdx_flag),
    .io_deq_3_bits_cf_waitForRobIdx_value(fpDq_io_deq_3_bits_cf_waitForRobIdx_value),
    .io_deq_3_bits_cf_loadWaitBit(fpDq_io_deq_3_bits_cf_loadWaitBit),
    .io_deq_3_bits_cf_loadWaitStrict(fpDq_io_deq_3_bits_cf_loadWaitStrict),
    .io_deq_3_bits_cf_ssid(fpDq_io_deq_3_bits_cf_ssid),
    .io_deq_3_bits_cf_ftqPtr_flag(fpDq_io_deq_3_bits_cf_ftqPtr_flag),
    .io_deq_3_bits_cf_ftqPtr_value(fpDq_io_deq_3_bits_cf_ftqPtr_value),
    .io_deq_3_bits_cf_ftqOffset(fpDq_io_deq_3_bits_cf_ftqOffset),
    .io_deq_3_bits_ctrl_srcType_0(fpDq_io_deq_3_bits_ctrl_srcType_0),
    .io_deq_3_bits_ctrl_srcType_1(fpDq_io_deq_3_bits_ctrl_srcType_1),
    .io_deq_3_bits_ctrl_fuType(fpDq_io_deq_3_bits_ctrl_fuType),
    .io_deq_3_bits_ctrl_fuOpType(fpDq_io_deq_3_bits_ctrl_fuOpType),
    .io_deq_3_bits_ctrl_rfWen(fpDq_io_deq_3_bits_ctrl_rfWen),
    .io_deq_3_bits_ctrl_fpWen(fpDq_io_deq_3_bits_ctrl_fpWen),
    .io_deq_3_bits_ctrl_flushPipe(fpDq_io_deq_3_bits_ctrl_flushPipe),
    .io_deq_3_bits_ctrl_imm(fpDq_io_deq_3_bits_ctrl_imm),
    .io_deq_3_bits_ctrl_replayInst(fpDq_io_deq_3_bits_ctrl_replayInst),
    .io_deq_3_bits_psrc_0(fpDq_io_deq_3_bits_psrc_0),
    .io_deq_3_bits_psrc_1(fpDq_io_deq_3_bits_psrc_1),
    .io_deq_3_bits_pdest(fpDq_io_deq_3_bits_pdest),
    .io_deq_3_bits_robIdx_flag(fpDq_io_deq_3_bits_robIdx_flag),
    .io_deq_3_bits_robIdx_value(fpDq_io_deq_3_bits_robIdx_value),
    .io_redirect_valid(fpDq_io_redirect_valid),
    .io_redirect_bits_robIdx_flag(fpDq_io_redirect_bits_robIdx_flag),
    .io_redirect_bits_robIdx_value(fpDq_io_redirect_bits_robIdx_value),
    .io_redirect_bits_level(fpDq_io_redirect_bits_level),
    .io_deqNext_0_cf_ftqPtr_value(fpDq_io_deqNext_0_cf_ftqPtr_value),
    .io_deqNext_0_cf_ftqOffset(fpDq_io_deqNext_0_cf_ftqOffset),
    .io_deqNext_0_ctrl_srcType_0(fpDq_io_deqNext_0_ctrl_srcType_0),
    .io_deqNext_0_ctrl_srcType_1(fpDq_io_deqNext_0_ctrl_srcType_1),
    .io_deqNext_0_ctrl_srcType_2(fpDq_io_deqNext_0_ctrl_srcType_2),
    .io_deqNext_0_ctrl_fuType(fpDq_io_deqNext_0_ctrl_fuType),
    .io_deqNext_0_ctrl_fuOpType(fpDq_io_deqNext_0_ctrl_fuOpType),
    .io_deqNext_0_ctrl_rfWen(fpDq_io_deqNext_0_ctrl_rfWen),
    .io_deqNext_0_ctrl_fpWen(fpDq_io_deqNext_0_ctrl_fpWen),
    .io_deqNext_0_ctrl_flushPipe(fpDq_io_deqNext_0_ctrl_flushPipe),
    .io_deqNext_0_ctrl_selImm(fpDq_io_deqNext_0_ctrl_selImm),
    .io_deqNext_0_ctrl_imm(fpDq_io_deqNext_0_ctrl_imm),
    .io_deqNext_0_ctrl_replayInst(fpDq_io_deqNext_0_ctrl_replayInst),
    .io_deqNext_0_psrc_0(fpDq_io_deqNext_0_psrc_0),
    .io_deqNext_0_psrc_1(fpDq_io_deqNext_0_psrc_1),
    .io_deqNext_0_psrc_2(fpDq_io_deqNext_0_psrc_2),
    .io_deqNext_0_pdest(fpDq_io_deqNext_0_pdest),
    .io_deqNext_0_robIdx_flag(fpDq_io_deqNext_0_robIdx_flag),
    .io_deqNext_0_robIdx_value(fpDq_io_deqNext_0_robIdx_value),
    .io_deqNext_0_lqIdx_flag(fpDq_io_deqNext_0_lqIdx_flag),
    .io_deqNext_0_lqIdx_value(fpDq_io_deqNext_0_lqIdx_value),
    .io_deqNext_0_sqIdx_flag(fpDq_io_deqNext_0_sqIdx_flag),
    .io_deqNext_0_sqIdx_value(fpDq_io_deqNext_0_sqIdx_value),
    .io_deqNext_1_cf_ftqPtr_value(fpDq_io_deqNext_1_cf_ftqPtr_value),
    .io_deqNext_1_cf_ftqOffset(fpDq_io_deqNext_1_cf_ftqOffset),
    .io_deqNext_1_ctrl_srcType_0(fpDq_io_deqNext_1_ctrl_srcType_0),
    .io_deqNext_1_ctrl_srcType_1(fpDq_io_deqNext_1_ctrl_srcType_1),
    .io_deqNext_1_ctrl_srcType_2(fpDq_io_deqNext_1_ctrl_srcType_2),
    .io_deqNext_1_ctrl_fuType(fpDq_io_deqNext_1_ctrl_fuType),
    .io_deqNext_1_ctrl_fuOpType(fpDq_io_deqNext_1_ctrl_fuOpType),
    .io_deqNext_1_ctrl_rfWen(fpDq_io_deqNext_1_ctrl_rfWen),
    .io_deqNext_1_ctrl_fpWen(fpDq_io_deqNext_1_ctrl_fpWen),
    .io_deqNext_1_ctrl_flushPipe(fpDq_io_deqNext_1_ctrl_flushPipe),
    .io_deqNext_1_ctrl_selImm(fpDq_io_deqNext_1_ctrl_selImm),
    .io_deqNext_1_ctrl_imm(fpDq_io_deqNext_1_ctrl_imm),
    .io_deqNext_1_ctrl_replayInst(fpDq_io_deqNext_1_ctrl_replayInst),
    .io_deqNext_1_psrc_0(fpDq_io_deqNext_1_psrc_0),
    .io_deqNext_1_psrc_1(fpDq_io_deqNext_1_psrc_1),
    .io_deqNext_1_psrc_2(fpDq_io_deqNext_1_psrc_2),
    .io_deqNext_1_pdest(fpDq_io_deqNext_1_pdest),
    .io_deqNext_1_robIdx_flag(fpDq_io_deqNext_1_robIdx_flag),
    .io_deqNext_1_robIdx_value(fpDq_io_deqNext_1_robIdx_value),
    .io_deqNext_1_lqIdx_flag(fpDq_io_deqNext_1_lqIdx_flag),
    .io_deqNext_1_lqIdx_value(fpDq_io_deqNext_1_lqIdx_value),
    .io_deqNext_1_sqIdx_flag(fpDq_io_deqNext_1_sqIdx_flag),
    .io_deqNext_1_sqIdx_value(fpDq_io_deqNext_1_sqIdx_value),
    .io_deqNext_2_cf_ftqPtr_value(fpDq_io_deqNext_2_cf_ftqPtr_value),
    .io_deqNext_2_cf_ftqOffset(fpDq_io_deqNext_2_cf_ftqOffset),
    .io_deqNext_2_ctrl_srcType_0(fpDq_io_deqNext_2_ctrl_srcType_0),
    .io_deqNext_2_ctrl_srcType_1(fpDq_io_deqNext_2_ctrl_srcType_1),
    .io_deqNext_2_ctrl_srcType_2(fpDq_io_deqNext_2_ctrl_srcType_2),
    .io_deqNext_2_ctrl_fuType(fpDq_io_deqNext_2_ctrl_fuType),
    .io_deqNext_2_ctrl_fuOpType(fpDq_io_deqNext_2_ctrl_fuOpType),
    .io_deqNext_2_ctrl_rfWen(fpDq_io_deqNext_2_ctrl_rfWen),
    .io_deqNext_2_ctrl_fpWen(fpDq_io_deqNext_2_ctrl_fpWen),
    .io_deqNext_2_ctrl_flushPipe(fpDq_io_deqNext_2_ctrl_flushPipe),
    .io_deqNext_2_ctrl_selImm(fpDq_io_deqNext_2_ctrl_selImm),
    .io_deqNext_2_ctrl_imm(fpDq_io_deqNext_2_ctrl_imm),
    .io_deqNext_2_ctrl_replayInst(fpDq_io_deqNext_2_ctrl_replayInst),
    .io_deqNext_2_psrc_0(fpDq_io_deqNext_2_psrc_0),
    .io_deqNext_2_psrc_1(fpDq_io_deqNext_2_psrc_1),
    .io_deqNext_2_psrc_2(fpDq_io_deqNext_2_psrc_2),
    .io_deqNext_2_pdest(fpDq_io_deqNext_2_pdest),
    .io_deqNext_2_robIdx_flag(fpDq_io_deqNext_2_robIdx_flag),
    .io_deqNext_2_robIdx_value(fpDq_io_deqNext_2_robIdx_value),
    .io_deqNext_2_lqIdx_flag(fpDq_io_deqNext_2_lqIdx_flag),
    .io_deqNext_2_lqIdx_value(fpDq_io_deqNext_2_lqIdx_value),
    .io_deqNext_2_sqIdx_flag(fpDq_io_deqNext_2_sqIdx_flag),
    .io_deqNext_2_sqIdx_value(fpDq_io_deqNext_2_sqIdx_value),
    .io_deqNext_3_cf_ftqPtr_value(fpDq_io_deqNext_3_cf_ftqPtr_value),
    .io_deqNext_3_cf_ftqOffset(fpDq_io_deqNext_3_cf_ftqOffset),
    .io_deqNext_3_ctrl_srcType_0(fpDq_io_deqNext_3_ctrl_srcType_0),
    .io_deqNext_3_ctrl_srcType_1(fpDq_io_deqNext_3_ctrl_srcType_1),
    .io_deqNext_3_ctrl_srcType_2(fpDq_io_deqNext_3_ctrl_srcType_2),
    .io_deqNext_3_ctrl_fuType(fpDq_io_deqNext_3_ctrl_fuType),
    .io_deqNext_3_ctrl_fuOpType(fpDq_io_deqNext_3_ctrl_fuOpType),
    .io_deqNext_3_ctrl_rfWen(fpDq_io_deqNext_3_ctrl_rfWen),
    .io_deqNext_3_ctrl_fpWen(fpDq_io_deqNext_3_ctrl_fpWen),
    .io_deqNext_3_ctrl_flushPipe(fpDq_io_deqNext_3_ctrl_flushPipe),
    .io_deqNext_3_ctrl_selImm(fpDq_io_deqNext_3_ctrl_selImm),
    .io_deqNext_3_ctrl_imm(fpDq_io_deqNext_3_ctrl_imm),
    .io_deqNext_3_ctrl_replayInst(fpDq_io_deqNext_3_ctrl_replayInst),
    .io_deqNext_3_psrc_0(fpDq_io_deqNext_3_psrc_0),
    .io_deqNext_3_psrc_1(fpDq_io_deqNext_3_psrc_1),
    .io_deqNext_3_psrc_2(fpDq_io_deqNext_3_psrc_2),
    .io_deqNext_3_pdest(fpDq_io_deqNext_3_pdest),
    .io_deqNext_3_robIdx_flag(fpDq_io_deqNext_3_robIdx_flag),
    .io_deqNext_3_robIdx_value(fpDq_io_deqNext_3_robIdx_value),
    .io_deqNext_3_lqIdx_flag(fpDq_io_deqNext_3_lqIdx_flag),
    .io_deqNext_3_lqIdx_value(fpDq_io_deqNext_3_lqIdx_value),
    .io_deqNext_3_sqIdx_flag(fpDq_io_deqNext_3_sqIdx_flag),
    .io_deqNext_3_sqIdx_value(fpDq_io_deqNext_3_sqIdx_value),
    .io_perf_0_value(fpDq_io_perf_0_value),
    .io_perf_1_value(fpDq_io_perf_1_value),
    .io_perf_2_value(fpDq_io_perf_2_value),
    .io_perf_3_value(fpDq_io_perf_3_value),
    .io_perf_4_value(fpDq_io_perf_4_value),
    .io_perf_5_value(fpDq_io_perf_5_value),
    .io_perf_6_value(fpDq_io_perf_6_value),
    .io_perf_7_value(fpDq_io_perf_7_value)
  );
  DispatchQueue lsDq ( // @[CtrlBlock.scala 272:20]
    .clock(lsDq_clock),
    .reset(lsDq_reset),
    .io_enq_canAccept(lsDq_io_enq_canAccept),
    .io_enq_needAlloc_0(lsDq_io_enq_needAlloc_0),
    .io_enq_needAlloc_1(lsDq_io_enq_needAlloc_1),
    .io_enq_req_0_valid(lsDq_io_enq_req_0_valid),
    .io_enq_req_0_bits_cf_foldpc(lsDq_io_enq_req_0_bits_cf_foldpc),
    .io_enq_req_0_bits_cf_trigger_backendEn_0(lsDq_io_enq_req_0_bits_cf_trigger_backendEn_0),
    .io_enq_req_0_bits_cf_trigger_backendEn_1(lsDq_io_enq_req_0_bits_cf_trigger_backendEn_1),
    .io_enq_req_0_bits_cf_pd_isRVC(lsDq_io_enq_req_0_bits_cf_pd_isRVC),
    .io_enq_req_0_bits_cf_pd_brType(lsDq_io_enq_req_0_bits_cf_pd_brType),
    .io_enq_req_0_bits_cf_pd_isCall(lsDq_io_enq_req_0_bits_cf_pd_isCall),
    .io_enq_req_0_bits_cf_pd_isRet(lsDq_io_enq_req_0_bits_cf_pd_isRet),
    .io_enq_req_0_bits_cf_pred_taken(lsDq_io_enq_req_0_bits_cf_pred_taken),
    .io_enq_req_0_bits_cf_storeSetHit(lsDq_io_enq_req_0_bits_cf_storeSetHit),
    .io_enq_req_0_bits_cf_waitForRobIdx_flag(lsDq_io_enq_req_0_bits_cf_waitForRobIdx_flag),
    .io_enq_req_0_bits_cf_waitForRobIdx_value(lsDq_io_enq_req_0_bits_cf_waitForRobIdx_value),
    .io_enq_req_0_bits_cf_loadWaitBit(lsDq_io_enq_req_0_bits_cf_loadWaitBit),
    .io_enq_req_0_bits_cf_loadWaitStrict(lsDq_io_enq_req_0_bits_cf_loadWaitStrict),
    .io_enq_req_0_bits_cf_ssid(lsDq_io_enq_req_0_bits_cf_ssid),
    .io_enq_req_0_bits_cf_ftqPtr_flag(lsDq_io_enq_req_0_bits_cf_ftqPtr_flag),
    .io_enq_req_0_bits_cf_ftqPtr_value(lsDq_io_enq_req_0_bits_cf_ftqPtr_value),
    .io_enq_req_0_bits_cf_ftqOffset(lsDq_io_enq_req_0_bits_cf_ftqOffset),
    .io_enq_req_0_bits_ctrl_srcType_0(lsDq_io_enq_req_0_bits_ctrl_srcType_0),
    .io_enq_req_0_bits_ctrl_srcType_1(lsDq_io_enq_req_0_bits_ctrl_srcType_1),
    .io_enq_req_0_bits_ctrl_srcType_2(lsDq_io_enq_req_0_bits_ctrl_srcType_2),
    .io_enq_req_0_bits_ctrl_fuType(lsDq_io_enq_req_0_bits_ctrl_fuType),
    .io_enq_req_0_bits_ctrl_fuOpType(lsDq_io_enq_req_0_bits_ctrl_fuOpType),
    .io_enq_req_0_bits_ctrl_rfWen(lsDq_io_enq_req_0_bits_ctrl_rfWen),
    .io_enq_req_0_bits_ctrl_fpWen(lsDq_io_enq_req_0_bits_ctrl_fpWen),
    .io_enq_req_0_bits_ctrl_flushPipe(lsDq_io_enq_req_0_bits_ctrl_flushPipe),
    .io_enq_req_0_bits_ctrl_selImm(lsDq_io_enq_req_0_bits_ctrl_selImm),
    .io_enq_req_0_bits_ctrl_imm(lsDq_io_enq_req_0_bits_ctrl_imm),
    .io_enq_req_0_bits_ctrl_fpu_isAddSub(lsDq_io_enq_req_0_bits_ctrl_fpu_isAddSub),
    .io_enq_req_0_bits_ctrl_fpu_typeTagIn(lsDq_io_enq_req_0_bits_ctrl_fpu_typeTagIn),
    .io_enq_req_0_bits_ctrl_fpu_typeTagOut(lsDq_io_enq_req_0_bits_ctrl_fpu_typeTagOut),
    .io_enq_req_0_bits_ctrl_fpu_fromInt(lsDq_io_enq_req_0_bits_ctrl_fpu_fromInt),
    .io_enq_req_0_bits_ctrl_fpu_wflags(lsDq_io_enq_req_0_bits_ctrl_fpu_wflags),
    .io_enq_req_0_bits_ctrl_fpu_fpWen(lsDq_io_enq_req_0_bits_ctrl_fpu_fpWen),
    .io_enq_req_0_bits_ctrl_fpu_fmaCmd(lsDq_io_enq_req_0_bits_ctrl_fpu_fmaCmd),
    .io_enq_req_0_bits_ctrl_fpu_div(lsDq_io_enq_req_0_bits_ctrl_fpu_div),
    .io_enq_req_0_bits_ctrl_fpu_sqrt(lsDq_io_enq_req_0_bits_ctrl_fpu_sqrt),
    .io_enq_req_0_bits_ctrl_fpu_fcvt(lsDq_io_enq_req_0_bits_ctrl_fpu_fcvt),
    .io_enq_req_0_bits_ctrl_fpu_typ(lsDq_io_enq_req_0_bits_ctrl_fpu_typ),
    .io_enq_req_0_bits_ctrl_fpu_fmt(lsDq_io_enq_req_0_bits_ctrl_fpu_fmt),
    .io_enq_req_0_bits_ctrl_fpu_ren3(lsDq_io_enq_req_0_bits_ctrl_fpu_ren3),
    .io_enq_req_0_bits_ctrl_fpu_rm(lsDq_io_enq_req_0_bits_ctrl_fpu_rm),
    .io_enq_req_0_bits_psrc_0(lsDq_io_enq_req_0_bits_psrc_0),
    .io_enq_req_0_bits_psrc_1(lsDq_io_enq_req_0_bits_psrc_1),
    .io_enq_req_0_bits_psrc_2(lsDq_io_enq_req_0_bits_psrc_2),
    .io_enq_req_0_bits_pdest(lsDq_io_enq_req_0_bits_pdest),
    .io_enq_req_0_bits_robIdx_flag(lsDq_io_enq_req_0_bits_robIdx_flag),
    .io_enq_req_0_bits_robIdx_value(lsDq_io_enq_req_0_bits_robIdx_value),
    .io_enq_req_1_valid(lsDq_io_enq_req_1_valid),
    .io_enq_req_1_bits_cf_foldpc(lsDq_io_enq_req_1_bits_cf_foldpc),
    .io_enq_req_1_bits_cf_trigger_backendEn_0(lsDq_io_enq_req_1_bits_cf_trigger_backendEn_0),
    .io_enq_req_1_bits_cf_trigger_backendEn_1(lsDq_io_enq_req_1_bits_cf_trigger_backendEn_1),
    .io_enq_req_1_bits_cf_pd_isRVC(lsDq_io_enq_req_1_bits_cf_pd_isRVC),
    .io_enq_req_1_bits_cf_pd_brType(lsDq_io_enq_req_1_bits_cf_pd_brType),
    .io_enq_req_1_bits_cf_pd_isCall(lsDq_io_enq_req_1_bits_cf_pd_isCall),
    .io_enq_req_1_bits_cf_pd_isRet(lsDq_io_enq_req_1_bits_cf_pd_isRet),
    .io_enq_req_1_bits_cf_pred_taken(lsDq_io_enq_req_1_bits_cf_pred_taken),
    .io_enq_req_1_bits_cf_storeSetHit(lsDq_io_enq_req_1_bits_cf_storeSetHit),
    .io_enq_req_1_bits_cf_waitForRobIdx_flag(lsDq_io_enq_req_1_bits_cf_waitForRobIdx_flag),
    .io_enq_req_1_bits_cf_waitForRobIdx_value(lsDq_io_enq_req_1_bits_cf_waitForRobIdx_value),
    .io_enq_req_1_bits_cf_loadWaitBit(lsDq_io_enq_req_1_bits_cf_loadWaitBit),
    .io_enq_req_1_bits_cf_loadWaitStrict(lsDq_io_enq_req_1_bits_cf_loadWaitStrict),
    .io_enq_req_1_bits_cf_ssid(lsDq_io_enq_req_1_bits_cf_ssid),
    .io_enq_req_1_bits_cf_ftqPtr_flag(lsDq_io_enq_req_1_bits_cf_ftqPtr_flag),
    .io_enq_req_1_bits_cf_ftqPtr_value(lsDq_io_enq_req_1_bits_cf_ftqPtr_value),
    .io_enq_req_1_bits_cf_ftqOffset(lsDq_io_enq_req_1_bits_cf_ftqOffset),
    .io_enq_req_1_bits_ctrl_srcType_0(lsDq_io_enq_req_1_bits_ctrl_srcType_0),
    .io_enq_req_1_bits_ctrl_srcType_1(lsDq_io_enq_req_1_bits_ctrl_srcType_1),
    .io_enq_req_1_bits_ctrl_srcType_2(lsDq_io_enq_req_1_bits_ctrl_srcType_2),
    .io_enq_req_1_bits_ctrl_fuType(lsDq_io_enq_req_1_bits_ctrl_fuType),
    .io_enq_req_1_bits_ctrl_fuOpType(lsDq_io_enq_req_1_bits_ctrl_fuOpType),
    .io_enq_req_1_bits_ctrl_rfWen(lsDq_io_enq_req_1_bits_ctrl_rfWen),
    .io_enq_req_1_bits_ctrl_fpWen(lsDq_io_enq_req_1_bits_ctrl_fpWen),
    .io_enq_req_1_bits_ctrl_flushPipe(lsDq_io_enq_req_1_bits_ctrl_flushPipe),
    .io_enq_req_1_bits_ctrl_selImm(lsDq_io_enq_req_1_bits_ctrl_selImm),
    .io_enq_req_1_bits_ctrl_imm(lsDq_io_enq_req_1_bits_ctrl_imm),
    .io_enq_req_1_bits_ctrl_fpu_isAddSub(lsDq_io_enq_req_1_bits_ctrl_fpu_isAddSub),
    .io_enq_req_1_bits_ctrl_fpu_typeTagIn(lsDq_io_enq_req_1_bits_ctrl_fpu_typeTagIn),
    .io_enq_req_1_bits_ctrl_fpu_typeTagOut(lsDq_io_enq_req_1_bits_ctrl_fpu_typeTagOut),
    .io_enq_req_1_bits_ctrl_fpu_fromInt(lsDq_io_enq_req_1_bits_ctrl_fpu_fromInt),
    .io_enq_req_1_bits_ctrl_fpu_wflags(lsDq_io_enq_req_1_bits_ctrl_fpu_wflags),
    .io_enq_req_1_bits_ctrl_fpu_fpWen(lsDq_io_enq_req_1_bits_ctrl_fpu_fpWen),
    .io_enq_req_1_bits_ctrl_fpu_fmaCmd(lsDq_io_enq_req_1_bits_ctrl_fpu_fmaCmd),
    .io_enq_req_1_bits_ctrl_fpu_div(lsDq_io_enq_req_1_bits_ctrl_fpu_div),
    .io_enq_req_1_bits_ctrl_fpu_sqrt(lsDq_io_enq_req_1_bits_ctrl_fpu_sqrt),
    .io_enq_req_1_bits_ctrl_fpu_fcvt(lsDq_io_enq_req_1_bits_ctrl_fpu_fcvt),
    .io_enq_req_1_bits_ctrl_fpu_typ(lsDq_io_enq_req_1_bits_ctrl_fpu_typ),
    .io_enq_req_1_bits_ctrl_fpu_fmt(lsDq_io_enq_req_1_bits_ctrl_fpu_fmt),
    .io_enq_req_1_bits_ctrl_fpu_ren3(lsDq_io_enq_req_1_bits_ctrl_fpu_ren3),
    .io_enq_req_1_bits_ctrl_fpu_rm(lsDq_io_enq_req_1_bits_ctrl_fpu_rm),
    .io_enq_req_1_bits_psrc_0(lsDq_io_enq_req_1_bits_psrc_0),
    .io_enq_req_1_bits_psrc_1(lsDq_io_enq_req_1_bits_psrc_1),
    .io_enq_req_1_bits_psrc_2(lsDq_io_enq_req_1_bits_psrc_2),
    .io_enq_req_1_bits_pdest(lsDq_io_enq_req_1_bits_pdest),
    .io_enq_req_1_bits_robIdx_flag(lsDq_io_enq_req_1_bits_robIdx_flag),
    .io_enq_req_1_bits_robIdx_value(lsDq_io_enq_req_1_bits_robIdx_value),
    .io_deq_0_ready(lsDq_io_deq_0_ready),
    .io_deq_0_valid(lsDq_io_deq_0_valid),
    .io_deq_0_bits_cf_foldpc(lsDq_io_deq_0_bits_cf_foldpc),
    .io_deq_0_bits_cf_trigger_backendEn_0(lsDq_io_deq_0_bits_cf_trigger_backendEn_0),
    .io_deq_0_bits_cf_trigger_backendEn_1(lsDq_io_deq_0_bits_cf_trigger_backendEn_1),
    .io_deq_0_bits_cf_pd_isRVC(lsDq_io_deq_0_bits_cf_pd_isRVC),
    .io_deq_0_bits_cf_pd_brType(lsDq_io_deq_0_bits_cf_pd_brType),
    .io_deq_0_bits_cf_pd_isCall(lsDq_io_deq_0_bits_cf_pd_isCall),
    .io_deq_0_bits_cf_pd_isRet(lsDq_io_deq_0_bits_cf_pd_isRet),
    .io_deq_0_bits_cf_pred_taken(lsDq_io_deq_0_bits_cf_pred_taken),
    .io_deq_0_bits_cf_storeSetHit(lsDq_io_deq_0_bits_cf_storeSetHit),
    .io_deq_0_bits_cf_waitForRobIdx_flag(lsDq_io_deq_0_bits_cf_waitForRobIdx_flag),
    .io_deq_0_bits_cf_waitForRobIdx_value(lsDq_io_deq_0_bits_cf_waitForRobIdx_value),
    .io_deq_0_bits_cf_loadWaitBit(lsDq_io_deq_0_bits_cf_loadWaitBit),
    .io_deq_0_bits_cf_loadWaitStrict(lsDq_io_deq_0_bits_cf_loadWaitStrict),
    .io_deq_0_bits_cf_ssid(lsDq_io_deq_0_bits_cf_ssid),
    .io_deq_0_bits_cf_ftqPtr_flag(lsDq_io_deq_0_bits_cf_ftqPtr_flag),
    .io_deq_0_bits_cf_ftqPtr_value(lsDq_io_deq_0_bits_cf_ftqPtr_value),
    .io_deq_0_bits_cf_ftqOffset(lsDq_io_deq_0_bits_cf_ftqOffset),
    .io_deq_0_bits_ctrl_srcType_0(lsDq_io_deq_0_bits_ctrl_srcType_0),
    .io_deq_0_bits_ctrl_srcType_1(lsDq_io_deq_0_bits_ctrl_srcType_1),
    .io_deq_0_bits_ctrl_srcType_2(lsDq_io_deq_0_bits_ctrl_srcType_2),
    .io_deq_0_bits_ctrl_fuType(lsDq_io_deq_0_bits_ctrl_fuType),
    .io_deq_0_bits_ctrl_fuOpType(lsDq_io_deq_0_bits_ctrl_fuOpType),
    .io_deq_0_bits_ctrl_rfWen(lsDq_io_deq_0_bits_ctrl_rfWen),
    .io_deq_0_bits_ctrl_fpWen(lsDq_io_deq_0_bits_ctrl_fpWen),
    .io_deq_0_bits_ctrl_flushPipe(lsDq_io_deq_0_bits_ctrl_flushPipe),
    .io_deq_0_bits_ctrl_selImm(lsDq_io_deq_0_bits_ctrl_selImm),
    .io_deq_0_bits_ctrl_imm(lsDq_io_deq_0_bits_ctrl_imm),
    .io_deq_0_bits_ctrl_fpu_isAddSub(lsDq_io_deq_0_bits_ctrl_fpu_isAddSub),
    .io_deq_0_bits_ctrl_fpu_typeTagIn(lsDq_io_deq_0_bits_ctrl_fpu_typeTagIn),
    .io_deq_0_bits_ctrl_fpu_typeTagOut(lsDq_io_deq_0_bits_ctrl_fpu_typeTagOut),
    .io_deq_0_bits_ctrl_fpu_fromInt(lsDq_io_deq_0_bits_ctrl_fpu_fromInt),
    .io_deq_0_bits_ctrl_fpu_wflags(lsDq_io_deq_0_bits_ctrl_fpu_wflags),
    .io_deq_0_bits_ctrl_fpu_fpWen(lsDq_io_deq_0_bits_ctrl_fpu_fpWen),
    .io_deq_0_bits_ctrl_fpu_fmaCmd(lsDq_io_deq_0_bits_ctrl_fpu_fmaCmd),
    .io_deq_0_bits_ctrl_fpu_div(lsDq_io_deq_0_bits_ctrl_fpu_div),
    .io_deq_0_bits_ctrl_fpu_sqrt(lsDq_io_deq_0_bits_ctrl_fpu_sqrt),
    .io_deq_0_bits_ctrl_fpu_fcvt(lsDq_io_deq_0_bits_ctrl_fpu_fcvt),
    .io_deq_0_bits_ctrl_fpu_typ(lsDq_io_deq_0_bits_ctrl_fpu_typ),
    .io_deq_0_bits_ctrl_fpu_fmt(lsDq_io_deq_0_bits_ctrl_fpu_fmt),
    .io_deq_0_bits_ctrl_fpu_ren3(lsDq_io_deq_0_bits_ctrl_fpu_ren3),
    .io_deq_0_bits_ctrl_fpu_rm(lsDq_io_deq_0_bits_ctrl_fpu_rm),
    .io_deq_0_bits_ctrl_replayInst(lsDq_io_deq_0_bits_ctrl_replayInst),
    .io_deq_0_bits_psrc_0(lsDq_io_deq_0_bits_psrc_0),
    .io_deq_0_bits_psrc_1(lsDq_io_deq_0_bits_psrc_1),
    .io_deq_0_bits_psrc_2(lsDq_io_deq_0_bits_psrc_2),
    .io_deq_0_bits_pdest(lsDq_io_deq_0_bits_pdest),
    .io_deq_0_bits_robIdx_flag(lsDq_io_deq_0_bits_robIdx_flag),
    .io_deq_0_bits_robIdx_value(lsDq_io_deq_0_bits_robIdx_value),
    .io_deq_0_bits_lqIdx_flag(lsDq_io_deq_0_bits_lqIdx_flag),
    .io_deq_0_bits_lqIdx_value(lsDq_io_deq_0_bits_lqIdx_value),
    .io_deq_0_bits_sqIdx_flag(lsDq_io_deq_0_bits_sqIdx_flag),
    .io_deq_0_bits_sqIdx_value(lsDq_io_deq_0_bits_sqIdx_value),
    .io_deq_1_ready(lsDq_io_deq_1_ready),
    .io_deq_1_valid(lsDq_io_deq_1_valid),
    .io_deq_1_bits_cf_foldpc(lsDq_io_deq_1_bits_cf_foldpc),
    .io_deq_1_bits_cf_trigger_backendEn_0(lsDq_io_deq_1_bits_cf_trigger_backendEn_0),
    .io_deq_1_bits_cf_trigger_backendEn_1(lsDq_io_deq_1_bits_cf_trigger_backendEn_1),
    .io_deq_1_bits_cf_pd_isRVC(lsDq_io_deq_1_bits_cf_pd_isRVC),
    .io_deq_1_bits_cf_pd_brType(lsDq_io_deq_1_bits_cf_pd_brType),
    .io_deq_1_bits_cf_pd_isCall(lsDq_io_deq_1_bits_cf_pd_isCall),
    .io_deq_1_bits_cf_pd_isRet(lsDq_io_deq_1_bits_cf_pd_isRet),
    .io_deq_1_bits_cf_pred_taken(lsDq_io_deq_1_bits_cf_pred_taken),
    .io_deq_1_bits_cf_storeSetHit(lsDq_io_deq_1_bits_cf_storeSetHit),
    .io_deq_1_bits_cf_waitForRobIdx_flag(lsDq_io_deq_1_bits_cf_waitForRobIdx_flag),
    .io_deq_1_bits_cf_waitForRobIdx_value(lsDq_io_deq_1_bits_cf_waitForRobIdx_value),
    .io_deq_1_bits_cf_loadWaitBit(lsDq_io_deq_1_bits_cf_loadWaitBit),
    .io_deq_1_bits_cf_loadWaitStrict(lsDq_io_deq_1_bits_cf_loadWaitStrict),
    .io_deq_1_bits_cf_ssid(lsDq_io_deq_1_bits_cf_ssid),
    .io_deq_1_bits_cf_ftqPtr_flag(lsDq_io_deq_1_bits_cf_ftqPtr_flag),
    .io_deq_1_bits_cf_ftqPtr_value(lsDq_io_deq_1_bits_cf_ftqPtr_value),
    .io_deq_1_bits_cf_ftqOffset(lsDq_io_deq_1_bits_cf_ftqOffset),
    .io_deq_1_bits_ctrl_srcType_0(lsDq_io_deq_1_bits_ctrl_srcType_0),
    .io_deq_1_bits_ctrl_srcType_1(lsDq_io_deq_1_bits_ctrl_srcType_1),
    .io_deq_1_bits_ctrl_fuType(lsDq_io_deq_1_bits_ctrl_fuType),
    .io_deq_1_bits_ctrl_fuOpType(lsDq_io_deq_1_bits_ctrl_fuOpType),
    .io_deq_1_bits_ctrl_rfWen(lsDq_io_deq_1_bits_ctrl_rfWen),
    .io_deq_1_bits_ctrl_fpWen(lsDq_io_deq_1_bits_ctrl_fpWen),
    .io_deq_1_bits_ctrl_flushPipe(lsDq_io_deq_1_bits_ctrl_flushPipe),
    .io_deq_1_bits_ctrl_selImm(lsDq_io_deq_1_bits_ctrl_selImm),
    .io_deq_1_bits_ctrl_imm(lsDq_io_deq_1_bits_ctrl_imm),
    .io_deq_1_bits_ctrl_replayInst(lsDq_io_deq_1_bits_ctrl_replayInst),
    .io_deq_1_bits_psrc_0(lsDq_io_deq_1_bits_psrc_0),
    .io_deq_1_bits_psrc_1(lsDq_io_deq_1_bits_psrc_1),
    .io_deq_1_bits_pdest(lsDq_io_deq_1_bits_pdest),
    .io_deq_1_bits_robIdx_flag(lsDq_io_deq_1_bits_robIdx_flag),
    .io_deq_1_bits_robIdx_value(lsDq_io_deq_1_bits_robIdx_value),
    .io_deq_1_bits_lqIdx_flag(lsDq_io_deq_1_bits_lqIdx_flag),
    .io_deq_1_bits_lqIdx_value(lsDq_io_deq_1_bits_lqIdx_value),
    .io_deq_1_bits_sqIdx_flag(lsDq_io_deq_1_bits_sqIdx_flag),
    .io_deq_1_bits_sqIdx_value(lsDq_io_deq_1_bits_sqIdx_value),
    .io_deq_2_ready(lsDq_io_deq_2_ready),
    .io_deq_2_valid(lsDq_io_deq_2_valid),
    .io_deq_2_bits_cf_foldpc(lsDq_io_deq_2_bits_cf_foldpc),
    .io_deq_2_bits_cf_trigger_backendEn_0(lsDq_io_deq_2_bits_cf_trigger_backendEn_0),
    .io_deq_2_bits_cf_trigger_backendEn_1(lsDq_io_deq_2_bits_cf_trigger_backendEn_1),
    .io_deq_2_bits_cf_pd_isRVC(lsDq_io_deq_2_bits_cf_pd_isRVC),
    .io_deq_2_bits_cf_pd_brType(lsDq_io_deq_2_bits_cf_pd_brType),
    .io_deq_2_bits_cf_pd_isCall(lsDq_io_deq_2_bits_cf_pd_isCall),
    .io_deq_2_bits_cf_pd_isRet(lsDq_io_deq_2_bits_cf_pd_isRet),
    .io_deq_2_bits_cf_pred_taken(lsDq_io_deq_2_bits_cf_pred_taken),
    .io_deq_2_bits_cf_storeSetHit(lsDq_io_deq_2_bits_cf_storeSetHit),
    .io_deq_2_bits_cf_waitForRobIdx_flag(lsDq_io_deq_2_bits_cf_waitForRobIdx_flag),
    .io_deq_2_bits_cf_waitForRobIdx_value(lsDq_io_deq_2_bits_cf_waitForRobIdx_value),
    .io_deq_2_bits_cf_loadWaitBit(lsDq_io_deq_2_bits_cf_loadWaitBit),
    .io_deq_2_bits_cf_loadWaitStrict(lsDq_io_deq_2_bits_cf_loadWaitStrict),
    .io_deq_2_bits_cf_ssid(lsDq_io_deq_2_bits_cf_ssid),
    .io_deq_2_bits_cf_ftqPtr_flag(lsDq_io_deq_2_bits_cf_ftqPtr_flag),
    .io_deq_2_bits_cf_ftqPtr_value(lsDq_io_deq_2_bits_cf_ftqPtr_value),
    .io_deq_2_bits_cf_ftqOffset(lsDq_io_deq_2_bits_cf_ftqOffset),
    .io_deq_2_bits_ctrl_srcType_0(lsDq_io_deq_2_bits_ctrl_srcType_0),
    .io_deq_2_bits_ctrl_srcType_1(lsDq_io_deq_2_bits_ctrl_srcType_1),
    .io_deq_2_bits_ctrl_fuType(lsDq_io_deq_2_bits_ctrl_fuType),
    .io_deq_2_bits_ctrl_fuOpType(lsDq_io_deq_2_bits_ctrl_fuOpType),
    .io_deq_2_bits_ctrl_rfWen(lsDq_io_deq_2_bits_ctrl_rfWen),
    .io_deq_2_bits_ctrl_fpWen(lsDq_io_deq_2_bits_ctrl_fpWen),
    .io_deq_2_bits_ctrl_flushPipe(lsDq_io_deq_2_bits_ctrl_flushPipe),
    .io_deq_2_bits_ctrl_imm(lsDq_io_deq_2_bits_ctrl_imm),
    .io_deq_2_bits_ctrl_replayInst(lsDq_io_deq_2_bits_ctrl_replayInst),
    .io_deq_2_bits_psrc_0(lsDq_io_deq_2_bits_psrc_0),
    .io_deq_2_bits_psrc_1(lsDq_io_deq_2_bits_psrc_1),
    .io_deq_2_bits_pdest(lsDq_io_deq_2_bits_pdest),
    .io_deq_2_bits_robIdx_flag(lsDq_io_deq_2_bits_robIdx_flag),
    .io_deq_2_bits_robIdx_value(lsDq_io_deq_2_bits_robIdx_value),
    .io_deq_3_ready(lsDq_io_deq_3_ready),
    .io_deq_3_valid(lsDq_io_deq_3_valid),
    .io_deq_3_bits_cf_foldpc(lsDq_io_deq_3_bits_cf_foldpc),
    .io_deq_3_bits_cf_trigger_backendEn_0(lsDq_io_deq_3_bits_cf_trigger_backendEn_0),
    .io_deq_3_bits_cf_trigger_backendEn_1(lsDq_io_deq_3_bits_cf_trigger_backendEn_1),
    .io_deq_3_bits_cf_pd_isRVC(lsDq_io_deq_3_bits_cf_pd_isRVC),
    .io_deq_3_bits_cf_pd_brType(lsDq_io_deq_3_bits_cf_pd_brType),
    .io_deq_3_bits_cf_pd_isCall(lsDq_io_deq_3_bits_cf_pd_isCall),
    .io_deq_3_bits_cf_pd_isRet(lsDq_io_deq_3_bits_cf_pd_isRet),
    .io_deq_3_bits_cf_pred_taken(lsDq_io_deq_3_bits_cf_pred_taken),
    .io_deq_3_bits_cf_storeSetHit(lsDq_io_deq_3_bits_cf_storeSetHit),
    .io_deq_3_bits_cf_waitForRobIdx_flag(lsDq_io_deq_3_bits_cf_waitForRobIdx_flag),
    .io_deq_3_bits_cf_waitForRobIdx_value(lsDq_io_deq_3_bits_cf_waitForRobIdx_value),
    .io_deq_3_bits_cf_loadWaitBit(lsDq_io_deq_3_bits_cf_loadWaitBit),
    .io_deq_3_bits_cf_loadWaitStrict(lsDq_io_deq_3_bits_cf_loadWaitStrict),
    .io_deq_3_bits_cf_ssid(lsDq_io_deq_3_bits_cf_ssid),
    .io_deq_3_bits_cf_ftqPtr_flag(lsDq_io_deq_3_bits_cf_ftqPtr_flag),
    .io_deq_3_bits_cf_ftqPtr_value(lsDq_io_deq_3_bits_cf_ftqPtr_value),
    .io_deq_3_bits_cf_ftqOffset(lsDq_io_deq_3_bits_cf_ftqOffset),
    .io_deq_3_bits_ctrl_srcType_0(lsDq_io_deq_3_bits_ctrl_srcType_0),
    .io_deq_3_bits_ctrl_srcType_1(lsDq_io_deq_3_bits_ctrl_srcType_1),
    .io_deq_3_bits_ctrl_fuType(lsDq_io_deq_3_bits_ctrl_fuType),
    .io_deq_3_bits_ctrl_fuOpType(lsDq_io_deq_3_bits_ctrl_fuOpType),
    .io_deq_3_bits_ctrl_rfWen(lsDq_io_deq_3_bits_ctrl_rfWen),
    .io_deq_3_bits_ctrl_fpWen(lsDq_io_deq_3_bits_ctrl_fpWen),
    .io_deq_3_bits_ctrl_flushPipe(lsDq_io_deq_3_bits_ctrl_flushPipe),
    .io_deq_3_bits_ctrl_imm(lsDq_io_deq_3_bits_ctrl_imm),
    .io_deq_3_bits_ctrl_replayInst(lsDq_io_deq_3_bits_ctrl_replayInst),
    .io_deq_3_bits_psrc_0(lsDq_io_deq_3_bits_psrc_0),
    .io_deq_3_bits_psrc_1(lsDq_io_deq_3_bits_psrc_1),
    .io_deq_3_bits_pdest(lsDq_io_deq_3_bits_pdest),
    .io_deq_3_bits_robIdx_flag(lsDq_io_deq_3_bits_robIdx_flag),
    .io_deq_3_bits_robIdx_value(lsDq_io_deq_3_bits_robIdx_value),
    .io_redirect_valid(lsDq_io_redirect_valid),
    .io_redirect_bits_robIdx_flag(lsDq_io_redirect_bits_robIdx_flag),
    .io_redirect_bits_robIdx_value(lsDq_io_redirect_bits_robIdx_value),
    .io_redirect_bits_level(lsDq_io_redirect_bits_level),
    .io_deqNext_0_cf_ftqPtr_value(lsDq_io_deqNext_0_cf_ftqPtr_value),
    .io_deqNext_0_cf_ftqOffset(lsDq_io_deqNext_0_cf_ftqOffset),
    .io_deqNext_0_ctrl_srcType_0(lsDq_io_deqNext_0_ctrl_srcType_0),
    .io_deqNext_0_ctrl_srcType_1(lsDq_io_deqNext_0_ctrl_srcType_1),
    .io_deqNext_0_ctrl_srcType_2(lsDq_io_deqNext_0_ctrl_srcType_2),
    .io_deqNext_0_ctrl_fuType(lsDq_io_deqNext_0_ctrl_fuType),
    .io_deqNext_0_ctrl_fuOpType(lsDq_io_deqNext_0_ctrl_fuOpType),
    .io_deqNext_0_ctrl_rfWen(lsDq_io_deqNext_0_ctrl_rfWen),
    .io_deqNext_0_ctrl_fpWen(lsDq_io_deqNext_0_ctrl_fpWen),
    .io_deqNext_0_ctrl_flushPipe(lsDq_io_deqNext_0_ctrl_flushPipe),
    .io_deqNext_0_ctrl_selImm(lsDq_io_deqNext_0_ctrl_selImm),
    .io_deqNext_0_ctrl_imm(lsDq_io_deqNext_0_ctrl_imm),
    .io_deqNext_0_ctrl_replayInst(lsDq_io_deqNext_0_ctrl_replayInst),
    .io_deqNext_0_psrc_0(lsDq_io_deqNext_0_psrc_0),
    .io_deqNext_0_psrc_1(lsDq_io_deqNext_0_psrc_1),
    .io_deqNext_0_psrc_2(lsDq_io_deqNext_0_psrc_2),
    .io_deqNext_0_pdest(lsDq_io_deqNext_0_pdest),
    .io_deqNext_0_robIdx_flag(lsDq_io_deqNext_0_robIdx_flag),
    .io_deqNext_0_robIdx_value(lsDq_io_deqNext_0_robIdx_value),
    .io_deqNext_0_lqIdx_flag(lsDq_io_deqNext_0_lqIdx_flag),
    .io_deqNext_0_lqIdx_value(lsDq_io_deqNext_0_lqIdx_value),
    .io_deqNext_0_sqIdx_flag(lsDq_io_deqNext_0_sqIdx_flag),
    .io_deqNext_0_sqIdx_value(lsDq_io_deqNext_0_sqIdx_value),
    .io_deqNext_1_cf_ftqPtr_value(lsDq_io_deqNext_1_cf_ftqPtr_value),
    .io_deqNext_1_cf_ftqOffset(lsDq_io_deqNext_1_cf_ftqOffset),
    .io_deqNext_1_ctrl_srcType_0(lsDq_io_deqNext_1_ctrl_srcType_0),
    .io_deqNext_1_ctrl_srcType_1(lsDq_io_deqNext_1_ctrl_srcType_1),
    .io_deqNext_1_ctrl_srcType_2(lsDq_io_deqNext_1_ctrl_srcType_2),
    .io_deqNext_1_ctrl_fuType(lsDq_io_deqNext_1_ctrl_fuType),
    .io_deqNext_1_ctrl_fuOpType(lsDq_io_deqNext_1_ctrl_fuOpType),
    .io_deqNext_1_ctrl_rfWen(lsDq_io_deqNext_1_ctrl_rfWen),
    .io_deqNext_1_ctrl_fpWen(lsDq_io_deqNext_1_ctrl_fpWen),
    .io_deqNext_1_ctrl_flushPipe(lsDq_io_deqNext_1_ctrl_flushPipe),
    .io_deqNext_1_ctrl_selImm(lsDq_io_deqNext_1_ctrl_selImm),
    .io_deqNext_1_ctrl_imm(lsDq_io_deqNext_1_ctrl_imm),
    .io_deqNext_1_ctrl_replayInst(lsDq_io_deqNext_1_ctrl_replayInst),
    .io_deqNext_1_psrc_0(lsDq_io_deqNext_1_psrc_0),
    .io_deqNext_1_psrc_1(lsDq_io_deqNext_1_psrc_1),
    .io_deqNext_1_psrc_2(lsDq_io_deqNext_1_psrc_2),
    .io_deqNext_1_pdest(lsDq_io_deqNext_1_pdest),
    .io_deqNext_1_robIdx_flag(lsDq_io_deqNext_1_robIdx_flag),
    .io_deqNext_1_robIdx_value(lsDq_io_deqNext_1_robIdx_value),
    .io_deqNext_1_lqIdx_flag(lsDq_io_deqNext_1_lqIdx_flag),
    .io_deqNext_1_lqIdx_value(lsDq_io_deqNext_1_lqIdx_value),
    .io_deqNext_1_sqIdx_flag(lsDq_io_deqNext_1_sqIdx_flag),
    .io_deqNext_1_sqIdx_value(lsDq_io_deqNext_1_sqIdx_value),
    .io_deqNext_2_cf_ftqPtr_value(lsDq_io_deqNext_2_cf_ftqPtr_value),
    .io_deqNext_2_cf_ftqOffset(lsDq_io_deqNext_2_cf_ftqOffset),
    .io_deqNext_2_ctrl_srcType_0(lsDq_io_deqNext_2_ctrl_srcType_0),
    .io_deqNext_2_ctrl_srcType_1(lsDq_io_deqNext_2_ctrl_srcType_1),
    .io_deqNext_2_ctrl_srcType_2(lsDq_io_deqNext_2_ctrl_srcType_2),
    .io_deqNext_2_ctrl_fuType(lsDq_io_deqNext_2_ctrl_fuType),
    .io_deqNext_2_ctrl_fuOpType(lsDq_io_deqNext_2_ctrl_fuOpType),
    .io_deqNext_2_ctrl_rfWen(lsDq_io_deqNext_2_ctrl_rfWen),
    .io_deqNext_2_ctrl_fpWen(lsDq_io_deqNext_2_ctrl_fpWen),
    .io_deqNext_2_ctrl_flushPipe(lsDq_io_deqNext_2_ctrl_flushPipe),
    .io_deqNext_2_ctrl_selImm(lsDq_io_deqNext_2_ctrl_selImm),
    .io_deqNext_2_ctrl_imm(lsDq_io_deqNext_2_ctrl_imm),
    .io_deqNext_2_ctrl_replayInst(lsDq_io_deqNext_2_ctrl_replayInst),
    .io_deqNext_2_psrc_0(lsDq_io_deqNext_2_psrc_0),
    .io_deqNext_2_psrc_1(lsDq_io_deqNext_2_psrc_1),
    .io_deqNext_2_psrc_2(lsDq_io_deqNext_2_psrc_2),
    .io_deqNext_2_pdest(lsDq_io_deqNext_2_pdest),
    .io_deqNext_2_robIdx_flag(lsDq_io_deqNext_2_robIdx_flag),
    .io_deqNext_2_robIdx_value(lsDq_io_deqNext_2_robIdx_value),
    .io_deqNext_2_lqIdx_flag(lsDq_io_deqNext_2_lqIdx_flag),
    .io_deqNext_2_lqIdx_value(lsDq_io_deqNext_2_lqIdx_value),
    .io_deqNext_2_sqIdx_flag(lsDq_io_deqNext_2_sqIdx_flag),
    .io_deqNext_2_sqIdx_value(lsDq_io_deqNext_2_sqIdx_value),
    .io_deqNext_3_cf_ftqPtr_value(lsDq_io_deqNext_3_cf_ftqPtr_value),
    .io_deqNext_3_cf_ftqOffset(lsDq_io_deqNext_3_cf_ftqOffset),
    .io_deqNext_3_ctrl_srcType_0(lsDq_io_deqNext_3_ctrl_srcType_0),
    .io_deqNext_3_ctrl_srcType_1(lsDq_io_deqNext_3_ctrl_srcType_1),
    .io_deqNext_3_ctrl_srcType_2(lsDq_io_deqNext_3_ctrl_srcType_2),
    .io_deqNext_3_ctrl_fuType(lsDq_io_deqNext_3_ctrl_fuType),
    .io_deqNext_3_ctrl_fuOpType(lsDq_io_deqNext_3_ctrl_fuOpType),
    .io_deqNext_3_ctrl_rfWen(lsDq_io_deqNext_3_ctrl_rfWen),
    .io_deqNext_3_ctrl_fpWen(lsDq_io_deqNext_3_ctrl_fpWen),
    .io_deqNext_3_ctrl_flushPipe(lsDq_io_deqNext_3_ctrl_flushPipe),
    .io_deqNext_3_ctrl_selImm(lsDq_io_deqNext_3_ctrl_selImm),
    .io_deqNext_3_ctrl_imm(lsDq_io_deqNext_3_ctrl_imm),
    .io_deqNext_3_ctrl_replayInst(lsDq_io_deqNext_3_ctrl_replayInst),
    .io_deqNext_3_psrc_0(lsDq_io_deqNext_3_psrc_0),
    .io_deqNext_3_psrc_1(lsDq_io_deqNext_3_psrc_1),
    .io_deqNext_3_psrc_2(lsDq_io_deqNext_3_psrc_2),
    .io_deqNext_3_pdest(lsDq_io_deqNext_3_pdest),
    .io_deqNext_3_robIdx_flag(lsDq_io_deqNext_3_robIdx_flag),
    .io_deqNext_3_robIdx_value(lsDq_io_deqNext_3_robIdx_value),
    .io_deqNext_3_lqIdx_flag(lsDq_io_deqNext_3_lqIdx_flag),
    .io_deqNext_3_lqIdx_value(lsDq_io_deqNext_3_lqIdx_value),
    .io_deqNext_3_sqIdx_flag(lsDq_io_deqNext_3_sqIdx_flag),
    .io_deqNext_3_sqIdx_value(lsDq_io_deqNext_3_sqIdx_value),
    .io_perf_0_value(lsDq_io_perf_0_value),
    .io_perf_1_value(lsDq_io_perf_1_value),
    .io_perf_2_value(lsDq_io_perf_2_value),
    .io_perf_3_value(lsDq_io_perf_3_value),
    .io_perf_4_value(lsDq_io_perf_4_value),
    .io_perf_5_value(lsDq_io_perf_5_value),
    .io_perf_6_value(lsDq_io_perf_6_value),
    .io_perf_7_value(lsDq_io_perf_7_value)
  );
  RedirectGenerator redirectGen ( // @[CtrlBlock.scala 273:27]
    .clock(redirectGen_clock),
    .reset(redirectGen_reset),
    .io_exuMispredict_0_valid(redirectGen_io_exuMispredict_0_valid),
    .io_exuMispredict_0_bits_uop_cf_pd_isRVC(redirectGen_io_exuMispredict_0_bits_uop_cf_pd_isRVC),
    .io_exuMispredict_0_bits_uop_cf_pd_brType(redirectGen_io_exuMispredict_0_bits_uop_cf_pd_brType),
    .io_exuMispredict_0_bits_uop_cf_pd_isCall(redirectGen_io_exuMispredict_0_bits_uop_cf_pd_isCall),
    .io_exuMispredict_0_bits_uop_cf_pd_isRet(redirectGen_io_exuMispredict_0_bits_uop_cf_pd_isRet),
    .io_exuMispredict_0_bits_uop_ctrl_imm(redirectGen_io_exuMispredict_0_bits_uop_ctrl_imm),
    .io_exuMispredict_0_bits_redirect_robIdx_flag(redirectGen_io_exuMispredict_0_bits_redirect_robIdx_flag),
    .io_exuMispredict_0_bits_redirect_robIdx_value(redirectGen_io_exuMispredict_0_bits_redirect_robIdx_value),
    .io_exuMispredict_0_bits_redirect_ftqIdx_flag(redirectGen_io_exuMispredict_0_bits_redirect_ftqIdx_flag),
    .io_exuMispredict_0_bits_redirect_ftqIdx_value(redirectGen_io_exuMispredict_0_bits_redirect_ftqIdx_value),
    .io_exuMispredict_0_bits_redirect_ftqOffset(redirectGen_io_exuMispredict_0_bits_redirect_ftqOffset),
    .io_exuMispredict_0_bits_redirect_cfiUpdate_target(redirectGen_io_exuMispredict_0_bits_redirect_cfiUpdate_target),
    .io_exuMispredict_0_bits_redirect_cfiUpdate_isMisPred(
      redirectGen_io_exuMispredict_0_bits_redirect_cfiUpdate_isMisPred),
    .io_exuMispredict_1_valid(redirectGen_io_exuMispredict_1_valid),
    .io_exuMispredict_1_bits_uop_cf_pd_isRVC(redirectGen_io_exuMispredict_1_bits_uop_cf_pd_isRVC),
    .io_exuMispredict_1_bits_uop_cf_pd_brType(redirectGen_io_exuMispredict_1_bits_uop_cf_pd_brType),
    .io_exuMispredict_1_bits_uop_cf_pd_isCall(redirectGen_io_exuMispredict_1_bits_uop_cf_pd_isCall),
    .io_exuMispredict_1_bits_uop_cf_pd_isRet(redirectGen_io_exuMispredict_1_bits_uop_cf_pd_isRet),
    .io_exuMispredict_1_bits_uop_ctrl_imm(redirectGen_io_exuMispredict_1_bits_uop_ctrl_imm),
    .io_exuMispredict_1_bits_redirect_robIdx_flag(redirectGen_io_exuMispredict_1_bits_redirect_robIdx_flag),
    .io_exuMispredict_1_bits_redirect_robIdx_value(redirectGen_io_exuMispredict_1_bits_redirect_robIdx_value),
    .io_exuMispredict_1_bits_redirect_ftqIdx_flag(redirectGen_io_exuMispredict_1_bits_redirect_ftqIdx_flag),
    .io_exuMispredict_1_bits_redirect_ftqIdx_value(redirectGen_io_exuMispredict_1_bits_redirect_ftqIdx_value),
    .io_exuMispredict_1_bits_redirect_ftqOffset(redirectGen_io_exuMispredict_1_bits_redirect_ftqOffset),
    .io_exuMispredict_1_bits_redirect_cfiUpdate_taken(redirectGen_io_exuMispredict_1_bits_redirect_cfiUpdate_taken),
    .io_exuMispredict_1_bits_redirect_cfiUpdate_isMisPred(
      redirectGen_io_exuMispredict_1_bits_redirect_cfiUpdate_isMisPred),
    .io_exuMispredict_2_valid(redirectGen_io_exuMispredict_2_valid),
    .io_exuMispredict_2_bits_uop_cf_pd_isRVC(redirectGen_io_exuMispredict_2_bits_uop_cf_pd_isRVC),
    .io_exuMispredict_2_bits_uop_cf_pd_brType(redirectGen_io_exuMispredict_2_bits_uop_cf_pd_brType),
    .io_exuMispredict_2_bits_uop_cf_pd_isCall(redirectGen_io_exuMispredict_2_bits_uop_cf_pd_isCall),
    .io_exuMispredict_2_bits_uop_cf_pd_isRet(redirectGen_io_exuMispredict_2_bits_uop_cf_pd_isRet),
    .io_exuMispredict_2_bits_uop_ctrl_imm(redirectGen_io_exuMispredict_2_bits_uop_ctrl_imm),
    .io_exuMispredict_2_bits_redirect_robIdx_flag(redirectGen_io_exuMispredict_2_bits_redirect_robIdx_flag),
    .io_exuMispredict_2_bits_redirect_robIdx_value(redirectGen_io_exuMispredict_2_bits_redirect_robIdx_value),
    .io_exuMispredict_2_bits_redirect_ftqIdx_flag(redirectGen_io_exuMispredict_2_bits_redirect_ftqIdx_flag),
    .io_exuMispredict_2_bits_redirect_ftqIdx_value(redirectGen_io_exuMispredict_2_bits_redirect_ftqIdx_value),
    .io_exuMispredict_2_bits_redirect_ftqOffset(redirectGen_io_exuMispredict_2_bits_redirect_ftqOffset),
    .io_exuMispredict_2_bits_redirect_cfiUpdate_taken(redirectGen_io_exuMispredict_2_bits_redirect_cfiUpdate_taken),
    .io_exuMispredict_2_bits_redirect_cfiUpdate_isMisPred(
      redirectGen_io_exuMispredict_2_bits_redirect_cfiUpdate_isMisPred),
    .io_loadReplay_valid(redirectGen_io_loadReplay_valid),
    .io_loadReplay_bits_robIdx_flag(redirectGen_io_loadReplay_bits_robIdx_flag),
    .io_loadReplay_bits_robIdx_value(redirectGen_io_loadReplay_bits_robIdx_value),
    .io_loadReplay_bits_ftqIdx_flag(redirectGen_io_loadReplay_bits_ftqIdx_flag),
    .io_loadReplay_bits_ftqIdx_value(redirectGen_io_loadReplay_bits_ftqIdx_value),
    .io_loadReplay_bits_ftqOffset(redirectGen_io_loadReplay_bits_ftqOffset),
    .io_loadReplay_bits_stFtqIdx_value(redirectGen_io_loadReplay_bits_stFtqIdx_value),
    .io_loadReplay_bits_stFtqOffset(redirectGen_io_loadReplay_bits_stFtqOffset),
    .io_flush(redirectGen_io_flush),
    .io_redirectPcRead_ptr_value(redirectGen_io_redirectPcRead_ptr_value),
    .io_redirectPcRead_offset(redirectGen_io_redirectPcRead_offset),
    .io_redirectPcRead_data(redirectGen_io_redirectPcRead_data),
    .io_stage2Redirect_valid(redirectGen_io_stage2Redirect_valid),
    .io_stage2Redirect_bits_robIdx_flag(redirectGen_io_stage2Redirect_bits_robIdx_flag),
    .io_stage2Redirect_bits_robIdx_value(redirectGen_io_stage2Redirect_bits_robIdx_value),
    .io_stage2Redirect_bits_ftqIdx_flag(redirectGen_io_stage2Redirect_bits_ftqIdx_flag),
    .io_stage2Redirect_bits_ftqIdx_value(redirectGen_io_stage2Redirect_bits_ftqIdx_value),
    .io_stage2Redirect_bits_ftqOffset(redirectGen_io_stage2Redirect_bits_ftqOffset),
    .io_stage2Redirect_bits_level(redirectGen_io_stage2Redirect_bits_level),
    .io_stage2Redirect_bits_cfiUpdate_pc(redirectGen_io_stage2Redirect_bits_cfiUpdate_pc),
    .io_stage2Redirect_bits_cfiUpdate_pd_isRVC(redirectGen_io_stage2Redirect_bits_cfiUpdate_pd_isRVC),
    .io_stage2Redirect_bits_cfiUpdate_pd_brType(redirectGen_io_stage2Redirect_bits_cfiUpdate_pd_brType),
    .io_stage2Redirect_bits_cfiUpdate_pd_isCall(redirectGen_io_stage2Redirect_bits_cfiUpdate_pd_isCall),
    .io_stage2Redirect_bits_cfiUpdate_pd_isRet(redirectGen_io_stage2Redirect_bits_cfiUpdate_pd_isRet),
    .io_stage2Redirect_bits_cfiUpdate_target(redirectGen_io_stage2Redirect_bits_cfiUpdate_target),
    .io_stage2Redirect_bits_cfiUpdate_taken(redirectGen_io_stage2Redirect_bits_cfiUpdate_taken),
    .io_stage2Redirect_bits_cfiUpdate_isMisPred(redirectGen_io_stage2Redirect_bits_cfiUpdate_isMisPred),
    .io_memPredUpdate_valid(redirectGen_io_memPredUpdate_valid),
    .io_memPredUpdate_ldpc(redirectGen_io_memPredUpdate_ldpc),
    .io_memPredUpdate_stpc(redirectGen_io_memPredUpdate_stpc),
    .io_memPredPcRead_ptr_value(redirectGen_io_memPredPcRead_ptr_value),
    .io_memPredPcRead_offset(redirectGen_io_memPredPcRead_offset),
    .io_memPredPcRead_data(redirectGen_io_memPredPcRead_data)
  );
  SyncDataModuleTemplate_CtrlPcMem_8entry pcMem ( // @[CtrlBlock.scala 283:21]
    .clock(pcMem_clock),
    .io_raddr_0(pcMem_io_raddr_0),
    .io_raddr_2(pcMem_io_raddr_2),
    .io_raddr_3(pcMem_io_raddr_3),
    .io_raddr_4(pcMem_io_raddr_4),
    .io_raddr_7(pcMem_io_raddr_7),
    .io_rdata_0_startAddr(pcMem_io_rdata_0_startAddr),
    .io_rdata_0_nextLineAddr(pcMem_io_rdata_0_nextLineAddr),
    .io_rdata_0_isNextMask_0(pcMem_io_rdata_0_isNextMask_0),
    .io_rdata_0_isNextMask_1(pcMem_io_rdata_0_isNextMask_1),
    .io_rdata_0_isNextMask_2(pcMem_io_rdata_0_isNextMask_2),
    .io_rdata_0_isNextMask_3(pcMem_io_rdata_0_isNextMask_3),
    .io_rdata_0_isNextMask_4(pcMem_io_rdata_0_isNextMask_4),
    .io_rdata_0_isNextMask_5(pcMem_io_rdata_0_isNextMask_5),
    .io_rdata_0_isNextMask_6(pcMem_io_rdata_0_isNextMask_6),
    .io_rdata_0_isNextMask_7(pcMem_io_rdata_0_isNextMask_7),
    .io_rdata_2_startAddr(pcMem_io_rdata_2_startAddr),
    .io_rdata_2_nextLineAddr(pcMem_io_rdata_2_nextLineAddr),
    .io_rdata_2_isNextMask_0(pcMem_io_rdata_2_isNextMask_0),
    .io_rdata_2_isNextMask_1(pcMem_io_rdata_2_isNextMask_1),
    .io_rdata_2_isNextMask_2(pcMem_io_rdata_2_isNextMask_2),
    .io_rdata_2_isNextMask_3(pcMem_io_rdata_2_isNextMask_3),
    .io_rdata_2_isNextMask_4(pcMem_io_rdata_2_isNextMask_4),
    .io_rdata_2_isNextMask_5(pcMem_io_rdata_2_isNextMask_5),
    .io_rdata_2_isNextMask_6(pcMem_io_rdata_2_isNextMask_6),
    .io_rdata_2_isNextMask_7(pcMem_io_rdata_2_isNextMask_7),
    .io_rdata_3_startAddr(pcMem_io_rdata_3_startAddr),
    .io_rdata_3_nextLineAddr(pcMem_io_rdata_3_nextLineAddr),
    .io_rdata_3_isNextMask_0(pcMem_io_rdata_3_isNextMask_0),
    .io_rdata_3_isNextMask_1(pcMem_io_rdata_3_isNextMask_1),
    .io_rdata_3_isNextMask_2(pcMem_io_rdata_3_isNextMask_2),
    .io_rdata_3_isNextMask_3(pcMem_io_rdata_3_isNextMask_3),
    .io_rdata_3_isNextMask_4(pcMem_io_rdata_3_isNextMask_4),
    .io_rdata_3_isNextMask_5(pcMem_io_rdata_3_isNextMask_5),
    .io_rdata_3_isNextMask_6(pcMem_io_rdata_3_isNextMask_6),
    .io_rdata_3_isNextMask_7(pcMem_io_rdata_3_isNextMask_7),
    .io_rdata_4_startAddr(pcMem_io_rdata_4_startAddr),
    .io_rdata_7_startAddr(pcMem_io_rdata_7_startAddr),
    .io_rdata_7_nextLineAddr(pcMem_io_rdata_7_nextLineAddr),
    .io_rdata_7_isNextMask_0(pcMem_io_rdata_7_isNextMask_0),
    .io_rdata_7_isNextMask_1(pcMem_io_rdata_7_isNextMask_1),
    .io_rdata_7_isNextMask_2(pcMem_io_rdata_7_isNextMask_2),
    .io_rdata_7_isNextMask_3(pcMem_io_rdata_7_isNextMask_3),
    .io_rdata_7_isNextMask_4(pcMem_io_rdata_7_isNextMask_4),
    .io_rdata_7_isNextMask_5(pcMem_io_rdata_7_isNextMask_5),
    .io_rdata_7_isNextMask_6(pcMem_io_rdata_7_isNextMask_6),
    .io_rdata_7_isNextMask_7(pcMem_io_rdata_7_isNextMask_7),
    .io_wen_0(pcMem_io_wen_0),
    .io_waddr_0(pcMem_io_waddr_0),
    .io_wdata_0_startAddr(pcMem_io_wdata_0_startAddr),
    .io_wdata_0_nextLineAddr(pcMem_io_wdata_0_nextLineAddr),
    .io_wdata_0_isNextMask_0(pcMem_io_wdata_0_isNextMask_0),
    .io_wdata_0_isNextMask_1(pcMem_io_wdata_0_isNextMask_1),
    .io_wdata_0_isNextMask_2(pcMem_io_wdata_0_isNextMask_2),
    .io_wdata_0_isNextMask_3(pcMem_io_wdata_0_isNextMask_3),
    .io_wdata_0_isNextMask_4(pcMem_io_wdata_0_isNextMask_4),
    .io_wdata_0_isNextMask_5(pcMem_io_wdata_0_isNextMask_5),
    .io_wdata_0_isNextMask_6(pcMem_io_wdata_0_isNextMask_6),
    .io_wdata_0_isNextMask_7(pcMem_io_wdata_0_isNextMask_7)
  );
  DelayN_26 frontendFlushValid_delay ( // @[Hold.scala 97:23]
    .clock(frontendFlushValid_delay_clock),
    .io_in(frontendFlushValid_delay_io_in),
    .io_out(frontendFlushValid_delay_io_out)
  );
  DelayN_248 pc_from_csr_delay ( // @[Hold.scala 97:23]
    .clock(pc_from_csr_delay_clock),
    .io_in(pc_from_csr_delay_io_in),
    .io_out(pc_from_csr_delay_io_out)
  );
  LFST lfst ( // @[CtrlBlock.scala 425:20]
    .clock(lfst_clock),
    .reset(lfst_reset),
    .io_redirect_valid(lfst_io_redirect_valid),
    .io_redirect_bits_robIdx_flag(lfst_io_redirect_bits_robIdx_flag),
    .io_redirect_bits_robIdx_value(lfst_io_redirect_bits_robIdx_value),
    .io_redirect_bits_level(lfst_io_redirect_bits_level),
    .io_dispatch_req_0_valid(lfst_io_dispatch_req_0_valid),
    .io_dispatch_req_0_bits_isstore(lfst_io_dispatch_req_0_bits_isstore),
    .io_dispatch_req_0_bits_ssid(lfst_io_dispatch_req_0_bits_ssid),
    .io_dispatch_req_0_bits_robIdx_flag(lfst_io_dispatch_req_0_bits_robIdx_flag),
    .io_dispatch_req_0_bits_robIdx_value(lfst_io_dispatch_req_0_bits_robIdx_value),
    .io_dispatch_req_1_valid(lfst_io_dispatch_req_1_valid),
    .io_dispatch_req_1_bits_isstore(lfst_io_dispatch_req_1_bits_isstore),
    .io_dispatch_req_1_bits_ssid(lfst_io_dispatch_req_1_bits_ssid),
    .io_dispatch_req_1_bits_robIdx_flag(lfst_io_dispatch_req_1_bits_robIdx_flag),
    .io_dispatch_req_1_bits_robIdx_value(lfst_io_dispatch_req_1_bits_robIdx_value),
    .io_dispatch_resp_0_bits_shouldWait(lfst_io_dispatch_resp_0_bits_shouldWait),
    .io_dispatch_resp_0_bits_robIdx_flag(lfst_io_dispatch_resp_0_bits_robIdx_flag),
    .io_dispatch_resp_0_bits_robIdx_value(lfst_io_dispatch_resp_0_bits_robIdx_value),
    .io_dispatch_resp_1_bits_shouldWait(lfst_io_dispatch_resp_1_bits_shouldWait),
    .io_dispatch_resp_1_bits_robIdx_flag(lfst_io_dispatch_resp_1_bits_robIdx_flag),
    .io_dispatch_resp_1_bits_robIdx_value(lfst_io_dispatch_resp_1_bits_robIdx_value),
    .io_storeIssue_0_valid(lfst_io_storeIssue_0_valid),
    .io_storeIssue_0_bits_uop_cf_storeSetHit(lfst_io_storeIssue_0_bits_uop_cf_storeSetHit),
    .io_storeIssue_0_bits_uop_cf_ssid(lfst_io_storeIssue_0_bits_uop_cf_ssid),
    .io_storeIssue_0_bits_uop_robIdx_value(lfst_io_storeIssue_0_bits_uop_robIdx_value),
    .io_storeIssue_1_valid(lfst_io_storeIssue_1_valid),
    .io_storeIssue_1_bits_uop_cf_storeSetHit(lfst_io_storeIssue_1_bits_uop_cf_storeSetHit),
    .io_storeIssue_1_bits_uop_cf_ssid(lfst_io_storeIssue_1_bits_uop_cf_ssid),
    .io_storeIssue_1_bits_uop_robIdx_value(lfst_io_storeIssue_1_bits_uop_robIdx_value),
    .io_csrCtrl_lvpred_disable(lfst_io_csrCtrl_lvpred_disable),
    .io_csrCtrl_no_spec_load(lfst_io_csrCtrl_no_spec_load),
    .io_csrCtrl_storeset_wait_store(lfst_io_csrCtrl_storeset_wait_store)
  );
  LsqEnqCtrl lsqCtrl ( // @[CtrlBlock.scala 519:27]
    .clock(lsqCtrl_clock),
    .reset(lsqCtrl_reset),
    .io_redirect_valid(lsqCtrl_io_redirect_valid),
    .io_enq_canAccept(lsqCtrl_io_enq_canAccept),
    .io_enq_needAlloc_0(lsqCtrl_io_enq_needAlloc_0),
    .io_enq_needAlloc_1(lsqCtrl_io_enq_needAlloc_1),
    .io_enq_needAlloc_2(lsqCtrl_io_enq_needAlloc_2),
    .io_enq_needAlloc_3(lsqCtrl_io_enq_needAlloc_3),
    .io_enq_req_0_valid(lsqCtrl_io_enq_req_0_valid),
    .io_enq_req_0_bits_cf_trigger_backendEn_0(lsqCtrl_io_enq_req_0_bits_cf_trigger_backendEn_0),
    .io_enq_req_0_bits_cf_trigger_backendEn_1(lsqCtrl_io_enq_req_0_bits_cf_trigger_backendEn_1),
    .io_enq_req_0_bits_ctrl_fuOpType(lsqCtrl_io_enq_req_0_bits_ctrl_fuOpType),
    .io_enq_req_0_bits_ctrl_rfWen(lsqCtrl_io_enq_req_0_bits_ctrl_rfWen),
    .io_enq_req_0_bits_ctrl_fpWen(lsqCtrl_io_enq_req_0_bits_ctrl_fpWen),
    .io_enq_req_0_bits_ctrl_flushPipe(lsqCtrl_io_enq_req_0_bits_ctrl_flushPipe),
    .io_enq_req_0_bits_ctrl_replayInst(lsqCtrl_io_enq_req_0_bits_ctrl_replayInst),
    .io_enq_req_0_bits_pdest(lsqCtrl_io_enq_req_0_bits_pdest),
    .io_enq_req_0_bits_robIdx_flag(lsqCtrl_io_enq_req_0_bits_robIdx_flag),
    .io_enq_req_0_bits_robIdx_value(lsqCtrl_io_enq_req_0_bits_robIdx_value),
    .io_enq_req_1_valid(lsqCtrl_io_enq_req_1_valid),
    .io_enq_req_1_bits_cf_trigger_backendEn_0(lsqCtrl_io_enq_req_1_bits_cf_trigger_backendEn_0),
    .io_enq_req_1_bits_cf_trigger_backendEn_1(lsqCtrl_io_enq_req_1_bits_cf_trigger_backendEn_1),
    .io_enq_req_1_bits_ctrl_fuOpType(lsqCtrl_io_enq_req_1_bits_ctrl_fuOpType),
    .io_enq_req_1_bits_ctrl_rfWen(lsqCtrl_io_enq_req_1_bits_ctrl_rfWen),
    .io_enq_req_1_bits_ctrl_fpWen(lsqCtrl_io_enq_req_1_bits_ctrl_fpWen),
    .io_enq_req_1_bits_ctrl_flushPipe(lsqCtrl_io_enq_req_1_bits_ctrl_flushPipe),
    .io_enq_req_1_bits_ctrl_replayInst(lsqCtrl_io_enq_req_1_bits_ctrl_replayInst),
    .io_enq_req_1_bits_pdest(lsqCtrl_io_enq_req_1_bits_pdest),
    .io_enq_req_1_bits_robIdx_flag(lsqCtrl_io_enq_req_1_bits_robIdx_flag),
    .io_enq_req_1_bits_robIdx_value(lsqCtrl_io_enq_req_1_bits_robIdx_value),
    .io_enq_req_2_valid(lsqCtrl_io_enq_req_2_valid),
    .io_enq_req_2_bits_cf_trigger_backendEn_0(lsqCtrl_io_enq_req_2_bits_cf_trigger_backendEn_0),
    .io_enq_req_2_bits_cf_trigger_backendEn_1(lsqCtrl_io_enq_req_2_bits_cf_trigger_backendEn_1),
    .io_enq_req_2_bits_ctrl_fuOpType(lsqCtrl_io_enq_req_2_bits_ctrl_fuOpType),
    .io_enq_req_2_bits_ctrl_rfWen(lsqCtrl_io_enq_req_2_bits_ctrl_rfWen),
    .io_enq_req_2_bits_ctrl_fpWen(lsqCtrl_io_enq_req_2_bits_ctrl_fpWen),
    .io_enq_req_2_bits_ctrl_flushPipe(lsqCtrl_io_enq_req_2_bits_ctrl_flushPipe),
    .io_enq_req_2_bits_ctrl_replayInst(lsqCtrl_io_enq_req_2_bits_ctrl_replayInst),
    .io_enq_req_2_bits_pdest(lsqCtrl_io_enq_req_2_bits_pdest),
    .io_enq_req_2_bits_robIdx_flag(lsqCtrl_io_enq_req_2_bits_robIdx_flag),
    .io_enq_req_2_bits_robIdx_value(lsqCtrl_io_enq_req_2_bits_robIdx_value),
    .io_enq_req_3_valid(lsqCtrl_io_enq_req_3_valid),
    .io_enq_req_3_bits_cf_trigger_backendEn_0(lsqCtrl_io_enq_req_3_bits_cf_trigger_backendEn_0),
    .io_enq_req_3_bits_cf_trigger_backendEn_1(lsqCtrl_io_enq_req_3_bits_cf_trigger_backendEn_1),
    .io_enq_req_3_bits_ctrl_fuOpType(lsqCtrl_io_enq_req_3_bits_ctrl_fuOpType),
    .io_enq_req_3_bits_ctrl_rfWen(lsqCtrl_io_enq_req_3_bits_ctrl_rfWen),
    .io_enq_req_3_bits_ctrl_fpWen(lsqCtrl_io_enq_req_3_bits_ctrl_fpWen),
    .io_enq_req_3_bits_ctrl_flushPipe(lsqCtrl_io_enq_req_3_bits_ctrl_flushPipe),
    .io_enq_req_3_bits_ctrl_replayInst(lsqCtrl_io_enq_req_3_bits_ctrl_replayInst),
    .io_enq_req_3_bits_pdest(lsqCtrl_io_enq_req_3_bits_pdest),
    .io_enq_req_3_bits_robIdx_flag(lsqCtrl_io_enq_req_3_bits_robIdx_flag),
    .io_enq_req_3_bits_robIdx_value(lsqCtrl_io_enq_req_3_bits_robIdx_value),
    .io_enq_resp_0_lqIdx_flag(lsqCtrl_io_enq_resp_0_lqIdx_flag),
    .io_enq_resp_0_lqIdx_value(lsqCtrl_io_enq_resp_0_lqIdx_value),
    .io_enq_resp_0_sqIdx_flag(lsqCtrl_io_enq_resp_0_sqIdx_flag),
    .io_enq_resp_0_sqIdx_value(lsqCtrl_io_enq_resp_0_sqIdx_value),
    .io_enq_resp_1_lqIdx_flag(lsqCtrl_io_enq_resp_1_lqIdx_flag),
    .io_enq_resp_1_lqIdx_value(lsqCtrl_io_enq_resp_1_lqIdx_value),
    .io_enq_resp_1_sqIdx_flag(lsqCtrl_io_enq_resp_1_sqIdx_flag),
    .io_enq_resp_1_sqIdx_value(lsqCtrl_io_enq_resp_1_sqIdx_value),
    .io_enq_resp_2_lqIdx_flag(lsqCtrl_io_enq_resp_2_lqIdx_flag),
    .io_enq_resp_2_lqIdx_value(lsqCtrl_io_enq_resp_2_lqIdx_value),
    .io_enq_resp_2_sqIdx_flag(lsqCtrl_io_enq_resp_2_sqIdx_flag),
    .io_enq_resp_2_sqIdx_value(lsqCtrl_io_enq_resp_2_sqIdx_value),
    .io_enq_resp_3_lqIdx_flag(lsqCtrl_io_enq_resp_3_lqIdx_flag),
    .io_enq_resp_3_lqIdx_value(lsqCtrl_io_enq_resp_3_lqIdx_value),
    .io_enq_resp_3_sqIdx_flag(lsqCtrl_io_enq_resp_3_sqIdx_flag),
    .io_enq_resp_3_sqIdx_value(lsqCtrl_io_enq_resp_3_sqIdx_value),
    .io_lcommit(lsqCtrl_io_lcommit),
    .io_scommit(lsqCtrl_io_scommit),
    .io_lqCancelCnt(lsqCtrl_io_lqCancelCnt),
    .io_sqCancelCnt(lsqCtrl_io_sqCancelCnt),
    .io_enqLsq_needAlloc_0(lsqCtrl_io_enqLsq_needAlloc_0),
    .io_enqLsq_needAlloc_1(lsqCtrl_io_enqLsq_needAlloc_1),
    .io_enqLsq_needAlloc_2(lsqCtrl_io_enqLsq_needAlloc_2),
    .io_enqLsq_needAlloc_3(lsqCtrl_io_enqLsq_needAlloc_3),
    .io_enqLsq_req_0_valid(lsqCtrl_io_enqLsq_req_0_valid),
    .io_enqLsq_req_0_bits_cf_trigger_backendEn_0(lsqCtrl_io_enqLsq_req_0_bits_cf_trigger_backendEn_0),
    .io_enqLsq_req_0_bits_cf_trigger_backendEn_1(lsqCtrl_io_enqLsq_req_0_bits_cf_trigger_backendEn_1),
    .io_enqLsq_req_0_bits_ctrl_fuOpType(lsqCtrl_io_enqLsq_req_0_bits_ctrl_fuOpType),
    .io_enqLsq_req_0_bits_ctrl_rfWen(lsqCtrl_io_enqLsq_req_0_bits_ctrl_rfWen),
    .io_enqLsq_req_0_bits_ctrl_fpWen(lsqCtrl_io_enqLsq_req_0_bits_ctrl_fpWen),
    .io_enqLsq_req_0_bits_ctrl_flushPipe(lsqCtrl_io_enqLsq_req_0_bits_ctrl_flushPipe),
    .io_enqLsq_req_0_bits_ctrl_replayInst(lsqCtrl_io_enqLsq_req_0_bits_ctrl_replayInst),
    .io_enqLsq_req_0_bits_pdest(lsqCtrl_io_enqLsq_req_0_bits_pdest),
    .io_enqLsq_req_0_bits_robIdx_flag(lsqCtrl_io_enqLsq_req_0_bits_robIdx_flag),
    .io_enqLsq_req_0_bits_robIdx_value(lsqCtrl_io_enqLsq_req_0_bits_robIdx_value),
    .io_enqLsq_req_0_bits_lqIdx_value(lsqCtrl_io_enqLsq_req_0_bits_lqIdx_value),
    .io_enqLsq_req_0_bits_sqIdx_value(lsqCtrl_io_enqLsq_req_0_bits_sqIdx_value),
    .io_enqLsq_req_1_valid(lsqCtrl_io_enqLsq_req_1_valid),
    .io_enqLsq_req_1_bits_cf_trigger_backendEn_0(lsqCtrl_io_enqLsq_req_1_bits_cf_trigger_backendEn_0),
    .io_enqLsq_req_1_bits_cf_trigger_backendEn_1(lsqCtrl_io_enqLsq_req_1_bits_cf_trigger_backendEn_1),
    .io_enqLsq_req_1_bits_ctrl_fuOpType(lsqCtrl_io_enqLsq_req_1_bits_ctrl_fuOpType),
    .io_enqLsq_req_1_bits_ctrl_rfWen(lsqCtrl_io_enqLsq_req_1_bits_ctrl_rfWen),
    .io_enqLsq_req_1_bits_ctrl_fpWen(lsqCtrl_io_enqLsq_req_1_bits_ctrl_fpWen),
    .io_enqLsq_req_1_bits_ctrl_flushPipe(lsqCtrl_io_enqLsq_req_1_bits_ctrl_flushPipe),
    .io_enqLsq_req_1_bits_ctrl_replayInst(lsqCtrl_io_enqLsq_req_1_bits_ctrl_replayInst),
    .io_enqLsq_req_1_bits_pdest(lsqCtrl_io_enqLsq_req_1_bits_pdest),
    .io_enqLsq_req_1_bits_robIdx_flag(lsqCtrl_io_enqLsq_req_1_bits_robIdx_flag),
    .io_enqLsq_req_1_bits_robIdx_value(lsqCtrl_io_enqLsq_req_1_bits_robIdx_value),
    .io_enqLsq_req_1_bits_lqIdx_value(lsqCtrl_io_enqLsq_req_1_bits_lqIdx_value),
    .io_enqLsq_req_1_bits_sqIdx_value(lsqCtrl_io_enqLsq_req_1_bits_sqIdx_value),
    .io_enqLsq_req_2_valid(lsqCtrl_io_enqLsq_req_2_valid),
    .io_enqLsq_req_2_bits_cf_trigger_backendEn_0(lsqCtrl_io_enqLsq_req_2_bits_cf_trigger_backendEn_0),
    .io_enqLsq_req_2_bits_cf_trigger_backendEn_1(lsqCtrl_io_enqLsq_req_2_bits_cf_trigger_backendEn_1),
    .io_enqLsq_req_2_bits_ctrl_fuOpType(lsqCtrl_io_enqLsq_req_2_bits_ctrl_fuOpType),
    .io_enqLsq_req_2_bits_ctrl_rfWen(lsqCtrl_io_enqLsq_req_2_bits_ctrl_rfWen),
    .io_enqLsq_req_2_bits_ctrl_fpWen(lsqCtrl_io_enqLsq_req_2_bits_ctrl_fpWen),
    .io_enqLsq_req_2_bits_ctrl_flushPipe(lsqCtrl_io_enqLsq_req_2_bits_ctrl_flushPipe),
    .io_enqLsq_req_2_bits_ctrl_replayInst(lsqCtrl_io_enqLsq_req_2_bits_ctrl_replayInst),
    .io_enqLsq_req_2_bits_pdest(lsqCtrl_io_enqLsq_req_2_bits_pdest),
    .io_enqLsq_req_2_bits_robIdx_flag(lsqCtrl_io_enqLsq_req_2_bits_robIdx_flag),
    .io_enqLsq_req_2_bits_robIdx_value(lsqCtrl_io_enqLsq_req_2_bits_robIdx_value),
    .io_enqLsq_req_2_bits_lqIdx_value(lsqCtrl_io_enqLsq_req_2_bits_lqIdx_value),
    .io_enqLsq_req_2_bits_sqIdx_value(lsqCtrl_io_enqLsq_req_2_bits_sqIdx_value),
    .io_enqLsq_req_3_valid(lsqCtrl_io_enqLsq_req_3_valid),
    .io_enqLsq_req_3_bits_cf_trigger_backendEn_0(lsqCtrl_io_enqLsq_req_3_bits_cf_trigger_backendEn_0),
    .io_enqLsq_req_3_bits_cf_trigger_backendEn_1(lsqCtrl_io_enqLsq_req_3_bits_cf_trigger_backendEn_1),
    .io_enqLsq_req_3_bits_ctrl_fuOpType(lsqCtrl_io_enqLsq_req_3_bits_ctrl_fuOpType),
    .io_enqLsq_req_3_bits_ctrl_rfWen(lsqCtrl_io_enqLsq_req_3_bits_ctrl_rfWen),
    .io_enqLsq_req_3_bits_ctrl_fpWen(lsqCtrl_io_enqLsq_req_3_bits_ctrl_fpWen),
    .io_enqLsq_req_3_bits_ctrl_flushPipe(lsqCtrl_io_enqLsq_req_3_bits_ctrl_flushPipe),
    .io_enqLsq_req_3_bits_ctrl_replayInst(lsqCtrl_io_enqLsq_req_3_bits_ctrl_replayInst),
    .io_enqLsq_req_3_bits_pdest(lsqCtrl_io_enqLsq_req_3_bits_pdest),
    .io_enqLsq_req_3_bits_robIdx_flag(lsqCtrl_io_enqLsq_req_3_bits_robIdx_flag),
    .io_enqLsq_req_3_bits_robIdx_value(lsqCtrl_io_enqLsq_req_3_bits_robIdx_value),
    .io_enqLsq_req_3_bits_lqIdx_value(lsqCtrl_io_enqLsq_req_3_bits_lqIdx_value),
    .io_enqLsq_req_3_bits_sqIdx_value(lsqCtrl_io_enqLsq_req_3_bits_sqIdx_value)
  );
  DelayN_26 io_cpu_halt_delay ( // @[Hold.scala 97:23]
    .clock(io_cpu_halt_delay_clock),
    .io_in(io_cpu_halt_delay_io_in),
    .io_out(io_cpu_halt_delay_io_out)
  );
  PFEvent pfevent ( // @[CtrlBlock.scala 585:23]
    .clock(pfevent_clock),
    .reset(pfevent_reset),
    .io_distribute_csr_wvalid(pfevent_io_distribute_csr_wvalid),
    .io_distribute_csr_waddr(pfevent_io_distribute_csr_waddr),
    .io_distribute_csr_wdata(pfevent_io_distribute_csr_wdata),
    .io_hpmevent_0(pfevent_io_hpmevent_0),
    .io_hpmevent_1(pfevent_io_hpmevent_1),
    .io_hpmevent_2(pfevent_io_hpmevent_2),
    .io_hpmevent_3(pfevent_io_hpmevent_3),
    .io_hpmevent_4(pfevent_io_hpmevent_4),
    .io_hpmevent_5(pfevent_io_hpmevent_5),
    .io_hpmevent_6(pfevent_io_hpmevent_6),
    .io_hpmevent_7(pfevent_io_hpmevent_7),
    .io_hpmevent_8(pfevent_io_hpmevent_8),
    .io_hpmevent_9(pfevent_io_hpmevent_9),
    .io_hpmevent_10(pfevent_io_hpmevent_10),
    .io_hpmevent_11(pfevent_io_hpmevent_11),
    .io_hpmevent_12(pfevent_io_hpmevent_12),
    .io_hpmevent_13(pfevent_io_hpmevent_13),
    .io_hpmevent_14(pfevent_io_hpmevent_14),
    .io_hpmevent_15(pfevent_io_hpmevent_15),
    .io_hpmevent_16(pfevent_io_hpmevent_16),
    .io_hpmevent_17(pfevent_io_hpmevent_17),
    .io_hpmevent_18(pfevent_io_hpmevent_18),
    .io_hpmevent_19(pfevent_io_hpmevent_19),
    .io_hpmevent_20(pfevent_io_hpmevent_20),
    .io_hpmevent_21(pfevent_io_hpmevent_21),
    .io_hpmevent_22(pfevent_io_hpmevent_22),
    .io_hpmevent_23(pfevent_io_hpmevent_23)
  );
  HPerfMonitor_3 hpm ( // @[PerfCounterUtils.scala 255:21]
    .clock(hpm_clock),
    .io_hpm_event_0(hpm_io_hpm_event_0),
    .io_hpm_event_1(hpm_io_hpm_event_1),
    .io_hpm_event_2(hpm_io_hpm_event_2),
    .io_hpm_event_3(hpm_io_hpm_event_3),
    .io_hpm_event_4(hpm_io_hpm_event_4),
    .io_hpm_event_5(hpm_io_hpm_event_5),
    .io_hpm_event_6(hpm_io_hpm_event_6),
    .io_hpm_event_7(hpm_io_hpm_event_7),
    .io_events_sets_0_value(hpm_io_events_sets_0_value),
    .io_events_sets_1_value(hpm_io_events_sets_1_value),
    .io_events_sets_2_value(hpm_io_events_sets_2_value),
    .io_events_sets_3_value(hpm_io_events_sets_3_value),
    .io_events_sets_4_value(hpm_io_events_sets_4_value),
    .io_events_sets_5_value(hpm_io_events_sets_5_value),
    .io_events_sets_6_value(hpm_io_events_sets_6_value),
    .io_events_sets_7_value(hpm_io_events_sets_7_value),
    .io_events_sets_8_value(hpm_io_events_sets_8_value),
    .io_events_sets_9_value(hpm_io_events_sets_9_value),
    .io_events_sets_10_value(hpm_io_events_sets_10_value),
    .io_events_sets_11_value(hpm_io_events_sets_11_value),
    .io_events_sets_12_value(hpm_io_events_sets_12_value),
    .io_events_sets_13_value(hpm_io_events_sets_13_value),
    .io_events_sets_14_value(hpm_io_events_sets_14_value),
    .io_events_sets_15_value(hpm_io_events_sets_15_value),
    .io_events_sets_16_value(hpm_io_events_sets_16_value),
    .io_events_sets_17_value(hpm_io_events_sets_17_value),
    .io_events_sets_18_value(hpm_io_events_sets_18_value),
    .io_events_sets_19_value(hpm_io_events_sets_19_value),
    .io_events_sets_20_value(hpm_io_events_sets_20_value),
    .io_events_sets_21_value(hpm_io_events_sets_21_value),
    .io_events_sets_23_value(hpm_io_events_sets_23_value),
    .io_events_sets_24_value(hpm_io_events_sets_24_value),
    .io_events_sets_25_value(hpm_io_events_sets_25_value),
    .io_events_sets_26_value(hpm_io_events_sets_26_value),
    .io_events_sets_27_value(hpm_io_events_sets_27_value),
    .io_events_sets_28_value(hpm_io_events_sets_28_value),
    .io_events_sets_29_value(hpm_io_events_sets_29_value),
    .io_events_sets_30_value(hpm_io_events_sets_30_value),
    .io_events_sets_31_value(hpm_io_events_sets_31_value),
    .io_events_sets_32_value(hpm_io_events_sets_32_value),
    .io_events_sets_33_value(hpm_io_events_sets_33_value),
    .io_events_sets_34_value(hpm_io_events_sets_34_value),
    .io_events_sets_35_value(hpm_io_events_sets_35_value),
    .io_events_sets_36_value(hpm_io_events_sets_36_value),
    .io_events_sets_37_value(hpm_io_events_sets_37_value),
    .io_events_sets_38_value(hpm_io_events_sets_38_value),
    .io_events_sets_39_value(hpm_io_events_sets_39_value),
    .io_events_sets_40_value(hpm_io_events_sets_40_value),
    .io_events_sets_41_value(hpm_io_events_sets_41_value),
    .io_events_sets_42_value(hpm_io_events_sets_42_value),
    .io_events_sets_43_value(hpm_io_events_sets_43_value),
    .io_events_sets_44_value(hpm_io_events_sets_44_value),
    .io_events_sets_45_value(hpm_io_events_sets_45_value),
    .io_events_sets_46_value(hpm_io_events_sets_46_value),
    .io_events_sets_47_value(hpm_io_events_sets_47_value),
    .io_events_sets_48_value(hpm_io_events_sets_48_value),
    .io_events_sets_49_value(hpm_io_events_sets_49_value),
    .io_events_sets_50_value(hpm_io_events_sets_50_value),
    .io_events_sets_51_value(hpm_io_events_sets_51_value),
    .io_events_sets_52_value(hpm_io_events_sets_52_value),
    .io_events_sets_53_value(hpm_io_events_sets_53_value),
    .io_events_sets_54_value(hpm_io_events_sets_54_value),
    .io_events_sets_55_value(hpm_io_events_sets_55_value),
    .io_events_sets_56_value(hpm_io_events_sets_56_value),
    .io_events_sets_57_value(hpm_io_events_sets_57_value),
    .io_events_sets_58_value(hpm_io_events_sets_58_value),
    .io_events_sets_59_value(hpm_io_events_sets_59_value),
    .io_events_sets_60_value(hpm_io_events_sets_60_value),
    .io_events_sets_61_value(hpm_io_events_sets_61_value),
    .io_events_sets_62_value(hpm_io_events_sets_62_value),
    .io_events_sets_63_value(hpm_io_events_sets_63_value),
    .io_events_sets_64_value(hpm_io_events_sets_64_value),
    .io_events_sets_65_value(hpm_io_events_sets_65_value),
    .io_events_sets_66_value(hpm_io_events_sets_66_value),
    .io_events_sets_67_value(hpm_io_events_sets_67_value),
    .io_events_sets_68_value(hpm_io_events_sets_68_value),
    .io_events_sets_69_value(hpm_io_events_sets_69_value),
    .io_events_sets_70_value(hpm_io_events_sets_70_value),
    .io_events_sets_71_value(hpm_io_events_sets_71_value),
    .io_events_sets_72_value(hpm_io_events_sets_72_value),
    .io_events_sets_73_value(hpm_io_events_sets_73_value),
    .io_events_sets_74_value(hpm_io_events_sets_74_value),
    .io_events_sets_75_value(hpm_io_events_sets_75_value),
    .io_events_sets_76_value(hpm_io_events_sets_76_value),
    .io_events_sets_77_value(hpm_io_events_sets_77_value),
    .io_events_sets_78_value(hpm_io_events_sets_78_value),
    .io_events_sets_79_value(hpm_io_events_sets_79_value),
    .io_events_sets_80_value(hpm_io_events_sets_80_value),
    .io_events_sets_81_value(hpm_io_events_sets_81_value),
    .io_events_sets_82_value(hpm_io_events_sets_82_value),
    .io_events_sets_83_value(hpm_io_events_sets_83_value),
    .io_events_sets_84_value(hpm_io_events_sets_84_value),
    .io_events_sets_85_value(hpm_io_events_sets_85_value),
    .io_events_sets_86_value(hpm_io_events_sets_86_value),
    .io_events_sets_87_value(hpm_io_events_sets_87_value),
    .io_events_sets_88_value(hpm_io_events_sets_88_value),
    .io_perf_0_value(hpm_io_perf_0_value),
    .io_perf_1_value(hpm_io_perf_1_value),
    .io_perf_2_value(hpm_io_perf_2_value),
    .io_perf_3_value(hpm_io_perf_3_value),
    .io_perf_4_value(hpm_io_perf_4_value),
    .io_perf_5_value(hpm_io_perf_5_value),
    .io_perf_6_value(hpm_io_perf_6_value),
    .io_perf_7_value(hpm_io_perf_7_value)
  );
  assign io_cpu_halt = io_cpu_halt_delay_io_out; // @[CtrlBlock.scala 560:15]
  assign io_frontend_cfVec_0_ready = decode_io_in_0_ready; // @[CtrlBlock.scala 402:16]
  assign io_frontend_cfVec_1_ready = decode_io_in_1_ready; // @[CtrlBlock.scala 402:16]
  assign io_frontend_toFtq_rob_commits_0_valid = io_frontend_toFtq_rob_commits_0_valid_REG; // @[CtrlBlock.scala 338:44]
  assign io_frontend_toFtq_rob_commits_0_bits_commitType = io_frontend_toFtq_rob_commits_0_bits_rcommitType; // @[CtrlBlock.scala 339:43]
  assign io_frontend_toFtq_rob_commits_0_bits_ftqIdx_flag = io_frontend_toFtq_rob_commits_0_bits_rftqIdx_flag; // @[CtrlBlock.scala 339:43]
  assign io_frontend_toFtq_rob_commits_0_bits_ftqIdx_value = io_frontend_toFtq_rob_commits_0_bits_rftqIdx_value; // @[CtrlBlock.scala 339:43]
  assign io_frontend_toFtq_rob_commits_0_bits_ftqOffset = io_frontend_toFtq_rob_commits_0_bits_rftqOffset; // @[CtrlBlock.scala 339:43]
  assign io_frontend_toFtq_rob_commits_1_valid = io_frontend_toFtq_rob_commits_1_valid_REG; // @[CtrlBlock.scala 338:44]
  assign io_frontend_toFtq_rob_commits_1_bits_commitType = io_frontend_toFtq_rob_commits_1_bits_rcommitType; // @[CtrlBlock.scala 339:43]
  assign io_frontend_toFtq_rob_commits_1_bits_ftqIdx_flag = io_frontend_toFtq_rob_commits_1_bits_rftqIdx_flag; // @[CtrlBlock.scala 339:43]
  assign io_frontend_toFtq_rob_commits_1_bits_ftqIdx_value = io_frontend_toFtq_rob_commits_1_bits_rftqIdx_value; // @[CtrlBlock.scala 339:43]
  assign io_frontend_toFtq_rob_commits_1_bits_ftqOffset = io_frontend_toFtq_rob_commits_1_bits_rftqOffset; // @[CtrlBlock.scala 339:43]
  assign io_frontend_toFtq_redirect_valid = frontendFlushValid_delay_io_out | redirectGen_io_stage2Redirect_valid; // @[CtrlBlock.scala 341:58]
  assign io_frontend_toFtq_redirect_bits_ftqIdx_flag = frontendFlushValid_delay_io_out ? frontendFlushBits_ftqIdx_flag
     : redirectGen_io_stage2Redirect_bits_ftqIdx_flag; // @[CtrlBlock.scala 342:41]
  assign io_frontend_toFtq_redirect_bits_ftqIdx_value = frontendFlushValid_delay_io_out ? frontendFlushBits_ftqIdx_value
     : redirectGen_io_stage2Redirect_bits_ftqIdx_value; // @[CtrlBlock.scala 342:41]
  assign io_frontend_toFtq_redirect_bits_ftqOffset = frontendFlushValid_delay_io_out ? frontendFlushBits_ftqOffset :
    redirectGen_io_stage2Redirect_bits_ftqOffset; // @[CtrlBlock.scala 342:41]
  assign io_frontend_toFtq_redirect_bits_level = frontendFlushValid_delay_io_out |
    _io_frontend_toFtq_redirect_bits_T_level; // @[CtrlBlock.scala 356:29 342:35 357:43]
  assign io_frontend_toFtq_redirect_bits_cfiUpdate_pc = frontendFlushValid_delay_io_out ? 39'h0 :
    redirectGen_io_stage2Redirect_bits_cfiUpdate_pc; // @[CtrlBlock.scala 342:41]
  assign io_frontend_toFtq_redirect_bits_cfiUpdate_pd_isRVC = frontendFlushValid_delay_io_out ? 1'h0 :
    redirectGen_io_stage2Redirect_bits_cfiUpdate_pd_isRVC; // @[CtrlBlock.scala 342:41]
  assign io_frontend_toFtq_redirect_bits_cfiUpdate_pd_brType = frontendFlushValid_delay_io_out ? 2'h0 :
    redirectGen_io_stage2Redirect_bits_cfiUpdate_pd_brType; // @[CtrlBlock.scala 342:41]
  assign io_frontend_toFtq_redirect_bits_cfiUpdate_pd_isCall = frontendFlushValid_delay_io_out ? 1'h0 :
    redirectGen_io_stage2Redirect_bits_cfiUpdate_pd_isCall; // @[CtrlBlock.scala 342:41]
  assign io_frontend_toFtq_redirect_bits_cfiUpdate_pd_isRet = frontendFlushValid_delay_io_out ? 1'h0 :
    redirectGen_io_stage2Redirect_bits_cfiUpdate_pd_isRet; // @[CtrlBlock.scala 342:41]
  assign io_frontend_toFtq_redirect_bits_cfiUpdate_target = frontendFlushValid_delay_io_out ?
    io_frontend_toFtq_redirect_bits_cfiUpdate_target_REG : _io_frontend_toFtq_redirect_bits_T_cfiUpdate_target; // @[CtrlBlock.scala 356:29 342:35 358:54]
  assign io_frontend_toFtq_redirect_bits_cfiUpdate_taken = frontendFlushValid_delay_io_out ? 1'h0 :
    redirectGen_io_stage2Redirect_bits_cfiUpdate_taken; // @[CtrlBlock.scala 342:41]
  assign io_frontend_toFtq_redirect_bits_cfiUpdate_isMisPred = frontendFlushValid_delay_io_out ? 1'h0 :
    redirectGen_io_stage2Redirect_bits_cfiUpdate_isMisPred; // @[CtrlBlock.scala 342:41]
  assign io_allocPregs_0_isInt = dispatch_io_allocPregs_0_isInt; // @[CtrlBlock.scala 500:26]
  assign io_allocPregs_0_isFp = dispatch_io_allocPregs_0_isFp; // @[CtrlBlock.scala 500:26]
  assign io_allocPregs_0_preg = dispatch_io_allocPregs_0_preg; // @[CtrlBlock.scala 500:26]
  assign io_allocPregs_1_isInt = dispatch_io_allocPregs_1_isInt; // @[CtrlBlock.scala 500:26]
  assign io_allocPregs_1_isFp = dispatch_io_allocPregs_1_isFp; // @[CtrlBlock.scala 500:26]
  assign io_allocPregs_1_preg = dispatch_io_allocPregs_1_preg; // @[CtrlBlock.scala 500:26]
  assign io_dispatch_0_valid = intDq_io_deq_0_valid; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_0_bits_cf_foldpc = intDq_io_deq_0_bits_cf_foldpc; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_0_bits_cf_trigger_backendEn_0 = intDq_io_deq_0_bits_cf_trigger_backendEn_0; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_0_bits_cf_trigger_backendEn_1 = intDq_io_deq_0_bits_cf_trigger_backendEn_1; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_0_bits_cf_pd_isRVC = intDq_io_deq_0_bits_cf_pd_isRVC; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_0_bits_cf_pd_brType = intDq_io_deq_0_bits_cf_pd_brType; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_0_bits_cf_pd_isCall = intDq_io_deq_0_bits_cf_pd_isCall; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_0_bits_cf_pd_isRet = intDq_io_deq_0_bits_cf_pd_isRet; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_0_bits_cf_pred_taken = intDq_io_deq_0_bits_cf_pred_taken; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_0_bits_cf_storeSetHit = intDq_io_deq_0_bits_cf_storeSetHit; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_0_bits_cf_waitForRobIdx_flag = intDq_io_deq_0_bits_cf_waitForRobIdx_flag; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_0_bits_cf_waitForRobIdx_value = intDq_io_deq_0_bits_cf_waitForRobIdx_value; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_0_bits_cf_loadWaitBit = intDq_io_deq_0_bits_cf_loadWaitBit; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_0_bits_cf_loadWaitStrict = intDq_io_deq_0_bits_cf_loadWaitStrict; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_0_bits_cf_ssid = intDq_io_deq_0_bits_cf_ssid; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_0_bits_cf_ftqPtr_flag = intDq_io_deq_0_bits_cf_ftqPtr_flag; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_0_bits_cf_ftqPtr_value = intDq_io_deq_0_bits_cf_ftqPtr_value; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_0_bits_cf_ftqOffset = intDq_io_deq_0_bits_cf_ftqOffset; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_0_bits_ctrl_srcType_0 = intDq_io_deq_0_bits_ctrl_srcType_0; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_0_bits_ctrl_srcType_1 = intDq_io_deq_0_bits_ctrl_srcType_1; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_0_bits_ctrl_fuType = intDq_io_deq_0_bits_ctrl_fuType; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_0_bits_ctrl_fuOpType = intDq_io_deq_0_bits_ctrl_fuOpType; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_0_bits_ctrl_rfWen = intDq_io_deq_0_bits_ctrl_rfWen; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_0_bits_ctrl_fpWen = intDq_io_deq_0_bits_ctrl_fpWen; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_0_bits_ctrl_selImm = intDq_io_deq_0_bits_ctrl_selImm; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_0_bits_ctrl_imm = intDq_io_deq_0_bits_ctrl_imm; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_0_bits_ctrl_fpu_isAddSub = intDq_io_deq_0_bits_ctrl_fpu_isAddSub; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_0_bits_ctrl_fpu_typeTagIn = intDq_io_deq_0_bits_ctrl_fpu_typeTagIn; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_0_bits_ctrl_fpu_typeTagOut = intDq_io_deq_0_bits_ctrl_fpu_typeTagOut; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_0_bits_ctrl_fpu_fromInt = intDq_io_deq_0_bits_ctrl_fpu_fromInt; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_0_bits_ctrl_fpu_wflags = intDq_io_deq_0_bits_ctrl_fpu_wflags; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_0_bits_ctrl_fpu_fpWen = intDq_io_deq_0_bits_ctrl_fpu_fpWen; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_0_bits_ctrl_fpu_fmaCmd = intDq_io_deq_0_bits_ctrl_fpu_fmaCmd; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_0_bits_ctrl_fpu_div = intDq_io_deq_0_bits_ctrl_fpu_div; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_0_bits_ctrl_fpu_sqrt = intDq_io_deq_0_bits_ctrl_fpu_sqrt; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_0_bits_ctrl_fpu_fcvt = intDq_io_deq_0_bits_ctrl_fpu_fcvt; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_0_bits_ctrl_fpu_typ = intDq_io_deq_0_bits_ctrl_fpu_typ; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_0_bits_ctrl_fpu_fmt = intDq_io_deq_0_bits_ctrl_fpu_fmt; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_0_bits_ctrl_fpu_ren3 = intDq_io_deq_0_bits_ctrl_fpu_ren3; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_0_bits_ctrl_fpu_rm = intDq_io_deq_0_bits_ctrl_fpu_rm; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_0_bits_psrc_0 = intDq_io_deq_0_bits_psrc_0; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_0_bits_psrc_1 = intDq_io_deq_0_bits_psrc_1; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_0_bits_pdest = intDq_io_deq_0_bits_pdest; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_0_bits_robIdx_flag = intDq_io_deq_0_bits_robIdx_flag; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_0_bits_robIdx_value = intDq_io_deq_0_bits_robIdx_value; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_0_bits_lqIdx_flag = intDq_io_deq_0_bits_lqIdx_flag; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_0_bits_lqIdx_value = intDq_io_deq_0_bits_lqIdx_value; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_0_bits_sqIdx_flag = intDq_io_deq_0_bits_sqIdx_flag; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_0_bits_sqIdx_value = intDq_io_deq_0_bits_sqIdx_value; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_1_valid = intDq_io_deq_1_valid; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_1_bits_cf_foldpc = intDq_io_deq_1_bits_cf_foldpc; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_1_bits_cf_trigger_backendEn_0 = intDq_io_deq_1_bits_cf_trigger_backendEn_0; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_1_bits_cf_trigger_backendEn_1 = intDq_io_deq_1_bits_cf_trigger_backendEn_1; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_1_bits_cf_pd_isRVC = intDq_io_deq_1_bits_cf_pd_isRVC; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_1_bits_cf_pd_brType = intDq_io_deq_1_bits_cf_pd_brType; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_1_bits_cf_pd_isCall = intDq_io_deq_1_bits_cf_pd_isCall; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_1_bits_cf_pd_isRet = intDq_io_deq_1_bits_cf_pd_isRet; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_1_bits_cf_pred_taken = intDq_io_deq_1_bits_cf_pred_taken; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_1_bits_cf_storeSetHit = intDq_io_deq_1_bits_cf_storeSetHit; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_1_bits_cf_waitForRobIdx_flag = intDq_io_deq_1_bits_cf_waitForRobIdx_flag; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_1_bits_cf_waitForRobIdx_value = intDq_io_deq_1_bits_cf_waitForRobIdx_value; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_1_bits_cf_loadWaitBit = intDq_io_deq_1_bits_cf_loadWaitBit; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_1_bits_cf_loadWaitStrict = intDq_io_deq_1_bits_cf_loadWaitStrict; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_1_bits_cf_ssid = intDq_io_deq_1_bits_cf_ssid; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_1_bits_cf_ftqPtr_flag = intDq_io_deq_1_bits_cf_ftqPtr_flag; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_1_bits_cf_ftqPtr_value = intDq_io_deq_1_bits_cf_ftqPtr_value; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_1_bits_cf_ftqOffset = intDq_io_deq_1_bits_cf_ftqOffset; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_1_bits_ctrl_srcType_0 = intDq_io_deq_1_bits_ctrl_srcType_0; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_1_bits_ctrl_srcType_1 = intDq_io_deq_1_bits_ctrl_srcType_1; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_1_bits_ctrl_fuType = intDq_io_deq_1_bits_ctrl_fuType; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_1_bits_ctrl_fuOpType = intDq_io_deq_1_bits_ctrl_fuOpType; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_1_bits_ctrl_rfWen = intDq_io_deq_1_bits_ctrl_rfWen; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_1_bits_ctrl_fpWen = intDq_io_deq_1_bits_ctrl_fpWen; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_1_bits_ctrl_selImm = intDq_io_deq_1_bits_ctrl_selImm; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_1_bits_ctrl_imm = intDq_io_deq_1_bits_ctrl_imm; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_1_bits_psrc_0 = intDq_io_deq_1_bits_psrc_0; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_1_bits_psrc_1 = intDq_io_deq_1_bits_psrc_1; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_1_bits_pdest = intDq_io_deq_1_bits_pdest; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_1_bits_robIdx_flag = intDq_io_deq_1_bits_robIdx_flag; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_1_bits_robIdx_value = intDq_io_deq_1_bits_robIdx_value; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_1_bits_lqIdx_flag = intDq_io_deq_1_bits_lqIdx_flag; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_1_bits_lqIdx_value = intDq_io_deq_1_bits_lqIdx_value; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_1_bits_sqIdx_flag = intDq_io_deq_1_bits_sqIdx_flag; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_1_bits_sqIdx_value = intDq_io_deq_1_bits_sqIdx_value; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_4_valid = lsDq_io_deq_0_valid; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_4_bits_cf_foldpc = lsDq_io_deq_0_bits_cf_foldpc; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_4_bits_cf_trigger_backendEn_0 = lsDq_io_deq_0_bits_cf_trigger_backendEn_0; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_4_bits_cf_trigger_backendEn_1 = lsDq_io_deq_0_bits_cf_trigger_backendEn_1; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_4_bits_cf_pd_isRVC = lsDq_io_deq_0_bits_cf_pd_isRVC; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_4_bits_cf_pd_brType = lsDq_io_deq_0_bits_cf_pd_brType; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_4_bits_cf_pd_isCall = lsDq_io_deq_0_bits_cf_pd_isCall; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_4_bits_cf_pd_isRet = lsDq_io_deq_0_bits_cf_pd_isRet; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_4_bits_cf_pred_taken = lsDq_io_deq_0_bits_cf_pred_taken; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_4_bits_cf_storeSetHit = lsDq_io_deq_0_bits_cf_storeSetHit; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_4_bits_cf_waitForRobIdx_flag = lsDq_io_deq_0_bits_cf_waitForRobIdx_flag; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_4_bits_cf_waitForRobIdx_value = lsDq_io_deq_0_bits_cf_waitForRobIdx_value; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_4_bits_cf_loadWaitBit = lsDq_io_deq_0_bits_cf_loadWaitBit; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_4_bits_cf_loadWaitStrict = lsDq_io_deq_0_bits_cf_loadWaitStrict; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_4_bits_cf_ssid = lsDq_io_deq_0_bits_cf_ssid; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_4_bits_cf_ftqPtr_flag = lsDq_io_deq_0_bits_cf_ftqPtr_flag; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_4_bits_cf_ftqPtr_value = lsDq_io_deq_0_bits_cf_ftqPtr_value; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_4_bits_cf_ftqOffset = lsDq_io_deq_0_bits_cf_ftqOffset; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_4_bits_ctrl_srcType_0 = lsDq_io_deq_0_bits_ctrl_srcType_0; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_4_bits_ctrl_srcType_1 = lsDq_io_deq_0_bits_ctrl_srcType_1; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_4_bits_ctrl_fuType = lsDq_io_deq_0_bits_ctrl_fuType; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_4_bits_ctrl_fuOpType = lsDq_io_deq_0_bits_ctrl_fuOpType; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_4_bits_ctrl_rfWen = lsDq_io_deq_0_bits_ctrl_rfWen; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_4_bits_ctrl_fpWen = lsDq_io_deq_0_bits_ctrl_fpWen; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_4_bits_ctrl_flushPipe = lsDq_io_deq_0_bits_ctrl_flushPipe; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_4_bits_ctrl_imm = lsDq_io_deq_0_bits_ctrl_imm; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_4_bits_ctrl_replayInst = lsDq_io_deq_0_bits_ctrl_replayInst; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_4_bits_psrc_0 = lsDq_io_deq_0_bits_psrc_0; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_4_bits_psrc_1 = lsDq_io_deq_0_bits_psrc_1; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_4_bits_pdest = lsDq_io_deq_0_bits_pdest; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_4_bits_robIdx_flag = lsDq_io_deq_0_bits_robIdx_flag; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_4_bits_robIdx_value = lsDq_io_deq_0_bits_robIdx_value; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_5_valid = lsDq_io_deq_1_valid; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_5_bits_cf_foldpc = lsDq_io_deq_1_bits_cf_foldpc; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_5_bits_cf_trigger_backendEn_0 = lsDq_io_deq_1_bits_cf_trigger_backendEn_0; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_5_bits_cf_trigger_backendEn_1 = lsDq_io_deq_1_bits_cf_trigger_backendEn_1; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_5_bits_cf_pd_isRVC = lsDq_io_deq_1_bits_cf_pd_isRVC; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_5_bits_cf_pd_brType = lsDq_io_deq_1_bits_cf_pd_brType; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_5_bits_cf_pd_isCall = lsDq_io_deq_1_bits_cf_pd_isCall; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_5_bits_cf_pd_isRet = lsDq_io_deq_1_bits_cf_pd_isRet; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_5_bits_cf_pred_taken = lsDq_io_deq_1_bits_cf_pred_taken; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_5_bits_cf_storeSetHit = lsDq_io_deq_1_bits_cf_storeSetHit; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_5_bits_cf_waitForRobIdx_flag = lsDq_io_deq_1_bits_cf_waitForRobIdx_flag; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_5_bits_cf_waitForRobIdx_value = lsDq_io_deq_1_bits_cf_waitForRobIdx_value; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_5_bits_cf_loadWaitBit = lsDq_io_deq_1_bits_cf_loadWaitBit; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_5_bits_cf_loadWaitStrict = lsDq_io_deq_1_bits_cf_loadWaitStrict; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_5_bits_cf_ssid = lsDq_io_deq_1_bits_cf_ssid; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_5_bits_cf_ftqPtr_flag = lsDq_io_deq_1_bits_cf_ftqPtr_flag; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_5_bits_cf_ftqPtr_value = lsDq_io_deq_1_bits_cf_ftqPtr_value; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_5_bits_cf_ftqOffset = lsDq_io_deq_1_bits_cf_ftqOffset; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_5_bits_ctrl_srcType_0 = lsDq_io_deq_1_bits_ctrl_srcType_0; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_5_bits_ctrl_srcType_1 = lsDq_io_deq_1_bits_ctrl_srcType_1; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_5_bits_ctrl_fuType = lsDq_io_deq_1_bits_ctrl_fuType; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_5_bits_ctrl_fuOpType = lsDq_io_deq_1_bits_ctrl_fuOpType; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_5_bits_ctrl_rfWen = lsDq_io_deq_1_bits_ctrl_rfWen; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_5_bits_ctrl_fpWen = lsDq_io_deq_1_bits_ctrl_fpWen; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_5_bits_ctrl_flushPipe = lsDq_io_deq_1_bits_ctrl_flushPipe; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_5_bits_ctrl_imm = lsDq_io_deq_1_bits_ctrl_imm; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_5_bits_ctrl_replayInst = lsDq_io_deq_1_bits_ctrl_replayInst; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_5_bits_psrc_0 = lsDq_io_deq_1_bits_psrc_0; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_5_bits_psrc_1 = lsDq_io_deq_1_bits_psrc_1; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_5_bits_pdest = lsDq_io_deq_1_bits_pdest; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_5_bits_robIdx_flag = lsDq_io_deq_1_bits_robIdx_flag; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_5_bits_robIdx_value = lsDq_io_deq_1_bits_robIdx_value; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_6_valid = lsDq_io_deq_2_valid; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_6_bits_cf_foldpc = lsDq_io_deq_2_bits_cf_foldpc; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_6_bits_cf_trigger_backendEn_0 = lsDq_io_deq_2_bits_cf_trigger_backendEn_0; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_6_bits_cf_trigger_backendEn_1 = lsDq_io_deq_2_bits_cf_trigger_backendEn_1; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_6_bits_cf_pd_isRVC = lsDq_io_deq_2_bits_cf_pd_isRVC; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_6_bits_cf_pd_brType = lsDq_io_deq_2_bits_cf_pd_brType; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_6_bits_cf_pd_isCall = lsDq_io_deq_2_bits_cf_pd_isCall; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_6_bits_cf_pd_isRet = lsDq_io_deq_2_bits_cf_pd_isRet; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_6_bits_cf_pred_taken = lsDq_io_deq_2_bits_cf_pred_taken; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_6_bits_cf_storeSetHit = lsDq_io_deq_2_bits_cf_storeSetHit; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_6_bits_cf_waitForRobIdx_flag = lsDq_io_deq_2_bits_cf_waitForRobIdx_flag; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_6_bits_cf_waitForRobIdx_value = lsDq_io_deq_2_bits_cf_waitForRobIdx_value; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_6_bits_cf_loadWaitBit = lsDq_io_deq_2_bits_cf_loadWaitBit; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_6_bits_cf_loadWaitStrict = lsDq_io_deq_2_bits_cf_loadWaitStrict; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_6_bits_cf_ssid = lsDq_io_deq_2_bits_cf_ssid; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_6_bits_cf_ftqPtr_flag = lsDq_io_deq_2_bits_cf_ftqPtr_flag; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_6_bits_cf_ftqPtr_value = lsDq_io_deq_2_bits_cf_ftqPtr_value; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_6_bits_cf_ftqOffset = lsDq_io_deq_2_bits_cf_ftqOffset; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_6_bits_ctrl_srcType_0 = lsDq_io_deq_2_bits_ctrl_srcType_0; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_6_bits_ctrl_srcType_1 = lsDq_io_deq_2_bits_ctrl_srcType_1; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_6_bits_ctrl_fuType = lsDq_io_deq_2_bits_ctrl_fuType; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_6_bits_ctrl_fuOpType = lsDq_io_deq_2_bits_ctrl_fuOpType; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_6_bits_ctrl_rfWen = lsDq_io_deq_2_bits_ctrl_rfWen; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_6_bits_ctrl_fpWen = lsDq_io_deq_2_bits_ctrl_fpWen; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_6_bits_ctrl_flushPipe = lsDq_io_deq_2_bits_ctrl_flushPipe; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_6_bits_ctrl_imm = lsDq_io_deq_2_bits_ctrl_imm; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_6_bits_ctrl_replayInst = lsDq_io_deq_2_bits_ctrl_replayInst; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_6_bits_psrc_0 = lsDq_io_deq_2_bits_psrc_0; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_6_bits_psrc_1 = lsDq_io_deq_2_bits_psrc_1; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_6_bits_pdest = lsDq_io_deq_2_bits_pdest; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_6_bits_robIdx_flag = lsDq_io_deq_2_bits_robIdx_flag; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_6_bits_robIdx_value = lsDq_io_deq_2_bits_robIdx_value; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_7_valid = lsDq_io_deq_3_valid; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_7_bits_cf_foldpc = lsDq_io_deq_3_bits_cf_foldpc; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_7_bits_cf_trigger_backendEn_0 = lsDq_io_deq_3_bits_cf_trigger_backendEn_0; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_7_bits_cf_trigger_backendEn_1 = lsDq_io_deq_3_bits_cf_trigger_backendEn_1; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_7_bits_cf_pd_isRVC = lsDq_io_deq_3_bits_cf_pd_isRVC; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_7_bits_cf_pd_brType = lsDq_io_deq_3_bits_cf_pd_brType; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_7_bits_cf_pd_isCall = lsDq_io_deq_3_bits_cf_pd_isCall; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_7_bits_cf_pd_isRet = lsDq_io_deq_3_bits_cf_pd_isRet; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_7_bits_cf_pred_taken = lsDq_io_deq_3_bits_cf_pred_taken; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_7_bits_cf_storeSetHit = lsDq_io_deq_3_bits_cf_storeSetHit; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_7_bits_cf_waitForRobIdx_flag = lsDq_io_deq_3_bits_cf_waitForRobIdx_flag; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_7_bits_cf_waitForRobIdx_value = lsDq_io_deq_3_bits_cf_waitForRobIdx_value; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_7_bits_cf_loadWaitBit = lsDq_io_deq_3_bits_cf_loadWaitBit; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_7_bits_cf_loadWaitStrict = lsDq_io_deq_3_bits_cf_loadWaitStrict; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_7_bits_cf_ssid = lsDq_io_deq_3_bits_cf_ssid; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_7_bits_cf_ftqPtr_flag = lsDq_io_deq_3_bits_cf_ftqPtr_flag; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_7_bits_cf_ftqPtr_value = lsDq_io_deq_3_bits_cf_ftqPtr_value; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_7_bits_cf_ftqOffset = lsDq_io_deq_3_bits_cf_ftqOffset; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_7_bits_ctrl_srcType_0 = lsDq_io_deq_3_bits_ctrl_srcType_0; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_7_bits_ctrl_srcType_1 = lsDq_io_deq_3_bits_ctrl_srcType_1; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_7_bits_ctrl_fuType = lsDq_io_deq_3_bits_ctrl_fuType; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_7_bits_ctrl_fuOpType = lsDq_io_deq_3_bits_ctrl_fuOpType; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_7_bits_ctrl_rfWen = lsDq_io_deq_3_bits_ctrl_rfWen; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_7_bits_ctrl_fpWen = lsDq_io_deq_3_bits_ctrl_fpWen; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_7_bits_ctrl_flushPipe = lsDq_io_deq_3_bits_ctrl_flushPipe; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_7_bits_ctrl_imm = lsDq_io_deq_3_bits_ctrl_imm; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_7_bits_ctrl_replayInst = lsDq_io_deq_3_bits_ctrl_replayInst; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_7_bits_psrc_0 = lsDq_io_deq_3_bits_psrc_0; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_7_bits_psrc_1 = lsDq_io_deq_3_bits_psrc_1; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_7_bits_pdest = lsDq_io_deq_3_bits_pdest; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_7_bits_robIdx_flag = lsDq_io_deq_3_bits_robIdx_flag; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_7_bits_robIdx_value = lsDq_io_deq_3_bits_robIdx_value; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_8_valid = fpDq_io_deq_0_valid; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_8_bits_cf_pd_isRVC = fpDq_io_deq_0_bits_cf_pd_isRVC; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_8_bits_cf_pd_brType = fpDq_io_deq_0_bits_cf_pd_brType; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_8_bits_cf_pd_isCall = fpDq_io_deq_0_bits_cf_pd_isCall; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_8_bits_cf_pd_isRet = fpDq_io_deq_0_bits_cf_pd_isRet; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_8_bits_cf_pred_taken = fpDq_io_deq_0_bits_cf_pred_taken; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_8_bits_cf_ftqPtr_flag = fpDq_io_deq_0_bits_cf_ftqPtr_flag; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_8_bits_cf_ftqPtr_value = fpDq_io_deq_0_bits_cf_ftqPtr_value; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_8_bits_cf_ftqOffset = fpDq_io_deq_0_bits_cf_ftqOffset; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_8_bits_ctrl_srcType_0 = fpDq_io_deq_0_bits_ctrl_srcType_0; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_8_bits_ctrl_srcType_1 = fpDq_io_deq_0_bits_ctrl_srcType_1; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_8_bits_ctrl_srcType_2 = fpDq_io_deq_0_bits_ctrl_srcType_2; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_8_bits_ctrl_fuType = fpDq_io_deq_0_bits_ctrl_fuType; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_8_bits_ctrl_fuOpType = fpDq_io_deq_0_bits_ctrl_fuOpType; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_8_bits_ctrl_rfWen = fpDq_io_deq_0_bits_ctrl_rfWen; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_8_bits_ctrl_fpWen = fpDq_io_deq_0_bits_ctrl_fpWen; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_8_bits_ctrl_imm = fpDq_io_deq_0_bits_ctrl_imm; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_8_bits_ctrl_fpu_isAddSub = fpDq_io_deq_0_bits_ctrl_fpu_isAddSub; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_8_bits_ctrl_fpu_typeTagIn = fpDq_io_deq_0_bits_ctrl_fpu_typeTagIn; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_8_bits_ctrl_fpu_typeTagOut = fpDq_io_deq_0_bits_ctrl_fpu_typeTagOut; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_8_bits_ctrl_fpu_fromInt = fpDq_io_deq_0_bits_ctrl_fpu_fromInt; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_8_bits_ctrl_fpu_wflags = fpDq_io_deq_0_bits_ctrl_fpu_wflags; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_8_bits_ctrl_fpu_fpWen = fpDq_io_deq_0_bits_ctrl_fpu_fpWen; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_8_bits_ctrl_fpu_fmaCmd = fpDq_io_deq_0_bits_ctrl_fpu_fmaCmd; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_8_bits_ctrl_fpu_div = fpDq_io_deq_0_bits_ctrl_fpu_div; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_8_bits_ctrl_fpu_sqrt = fpDq_io_deq_0_bits_ctrl_fpu_sqrt; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_8_bits_ctrl_fpu_fcvt = fpDq_io_deq_0_bits_ctrl_fpu_fcvt; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_8_bits_ctrl_fpu_typ = fpDq_io_deq_0_bits_ctrl_fpu_typ; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_8_bits_ctrl_fpu_fmt = fpDq_io_deq_0_bits_ctrl_fpu_fmt; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_8_bits_ctrl_fpu_ren3 = fpDq_io_deq_0_bits_ctrl_fpu_ren3; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_8_bits_ctrl_fpu_rm = fpDq_io_deq_0_bits_ctrl_fpu_rm; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_8_bits_psrc_0 = fpDq_io_deq_0_bits_psrc_0; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_8_bits_psrc_1 = fpDq_io_deq_0_bits_psrc_1; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_8_bits_psrc_2 = fpDq_io_deq_0_bits_psrc_2; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_8_bits_pdest = fpDq_io_deq_0_bits_pdest; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_8_bits_robIdx_flag = fpDq_io_deq_0_bits_robIdx_flag; // @[CtrlBlock.scala 508:15]
  assign io_dispatch_8_bits_robIdx_value = fpDq_io_deq_0_bits_robIdx_value; // @[CtrlBlock.scala 508:15]
  assign io_enqLsq_needAlloc_0 = lsqCtrl_io_enqLsq_needAlloc_0; // @[CtrlBlock.scala 526:17]
  assign io_enqLsq_needAlloc_1 = lsqCtrl_io_enqLsq_needAlloc_1; // @[CtrlBlock.scala 526:17]
  assign io_enqLsq_needAlloc_2 = lsqCtrl_io_enqLsq_needAlloc_2; // @[CtrlBlock.scala 526:17]
  assign io_enqLsq_needAlloc_3 = lsqCtrl_io_enqLsq_needAlloc_3; // @[CtrlBlock.scala 526:17]
  assign io_enqLsq_req_0_valid = lsqCtrl_io_enqLsq_req_0_valid; // @[CtrlBlock.scala 526:17]
  assign io_enqLsq_req_0_bits_cf_trigger_backendEn_0 = lsqCtrl_io_enqLsq_req_0_bits_cf_trigger_backendEn_0; // @[CtrlBlock.scala 526:17]
  assign io_enqLsq_req_0_bits_cf_trigger_backendEn_1 = lsqCtrl_io_enqLsq_req_0_bits_cf_trigger_backendEn_1; // @[CtrlBlock.scala 526:17]
  assign io_enqLsq_req_0_bits_ctrl_fuOpType = lsqCtrl_io_enqLsq_req_0_bits_ctrl_fuOpType; // @[CtrlBlock.scala 526:17]
  assign io_enqLsq_req_0_bits_ctrl_rfWen = lsqCtrl_io_enqLsq_req_0_bits_ctrl_rfWen; // @[CtrlBlock.scala 526:17]
  assign io_enqLsq_req_0_bits_ctrl_fpWen = lsqCtrl_io_enqLsq_req_0_bits_ctrl_fpWen; // @[CtrlBlock.scala 526:17]
  assign io_enqLsq_req_0_bits_ctrl_flushPipe = lsqCtrl_io_enqLsq_req_0_bits_ctrl_flushPipe; // @[CtrlBlock.scala 526:17]
  assign io_enqLsq_req_0_bits_ctrl_replayInst = lsqCtrl_io_enqLsq_req_0_bits_ctrl_replayInst; // @[CtrlBlock.scala 526:17]
  assign io_enqLsq_req_0_bits_pdest = lsqCtrl_io_enqLsq_req_0_bits_pdest; // @[CtrlBlock.scala 526:17]
  assign io_enqLsq_req_0_bits_robIdx_flag = lsqCtrl_io_enqLsq_req_0_bits_robIdx_flag; // @[CtrlBlock.scala 526:17]
  assign io_enqLsq_req_0_bits_robIdx_value = lsqCtrl_io_enqLsq_req_0_bits_robIdx_value; // @[CtrlBlock.scala 526:17]
  assign io_enqLsq_req_0_bits_lqIdx_value = lsqCtrl_io_enqLsq_req_0_bits_lqIdx_value; // @[CtrlBlock.scala 526:17]
  assign io_enqLsq_req_0_bits_sqIdx_value = lsqCtrl_io_enqLsq_req_0_bits_sqIdx_value; // @[CtrlBlock.scala 526:17]
  assign io_enqLsq_req_1_valid = lsqCtrl_io_enqLsq_req_1_valid; // @[CtrlBlock.scala 526:17]
  assign io_enqLsq_req_1_bits_cf_trigger_backendEn_0 = lsqCtrl_io_enqLsq_req_1_bits_cf_trigger_backendEn_0; // @[CtrlBlock.scala 526:17]
  assign io_enqLsq_req_1_bits_cf_trigger_backendEn_1 = lsqCtrl_io_enqLsq_req_1_bits_cf_trigger_backendEn_1; // @[CtrlBlock.scala 526:17]
  assign io_enqLsq_req_1_bits_ctrl_fuOpType = lsqCtrl_io_enqLsq_req_1_bits_ctrl_fuOpType; // @[CtrlBlock.scala 526:17]
  assign io_enqLsq_req_1_bits_ctrl_rfWen = lsqCtrl_io_enqLsq_req_1_bits_ctrl_rfWen; // @[CtrlBlock.scala 526:17]
  assign io_enqLsq_req_1_bits_ctrl_fpWen = lsqCtrl_io_enqLsq_req_1_bits_ctrl_fpWen; // @[CtrlBlock.scala 526:17]
  assign io_enqLsq_req_1_bits_ctrl_flushPipe = lsqCtrl_io_enqLsq_req_1_bits_ctrl_flushPipe; // @[CtrlBlock.scala 526:17]
  assign io_enqLsq_req_1_bits_ctrl_replayInst = lsqCtrl_io_enqLsq_req_1_bits_ctrl_replayInst; // @[CtrlBlock.scala 526:17]
  assign io_enqLsq_req_1_bits_pdest = lsqCtrl_io_enqLsq_req_1_bits_pdest; // @[CtrlBlock.scala 526:17]
  assign io_enqLsq_req_1_bits_robIdx_flag = lsqCtrl_io_enqLsq_req_1_bits_robIdx_flag; // @[CtrlBlock.scala 526:17]
  assign io_enqLsq_req_1_bits_robIdx_value = lsqCtrl_io_enqLsq_req_1_bits_robIdx_value; // @[CtrlBlock.scala 526:17]
  assign io_enqLsq_req_1_bits_lqIdx_value = lsqCtrl_io_enqLsq_req_1_bits_lqIdx_value; // @[CtrlBlock.scala 526:17]
  assign io_enqLsq_req_1_bits_sqIdx_value = lsqCtrl_io_enqLsq_req_1_bits_sqIdx_value; // @[CtrlBlock.scala 526:17]
  assign io_enqLsq_req_2_valid = lsqCtrl_io_enqLsq_req_2_valid; // @[CtrlBlock.scala 526:17]
  assign io_enqLsq_req_2_bits_cf_trigger_backendEn_0 = lsqCtrl_io_enqLsq_req_2_bits_cf_trigger_backendEn_0; // @[CtrlBlock.scala 526:17]
  assign io_enqLsq_req_2_bits_cf_trigger_backendEn_1 = lsqCtrl_io_enqLsq_req_2_bits_cf_trigger_backendEn_1; // @[CtrlBlock.scala 526:17]
  assign io_enqLsq_req_2_bits_ctrl_fuOpType = lsqCtrl_io_enqLsq_req_2_bits_ctrl_fuOpType; // @[CtrlBlock.scala 526:17]
  assign io_enqLsq_req_2_bits_ctrl_rfWen = lsqCtrl_io_enqLsq_req_2_bits_ctrl_rfWen; // @[CtrlBlock.scala 526:17]
  assign io_enqLsq_req_2_bits_ctrl_fpWen = lsqCtrl_io_enqLsq_req_2_bits_ctrl_fpWen; // @[CtrlBlock.scala 526:17]
  assign io_enqLsq_req_2_bits_ctrl_flushPipe = lsqCtrl_io_enqLsq_req_2_bits_ctrl_flushPipe; // @[CtrlBlock.scala 526:17]
  assign io_enqLsq_req_2_bits_ctrl_replayInst = lsqCtrl_io_enqLsq_req_2_bits_ctrl_replayInst; // @[CtrlBlock.scala 526:17]
  assign io_enqLsq_req_2_bits_pdest = lsqCtrl_io_enqLsq_req_2_bits_pdest; // @[CtrlBlock.scala 526:17]
  assign io_enqLsq_req_2_bits_robIdx_flag = lsqCtrl_io_enqLsq_req_2_bits_robIdx_flag; // @[CtrlBlock.scala 526:17]
  assign io_enqLsq_req_2_bits_robIdx_value = lsqCtrl_io_enqLsq_req_2_bits_robIdx_value; // @[CtrlBlock.scala 526:17]
  assign io_enqLsq_req_2_bits_lqIdx_value = lsqCtrl_io_enqLsq_req_2_bits_lqIdx_value; // @[CtrlBlock.scala 526:17]
  assign io_enqLsq_req_2_bits_sqIdx_value = lsqCtrl_io_enqLsq_req_2_bits_sqIdx_value; // @[CtrlBlock.scala 526:17]
  assign io_enqLsq_req_3_valid = lsqCtrl_io_enqLsq_req_3_valid; // @[CtrlBlock.scala 526:17]
  assign io_enqLsq_req_3_bits_cf_trigger_backendEn_0 = lsqCtrl_io_enqLsq_req_3_bits_cf_trigger_backendEn_0; // @[CtrlBlock.scala 526:17]
  assign io_enqLsq_req_3_bits_cf_trigger_backendEn_1 = lsqCtrl_io_enqLsq_req_3_bits_cf_trigger_backendEn_1; // @[CtrlBlock.scala 526:17]
  assign io_enqLsq_req_3_bits_ctrl_fuOpType = lsqCtrl_io_enqLsq_req_3_bits_ctrl_fuOpType; // @[CtrlBlock.scala 526:17]
  assign io_enqLsq_req_3_bits_ctrl_rfWen = lsqCtrl_io_enqLsq_req_3_bits_ctrl_rfWen; // @[CtrlBlock.scala 526:17]
  assign io_enqLsq_req_3_bits_ctrl_fpWen = lsqCtrl_io_enqLsq_req_3_bits_ctrl_fpWen; // @[CtrlBlock.scala 526:17]
  assign io_enqLsq_req_3_bits_ctrl_flushPipe = lsqCtrl_io_enqLsq_req_3_bits_ctrl_flushPipe; // @[CtrlBlock.scala 526:17]
  assign io_enqLsq_req_3_bits_ctrl_replayInst = lsqCtrl_io_enqLsq_req_3_bits_ctrl_replayInst; // @[CtrlBlock.scala 526:17]
  assign io_enqLsq_req_3_bits_pdest = lsqCtrl_io_enqLsq_req_3_bits_pdest; // @[CtrlBlock.scala 526:17]
  assign io_enqLsq_req_3_bits_robIdx_flag = lsqCtrl_io_enqLsq_req_3_bits_robIdx_flag; // @[CtrlBlock.scala 526:17]
  assign io_enqLsq_req_3_bits_robIdx_value = lsqCtrl_io_enqLsq_req_3_bits_robIdx_value; // @[CtrlBlock.scala 526:17]
  assign io_enqLsq_req_3_bits_lqIdx_value = lsqCtrl_io_enqLsq_req_3_bits_lqIdx_value; // @[CtrlBlock.scala 526:17]
  assign io_enqLsq_req_3_bits_sqIdx_value = lsqCtrl_io_enqLsq_req_3_bits_sqIdx_value; // @[CtrlBlock.scala 526:17]
  assign io_jumpPc = {jumpPcRead0_hi,1'h0}; // @[Cat.scala 31:58]
  assign io_jalr_target = read_from_newest_entry ? io_jalr_target_REG : pcMem_io_rdata_4_startAddr; // @[CtrlBlock.scala 552:24]
  assign io_robio_toCSR_fflags_valid = rob_io_csr_fflags_valid; // @[CtrlBlock.scala 567:18]
  assign io_robio_toCSR_fflags_bits = rob_io_csr_fflags_bits; // @[CtrlBlock.scala 567:18]
  assign io_robio_toCSR_dirty_fs = rob_io_csr_dirty_fs; // @[CtrlBlock.scala 567:18]
  assign io_robio_toCSR_perfinfo_retiredInstr = io_robio_toCSR_perfinfo_retiredInstr_REG; // @[CtrlBlock.scala 571:40]
  assign io_robio_exception_valid = rob_io_exception_valid; // @[CtrlBlock.scala 572:22]
  assign io_robio_exception_bits_uop_cf_pc = {flushPC_hi,1'h0}; // @[Cat.scala 31:58]
  assign io_robio_exception_bits_uop_cf_exceptionVec_0 = rob_io_exception_bits_uop_cf_exceptionVec_0; // @[CtrlBlock.scala 572:22]
  assign io_robio_exception_bits_uop_cf_exceptionVec_1 = rob_io_exception_bits_uop_cf_exceptionVec_1; // @[CtrlBlock.scala 572:22]
  assign io_robio_exception_bits_uop_cf_exceptionVec_2 = rob_io_exception_bits_uop_cf_exceptionVec_2; // @[CtrlBlock.scala 572:22]
  assign io_robio_exception_bits_uop_cf_exceptionVec_3 = rob_io_exception_bits_uop_cf_exceptionVec_3; // @[CtrlBlock.scala 572:22]
  assign io_robio_exception_bits_uop_cf_exceptionVec_4 = rob_io_exception_bits_uop_cf_exceptionVec_4; // @[CtrlBlock.scala 572:22]
  assign io_robio_exception_bits_uop_cf_exceptionVec_5 = rob_io_exception_bits_uop_cf_exceptionVec_5; // @[CtrlBlock.scala 572:22]
  assign io_robio_exception_bits_uop_cf_exceptionVec_6 = rob_io_exception_bits_uop_cf_exceptionVec_6; // @[CtrlBlock.scala 572:22]
  assign io_robio_exception_bits_uop_cf_exceptionVec_7 = rob_io_exception_bits_uop_cf_exceptionVec_7; // @[CtrlBlock.scala 572:22]
  assign io_robio_exception_bits_uop_cf_exceptionVec_8 = rob_io_exception_bits_uop_cf_exceptionVec_8; // @[CtrlBlock.scala 572:22]
  assign io_robio_exception_bits_uop_cf_exceptionVec_9 = rob_io_exception_bits_uop_cf_exceptionVec_9; // @[CtrlBlock.scala 572:22]
  assign io_robio_exception_bits_uop_cf_exceptionVec_11 = rob_io_exception_bits_uop_cf_exceptionVec_11; // @[CtrlBlock.scala 572:22]
  assign io_robio_exception_bits_uop_cf_exceptionVec_12 = rob_io_exception_bits_uop_cf_exceptionVec_12; // @[CtrlBlock.scala 572:22]
  assign io_robio_exception_bits_uop_cf_exceptionVec_13 = rob_io_exception_bits_uop_cf_exceptionVec_13; // @[CtrlBlock.scala 572:22]
  assign io_robio_exception_bits_uop_cf_exceptionVec_15 = rob_io_exception_bits_uop_cf_exceptionVec_15; // @[CtrlBlock.scala 572:22]
  assign io_robio_exception_bits_uop_cf_trigger_frontendHit_0 = rob_io_exception_bits_uop_cf_trigger_frontendHit_0; // @[CtrlBlock.scala 572:22]
  assign io_robio_exception_bits_uop_cf_trigger_frontendHit_1 = rob_io_exception_bits_uop_cf_trigger_frontendHit_1; // @[CtrlBlock.scala 572:22]
  assign io_robio_exception_bits_uop_cf_trigger_frontendHit_2 = rob_io_exception_bits_uop_cf_trigger_frontendHit_2; // @[CtrlBlock.scala 572:22]
  assign io_robio_exception_bits_uop_cf_trigger_frontendHit_3 = rob_io_exception_bits_uop_cf_trigger_frontendHit_3; // @[CtrlBlock.scala 572:22]
  assign io_robio_exception_bits_uop_cf_trigger_backendHit_0 = rob_io_exception_bits_uop_cf_trigger_backendHit_0; // @[CtrlBlock.scala 572:22]
  assign io_robio_exception_bits_uop_cf_trigger_backendHit_1 = rob_io_exception_bits_uop_cf_trigger_backendHit_1; // @[CtrlBlock.scala 572:22]
  assign io_robio_exception_bits_uop_cf_trigger_backendHit_2 = rob_io_exception_bits_uop_cf_trigger_backendHit_2; // @[CtrlBlock.scala 572:22]
  assign io_robio_exception_bits_uop_cf_trigger_backendHit_3 = rob_io_exception_bits_uop_cf_trigger_backendHit_3; // @[CtrlBlock.scala 572:22]
  assign io_robio_exception_bits_uop_cf_trigger_backendHit_4 = rob_io_exception_bits_uop_cf_trigger_backendHit_4; // @[CtrlBlock.scala 572:22]
  assign io_robio_exception_bits_uop_cf_trigger_backendHit_5 = rob_io_exception_bits_uop_cf_trigger_backendHit_5; // @[CtrlBlock.scala 572:22]
  assign io_robio_exception_bits_uop_cf_crossPageIPFFix = rob_io_exception_bits_uop_cf_crossPageIPFFix; // @[CtrlBlock.scala 572:22]
  assign io_robio_exception_bits_uop_ctrl_commitType = rob_io_exception_bits_uop_ctrl_commitType; // @[CtrlBlock.scala 572:22]
  assign io_robio_exception_bits_uop_ctrl_singleStep = rob_io_exception_bits_uop_ctrl_singleStep; // @[CtrlBlock.scala 572:22]
  assign io_robio_exception_bits_isInterrupt = rob_io_exception_bits_isInterrupt; // @[CtrlBlock.scala 572:22]
  assign io_robio_lsq_scommit = rob_io_lsq_scommit; // @[CtrlBlock.scala 576:16]
  assign io_robio_lsq_pendingld = rob_io_lsq_pendingld; // @[CtrlBlock.scala 576:16]
  assign io_robio_lsq_pendingst = rob_io_lsq_pendingst; // @[CtrlBlock.scala 576:16]
  assign io_robio_lsq_commit = rob_io_lsq_commit; // @[CtrlBlock.scala 576:16]
  assign io_redirect_valid = flushRedirect_valid_REG ? flushRedirect_valid_REG : redirectGen_io_stage2Redirect_valid; // @[CtrlBlock.scala 302:27]
  assign io_redirect_bits_robIdx_flag = flushRedirect_valid_REG ? flushRedirect_bits_rrobIdx_flag :
    redirectGen_io_stage2Redirect_bits_robIdx_flag; // @[CtrlBlock.scala 302:27]
  assign io_redirect_bits_robIdx_value = flushRedirect_valid_REG ? flushRedirect_bits_rrobIdx_value :
    redirectGen_io_stage2Redirect_bits_robIdx_value; // @[CtrlBlock.scala 302:27]
  assign io_redirect_bits_level = flushRedirect_valid_REG ? flushRedirect_bits_rlevel :
    redirectGen_io_stage2Redirect_bits_level; // @[CtrlBlock.scala 302:27]
  assign io_debug_int_rat_0 = rat_io_debug_int_rat_0; // @[CtrlBlock.scala 435:24]
  assign io_debug_int_rat_1 = rat_io_debug_int_rat_1; // @[CtrlBlock.scala 435:24]
  assign io_debug_int_rat_2 = rat_io_debug_int_rat_2; // @[CtrlBlock.scala 435:24]
  assign io_debug_int_rat_3 = rat_io_debug_int_rat_3; // @[CtrlBlock.scala 435:24]
  assign io_debug_int_rat_4 = rat_io_debug_int_rat_4; // @[CtrlBlock.scala 435:24]
  assign io_debug_int_rat_5 = rat_io_debug_int_rat_5; // @[CtrlBlock.scala 435:24]
  assign io_debug_int_rat_6 = rat_io_debug_int_rat_6; // @[CtrlBlock.scala 435:24]
  assign io_debug_int_rat_7 = rat_io_debug_int_rat_7; // @[CtrlBlock.scala 435:24]
  assign io_debug_int_rat_8 = rat_io_debug_int_rat_8; // @[CtrlBlock.scala 435:24]
  assign io_debug_int_rat_9 = rat_io_debug_int_rat_9; // @[CtrlBlock.scala 435:24]
  assign io_debug_int_rat_10 = rat_io_debug_int_rat_10; // @[CtrlBlock.scala 435:24]
  assign io_debug_int_rat_11 = rat_io_debug_int_rat_11; // @[CtrlBlock.scala 435:24]
  assign io_debug_int_rat_12 = rat_io_debug_int_rat_12; // @[CtrlBlock.scala 435:24]
  assign io_debug_int_rat_13 = rat_io_debug_int_rat_13; // @[CtrlBlock.scala 435:24]
  assign io_debug_int_rat_14 = rat_io_debug_int_rat_14; // @[CtrlBlock.scala 435:24]
  assign io_debug_int_rat_15 = rat_io_debug_int_rat_15; // @[CtrlBlock.scala 435:24]
  assign io_debug_int_rat_16 = rat_io_debug_int_rat_16; // @[CtrlBlock.scala 435:24]
  assign io_debug_int_rat_17 = rat_io_debug_int_rat_17; // @[CtrlBlock.scala 435:24]
  assign io_debug_int_rat_18 = rat_io_debug_int_rat_18; // @[CtrlBlock.scala 435:24]
  assign io_debug_int_rat_19 = rat_io_debug_int_rat_19; // @[CtrlBlock.scala 435:24]
  assign io_debug_int_rat_20 = rat_io_debug_int_rat_20; // @[CtrlBlock.scala 435:24]
  assign io_debug_int_rat_21 = rat_io_debug_int_rat_21; // @[CtrlBlock.scala 435:24]
  assign io_debug_int_rat_22 = rat_io_debug_int_rat_22; // @[CtrlBlock.scala 435:24]
  assign io_debug_int_rat_23 = rat_io_debug_int_rat_23; // @[CtrlBlock.scala 435:24]
  assign io_debug_int_rat_24 = rat_io_debug_int_rat_24; // @[CtrlBlock.scala 435:24]
  assign io_debug_int_rat_25 = rat_io_debug_int_rat_25; // @[CtrlBlock.scala 435:24]
  assign io_debug_int_rat_26 = rat_io_debug_int_rat_26; // @[CtrlBlock.scala 435:24]
  assign io_debug_int_rat_27 = rat_io_debug_int_rat_27; // @[CtrlBlock.scala 435:24]
  assign io_debug_int_rat_28 = rat_io_debug_int_rat_28; // @[CtrlBlock.scala 435:24]
  assign io_debug_int_rat_29 = rat_io_debug_int_rat_29; // @[CtrlBlock.scala 435:24]
  assign io_debug_int_rat_30 = rat_io_debug_int_rat_30; // @[CtrlBlock.scala 435:24]
  assign io_debug_int_rat_31 = rat_io_debug_int_rat_31; // @[CtrlBlock.scala 435:24]
  assign io_debug_fp_rat_0 = rat_io_debug_fp_rat_0; // @[CtrlBlock.scala 436:23]
  assign io_debug_fp_rat_1 = rat_io_debug_fp_rat_1; // @[CtrlBlock.scala 436:23]
  assign io_debug_fp_rat_2 = rat_io_debug_fp_rat_2; // @[CtrlBlock.scala 436:23]
  assign io_debug_fp_rat_3 = rat_io_debug_fp_rat_3; // @[CtrlBlock.scala 436:23]
  assign io_debug_fp_rat_4 = rat_io_debug_fp_rat_4; // @[CtrlBlock.scala 436:23]
  assign io_debug_fp_rat_5 = rat_io_debug_fp_rat_5; // @[CtrlBlock.scala 436:23]
  assign io_debug_fp_rat_6 = rat_io_debug_fp_rat_6; // @[CtrlBlock.scala 436:23]
  assign io_debug_fp_rat_7 = rat_io_debug_fp_rat_7; // @[CtrlBlock.scala 436:23]
  assign io_debug_fp_rat_8 = rat_io_debug_fp_rat_8; // @[CtrlBlock.scala 436:23]
  assign io_debug_fp_rat_9 = rat_io_debug_fp_rat_9; // @[CtrlBlock.scala 436:23]
  assign io_debug_fp_rat_10 = rat_io_debug_fp_rat_10; // @[CtrlBlock.scala 436:23]
  assign io_debug_fp_rat_11 = rat_io_debug_fp_rat_11; // @[CtrlBlock.scala 436:23]
  assign io_debug_fp_rat_12 = rat_io_debug_fp_rat_12; // @[CtrlBlock.scala 436:23]
  assign io_debug_fp_rat_13 = rat_io_debug_fp_rat_13; // @[CtrlBlock.scala 436:23]
  assign io_debug_fp_rat_14 = rat_io_debug_fp_rat_14; // @[CtrlBlock.scala 436:23]
  assign io_debug_fp_rat_15 = rat_io_debug_fp_rat_15; // @[CtrlBlock.scala 436:23]
  assign io_debug_fp_rat_16 = rat_io_debug_fp_rat_16; // @[CtrlBlock.scala 436:23]
  assign io_debug_fp_rat_17 = rat_io_debug_fp_rat_17; // @[CtrlBlock.scala 436:23]
  assign io_debug_fp_rat_18 = rat_io_debug_fp_rat_18; // @[CtrlBlock.scala 436:23]
  assign io_debug_fp_rat_19 = rat_io_debug_fp_rat_19; // @[CtrlBlock.scala 436:23]
  assign io_debug_fp_rat_20 = rat_io_debug_fp_rat_20; // @[CtrlBlock.scala 436:23]
  assign io_debug_fp_rat_21 = rat_io_debug_fp_rat_21; // @[CtrlBlock.scala 436:23]
  assign io_debug_fp_rat_22 = rat_io_debug_fp_rat_22; // @[CtrlBlock.scala 436:23]
  assign io_debug_fp_rat_23 = rat_io_debug_fp_rat_23; // @[CtrlBlock.scala 436:23]
  assign io_debug_fp_rat_24 = rat_io_debug_fp_rat_24; // @[CtrlBlock.scala 436:23]
  assign io_debug_fp_rat_25 = rat_io_debug_fp_rat_25; // @[CtrlBlock.scala 436:23]
  assign io_debug_fp_rat_26 = rat_io_debug_fp_rat_26; // @[CtrlBlock.scala 436:23]
  assign io_debug_fp_rat_27 = rat_io_debug_fp_rat_27; // @[CtrlBlock.scala 436:23]
  assign io_debug_fp_rat_28 = rat_io_debug_fp_rat_28; // @[CtrlBlock.scala 436:23]
  assign io_debug_fp_rat_29 = rat_io_debug_fp_rat_29; // @[CtrlBlock.scala 436:23]
  assign io_debug_fp_rat_30 = rat_io_debug_fp_rat_30; // @[CtrlBlock.scala 436:23]
  assign io_debug_fp_rat_31 = rat_io_debug_fp_rat_31; // @[CtrlBlock.scala 436:23]
  assign io_perf_0_value = io_perf_0_value_REG_1; // @[PerfCounterUtils.scala 188:17]
  assign io_perf_1_value = io_perf_1_value_REG_1; // @[PerfCounterUtils.scala 188:17]
  assign io_perf_2_value = io_perf_2_value_REG_1; // @[PerfCounterUtils.scala 188:17]
  assign io_perf_3_value = io_perf_3_value_REG_1; // @[PerfCounterUtils.scala 188:17]
  assign io_perf_4_value = io_perf_4_value_REG_1; // @[PerfCounterUtils.scala 188:17]
  assign io_perf_5_value = io_perf_5_value_REG_1; // @[PerfCounterUtils.scala 188:17]
  assign io_perf_6_value = io_perf_6_value_REG_1; // @[PerfCounterUtils.scala 188:17]
  assign io_perf_7_value = io_perf_7_value_REG_1; // @[PerfCounterUtils.scala 188:17]
  assign rob_clock = clock;
  assign rob_reset = reset;
  assign rob_io_hartId = io_hartId; // @[CtrlBlock.scala 559:17]
  assign rob_io_redirect_valid = flushRedirect_valid_REG ? flushRedirect_valid_REG : redirectGen_io_stage2Redirect_valid
    ; // @[CtrlBlock.scala 302:27]
  assign rob_io_redirect_bits_robIdx_flag = flushRedirect_valid_REG ? flushRedirect_bits_rrobIdx_flag :
    redirectGen_io_stage2Redirect_bits_robIdx_flag; // @[CtrlBlock.scala 302:27]
  assign rob_io_redirect_bits_robIdx_value = flushRedirect_valid_REG ? flushRedirect_bits_rrobIdx_value :
    redirectGen_io_stage2Redirect_bits_robIdx_value; // @[CtrlBlock.scala 302:27]
  assign rob_io_redirect_bits_level = flushRedirect_valid_REG ? flushRedirect_bits_rlevel :
    redirectGen_io_stage2Redirect_bits_level; // @[CtrlBlock.scala 302:27]
  assign rob_io_enq_needAlloc_0 = dispatch_io_enqRob_needAlloc_0; // @[CtrlBlock.scala 496:22]
  assign rob_io_enq_req_0_valid = dispatch_io_enqRob_req_0_valid; // @[CtrlBlock.scala 496:22]
  assign rob_io_enq_req_0_bits_cf_exceptionVec_1 = dispatch_io_enqRob_req_0_bits_cf_exceptionVec_1; // @[CtrlBlock.scala 496:22]
  assign rob_io_enq_req_0_bits_cf_exceptionVec_2 = dispatch_io_enqRob_req_0_bits_cf_exceptionVec_2; // @[CtrlBlock.scala 496:22]
  assign rob_io_enq_req_0_bits_cf_exceptionVec_12 = dispatch_io_enqRob_req_0_bits_cf_exceptionVec_12; // @[CtrlBlock.scala 496:22]
  assign rob_io_enq_req_0_bits_cf_trigger_frontendHit_0 = dispatch_io_enqRob_req_0_bits_cf_trigger_frontendHit_0; // @[CtrlBlock.scala 496:22]
  assign rob_io_enq_req_0_bits_cf_trigger_frontendHit_1 = dispatch_io_enqRob_req_0_bits_cf_trigger_frontendHit_1; // @[CtrlBlock.scala 496:22]
  assign rob_io_enq_req_0_bits_cf_trigger_frontendHit_2 = dispatch_io_enqRob_req_0_bits_cf_trigger_frontendHit_2; // @[CtrlBlock.scala 496:22]
  assign rob_io_enq_req_0_bits_cf_trigger_frontendHit_3 = dispatch_io_enqRob_req_0_bits_cf_trigger_frontendHit_3; // @[CtrlBlock.scala 496:22]
  assign rob_io_enq_req_0_bits_cf_pd_isRVC = dispatch_io_enqRob_req_0_bits_cf_pd_isRVC; // @[CtrlBlock.scala 496:22]
  assign rob_io_enq_req_0_bits_cf_crossPageIPFFix = dispatch_io_enqRob_req_0_bits_cf_crossPageIPFFix; // @[CtrlBlock.scala 496:22]
  assign rob_io_enq_req_0_bits_cf_loadWaitBit = dispatch_io_enqRob_req_0_bits_cf_loadWaitBit; // @[CtrlBlock.scala 496:22]
  assign rob_io_enq_req_0_bits_cf_ftqPtr_flag = dispatch_io_enqRob_req_0_bits_cf_ftqPtr_flag; // @[CtrlBlock.scala 496:22]
  assign rob_io_enq_req_0_bits_cf_ftqPtr_value = dispatch_io_enqRob_req_0_bits_cf_ftqPtr_value; // @[CtrlBlock.scala 496:22]
  assign rob_io_enq_req_0_bits_cf_ftqOffset = dispatch_io_enqRob_req_0_bits_cf_ftqOffset; // @[CtrlBlock.scala 496:22]
  assign rob_io_enq_req_0_bits_ctrl_ldest = dispatch_io_enqRob_req_0_bits_ctrl_ldest; // @[CtrlBlock.scala 496:22]
  assign rob_io_enq_req_0_bits_ctrl_fuType = dispatch_io_enqRob_req_0_bits_ctrl_fuType; // @[CtrlBlock.scala 496:22]
  assign rob_io_enq_req_0_bits_ctrl_fuOpType = dispatch_io_enqRob_req_0_bits_ctrl_fuOpType; // @[CtrlBlock.scala 496:22]
  assign rob_io_enq_req_0_bits_ctrl_rfWen = dispatch_io_enqRob_req_0_bits_ctrl_rfWen; // @[CtrlBlock.scala 496:22]
  assign rob_io_enq_req_0_bits_ctrl_fpWen = dispatch_io_enqRob_req_0_bits_ctrl_fpWen; // @[CtrlBlock.scala 496:22]
  assign rob_io_enq_req_0_bits_ctrl_isXSTrap = dispatch_io_enqRob_req_0_bits_ctrl_isXSTrap; // @[CtrlBlock.scala 496:22]
  assign rob_io_enq_req_0_bits_ctrl_noSpecExec = dispatch_io_enqRob_req_0_bits_ctrl_noSpecExec; // @[CtrlBlock.scala 496:22]
  assign rob_io_enq_req_0_bits_ctrl_blockBackward = dispatch_io_enqRob_req_0_bits_ctrl_blockBackward; // @[CtrlBlock.scala 496:22]
  assign rob_io_enq_req_0_bits_ctrl_flushPipe = dispatch_io_enqRob_req_0_bits_ctrl_flushPipe; // @[CtrlBlock.scala 496:22]
  assign rob_io_enq_req_0_bits_ctrl_commitType = dispatch_io_enqRob_req_0_bits_ctrl_commitType; // @[CtrlBlock.scala 496:22]
  assign rob_io_enq_req_0_bits_ctrl_fpu_wflags = dispatch_io_enqRob_req_0_bits_ctrl_fpu_wflags; // @[CtrlBlock.scala 496:22]
  assign rob_io_enq_req_0_bits_ctrl_isMove = dispatch_io_enqRob_req_0_bits_ctrl_isMove; // @[CtrlBlock.scala 496:22]
  assign rob_io_enq_req_0_bits_ctrl_singleStep = dispatch_io_enqRob_req_0_bits_ctrl_singleStep; // @[CtrlBlock.scala 496:22]
  assign rob_io_enq_req_0_bits_pdest = dispatch_io_enqRob_req_0_bits_pdest; // @[CtrlBlock.scala 496:22]
  assign rob_io_enq_req_0_bits_old_pdest = dispatch_io_enqRob_req_0_bits_old_pdest; // @[CtrlBlock.scala 496:22]
  assign rob_io_enq_req_0_bits_robIdx_flag = dispatch_io_enqRob_req_0_bits_robIdx_flag; // @[CtrlBlock.scala 496:22]
  assign rob_io_enq_req_0_bits_robIdx_value = dispatch_io_enqRob_req_0_bits_robIdx_value; // @[CtrlBlock.scala 496:22]
  assign rob_io_enq_req_0_bits_eliminatedMove = dispatch_io_enqRob_req_0_bits_eliminatedMove; // @[CtrlBlock.scala 496:22]
  assign rob_io_enq_req_1_valid = dispatch_io_enqRob_req_1_valid; // @[CtrlBlock.scala 496:22]
  assign rob_io_enq_req_1_bits_cf_exceptionVec_1 = dispatch_io_enqRob_req_1_bits_cf_exceptionVec_1; // @[CtrlBlock.scala 496:22]
  assign rob_io_enq_req_1_bits_cf_exceptionVec_2 = dispatch_io_enqRob_req_1_bits_cf_exceptionVec_2; // @[CtrlBlock.scala 496:22]
  assign rob_io_enq_req_1_bits_cf_exceptionVec_12 = dispatch_io_enqRob_req_1_bits_cf_exceptionVec_12; // @[CtrlBlock.scala 496:22]
  assign rob_io_enq_req_1_bits_cf_trigger_frontendHit_0 = dispatch_io_enqRob_req_1_bits_cf_trigger_frontendHit_0; // @[CtrlBlock.scala 496:22]
  assign rob_io_enq_req_1_bits_cf_trigger_frontendHit_1 = dispatch_io_enqRob_req_1_bits_cf_trigger_frontendHit_1; // @[CtrlBlock.scala 496:22]
  assign rob_io_enq_req_1_bits_cf_trigger_frontendHit_2 = dispatch_io_enqRob_req_1_bits_cf_trigger_frontendHit_2; // @[CtrlBlock.scala 496:22]
  assign rob_io_enq_req_1_bits_cf_trigger_frontendHit_3 = dispatch_io_enqRob_req_1_bits_cf_trigger_frontendHit_3; // @[CtrlBlock.scala 496:22]
  assign rob_io_enq_req_1_bits_cf_pd_isRVC = dispatch_io_enqRob_req_1_bits_cf_pd_isRVC; // @[CtrlBlock.scala 496:22]
  assign rob_io_enq_req_1_bits_cf_crossPageIPFFix = dispatch_io_enqRob_req_1_bits_cf_crossPageIPFFix; // @[CtrlBlock.scala 496:22]
  assign rob_io_enq_req_1_bits_cf_loadWaitBit = dispatch_io_enqRob_req_1_bits_cf_loadWaitBit; // @[CtrlBlock.scala 496:22]
  assign rob_io_enq_req_1_bits_cf_ftqPtr_flag = dispatch_io_enqRob_req_1_bits_cf_ftqPtr_flag; // @[CtrlBlock.scala 496:22]
  assign rob_io_enq_req_1_bits_cf_ftqPtr_value = dispatch_io_enqRob_req_1_bits_cf_ftqPtr_value; // @[CtrlBlock.scala 496:22]
  assign rob_io_enq_req_1_bits_cf_ftqOffset = dispatch_io_enqRob_req_1_bits_cf_ftqOffset; // @[CtrlBlock.scala 496:22]
  assign rob_io_enq_req_1_bits_ctrl_ldest = dispatch_io_enqRob_req_1_bits_ctrl_ldest; // @[CtrlBlock.scala 496:22]
  assign rob_io_enq_req_1_bits_ctrl_fuType = dispatch_io_enqRob_req_1_bits_ctrl_fuType; // @[CtrlBlock.scala 496:22]
  assign rob_io_enq_req_1_bits_ctrl_fuOpType = dispatch_io_enqRob_req_1_bits_ctrl_fuOpType; // @[CtrlBlock.scala 496:22]
  assign rob_io_enq_req_1_bits_ctrl_rfWen = dispatch_io_enqRob_req_1_bits_ctrl_rfWen; // @[CtrlBlock.scala 496:22]
  assign rob_io_enq_req_1_bits_ctrl_fpWen = dispatch_io_enqRob_req_1_bits_ctrl_fpWen; // @[CtrlBlock.scala 496:22]
  assign rob_io_enq_req_1_bits_ctrl_isXSTrap = dispatch_io_enqRob_req_1_bits_ctrl_isXSTrap; // @[CtrlBlock.scala 496:22]
  assign rob_io_enq_req_1_bits_ctrl_noSpecExec = dispatch_io_enqRob_req_1_bits_ctrl_noSpecExec; // @[CtrlBlock.scala 496:22]
  assign rob_io_enq_req_1_bits_ctrl_blockBackward = dispatch_io_enqRob_req_1_bits_ctrl_blockBackward; // @[CtrlBlock.scala 496:22]
  assign rob_io_enq_req_1_bits_ctrl_flushPipe = dispatch_io_enqRob_req_1_bits_ctrl_flushPipe; // @[CtrlBlock.scala 496:22]
  assign rob_io_enq_req_1_bits_ctrl_commitType = dispatch_io_enqRob_req_1_bits_ctrl_commitType; // @[CtrlBlock.scala 496:22]
  assign rob_io_enq_req_1_bits_ctrl_fpu_wflags = dispatch_io_enqRob_req_1_bits_ctrl_fpu_wflags; // @[CtrlBlock.scala 496:22]
  assign rob_io_enq_req_1_bits_ctrl_isMove = dispatch_io_enqRob_req_1_bits_ctrl_isMove; // @[CtrlBlock.scala 496:22]
  assign rob_io_enq_req_1_bits_ctrl_singleStep = dispatch_io_enqRob_req_1_bits_ctrl_singleStep; // @[CtrlBlock.scala 496:22]
  assign rob_io_enq_req_1_bits_pdest = dispatch_io_enqRob_req_1_bits_pdest; // @[CtrlBlock.scala 496:22]
  assign rob_io_enq_req_1_bits_old_pdest = dispatch_io_enqRob_req_1_bits_old_pdest; // @[CtrlBlock.scala 496:22]
  assign rob_io_enq_req_1_bits_robIdx_flag = dispatch_io_enqRob_req_1_bits_robIdx_flag; // @[CtrlBlock.scala 496:22]
  assign rob_io_enq_req_1_bits_robIdx_value = dispatch_io_enqRob_req_1_bits_robIdx_value; // @[CtrlBlock.scala 496:22]
  assign rob_io_enq_req_1_bits_eliminatedMove = dispatch_io_enqRob_req_1_bits_eliminatedMove; // @[CtrlBlock.scala 496:22]
  assign rob_io_writeback_1_0_valid = sources_source_exuOutput_0_valid_REG_3; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_0_bits_uop_robIdx_value = sources_source_exuOutput_0_bits_REG_3_uop_robIdx_value; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_0_bits_redirectValid = sources_source_exuOutput_0_bits_REG_3_redirectValid; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_0_bits_redirect_cfiUpdate_isMisPred =
    sources_source_exuOutput_0_bits_REG_3_redirect_cfiUpdate_isMisPred; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_1_valid = sources_source_exuOutput_1_valid_REG_3; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_1_bits_uop_robIdx_value = sources_source_exuOutput_1_bits_REG_3_uop_robIdx_value; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_1_bits_redirectValid = sources_source_exuOutput_1_bits_REG_3_redirectValid; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_1_bits_redirect_cfiUpdate_isMisPred =
    sources_source_exuOutput_1_bits_REG_3_redirect_cfiUpdate_isMisPred; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_2_valid = sources_source_exuOutput_2_valid_REG_3; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_2_bits_uop_cf_exceptionVec_4 = sources_source_exuOutput_2_bits_REG_3_uop_cf_exceptionVec_4; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_2_bits_uop_cf_exceptionVec_5 = sources_source_exuOutput_2_bits_REG_3_uop_cf_exceptionVec_5; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_2_bits_uop_cf_exceptionVec_13 = sources_source_exuOutput_2_bits_REG_3_uop_cf_exceptionVec_13
    ; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_2_bits_uop_cf_trigger_backendHit_0 =
    sources_source_exuOutput_2_bits_REG_3_uop_cf_trigger_backendHit_0; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_2_bits_uop_cf_trigger_backendHit_1 =
    sources_source_exuOutput_2_bits_REG_3_uop_cf_trigger_backendHit_1; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_2_bits_uop_cf_trigger_backendHit_2 =
    sources_source_exuOutput_2_bits_REG_3_uop_cf_trigger_backendHit_2; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_2_bits_uop_cf_trigger_backendHit_3 =
    sources_source_exuOutput_2_bits_REG_3_uop_cf_trigger_backendHit_3; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_2_bits_uop_cf_trigger_backendHit_4 =
    sources_source_exuOutput_2_bits_REG_3_uop_cf_trigger_backendHit_4; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_2_bits_uop_cf_trigger_backendHit_5 =
    sources_source_exuOutput_2_bits_REG_3_uop_cf_trigger_backendHit_5; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_2_bits_uop_ctrl_flushPipe = sources_source_exuOutput_2_bits_REG_3_uop_ctrl_flushPipe; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_2_bits_uop_ctrl_replayInst = sources_source_exuOutput_2_bits_REG_3_uop_ctrl_replayInst; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_2_bits_uop_robIdx_value = sources_source_exuOutput_2_bits_REG_3_uop_robIdx_value; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_2_bits_debug_isMMIO = sources_source_exuOutput_2_bits_REG_3_debug_isMMIO; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_3_valid = sources_source_exuOutput_3_valid_REG_3; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_3_bits_uop_cf_exceptionVec_4 = sources_source_exuOutput_3_bits_REG_3_uop_cf_exceptionVec_4; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_3_bits_uop_cf_exceptionVec_5 = sources_source_exuOutput_3_bits_REG_3_uop_cf_exceptionVec_5; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_3_bits_uop_cf_exceptionVec_13 = sources_source_exuOutput_3_bits_REG_3_uop_cf_exceptionVec_13
    ; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_3_bits_uop_cf_trigger_backendHit_0 =
    sources_source_exuOutput_3_bits_REG_3_uop_cf_trigger_backendHit_0; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_3_bits_uop_cf_trigger_backendHit_1 =
    sources_source_exuOutput_3_bits_REG_3_uop_cf_trigger_backendHit_1; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_3_bits_uop_cf_trigger_backendHit_2 =
    sources_source_exuOutput_3_bits_REG_3_uop_cf_trigger_backendHit_2; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_3_bits_uop_cf_trigger_backendHit_3 =
    sources_source_exuOutput_3_bits_REG_3_uop_cf_trigger_backendHit_3; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_3_bits_uop_cf_trigger_backendHit_4 =
    sources_source_exuOutput_3_bits_REG_3_uop_cf_trigger_backendHit_4; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_3_bits_uop_cf_trigger_backendHit_5 =
    sources_source_exuOutput_3_bits_REG_3_uop_cf_trigger_backendHit_5; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_3_bits_uop_ctrl_flushPipe = sources_source_exuOutput_3_bits_REG_3_uop_ctrl_flushPipe; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_3_bits_uop_ctrl_replayInst = sources_source_exuOutput_3_bits_REG_3_uop_ctrl_replayInst; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_3_bits_uop_robIdx_value = sources_source_exuOutput_3_bits_REG_3_uop_robIdx_value; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_3_bits_debug_isMMIO = sources_source_exuOutput_3_bits_REG_3_debug_isMMIO; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_4_valid = sources_source_exuOutput_4_valid_REG_3; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_4_bits_uop_cf_exceptionVec_2 = sources_source_exuOutput_4_bits_REG_3_uop_cf_exceptionVec_2; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_4_bits_uop_cf_exceptionVec_3 = sources_source_exuOutput_4_bits_REG_3_uop_cf_exceptionVec_3; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_4_bits_uop_cf_exceptionVec_8 = sources_source_exuOutput_4_bits_REG_3_uop_cf_exceptionVec_8; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_4_bits_uop_cf_exceptionVec_9 = sources_source_exuOutput_4_bits_REG_3_uop_cf_exceptionVec_9; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_4_bits_uop_cf_exceptionVec_11 = sources_source_exuOutput_4_bits_REG_3_uop_cf_exceptionVec_11
    ; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_4_bits_uop_ctrl_flushPipe = sources_source_exuOutput_4_bits_REG_3_uop_ctrl_flushPipe; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_4_bits_uop_robIdx_value = sources_source_exuOutput_4_bits_REG_3_uop_robIdx_value; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_4_bits_redirectValid = sources_source_exuOutput_4_bits_REG_3_redirectValid; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_4_bits_redirect_cfiUpdate_isMisPred =
    sources_source_exuOutput_4_bits_REG_3_redirect_cfiUpdate_isMisPred; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_4_bits_debug_isPerfCnt = sources_source_exuOutput_4_bits_REG_3_debug_isPerfCnt; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_5_valid = sources_source_exuOutput_5_valid_REG_3; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_5_bits_uop_cf_trigger_backendHit_0 =
    sources_source_exuOutput_5_bits_REG_3_uop_cf_trigger_backendHit_0; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_5_bits_uop_cf_trigger_backendHit_1 =
    sources_source_exuOutput_5_bits_REG_3_uop_cf_trigger_backendHit_1; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_5_bits_uop_cf_trigger_backendHit_2 =
    sources_source_exuOutput_5_bits_REG_3_uop_cf_trigger_backendHit_2; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_5_bits_uop_cf_trigger_backendHit_3 =
    sources_source_exuOutput_5_bits_REG_3_uop_cf_trigger_backendHit_3; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_5_bits_uop_cf_trigger_backendHit_4 =
    sources_source_exuOutput_5_bits_REG_3_uop_cf_trigger_backendHit_4; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_5_bits_uop_cf_trigger_backendHit_5 =
    sources_source_exuOutput_5_bits_REG_3_uop_cf_trigger_backendHit_5; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_5_bits_uop_robIdx_value = sources_source_exuOutput_5_bits_REG_3_uop_robIdx_value; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_6_valid = sources_source_exuOutput_6_valid_REG_3; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_6_bits_uop_cf_exceptionVec_2 = sources_source_exuOutput_6_bits_REG_3_uop_cf_exceptionVec_2; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_6_bits_uop_cf_exceptionVec_3 = sources_source_exuOutput_6_bits_REG_3_uop_cf_exceptionVec_3; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_6_bits_uop_cf_exceptionVec_8 = sources_source_exuOutput_6_bits_REG_3_uop_cf_exceptionVec_8; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_6_bits_uop_cf_exceptionVec_9 = sources_source_exuOutput_6_bits_REG_3_uop_cf_exceptionVec_9; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_6_bits_uop_cf_exceptionVec_11 = sources_source_exuOutput_6_bits_REG_3_uop_cf_exceptionVec_11
    ; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_6_bits_uop_ctrl_flushPipe = sources_source_exuOutput_6_bits_REG_3_uop_ctrl_flushPipe; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_6_bits_uop_robIdx_value = sources_source_exuOutput_6_bits_REG_3_uop_robIdx_value; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_6_bits_redirectValid = sources_source_exuOutput_6_bits_REG_3_redirectValid; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_6_bits_redirect_cfiUpdate_isMisPred =
    sources_source_exuOutput_6_bits_REG_3_redirect_cfiUpdate_isMisPred; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_6_bits_debug_isPerfCnt = sources_source_exuOutput_6_bits_REG_3_debug_isPerfCnt; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_7_valid = sources_source_exuOutput_7_valid_REG_3; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_7_bits_uop_cf_exceptionVec_4 = sources_source_exuOutput_7_bits_REG_3_uop_cf_exceptionVec_4; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_7_bits_uop_cf_exceptionVec_5 = sources_source_exuOutput_7_bits_REG_3_uop_cf_exceptionVec_5; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_7_bits_uop_cf_exceptionVec_6 = sources_source_exuOutput_7_bits_REG_3_uop_cf_exceptionVec_6; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_7_bits_uop_cf_exceptionVec_7 = sources_source_exuOutput_7_bits_REG_3_uop_cf_exceptionVec_7; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_7_bits_uop_cf_exceptionVec_13 = sources_source_exuOutput_7_bits_REG_3_uop_cf_exceptionVec_13
    ; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_7_bits_uop_cf_exceptionVec_15 = sources_source_exuOutput_7_bits_REG_3_uop_cf_exceptionVec_15
    ; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_7_bits_uop_cf_trigger_backendHit_0 =
    sources_source_exuOutput_7_bits_REG_3_uop_cf_trigger_backendHit_0; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_7_bits_uop_cf_trigger_backendHit_1 =
    sources_source_exuOutput_7_bits_REG_3_uop_cf_trigger_backendHit_1; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_7_bits_uop_cf_trigger_backendHit_2 =
    sources_source_exuOutput_7_bits_REG_3_uop_cf_trigger_backendHit_2; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_7_bits_uop_cf_trigger_backendHit_3 =
    sources_source_exuOutput_7_bits_REG_3_uop_cf_trigger_backendHit_3; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_7_bits_uop_cf_trigger_backendHit_4 =
    sources_source_exuOutput_7_bits_REG_3_uop_cf_trigger_backendHit_4; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_7_bits_uop_cf_trigger_backendHit_5 =
    sources_source_exuOutput_7_bits_REG_3_uop_cf_trigger_backendHit_5; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_7_bits_uop_robIdx_value = sources_source_exuOutput_7_bits_REG_3_uop_robIdx_value; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_7_bits_redirectValid = sources_source_exuOutput_7_bits_REG_3_redirectValid; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_7_bits_redirect_cfiUpdate_isMisPred =
    sources_source_exuOutput_7_bits_REG_3_redirect_cfiUpdate_isMisPred; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_7_bits_debug_isMMIO = sources_source_exuOutput_7_bits_REG_3_debug_isMMIO; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_7_bits_debug_isPerfCnt = sources_source_exuOutput_7_bits_REG_3_debug_isPerfCnt; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_8_valid = sources_source_exuOutput_8_valid_REG_3; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_8_bits_uop_cf_exceptionVec_4 = sources_source_exuOutput_8_bits_REG_3_uop_cf_exceptionVec_4; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_8_bits_uop_cf_exceptionVec_5 = sources_source_exuOutput_8_bits_REG_3_uop_cf_exceptionVec_5; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_8_bits_uop_cf_exceptionVec_6 = sources_source_exuOutput_8_bits_REG_3_uop_cf_exceptionVec_6; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_8_bits_uop_cf_exceptionVec_7 = sources_source_exuOutput_8_bits_REG_3_uop_cf_exceptionVec_7; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_8_bits_uop_cf_exceptionVec_13 = sources_source_exuOutput_8_bits_REG_3_uop_cf_exceptionVec_13
    ; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_8_bits_uop_cf_exceptionVec_15 = sources_source_exuOutput_8_bits_REG_3_uop_cf_exceptionVec_15
    ; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_8_bits_uop_cf_trigger_backendHit_0 =
    sources_source_exuOutput_8_bits_REG_3_uop_cf_trigger_backendHit_0; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_8_bits_uop_cf_trigger_backendHit_1 =
    sources_source_exuOutput_8_bits_REG_3_uop_cf_trigger_backendHit_1; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_8_bits_uop_cf_trigger_backendHit_2 =
    sources_source_exuOutput_8_bits_REG_3_uop_cf_trigger_backendHit_2; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_8_bits_uop_cf_trigger_backendHit_3 =
    sources_source_exuOutput_8_bits_REG_3_uop_cf_trigger_backendHit_3; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_8_bits_uop_cf_trigger_backendHit_4 =
    sources_source_exuOutput_8_bits_REG_3_uop_cf_trigger_backendHit_4; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_8_bits_uop_cf_trigger_backendHit_5 =
    sources_source_exuOutput_8_bits_REG_3_uop_cf_trigger_backendHit_5; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_8_bits_uop_robIdx_value = sources_source_exuOutput_8_bits_REG_3_uop_robIdx_value; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_8_bits_redirectValid = sources_source_exuOutput_8_bits_REG_3_redirectValid; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_8_bits_redirect_cfiUpdate_isMisPred =
    sources_source_exuOutput_8_bits_REG_3_redirect_cfiUpdate_isMisPred; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_8_bits_debug_isMMIO = sources_source_exuOutput_8_bits_REG_3_debug_isMMIO; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_8_bits_debug_isPerfCnt = sources_source_exuOutput_8_bits_REG_3_debug_isPerfCnt; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_9_valid = sources_source_exuOutput_9_valid_REG_3; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_9_bits_uop_robIdx_value = sources_source_exuOutput_9_bits_REG_3_uop_robIdx_value; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_10_valid = sources_source_exuOutput_10_valid_REG_3; // @[Rob.scala 379:56]
  assign rob_io_writeback_1_10_bits_uop_robIdx_value = sources_source_exuOutput_10_bits_REG_3_uop_robIdx_value; // @[Rob.scala 379:56]
  assign rob_io_writeback_0_3_valid = sources_source_exuOutput_3_valid_REG; // @[Rob.scala 379:56]
  assign rob_io_writeback_0_3_bits_uop_cf_exceptionVec_2 = sources_source_exuOutput_3_bits_REG_uop_cf_exceptionVec_2; // @[Rob.scala 379:56]
  assign rob_io_writeback_0_3_bits_uop_cf_exceptionVec_3 = sources_source_exuOutput_3_bits_REG_uop_cf_exceptionVec_3; // @[Rob.scala 379:56]
  assign rob_io_writeback_0_3_bits_uop_cf_exceptionVec_8 = sources_source_exuOutput_3_bits_REG_uop_cf_exceptionVec_8; // @[Rob.scala 379:56]
  assign rob_io_writeback_0_3_bits_uop_cf_exceptionVec_9 = sources_source_exuOutput_3_bits_REG_uop_cf_exceptionVec_9; // @[Rob.scala 379:56]
  assign rob_io_writeback_0_3_bits_uop_cf_exceptionVec_11 = sources_source_exuOutput_3_bits_REG_uop_cf_exceptionVec_11; // @[Rob.scala 379:56]
  assign rob_io_writeback_0_3_bits_uop_ctrl_flushPipe = sources_source_exuOutput_3_bits_REG_uop_ctrl_flushPipe; // @[Rob.scala 379:56]
  assign rob_io_writeback_0_3_bits_uop_robIdx_flag = sources_source_exuOutput_3_bits_REG_uop_robIdx_flag; // @[Rob.scala 379:56]
  assign rob_io_writeback_0_3_bits_uop_robIdx_value = sources_source_exuOutput_3_bits_REG_uop_robIdx_value; // @[Rob.scala 379:56]
  assign rob_io_writeback_0_3_bits_fflags = sources_source_exuOutput_3_bits_REG_fflags; // @[Rob.scala 379:56]
  assign rob_io_writeback_0_4_valid = sources_source_exuOutput_4_valid_REG; // @[Rob.scala 379:56]
  assign rob_io_writeback_0_4_bits_uop_robIdx_value = sources_source_exuOutput_4_bits_REG_uop_robIdx_value; // @[Rob.scala 379:56]
  assign rob_io_writeback_0_4_bits_fflags = sources_source_exuOutput_4_bits_REG_fflags; // @[Rob.scala 379:56]
  assign rob_io_writeback_0_5_valid = sources_source_exuOutput_5_valid_REG; // @[Rob.scala 379:56]
  assign rob_io_writeback_0_5_bits_uop_robIdx_value = sources_source_exuOutput_5_bits_REG_uop_robIdx_value; // @[Rob.scala 379:56]
  assign rob_io_writeback_0_5_bits_fflags = sources_source_exuOutput_5_bits_REG_fflags; // @[Rob.scala 379:56]
  assign rob_io_writeback_0_6_valid = sources_source_exuOutput_6_valid_REG; // @[Rob.scala 379:56]
  assign rob_io_writeback_0_6_bits_uop_cf_exceptionVec_4 = sources_source_exuOutput_6_bits_REG_uop_cf_exceptionVec_4; // @[Rob.scala 379:56]
  assign rob_io_writeback_0_6_bits_uop_cf_exceptionVec_5 = sources_source_exuOutput_6_bits_REG_uop_cf_exceptionVec_5; // @[Rob.scala 379:56]
  assign rob_io_writeback_0_6_bits_uop_cf_exceptionVec_13 = sources_source_exuOutput_6_bits_REG_uop_cf_exceptionVec_13; // @[Rob.scala 379:56]
  assign rob_io_writeback_0_6_bits_uop_cf_trigger_backendHit_0 =
    sources_source_exuOutput_6_bits_REG_uop_cf_trigger_backendHit_0; // @[Rob.scala 379:56]
  assign rob_io_writeback_0_6_bits_uop_cf_trigger_backendHit_1 =
    sources_source_exuOutput_6_bits_REG_uop_cf_trigger_backendHit_1; // @[Rob.scala 379:56]
  assign rob_io_writeback_0_6_bits_uop_cf_trigger_backendHit_2 =
    sources_source_exuOutput_6_bits_REG_uop_cf_trigger_backendHit_2; // @[Rob.scala 379:56]
  assign rob_io_writeback_0_6_bits_uop_cf_trigger_backendHit_3 =
    sources_source_exuOutput_6_bits_REG_uop_cf_trigger_backendHit_3; // @[Rob.scala 379:56]
  assign rob_io_writeback_0_6_bits_uop_cf_trigger_backendHit_4 =
    sources_source_exuOutput_6_bits_REG_uop_cf_trigger_backendHit_4; // @[Rob.scala 379:56]
  assign rob_io_writeback_0_6_bits_uop_cf_trigger_backendHit_5 =
    sources_source_exuOutput_6_bits_REG_uop_cf_trigger_backendHit_5; // @[Rob.scala 379:56]
  assign rob_io_writeback_0_6_bits_uop_ctrl_flushPipe = sources_source_exuOutput_6_bits_REG_uop_ctrl_flushPipe; // @[Rob.scala 379:56]
  assign rob_io_writeback_0_6_bits_uop_ctrl_replayInst = sources_source_exuOutput_6_bits_REG_uop_ctrl_replayInst; // @[Rob.scala 379:56]
  assign rob_io_writeback_0_6_bits_uop_robIdx_flag = sources_source_exuOutput_6_bits_REG_uop_robIdx_flag; // @[Rob.scala 379:56]
  assign rob_io_writeback_0_6_bits_uop_robIdx_value = sources_source_exuOutput_6_bits_REG_uop_robIdx_value; // @[Rob.scala 379:56]
  assign rob_io_writeback_0_7_valid = sources_source_exuOutput_7_valid_REG; // @[Rob.scala 379:56]
  assign rob_io_writeback_0_7_bits_uop_cf_exceptionVec_4 = sources_source_exuOutput_7_bits_REG_uop_cf_exceptionVec_4; // @[Rob.scala 379:56]
  assign rob_io_writeback_0_7_bits_uop_cf_exceptionVec_5 = sources_source_exuOutput_7_bits_REG_uop_cf_exceptionVec_5; // @[Rob.scala 379:56]
  assign rob_io_writeback_0_7_bits_uop_cf_exceptionVec_13 = sources_source_exuOutput_7_bits_REG_uop_cf_exceptionVec_13; // @[Rob.scala 379:56]
  assign rob_io_writeback_0_7_bits_uop_cf_trigger_backendHit_0 =
    sources_source_exuOutput_7_bits_REG_uop_cf_trigger_backendHit_0; // @[Rob.scala 379:56]
  assign rob_io_writeback_0_7_bits_uop_cf_trigger_backendHit_1 =
    sources_source_exuOutput_7_bits_REG_uop_cf_trigger_backendHit_1; // @[Rob.scala 379:56]
  assign rob_io_writeback_0_7_bits_uop_cf_trigger_backendHit_2 =
    sources_source_exuOutput_7_bits_REG_uop_cf_trigger_backendHit_2; // @[Rob.scala 379:56]
  assign rob_io_writeback_0_7_bits_uop_cf_trigger_backendHit_3 =
    sources_source_exuOutput_7_bits_REG_uop_cf_trigger_backendHit_3; // @[Rob.scala 379:56]
  assign rob_io_writeback_0_7_bits_uop_cf_trigger_backendHit_4 =
    sources_source_exuOutput_7_bits_REG_uop_cf_trigger_backendHit_4; // @[Rob.scala 379:56]
  assign rob_io_writeback_0_7_bits_uop_cf_trigger_backendHit_5 =
    sources_source_exuOutput_7_bits_REG_uop_cf_trigger_backendHit_5; // @[Rob.scala 379:56]
  assign rob_io_writeback_0_7_bits_uop_ctrl_flushPipe = sources_source_exuOutput_7_bits_REG_uop_ctrl_flushPipe; // @[Rob.scala 379:56]
  assign rob_io_writeback_0_7_bits_uop_ctrl_replayInst = sources_source_exuOutput_7_bits_REG_uop_ctrl_replayInst; // @[Rob.scala 379:56]
  assign rob_io_writeback_0_7_bits_uop_robIdx_flag = sources_source_exuOutput_7_bits_REG_uop_robIdx_flag; // @[Rob.scala 379:56]
  assign rob_io_writeback_0_7_bits_uop_robIdx_value = sources_source_exuOutput_7_bits_REG_uop_robIdx_value; // @[Rob.scala 379:56]
  assign rob_io_writeback_0_8_valid = sources_source_exuOutput_8_valid_REG; // @[Rob.scala 379:56]
  assign rob_io_writeback_0_8_bits_uop_cf_exceptionVec_4 = sources_source_exuOutput_8_bits_REG_uop_cf_exceptionVec_4; // @[Rob.scala 379:56]
  assign rob_io_writeback_0_8_bits_uop_cf_exceptionVec_5 = sources_source_exuOutput_8_bits_REG_uop_cf_exceptionVec_5; // @[Rob.scala 379:56]
  assign rob_io_writeback_0_8_bits_uop_cf_exceptionVec_6 = sources_source_exuOutput_8_bits_REG_uop_cf_exceptionVec_6; // @[Rob.scala 379:56]
  assign rob_io_writeback_0_8_bits_uop_cf_exceptionVec_7 = sources_source_exuOutput_8_bits_REG_uop_cf_exceptionVec_7; // @[Rob.scala 379:56]
  assign rob_io_writeback_0_8_bits_uop_cf_exceptionVec_13 = sources_source_exuOutput_8_bits_REG_uop_cf_exceptionVec_13; // @[Rob.scala 379:56]
  assign rob_io_writeback_0_8_bits_uop_cf_exceptionVec_15 = sources_source_exuOutput_8_bits_REG_uop_cf_exceptionVec_15; // @[Rob.scala 379:56]
  assign rob_io_writeback_0_8_bits_uop_cf_trigger_backendHit_0 =
    sources_source_exuOutput_8_bits_REG_uop_cf_trigger_backendHit_0; // @[Rob.scala 379:56]
  assign rob_io_writeback_0_8_bits_uop_cf_trigger_backendHit_1 =
    sources_source_exuOutput_8_bits_REG_uop_cf_trigger_backendHit_1; // @[Rob.scala 379:56]
  assign rob_io_writeback_0_8_bits_uop_cf_trigger_backendHit_2 =
    sources_source_exuOutput_8_bits_REG_uop_cf_trigger_backendHit_2; // @[Rob.scala 379:56]
  assign rob_io_writeback_0_8_bits_uop_cf_trigger_backendHit_3 =
    sources_source_exuOutput_8_bits_REG_uop_cf_trigger_backendHit_3; // @[Rob.scala 379:56]
  assign rob_io_writeback_0_8_bits_uop_cf_trigger_backendHit_4 =
    sources_source_exuOutput_8_bits_REG_uop_cf_trigger_backendHit_4; // @[Rob.scala 379:56]
  assign rob_io_writeback_0_8_bits_uop_cf_trigger_backendHit_5 =
    sources_source_exuOutput_8_bits_REG_uop_cf_trigger_backendHit_5; // @[Rob.scala 379:56]
  assign rob_io_writeback_0_8_bits_uop_robIdx_flag = sources_source_exuOutput_8_bits_REG_uop_robIdx_flag; // @[Rob.scala 379:56]
  assign rob_io_writeback_0_8_bits_uop_robIdx_value = sources_source_exuOutput_8_bits_REG_uop_robIdx_value; // @[Rob.scala 379:56]
  assign rob_io_writeback_0_9_valid = sources_source_exuOutput_9_valid_REG; // @[Rob.scala 379:56]
  assign rob_io_writeback_0_9_bits_uop_cf_exceptionVec_6 = sources_source_exuOutput_9_bits_REG_uop_cf_exceptionVec_6; // @[Rob.scala 379:56]
  assign rob_io_writeback_0_9_bits_uop_cf_exceptionVec_7 = sources_source_exuOutput_9_bits_REG_uop_cf_exceptionVec_7; // @[Rob.scala 379:56]
  assign rob_io_writeback_0_9_bits_uop_cf_exceptionVec_15 = sources_source_exuOutput_9_bits_REG_uop_cf_exceptionVec_15; // @[Rob.scala 379:56]
  assign rob_io_writeback_0_9_bits_uop_cf_trigger_backendHit_0 =
    sources_source_exuOutput_9_bits_REG_uop_cf_trigger_backendHit_0; // @[Rob.scala 379:56]
  assign rob_io_writeback_0_9_bits_uop_cf_trigger_backendHit_1 =
    sources_source_exuOutput_9_bits_REG_uop_cf_trigger_backendHit_1; // @[Rob.scala 379:56]
  assign rob_io_writeback_0_9_bits_uop_cf_trigger_backendHit_4 =
    sources_source_exuOutput_9_bits_REG_uop_cf_trigger_backendHit_4; // @[Rob.scala 379:56]
  assign rob_io_writeback_0_9_bits_uop_robIdx_flag = sources_source_exuOutput_9_bits_REG_uop_robIdx_flag; // @[Rob.scala 379:56]
  assign rob_io_writeback_0_9_bits_uop_robIdx_value = sources_source_exuOutput_9_bits_REG_uop_robIdx_value; // @[Rob.scala 379:56]
  assign rob_io_lsq_isMMIO_0 = io_robio_lsq_isMMIO_0; // @[CtrlBlock.scala 576:16]
  assign rob_io_lsq_isMMIO_1 = io_robio_lsq_isMMIO_1; // @[CtrlBlock.scala 576:16]
  assign rob_io_lsq_uop_0_robIdx_value = io_robio_lsq_uop_0_robIdx_value; // @[CtrlBlock.scala 576:16]
  assign rob_io_lsq_uop_1_robIdx_value = io_robio_lsq_uop_1_robIdx_value; // @[CtrlBlock.scala 576:16]
  assign rob_io_csr_intrBitSet = io_robio_toCSR_intrBitSet; // @[CtrlBlock.scala 567:18]
  assign rob_io_csr_wfiEvent = io_robio_toCSR_wfiEvent; // @[CtrlBlock.scala 569:23]
  assign rob_io_wfi_enable = decode_io_csrCtrl_wfi_enable; // @[CtrlBlock.scala 570:21]
  assign dispatch2_io_in_1_bits_ctrl_fuType = intDq_io_deq_1_bits_ctrl_fuType; // @[CtrlBlock.scala 531:16]
  assign dispatch2_io_out_0_ready = io_rsReady_0; // @[CtrlBlock.scala 536:18]
  assign dispatch2_io_out_1_ready = io_rsReady_1; // @[CtrlBlock.scala 536:18]
  assign dispatch2_1_clock = clock;
  assign dispatch2_1_reset = reset;
  assign dispatch2_1_io_redirect_valid = redirectForExu_next_valid_REG; // @[BitUtils.scala 26:20 28:18]
  assign dispatch2_1_io_redirect_bits_robIdx_flag = redirectForExu_next_bits_rrobIdx_flag; // @[BitUtils.scala 26:20 33:15]
  assign dispatch2_1_io_redirect_bits_robIdx_value = redirectForExu_next_bits_rrobIdx_value; // @[BitUtils.scala 26:20 33:15]
  assign dispatch2_1_io_redirect_bits_level = redirectForExu_next_bits_rlevel; // @[BitUtils.scala 26:20 33:15]
  assign dispatch2_1_io_in_0_valid = lsDq_io_deq_0_valid; // @[CtrlBlock.scala 530:17]
  assign dispatch2_1_io_in_0_bits_cf_foldpc = lsDq_io_deq_0_bits_cf_foldpc; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_0_bits_cf_trigger_backendEn_0 = lsDq_io_deq_0_bits_cf_trigger_backendEn_0; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_0_bits_cf_trigger_backendEn_1 = lsDq_io_deq_0_bits_cf_trigger_backendEn_1; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_0_bits_cf_pd_isRVC = lsDq_io_deq_0_bits_cf_pd_isRVC; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_0_bits_cf_pd_brType = lsDq_io_deq_0_bits_cf_pd_brType; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_0_bits_cf_pd_isCall = lsDq_io_deq_0_bits_cf_pd_isCall; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_0_bits_cf_pd_isRet = lsDq_io_deq_0_bits_cf_pd_isRet; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_0_bits_cf_pred_taken = lsDq_io_deq_0_bits_cf_pred_taken; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_0_bits_cf_storeSetHit = lsDq_io_deq_0_bits_cf_storeSetHit; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_0_bits_cf_waitForRobIdx_flag = lsDq_io_deq_0_bits_cf_waitForRobIdx_flag; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_0_bits_cf_waitForRobIdx_value = lsDq_io_deq_0_bits_cf_waitForRobIdx_value; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_0_bits_cf_loadWaitBit = lsDq_io_deq_0_bits_cf_loadWaitBit; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_0_bits_cf_loadWaitStrict = lsDq_io_deq_0_bits_cf_loadWaitStrict; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_0_bits_cf_ssid = lsDq_io_deq_0_bits_cf_ssid; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_0_bits_cf_ftqPtr_flag = lsDq_io_deq_0_bits_cf_ftqPtr_flag; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_0_bits_cf_ftqPtr_value = lsDq_io_deq_0_bits_cf_ftqPtr_value; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_0_bits_cf_ftqOffset = lsDq_io_deq_0_bits_cf_ftqOffset; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_0_bits_ctrl_srcType_0 = lsDq_io_deq_0_bits_ctrl_srcType_0; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_0_bits_ctrl_srcType_1 = lsDq_io_deq_0_bits_ctrl_srcType_1; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_0_bits_ctrl_fuType = lsDq_io_deq_0_bits_ctrl_fuType; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_0_bits_ctrl_fuOpType = lsDq_io_deq_0_bits_ctrl_fuOpType; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_0_bits_ctrl_rfWen = lsDq_io_deq_0_bits_ctrl_rfWen; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_0_bits_ctrl_fpWen = lsDq_io_deq_0_bits_ctrl_fpWen; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_0_bits_ctrl_flushPipe = lsDq_io_deq_0_bits_ctrl_flushPipe; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_0_bits_ctrl_imm = lsDq_io_deq_0_bits_ctrl_imm; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_0_bits_ctrl_replayInst = lsDq_io_deq_0_bits_ctrl_replayInst; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_0_bits_psrc_0 = lsDq_io_deq_0_bits_psrc_0; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_0_bits_psrc_1 = lsDq_io_deq_0_bits_psrc_1; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_0_bits_pdest = lsDq_io_deq_0_bits_pdest; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_0_bits_robIdx_flag = lsDq_io_deq_0_bits_robIdx_flag; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_0_bits_robIdx_value = lsDq_io_deq_0_bits_robIdx_value; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_1_valid = lsDq_io_deq_1_valid; // @[CtrlBlock.scala 530:17]
  assign dispatch2_1_io_in_1_bits_cf_foldpc = lsDq_io_deq_1_bits_cf_foldpc; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_1_bits_cf_trigger_backendEn_0 = lsDq_io_deq_1_bits_cf_trigger_backendEn_0; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_1_bits_cf_trigger_backendEn_1 = lsDq_io_deq_1_bits_cf_trigger_backendEn_1; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_1_bits_cf_pd_isRVC = lsDq_io_deq_1_bits_cf_pd_isRVC; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_1_bits_cf_pd_brType = lsDq_io_deq_1_bits_cf_pd_brType; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_1_bits_cf_pd_isCall = lsDq_io_deq_1_bits_cf_pd_isCall; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_1_bits_cf_pd_isRet = lsDq_io_deq_1_bits_cf_pd_isRet; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_1_bits_cf_pred_taken = lsDq_io_deq_1_bits_cf_pred_taken; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_1_bits_cf_storeSetHit = lsDq_io_deq_1_bits_cf_storeSetHit; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_1_bits_cf_waitForRobIdx_flag = lsDq_io_deq_1_bits_cf_waitForRobIdx_flag; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_1_bits_cf_waitForRobIdx_value = lsDq_io_deq_1_bits_cf_waitForRobIdx_value; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_1_bits_cf_loadWaitBit = lsDq_io_deq_1_bits_cf_loadWaitBit; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_1_bits_cf_loadWaitStrict = lsDq_io_deq_1_bits_cf_loadWaitStrict; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_1_bits_cf_ssid = lsDq_io_deq_1_bits_cf_ssid; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_1_bits_cf_ftqPtr_flag = lsDq_io_deq_1_bits_cf_ftqPtr_flag; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_1_bits_cf_ftqPtr_value = lsDq_io_deq_1_bits_cf_ftqPtr_value; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_1_bits_cf_ftqOffset = lsDq_io_deq_1_bits_cf_ftqOffset; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_1_bits_ctrl_srcType_0 = lsDq_io_deq_1_bits_ctrl_srcType_0; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_1_bits_ctrl_srcType_1 = lsDq_io_deq_1_bits_ctrl_srcType_1; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_1_bits_ctrl_fuType = lsDq_io_deq_1_bits_ctrl_fuType; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_1_bits_ctrl_fuOpType = lsDq_io_deq_1_bits_ctrl_fuOpType; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_1_bits_ctrl_rfWen = lsDq_io_deq_1_bits_ctrl_rfWen; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_1_bits_ctrl_fpWen = lsDq_io_deq_1_bits_ctrl_fpWen; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_1_bits_ctrl_flushPipe = lsDq_io_deq_1_bits_ctrl_flushPipe; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_1_bits_ctrl_imm = lsDq_io_deq_1_bits_ctrl_imm; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_1_bits_ctrl_replayInst = lsDq_io_deq_1_bits_ctrl_replayInst; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_1_bits_psrc_0 = lsDq_io_deq_1_bits_psrc_0; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_1_bits_psrc_1 = lsDq_io_deq_1_bits_psrc_1; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_1_bits_pdest = lsDq_io_deq_1_bits_pdest; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_1_bits_robIdx_flag = lsDq_io_deq_1_bits_robIdx_flag; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_1_bits_robIdx_value = lsDq_io_deq_1_bits_robIdx_value; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_2_valid = lsDq_io_deq_2_valid; // @[CtrlBlock.scala 530:17]
  assign dispatch2_1_io_in_2_bits_cf_foldpc = lsDq_io_deq_2_bits_cf_foldpc; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_2_bits_cf_trigger_backendEn_0 = lsDq_io_deq_2_bits_cf_trigger_backendEn_0; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_2_bits_cf_trigger_backendEn_1 = lsDq_io_deq_2_bits_cf_trigger_backendEn_1; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_2_bits_cf_pd_isRVC = lsDq_io_deq_2_bits_cf_pd_isRVC; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_2_bits_cf_pd_brType = lsDq_io_deq_2_bits_cf_pd_brType; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_2_bits_cf_pd_isCall = lsDq_io_deq_2_bits_cf_pd_isCall; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_2_bits_cf_pd_isRet = lsDq_io_deq_2_bits_cf_pd_isRet; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_2_bits_cf_pred_taken = lsDq_io_deq_2_bits_cf_pred_taken; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_2_bits_cf_storeSetHit = lsDq_io_deq_2_bits_cf_storeSetHit; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_2_bits_cf_waitForRobIdx_flag = lsDq_io_deq_2_bits_cf_waitForRobIdx_flag; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_2_bits_cf_waitForRobIdx_value = lsDq_io_deq_2_bits_cf_waitForRobIdx_value; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_2_bits_cf_loadWaitBit = lsDq_io_deq_2_bits_cf_loadWaitBit; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_2_bits_cf_loadWaitStrict = lsDq_io_deq_2_bits_cf_loadWaitStrict; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_2_bits_cf_ssid = lsDq_io_deq_2_bits_cf_ssid; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_2_bits_cf_ftqPtr_flag = lsDq_io_deq_2_bits_cf_ftqPtr_flag; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_2_bits_cf_ftqPtr_value = lsDq_io_deq_2_bits_cf_ftqPtr_value; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_2_bits_cf_ftqOffset = lsDq_io_deq_2_bits_cf_ftqOffset; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_2_bits_ctrl_srcType_0 = lsDq_io_deq_2_bits_ctrl_srcType_0; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_2_bits_ctrl_srcType_1 = lsDq_io_deq_2_bits_ctrl_srcType_1; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_2_bits_ctrl_fuType = lsDq_io_deq_2_bits_ctrl_fuType; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_2_bits_ctrl_fuOpType = lsDq_io_deq_2_bits_ctrl_fuOpType; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_2_bits_ctrl_rfWen = lsDq_io_deq_2_bits_ctrl_rfWen; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_2_bits_ctrl_fpWen = lsDq_io_deq_2_bits_ctrl_fpWen; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_2_bits_ctrl_flushPipe = lsDq_io_deq_2_bits_ctrl_flushPipe; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_2_bits_ctrl_imm = lsDq_io_deq_2_bits_ctrl_imm; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_2_bits_ctrl_replayInst = lsDq_io_deq_2_bits_ctrl_replayInst; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_2_bits_psrc_0 = lsDq_io_deq_2_bits_psrc_0; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_2_bits_psrc_1 = lsDq_io_deq_2_bits_psrc_1; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_2_bits_pdest = lsDq_io_deq_2_bits_pdest; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_2_bits_robIdx_flag = lsDq_io_deq_2_bits_robIdx_flag; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_2_bits_robIdx_value = lsDq_io_deq_2_bits_robIdx_value; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_3_valid = lsDq_io_deq_3_valid; // @[CtrlBlock.scala 530:17]
  assign dispatch2_1_io_in_3_bits_cf_foldpc = lsDq_io_deq_3_bits_cf_foldpc; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_3_bits_cf_trigger_backendEn_0 = lsDq_io_deq_3_bits_cf_trigger_backendEn_0; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_3_bits_cf_trigger_backendEn_1 = lsDq_io_deq_3_bits_cf_trigger_backendEn_1; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_3_bits_cf_pd_isRVC = lsDq_io_deq_3_bits_cf_pd_isRVC; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_3_bits_cf_pd_brType = lsDq_io_deq_3_bits_cf_pd_brType; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_3_bits_cf_pd_isCall = lsDq_io_deq_3_bits_cf_pd_isCall; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_3_bits_cf_pd_isRet = lsDq_io_deq_3_bits_cf_pd_isRet; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_3_bits_cf_pred_taken = lsDq_io_deq_3_bits_cf_pred_taken; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_3_bits_cf_storeSetHit = lsDq_io_deq_3_bits_cf_storeSetHit; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_3_bits_cf_waitForRobIdx_flag = lsDq_io_deq_3_bits_cf_waitForRobIdx_flag; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_3_bits_cf_waitForRobIdx_value = lsDq_io_deq_3_bits_cf_waitForRobIdx_value; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_3_bits_cf_loadWaitBit = lsDq_io_deq_3_bits_cf_loadWaitBit; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_3_bits_cf_loadWaitStrict = lsDq_io_deq_3_bits_cf_loadWaitStrict; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_3_bits_cf_ssid = lsDq_io_deq_3_bits_cf_ssid; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_3_bits_cf_ftqPtr_flag = lsDq_io_deq_3_bits_cf_ftqPtr_flag; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_3_bits_cf_ftqPtr_value = lsDq_io_deq_3_bits_cf_ftqPtr_value; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_3_bits_cf_ftqOffset = lsDq_io_deq_3_bits_cf_ftqOffset; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_3_bits_ctrl_srcType_0 = lsDq_io_deq_3_bits_ctrl_srcType_0; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_3_bits_ctrl_srcType_1 = lsDq_io_deq_3_bits_ctrl_srcType_1; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_3_bits_ctrl_fuType = lsDq_io_deq_3_bits_ctrl_fuType; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_3_bits_ctrl_fuOpType = lsDq_io_deq_3_bits_ctrl_fuOpType; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_3_bits_ctrl_rfWen = lsDq_io_deq_3_bits_ctrl_rfWen; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_3_bits_ctrl_fpWen = lsDq_io_deq_3_bits_ctrl_fpWen; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_3_bits_ctrl_flushPipe = lsDq_io_deq_3_bits_ctrl_flushPipe; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_3_bits_ctrl_imm = lsDq_io_deq_3_bits_ctrl_imm; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_3_bits_ctrl_replayInst = lsDq_io_deq_3_bits_ctrl_replayInst; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_3_bits_psrc_0 = lsDq_io_deq_3_bits_psrc_0; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_3_bits_psrc_1 = lsDq_io_deq_3_bits_psrc_1; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_3_bits_pdest = lsDq_io_deq_3_bits_pdest; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_3_bits_robIdx_flag = lsDq_io_deq_3_bits_robIdx_flag; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_in_3_bits_robIdx_value = lsDq_io_deq_3_bits_robIdx_value; // @[CtrlBlock.scala 531:16]
  assign dispatch2_1_io_readIntState_0_resp = 1'h0;
  assign dispatch2_1_io_readIntState_1_resp = 1'h0;
  assign dispatch2_1_io_readIntState_2_resp = 1'h0;
  assign dispatch2_1_io_readIntState_3_resp = 1'h0;
  assign dispatch2_1_io_readIntState_4_resp = 1'h0;
  assign dispatch2_1_io_readIntState_5_resp = 1'h0;
  assign dispatch2_1_io_readFpState_0_resp = 1'h0;
  assign dispatch2_1_io_readFpState_1_resp = 1'h0;
  assign dispatch2_1_io_out_0_ready = io_rsReady_2; // @[CtrlBlock.scala 536:18]
  assign dispatch2_1_io_out_1_ready = io_rsReady_3; // @[CtrlBlock.scala 536:18]
  assign dispatch2_1_io_out_2_ready = io_rsReady_4; // @[CtrlBlock.scala 536:18]
  assign dispatch2_1_io_out_3_ready = io_rsReady_5; // @[CtrlBlock.scala 536:18]
  assign dispatch2_1_io_out_4_ready = io_rsReady_6; // @[CtrlBlock.scala 536:18]
  assign dispatch2_1_io_out_5_ready = io_rsReady_7; // @[CtrlBlock.scala 536:18]
  assign dispatch2_1_io_enqLsq_canAccept = lsqCtrl_io_enq_canAccept; // @[CtrlBlock.scala 521:22]
  assign dispatch2_1_io_enqLsq_resp_0_lqIdx_flag = lsqCtrl_io_enq_resp_0_lqIdx_flag; // @[CtrlBlock.scala 521:22]
  assign dispatch2_1_io_enqLsq_resp_0_lqIdx_value = lsqCtrl_io_enq_resp_0_lqIdx_value; // @[CtrlBlock.scala 521:22]
  assign dispatch2_1_io_enqLsq_resp_0_sqIdx_flag = lsqCtrl_io_enq_resp_0_sqIdx_flag; // @[CtrlBlock.scala 521:22]
  assign dispatch2_1_io_enqLsq_resp_0_sqIdx_value = lsqCtrl_io_enq_resp_0_sqIdx_value; // @[CtrlBlock.scala 521:22]
  assign dispatch2_1_io_enqLsq_resp_1_lqIdx_flag = lsqCtrl_io_enq_resp_1_lqIdx_flag; // @[CtrlBlock.scala 521:22]
  assign dispatch2_1_io_enqLsq_resp_1_lqIdx_value = lsqCtrl_io_enq_resp_1_lqIdx_value; // @[CtrlBlock.scala 521:22]
  assign dispatch2_1_io_enqLsq_resp_1_sqIdx_flag = lsqCtrl_io_enq_resp_1_sqIdx_flag; // @[CtrlBlock.scala 521:22]
  assign dispatch2_1_io_enqLsq_resp_1_sqIdx_value = lsqCtrl_io_enq_resp_1_sqIdx_value; // @[CtrlBlock.scala 521:22]
  assign dispatch2_1_io_enqLsq_resp_2_lqIdx_flag = lsqCtrl_io_enq_resp_2_lqIdx_flag; // @[CtrlBlock.scala 521:22]
  assign dispatch2_1_io_enqLsq_resp_2_lqIdx_value = lsqCtrl_io_enq_resp_2_lqIdx_value; // @[CtrlBlock.scala 521:22]
  assign dispatch2_1_io_enqLsq_resp_2_sqIdx_flag = lsqCtrl_io_enq_resp_2_sqIdx_flag; // @[CtrlBlock.scala 521:22]
  assign dispatch2_1_io_enqLsq_resp_2_sqIdx_value = lsqCtrl_io_enq_resp_2_sqIdx_value; // @[CtrlBlock.scala 521:22]
  assign dispatch2_1_io_enqLsq_resp_3_lqIdx_flag = lsqCtrl_io_enq_resp_3_lqIdx_flag; // @[CtrlBlock.scala 521:22]
  assign dispatch2_1_io_enqLsq_resp_3_lqIdx_value = lsqCtrl_io_enq_resp_3_lqIdx_value; // @[CtrlBlock.scala 521:22]
  assign dispatch2_1_io_enqLsq_resp_3_sqIdx_flag = lsqCtrl_io_enq_resp_3_sqIdx_flag; // @[CtrlBlock.scala 521:22]
  assign dispatch2_1_io_enqLsq_resp_3_sqIdx_value = lsqCtrl_io_enq_resp_3_sqIdx_value; // @[CtrlBlock.scala 521:22]
  assign dispatch2_2_io_out_0_ready = io_rsReady_8; // @[CtrlBlock.scala 536:18]
  assign decode_clock = clock;
  assign decode_io_in_0_valid = io_frontend_cfVec_0_valid; // @[CtrlBlock.scala 402:16]
  assign decode_io_in_0_bits_instr = io_frontend_cfVec_0_bits_instr; // @[CtrlBlock.scala 402:16]
  assign decode_io_in_0_bits_foldpc = io_frontend_cfVec_0_bits_foldpc; // @[CtrlBlock.scala 402:16]
  assign decode_io_in_0_bits_exceptionVec_1 = io_frontend_cfVec_0_bits_exceptionVec_1; // @[CtrlBlock.scala 402:16]
  assign decode_io_in_0_bits_exceptionVec_12 = io_frontend_cfVec_0_bits_exceptionVec_12; // @[CtrlBlock.scala 402:16]
  assign decode_io_in_0_bits_trigger_frontendHit_0 = io_frontend_cfVec_0_bits_trigger_frontendHit_0; // @[CtrlBlock.scala 402:16]
  assign decode_io_in_0_bits_trigger_frontendHit_1 = io_frontend_cfVec_0_bits_trigger_frontendHit_1; // @[CtrlBlock.scala 402:16]
  assign decode_io_in_0_bits_trigger_frontendHit_2 = io_frontend_cfVec_0_bits_trigger_frontendHit_2; // @[CtrlBlock.scala 402:16]
  assign decode_io_in_0_bits_trigger_frontendHit_3 = io_frontend_cfVec_0_bits_trigger_frontendHit_3; // @[CtrlBlock.scala 402:16]
  assign decode_io_in_0_bits_trigger_backendEn_0 = io_frontend_cfVec_0_bits_trigger_backendEn_0; // @[CtrlBlock.scala 402:16]
  assign decode_io_in_0_bits_trigger_backendEn_1 = io_frontend_cfVec_0_bits_trigger_backendEn_1; // @[CtrlBlock.scala 402:16]
  assign decode_io_in_0_bits_pd_isRVC = io_frontend_cfVec_0_bits_pd_isRVC; // @[CtrlBlock.scala 402:16]
  assign decode_io_in_0_bits_pd_brType = io_frontend_cfVec_0_bits_pd_brType; // @[CtrlBlock.scala 402:16]
  assign decode_io_in_0_bits_pd_isCall = io_frontend_cfVec_0_bits_pd_isCall; // @[CtrlBlock.scala 402:16]
  assign decode_io_in_0_bits_pd_isRet = io_frontend_cfVec_0_bits_pd_isRet; // @[CtrlBlock.scala 402:16]
  assign decode_io_in_0_bits_pred_taken = io_frontend_cfVec_0_bits_pred_taken; // @[CtrlBlock.scala 402:16]
  assign decode_io_in_0_bits_crossPageIPFFix = io_frontend_cfVec_0_bits_crossPageIPFFix; // @[CtrlBlock.scala 402:16]
  assign decode_io_in_0_bits_ftqPtr_flag = io_frontend_cfVec_0_bits_ftqPtr_flag; // @[CtrlBlock.scala 402:16]
  assign decode_io_in_0_bits_ftqPtr_value = io_frontend_cfVec_0_bits_ftqPtr_value; // @[CtrlBlock.scala 402:16]
  assign decode_io_in_0_bits_ftqOffset = io_frontend_cfVec_0_bits_ftqOffset; // @[CtrlBlock.scala 402:16]
  assign decode_io_in_1_valid = io_frontend_cfVec_1_valid; // @[CtrlBlock.scala 402:16]
  assign decode_io_in_1_bits_instr = io_frontend_cfVec_1_bits_instr; // @[CtrlBlock.scala 402:16]
  assign decode_io_in_1_bits_foldpc = io_frontend_cfVec_1_bits_foldpc; // @[CtrlBlock.scala 402:16]
  assign decode_io_in_1_bits_exceptionVec_1 = io_frontend_cfVec_1_bits_exceptionVec_1; // @[CtrlBlock.scala 402:16]
  assign decode_io_in_1_bits_exceptionVec_12 = io_frontend_cfVec_1_bits_exceptionVec_12; // @[CtrlBlock.scala 402:16]
  assign decode_io_in_1_bits_trigger_frontendHit_0 = io_frontend_cfVec_1_bits_trigger_frontendHit_0; // @[CtrlBlock.scala 402:16]
  assign decode_io_in_1_bits_trigger_frontendHit_1 = io_frontend_cfVec_1_bits_trigger_frontendHit_1; // @[CtrlBlock.scala 402:16]
  assign decode_io_in_1_bits_trigger_frontendHit_2 = io_frontend_cfVec_1_bits_trigger_frontendHit_2; // @[CtrlBlock.scala 402:16]
  assign decode_io_in_1_bits_trigger_frontendHit_3 = io_frontend_cfVec_1_bits_trigger_frontendHit_3; // @[CtrlBlock.scala 402:16]
  assign decode_io_in_1_bits_trigger_backendEn_0 = io_frontend_cfVec_1_bits_trigger_backendEn_0; // @[CtrlBlock.scala 402:16]
  assign decode_io_in_1_bits_trigger_backendEn_1 = io_frontend_cfVec_1_bits_trigger_backendEn_1; // @[CtrlBlock.scala 402:16]
  assign decode_io_in_1_bits_pd_isRVC = io_frontend_cfVec_1_bits_pd_isRVC; // @[CtrlBlock.scala 402:16]
  assign decode_io_in_1_bits_pd_brType = io_frontend_cfVec_1_bits_pd_brType; // @[CtrlBlock.scala 402:16]
  assign decode_io_in_1_bits_pd_isCall = io_frontend_cfVec_1_bits_pd_isCall; // @[CtrlBlock.scala 402:16]
  assign decode_io_in_1_bits_pd_isRet = io_frontend_cfVec_1_bits_pd_isRet; // @[CtrlBlock.scala 402:16]
  assign decode_io_in_1_bits_pred_taken = io_frontend_cfVec_1_bits_pred_taken; // @[CtrlBlock.scala 402:16]
  assign decode_io_in_1_bits_crossPageIPFFix = io_frontend_cfVec_1_bits_crossPageIPFFix; // @[CtrlBlock.scala 402:16]
  assign decode_io_in_1_bits_ftqPtr_flag = io_frontend_cfVec_1_bits_ftqPtr_flag; // @[CtrlBlock.scala 402:16]
  assign decode_io_in_1_bits_ftqPtr_value = io_frontend_cfVec_1_bits_ftqPtr_value; // @[CtrlBlock.scala 402:16]
  assign decode_io_in_1_bits_ftqOffset = io_frontend_cfVec_1_bits_ftqOffset; // @[CtrlBlock.scala 402:16]
  assign decode_io_out_0_ready = rename_io_in_0_ready; // @[PipelineConnect.scala 182:21 CtrlBlock.scala 452:22]
  assign decode_io_out_1_ready = rename_io_in_1_ready; // @[PipelineConnect.scala 182:21 CtrlBlock.scala 452:22]
  assign decode_io_csrCtrl_fusion_enable = decode_io_csrCtrl_REG_fusion_enable; // @[CtrlBlock.scala 403:21]
  assign decode_io_csrCtrl_wfi_enable = decode_io_csrCtrl_REG_wfi_enable; // @[CtrlBlock.scala 403:21]
  assign decode_io_csrCtrl_svinval_enable = decode_io_csrCtrl_REG_svinval_enable; // @[CtrlBlock.scala 403:21]
  assign decode_io_csrCtrl_singlestep = decode_io_csrCtrl_REG_singlestep; // @[CtrlBlock.scala 403:21]
  assign decode_io_fusion_0 = fusionDecoder_io_out_0_valid & _decode_io_fusion_0_T; // @[CtrlBlock.scala 465:60]
  assign fusionDecoder_clock = clock;
  assign fusionDecoder_reset = reset;
  assign fusionDecoder_io_in_0_valid = io_frontend_cfVec_0_valid & ~(decodeHasException | disableFusion); // @[CtrlBlock.scala 443:64]
  assign fusionDecoder_io_in_0_bits = io_frontend_cfVec_0_bits_instr; // @[CtrlBlock.scala 444:33]
  assign fusionDecoder_io_in_1_valid = io_frontend_cfVec_1_valid & ~(decodeHasException_1 | disableFusion); // @[CtrlBlock.scala 443:64]
  assign fusionDecoder_io_in_1_bits = io_frontend_cfVec_1_bits_instr; // @[CtrlBlock.scala 444:33]
  assign fusionDecoder_io_inReady_0 = decode_io_out_1_ready; // @[CtrlBlock.scala 446:39]
  assign fusionDecoder_io_dec_0_fuOpType = renamePipe_data_ctrl_fuOpType; // @[PipelineConnect.scala 116:16 182:21]
  assign rat_clock = clock;
  assign rat_reset = reset;
  assign rat_io_redirect = flushRedirect_valid_REG ? flushRedirect_valid_REG : redirectGen_io_stage2Redirect_valid; // @[CtrlBlock.scala 302:27]
  assign rat_io_robCommits_isCommit = rob_io_commits_isCommit; // @[CtrlBlock.scala 432:21]
  assign rat_io_robCommits_commitValid_0 = rob_io_commits_commitValid_0; // @[CtrlBlock.scala 432:21]
  assign rat_io_robCommits_commitValid_1 = rob_io_commits_commitValid_1; // @[CtrlBlock.scala 432:21]
  assign rat_io_robCommits_isWalk = rob_io_commits_isWalk; // @[CtrlBlock.scala 432:21]
  assign rat_io_robCommits_walkValid_0 = rob_io_commits_walkValid_0; // @[CtrlBlock.scala 432:21]
  assign rat_io_robCommits_walkValid_1 = rob_io_commits_walkValid_1; // @[CtrlBlock.scala 432:21]
  assign rat_io_robCommits_info_0_ldest = rob_io_commits_info_0_ldest; // @[CtrlBlock.scala 432:21]
  assign rat_io_robCommits_info_0_rfWen = rob_io_commits_info_0_rfWen; // @[CtrlBlock.scala 432:21]
  assign rat_io_robCommits_info_0_fpWen = rob_io_commits_info_0_fpWen; // @[CtrlBlock.scala 432:21]
  assign rat_io_robCommits_info_0_pdest = rob_io_commits_info_0_pdest; // @[CtrlBlock.scala 432:21]
  assign rat_io_robCommits_info_1_ldest = rob_io_commits_info_1_ldest; // @[CtrlBlock.scala 432:21]
  assign rat_io_robCommits_info_1_rfWen = rob_io_commits_info_1_rfWen; // @[CtrlBlock.scala 432:21]
  assign rat_io_robCommits_info_1_fpWen = rob_io_commits_info_1_fpWen; // @[CtrlBlock.scala 432:21]
  assign rat_io_robCommits_info_1_pdest = rob_io_commits_info_1_pdest; // @[CtrlBlock.scala 432:21]
  assign rat_io_intReadPorts_0_0_hold = decode_io_intRat_0_0_hold; // @[CtrlBlock.scala 404:20]
  assign rat_io_intReadPorts_0_0_addr = decode_io_intRat_0_0_addr; // @[CtrlBlock.scala 404:20]
  assign rat_io_intReadPorts_0_1_hold = decode_io_intRat_0_1_hold; // @[CtrlBlock.scala 404:20]
  assign rat_io_intReadPorts_0_1_addr = decode_io_intRat_0_1_addr; // @[CtrlBlock.scala 404:20]
  assign rat_io_intReadPorts_0_2_hold = decode_io_intRat_0_2_hold; // @[CtrlBlock.scala 404:20]
  assign rat_io_intReadPorts_0_2_addr = decode_io_intRat_0_2_addr; // @[CtrlBlock.scala 404:20]
  assign rat_io_intReadPorts_1_0_hold = decode_io_intRat_1_0_hold; // @[CtrlBlock.scala 404:20]
  assign rat_io_intReadPorts_1_0_addr = decode_io_intRat_1_0_addr; // @[CtrlBlock.scala 404:20]
  assign rat_io_intReadPorts_1_1_hold = decode_io_intRat_1_1_hold; // @[CtrlBlock.scala 404:20]
  assign rat_io_intReadPorts_1_1_addr = decode_io_intRat_1_1_addr; // @[CtrlBlock.scala 404:20]
  assign rat_io_intReadPorts_1_2_hold = decode_io_intRat_1_2_hold; // @[CtrlBlock.scala 404:20]
  assign rat_io_intReadPorts_1_2_addr = decode_io_intRat_1_2_addr; // @[CtrlBlock.scala 404:20]
  assign rat_io_intRenamePorts_0_wen = rename_io_intRenamePorts_0_wen; // @[CtrlBlock.scala 433:25]
  assign rat_io_intRenamePorts_0_addr = rename_io_intRenamePorts_0_addr; // @[CtrlBlock.scala 433:25]
  assign rat_io_intRenamePorts_0_data = rename_io_intRenamePorts_0_data; // @[CtrlBlock.scala 433:25]
  assign rat_io_intRenamePorts_1_wen = rename_io_intRenamePorts_1_wen; // @[CtrlBlock.scala 433:25]
  assign rat_io_intRenamePorts_1_addr = rename_io_intRenamePorts_1_addr; // @[CtrlBlock.scala 433:25]
  assign rat_io_intRenamePorts_1_data = rename_io_intRenamePorts_1_data; // @[CtrlBlock.scala 433:25]
  assign rat_io_fpReadPorts_0_0_hold = decode_io_fpRat_0_0_hold; // @[CtrlBlock.scala 405:19]
  assign rat_io_fpReadPorts_0_0_addr = decode_io_fpRat_0_0_addr; // @[CtrlBlock.scala 405:19]
  assign rat_io_fpReadPorts_0_1_hold = decode_io_fpRat_0_1_hold; // @[CtrlBlock.scala 405:19]
  assign rat_io_fpReadPorts_0_1_addr = decode_io_fpRat_0_1_addr; // @[CtrlBlock.scala 405:19]
  assign rat_io_fpReadPorts_0_2_hold = decode_io_fpRat_0_2_hold; // @[CtrlBlock.scala 405:19]
  assign rat_io_fpReadPorts_0_2_addr = decode_io_fpRat_0_2_addr; // @[CtrlBlock.scala 405:19]
  assign rat_io_fpReadPorts_0_3_hold = decode_io_fpRat_0_3_hold; // @[CtrlBlock.scala 405:19]
  assign rat_io_fpReadPorts_0_3_addr = decode_io_fpRat_0_3_addr; // @[CtrlBlock.scala 405:19]
  assign rat_io_fpReadPorts_1_0_hold = decode_io_fpRat_1_0_hold; // @[CtrlBlock.scala 405:19]
  assign rat_io_fpReadPorts_1_0_addr = decode_io_fpRat_1_0_addr; // @[CtrlBlock.scala 405:19]
  assign rat_io_fpReadPorts_1_1_hold = decode_io_fpRat_1_1_hold; // @[CtrlBlock.scala 405:19]
  assign rat_io_fpReadPorts_1_1_addr = decode_io_fpRat_1_1_addr; // @[CtrlBlock.scala 405:19]
  assign rat_io_fpReadPorts_1_2_hold = decode_io_fpRat_1_2_hold; // @[CtrlBlock.scala 405:19]
  assign rat_io_fpReadPorts_1_2_addr = decode_io_fpRat_1_2_addr; // @[CtrlBlock.scala 405:19]
  assign rat_io_fpReadPorts_1_3_hold = decode_io_fpRat_1_3_hold; // @[CtrlBlock.scala 405:19]
  assign rat_io_fpReadPorts_1_3_addr = decode_io_fpRat_1_3_addr; // @[CtrlBlock.scala 405:19]
  assign rat_io_fpRenamePorts_0_wen = rename_io_fpRenamePorts_0_wen; // @[CtrlBlock.scala 434:24]
  assign rat_io_fpRenamePorts_0_addr = rename_io_fpRenamePorts_0_addr; // @[CtrlBlock.scala 434:24]
  assign rat_io_fpRenamePorts_0_data = rename_io_fpRenamePorts_0_data; // @[CtrlBlock.scala 434:24]
  assign rat_io_fpRenamePorts_1_wen = rename_io_fpRenamePorts_1_wen; // @[CtrlBlock.scala 434:24]
  assign rat_io_fpRenamePorts_1_addr = rename_io_fpRenamePorts_1_addr; // @[CtrlBlock.scala 434:24]
  assign rat_io_fpRenamePorts_1_data = rename_io_fpRenamePorts_1_data; // @[CtrlBlock.scala 434:24]
  assign ssit_clock = clock;
  assign ssit_reset = reset;
  assign ssit_io_raddr_0 = _mdp_foldpc_T ? decode_io_in_0_bits_foldpc : rename_io_in_0_bits_cf_foldpc; // @[CtrlBlock.scala 410:25]
  assign ssit_io_raddr_1 = _mdp_foldpc_T_1 ? decode_io_in_1_bits_foldpc : rename_io_in_1_bits_cf_foldpc; // @[CtrlBlock.scala 410:25]
  assign ssit_io_update_valid = ssit_io_update_REG_valid; // @[CtrlBlock.scala 419:18]
  assign ssit_io_update_ldpc = ssit_io_update_REG_ldpc; // @[CtrlBlock.scala 419:18]
  assign ssit_io_update_stpc = ssit_io_update_REG_stpc; // @[CtrlBlock.scala 419:18]
  assign ssit_io_csrCtrl_lvpred_timeout = ssit_io_csrCtrl_REG_lvpred_timeout; // @[CtrlBlock.scala 420:19]
  assign rename_clock = clock;
  assign rename_reset = reset;
  assign rename_io_redirect_valid = flushRedirect_valid_REG ? flushRedirect_valid_REG :
    redirectGen_io_stage2Redirect_valid; // @[CtrlBlock.scala 302:27]
  assign rename_io_redirect_bits_robIdx_flag = flushRedirect_valid_REG ? flushRedirect_bits_rrobIdx_flag :
    redirectGen_io_stage2Redirect_bits_robIdx_flag; // @[CtrlBlock.scala 302:27]
  assign rename_io_redirect_bits_robIdx_value = flushRedirect_valid_REG ? flushRedirect_bits_rrobIdx_value :
    redirectGen_io_stage2Redirect_bits_robIdx_value; // @[CtrlBlock.scala 302:27]
  assign rename_io_redirect_bits_level = flushRedirect_valid_REG ? flushRedirect_bits_rlevel :
    redirectGen_io_stage2Redirect_bits_level; // @[CtrlBlock.scala 302:27]
  assign rename_io_robCommits_isCommit = rob_io_commits_isCommit; // @[CtrlBlock.scala 484:24]
  assign rename_io_robCommits_commitValid_0 = rob_io_commits_commitValid_0; // @[CtrlBlock.scala 484:24]
  assign rename_io_robCommits_commitValid_1 = rob_io_commits_commitValid_1; // @[CtrlBlock.scala 484:24]
  assign rename_io_robCommits_isWalk = rob_io_commits_isWalk; // @[CtrlBlock.scala 484:24]
  assign rename_io_robCommits_walkValid_0 = rob_io_commits_walkValid_0; // @[CtrlBlock.scala 484:24]
  assign rename_io_robCommits_walkValid_1 = rob_io_commits_walkValid_1; // @[CtrlBlock.scala 484:24]
  assign rename_io_robCommits_info_0_ldest = rob_io_commits_info_0_ldest; // @[CtrlBlock.scala 484:24]
  assign rename_io_robCommits_info_0_rfWen = rob_io_commits_info_0_rfWen; // @[CtrlBlock.scala 484:24]
  assign rename_io_robCommits_info_0_fpWen = rob_io_commits_info_0_fpWen; // @[CtrlBlock.scala 484:24]
  assign rename_io_robCommits_info_0_pdest = rob_io_commits_info_0_pdest; // @[CtrlBlock.scala 484:24]
  assign rename_io_robCommits_info_0_old_pdest = rob_io_commits_info_0_old_pdest; // @[CtrlBlock.scala 484:24]
  assign rename_io_robCommits_info_0_isMove = rob_io_commits_info_0_isMove; // @[CtrlBlock.scala 484:24]
  assign rename_io_robCommits_info_1_ldest = rob_io_commits_info_1_ldest; // @[CtrlBlock.scala 484:24]
  assign rename_io_robCommits_info_1_rfWen = rob_io_commits_info_1_rfWen; // @[CtrlBlock.scala 484:24]
  assign rename_io_robCommits_info_1_fpWen = rob_io_commits_info_1_fpWen; // @[CtrlBlock.scala 484:24]
  assign rename_io_robCommits_info_1_pdest = rob_io_commits_info_1_pdest; // @[CtrlBlock.scala 484:24]
  assign rename_io_robCommits_info_1_old_pdest = rob_io_commits_info_1_old_pdest; // @[CtrlBlock.scala 484:24]
  assign rename_io_robCommits_info_1_isMove = rob_io_commits_info_1_isMove; // @[CtrlBlock.scala 484:24]
  assign rename_io_in_0_valid = renamePipe_valid; // @[CtrlBlock.scala 453:47]
  assign rename_io_in_0_bits_cf_foldpc = renamePipe_data_cf_foldpc; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_0_bits_cf_exceptionVec_1 = renamePipe_data_cf_exceptionVec_1; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_0_bits_cf_exceptionVec_2 = renamePipe_data_cf_exceptionVec_2; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_0_bits_cf_exceptionVec_12 = renamePipe_data_cf_exceptionVec_12; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_0_bits_cf_trigger_frontendHit_0 = renamePipe_data_cf_trigger_frontendHit_0; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_0_bits_cf_trigger_frontendHit_1 = renamePipe_data_cf_trigger_frontendHit_1; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_0_bits_cf_trigger_frontendHit_2 = renamePipe_data_cf_trigger_frontendHit_2; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_0_bits_cf_trigger_frontendHit_3 = renamePipe_data_cf_trigger_frontendHit_3; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_0_bits_cf_trigger_backendEn_0 = renamePipe_data_cf_trigger_backendEn_0; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_0_bits_cf_trigger_backendEn_1 = renamePipe_data_cf_trigger_backendEn_1; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_0_bits_cf_pd_isRVC = renamePipe_data_cf_pd_isRVC; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_0_bits_cf_pd_brType = renamePipe_data_cf_pd_brType; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_0_bits_cf_pd_isCall = renamePipe_data_cf_pd_isCall; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_0_bits_cf_pd_isRet = renamePipe_data_cf_pd_isRet; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_0_bits_cf_pred_taken = renamePipe_data_cf_pred_taken; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_0_bits_cf_crossPageIPFFix = renamePipe_data_cf_crossPageIPFFix; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_0_bits_cf_ftqPtr_flag = renamePipe_data_cf_ftqPtr_flag; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_0_bits_cf_ftqPtr_value = renamePipe_data_cf_ftqPtr_value; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_0_bits_cf_ftqOffset = renamePipe_data_cf_ftqOffset; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_0_bits_ctrl_srcType_0 = renamePipe_data_ctrl_srcType_0; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_0_bits_ctrl_srcType_1 = fusionDecoder_io_out_0_valid ? _GEN_1088 : renamePipe_data_ctrl_srcType_1; // @[CtrlBlock.scala 454:26 466:44]
  assign rename_io_in_0_bits_ctrl_srcType_2 = renamePipe_data_ctrl_srcType_2; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_0_bits_ctrl_lsrc_0 = renamePipe_data_ctrl_lsrc_0; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_0_bits_ctrl_lsrc_1 = fusionDecoder_io_out_0_valid ? _GEN_1087 : renamePipe_data_ctrl_lsrc_1; // @[CtrlBlock.scala 454:26 466:44]
  assign rename_io_in_0_bits_ctrl_ldest = renamePipe_data_ctrl_ldest; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_0_bits_ctrl_fuType = fusionDecoder_io_out_0_valid ? _GEN_1085 : renamePipe_data_ctrl_fuType; // @[CtrlBlock.scala 454:26 466:44]
  assign rename_io_in_0_bits_ctrl_fuOpType = fusionDecoder_io_out_0_valid ? _GEN_1086 : renamePipe_data_ctrl_fuOpType; // @[CtrlBlock.scala 454:26 466:44]
  assign rename_io_in_0_bits_ctrl_rfWen = renamePipe_data_ctrl_rfWen; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_0_bits_ctrl_fpWen = renamePipe_data_ctrl_fpWen; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_0_bits_ctrl_isXSTrap = renamePipe_data_ctrl_isXSTrap; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_0_bits_ctrl_noSpecExec = renamePipe_data_ctrl_noSpecExec; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_0_bits_ctrl_blockBackward = renamePipe_data_ctrl_blockBackward; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_0_bits_ctrl_flushPipe = renamePipe_data_ctrl_flushPipe; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_0_bits_ctrl_selImm = renamePipe_data_ctrl_selImm; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_0_bits_ctrl_imm = renamePipe_data_ctrl_imm; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_0_bits_ctrl_commitType = fusionDecoder_io_out_0_valid ? _rename_io_in_0_bits_ctrl_commitType_T_2
     : 3'h0; // @[CtrlBlock.scala 454:26 466:44 477:46]
  assign rename_io_in_0_bits_ctrl_fpu_isAddSub = renamePipe_data_ctrl_fpu_isAddSub; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_0_bits_ctrl_fpu_typeTagIn = renamePipe_data_ctrl_fpu_typeTagIn; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_0_bits_ctrl_fpu_typeTagOut = renamePipe_data_ctrl_fpu_typeTagOut; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_0_bits_ctrl_fpu_fromInt = renamePipe_data_ctrl_fpu_fromInt; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_0_bits_ctrl_fpu_wflags = renamePipe_data_ctrl_fpu_wflags; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_0_bits_ctrl_fpu_fpWen = renamePipe_data_ctrl_fpu_fpWen; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_0_bits_ctrl_fpu_fmaCmd = renamePipe_data_ctrl_fpu_fmaCmd; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_0_bits_ctrl_fpu_div = renamePipe_data_ctrl_fpu_div; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_0_bits_ctrl_fpu_sqrt = renamePipe_data_ctrl_fpu_sqrt; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_0_bits_ctrl_fpu_fcvt = renamePipe_data_ctrl_fpu_fcvt; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_0_bits_ctrl_fpu_typ = renamePipe_data_ctrl_fpu_typ; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_0_bits_ctrl_fpu_fmt = renamePipe_data_ctrl_fpu_fmt; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_0_bits_ctrl_fpu_ren3 = renamePipe_data_ctrl_fpu_ren3; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_0_bits_ctrl_fpu_rm = renamePipe_data_ctrl_fpu_rm; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_0_bits_ctrl_isMove = renamePipe_data_ctrl_isMove; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_1_valid = renamePipe_valid_1 & ~fusionDecoder_io_clear_1; // @[CtrlBlock.scala 453:47]
  assign rename_io_in_1_bits_cf_foldpc = renamePipe_data_1_cf_foldpc; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_1_bits_cf_exceptionVec_1 = renamePipe_data_1_cf_exceptionVec_1; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_1_bits_cf_exceptionVec_2 = renamePipe_data_1_cf_exceptionVec_2; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_1_bits_cf_exceptionVec_12 = renamePipe_data_1_cf_exceptionVec_12; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_1_bits_cf_trigger_frontendHit_0 = renamePipe_data_1_cf_trigger_frontendHit_0; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_1_bits_cf_trigger_frontendHit_1 = renamePipe_data_1_cf_trigger_frontendHit_1; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_1_bits_cf_trigger_frontendHit_2 = renamePipe_data_1_cf_trigger_frontendHit_2; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_1_bits_cf_trigger_frontendHit_3 = renamePipe_data_1_cf_trigger_frontendHit_3; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_1_bits_cf_trigger_backendEn_0 = renamePipe_data_1_cf_trigger_backendEn_0; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_1_bits_cf_trigger_backendEn_1 = renamePipe_data_1_cf_trigger_backendEn_1; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_1_bits_cf_pd_isRVC = renamePipe_data_1_cf_pd_isRVC; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_1_bits_cf_pd_brType = renamePipe_data_1_cf_pd_brType; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_1_bits_cf_pd_isCall = renamePipe_data_1_cf_pd_isCall; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_1_bits_cf_pd_isRet = renamePipe_data_1_cf_pd_isRet; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_1_bits_cf_pred_taken = renamePipe_data_1_cf_pred_taken; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_1_bits_cf_crossPageIPFFix = renamePipe_data_1_cf_crossPageIPFFix; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_1_bits_cf_ftqPtr_flag = renamePipe_data_1_cf_ftqPtr_flag; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_1_bits_cf_ftqPtr_value = renamePipe_data_1_cf_ftqPtr_value; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_1_bits_cf_ftqOffset = renamePipe_data_1_cf_ftqOffset; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_1_bits_ctrl_srcType_0 = renamePipe_data_1_ctrl_srcType_0; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_1_bits_ctrl_srcType_1 = renamePipe_data_1_ctrl_srcType_1; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_1_bits_ctrl_srcType_2 = renamePipe_data_1_ctrl_srcType_2; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_1_bits_ctrl_lsrc_0 = renamePipe_data_1_ctrl_lsrc_0; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_1_bits_ctrl_lsrc_1 = renamePipe_data_1_ctrl_lsrc_1; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_1_bits_ctrl_lsrc_2 = renamePipe_data_1_ctrl_lsrc_2; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_1_bits_ctrl_ldest = renamePipe_data_1_ctrl_ldest; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_1_bits_ctrl_fuType = renamePipe_data_1_ctrl_fuType; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_1_bits_ctrl_fuOpType = renamePipe_data_1_ctrl_fuOpType; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_1_bits_ctrl_rfWen = renamePipe_data_1_ctrl_rfWen; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_1_bits_ctrl_fpWen = renamePipe_data_1_ctrl_fpWen; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_1_bits_ctrl_isXSTrap = renamePipe_data_1_ctrl_isXSTrap; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_1_bits_ctrl_noSpecExec = renamePipe_data_1_ctrl_noSpecExec; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_1_bits_ctrl_blockBackward = renamePipe_data_1_ctrl_blockBackward; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_1_bits_ctrl_flushPipe = renamePipe_data_1_ctrl_flushPipe; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_1_bits_ctrl_selImm = renamePipe_data_1_ctrl_selImm; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_1_bits_ctrl_imm = renamePipe_data_1_ctrl_imm; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_1_bits_ctrl_fpu_isAddSub = renamePipe_data_1_ctrl_fpu_isAddSub; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_1_bits_ctrl_fpu_typeTagIn = renamePipe_data_1_ctrl_fpu_typeTagIn; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_1_bits_ctrl_fpu_typeTagOut = renamePipe_data_1_ctrl_fpu_typeTagOut; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_1_bits_ctrl_fpu_fromInt = renamePipe_data_1_ctrl_fpu_fromInt; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_1_bits_ctrl_fpu_wflags = renamePipe_data_1_ctrl_fpu_wflags; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_1_bits_ctrl_fpu_fpWen = renamePipe_data_1_ctrl_fpu_fpWen; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_1_bits_ctrl_fpu_fmaCmd = renamePipe_data_1_ctrl_fpu_fmaCmd; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_1_bits_ctrl_fpu_div = renamePipe_data_1_ctrl_fpu_div; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_1_bits_ctrl_fpu_sqrt = renamePipe_data_1_ctrl_fpu_sqrt; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_1_bits_ctrl_fpu_fcvt = renamePipe_data_1_ctrl_fpu_fcvt; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_1_bits_ctrl_fpu_typ = renamePipe_data_1_ctrl_fpu_typ; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_1_bits_ctrl_fpu_fmt = renamePipe_data_1_ctrl_fpu_fmt; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_1_bits_ctrl_fpu_ren3 = renamePipe_data_1_ctrl_fpu_ren3; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_1_bits_ctrl_fpu_rm = renamePipe_data_1_ctrl_fpu_rm; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_in_1_bits_ctrl_isMove = renamePipe_data_1_ctrl_isMove; // @[PipelineConnect.scala 116:16 182:21]
  assign rename_io_fusionInfo_0_rs2FromRs1 = fusionDecoder_io_info_0_rs2FromRs1; // @[CtrlBlock.scala 462:31]
  assign rename_io_fusionInfo_0_rs2FromRs2 = fusionDecoder_io_info_0_rs2FromRs2; // @[CtrlBlock.scala 462:31]
  assign rename_io_fusionInfo_0_rs2FromZero = fusionDecoder_io_info_0_rs2FromZero; // @[CtrlBlock.scala 462:31]
  assign rename_io_ssit_0_valid = ssit_io_rdata_0_valid; // @[CtrlBlock.scala 485:18]
  assign rename_io_ssit_0_ssid = ssit_io_rdata_0_ssid; // @[CtrlBlock.scala 485:18]
  assign rename_io_ssit_0_strict = ssit_io_rdata_0_strict; // @[CtrlBlock.scala 485:18]
  assign rename_io_ssit_1_valid = ssit_io_rdata_1_valid; // @[CtrlBlock.scala 485:18]
  assign rename_io_ssit_1_ssid = ssit_io_rdata_1_ssid; // @[CtrlBlock.scala 485:18]
  assign rename_io_ssit_1_strict = ssit_io_rdata_1_strict; // @[CtrlBlock.scala 485:18]
  assign rename_io_intReadPorts_0_0 = rat_io_intReadPorts_0_0_data; // @[CtrlBlock.scala 455:31]
  assign rename_io_intReadPorts_0_1 = rat_io_intReadPorts_0_1_data; // @[CtrlBlock.scala 455:31]
  assign rename_io_intReadPorts_0_2 = rat_io_intReadPorts_0_2_data; // @[CtrlBlock.scala 455:31]
  assign rename_io_intReadPorts_1_0 = rat_io_intReadPorts_1_0_data; // @[CtrlBlock.scala 455:31]
  assign rename_io_intReadPorts_1_1 = rat_io_intReadPorts_1_1_data; // @[CtrlBlock.scala 455:31]
  assign rename_io_intReadPorts_1_2 = rat_io_intReadPorts_1_2_data; // @[CtrlBlock.scala 455:31]
  assign rename_io_fpReadPorts_0_0 = rat_io_fpReadPorts_0_0_data; // @[CtrlBlock.scala 456:30]
  assign rename_io_fpReadPorts_0_1 = rat_io_fpReadPorts_0_1_data; // @[CtrlBlock.scala 456:30]
  assign rename_io_fpReadPorts_0_2 = rat_io_fpReadPorts_0_2_data; // @[CtrlBlock.scala 456:30]
  assign rename_io_fpReadPorts_0_3 = rat_io_fpReadPorts_0_3_data; // @[CtrlBlock.scala 456:30]
  assign rename_io_fpReadPorts_1_0 = rat_io_fpReadPorts_1_0_data; // @[CtrlBlock.scala 456:30]
  assign rename_io_fpReadPorts_1_1 = rat_io_fpReadPorts_1_1_data; // @[CtrlBlock.scala 456:30]
  assign rename_io_fpReadPorts_1_2 = rat_io_fpReadPorts_1_2_data; // @[CtrlBlock.scala 456:30]
  assign rename_io_fpReadPorts_1_3 = rat_io_fpReadPorts_1_3_data; // @[CtrlBlock.scala 456:30]
  assign rename_io_out_0_ready = dispatch_io_fromRename_0_ready; // @[PipelineConnect.scala 114:31]
  assign dispatch_clock = clock;
  assign dispatch_reset = reset;
  assign dispatch_io_fromRename_0_valid = valid; // @[PipelineConnect.scala 117:17]
  assign dispatch_io_fromRename_0_bits_cf_foldpc = data_cf_foldpc; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_0_bits_cf_exceptionVec_1 = data_cf_exceptionVec_1; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_0_bits_cf_exceptionVec_2 = data_cf_exceptionVec_2; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_0_bits_cf_exceptionVec_12 = data_cf_exceptionVec_12; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_0_bits_cf_trigger_frontendHit_0 = data_cf_trigger_frontendHit_0; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_0_bits_cf_trigger_frontendHit_1 = data_cf_trigger_frontendHit_1; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_0_bits_cf_trigger_frontendHit_2 = data_cf_trigger_frontendHit_2; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_0_bits_cf_trigger_frontendHit_3 = data_cf_trigger_frontendHit_3; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_0_bits_cf_trigger_backendEn_0 = data_cf_trigger_backendEn_0; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_0_bits_cf_trigger_backendEn_1 = data_cf_trigger_backendEn_1; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_0_bits_cf_pd_isRVC = data_cf_pd_isRVC; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_0_bits_cf_pd_brType = data_cf_pd_brType; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_0_bits_cf_pd_isCall = data_cf_pd_isCall; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_0_bits_cf_pd_isRet = data_cf_pd_isRet; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_0_bits_cf_pred_taken = data_cf_pred_taken; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_0_bits_cf_crossPageIPFFix = data_cf_crossPageIPFFix; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_0_bits_cf_storeSetHit = data_cf_storeSetHit; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_0_bits_cf_loadWaitStrict = data_cf_loadWaitStrict; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_0_bits_cf_ssid = data_cf_ssid; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_0_bits_cf_ftqPtr_flag = data_cf_ftqPtr_flag; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_0_bits_cf_ftqPtr_value = data_cf_ftqPtr_value; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_0_bits_cf_ftqOffset = data_cf_ftqOffset; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_0_bits_ctrl_srcType_0 = data_ctrl_srcType_0; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_0_bits_ctrl_srcType_1 = data_ctrl_srcType_1; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_0_bits_ctrl_srcType_2 = data_ctrl_srcType_2; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_0_bits_ctrl_ldest = data_ctrl_ldest; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_0_bits_ctrl_fuType = data_ctrl_fuType; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_0_bits_ctrl_fuOpType = data_ctrl_fuOpType; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_0_bits_ctrl_rfWen = data_ctrl_rfWen; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_0_bits_ctrl_fpWen = data_ctrl_fpWen; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_0_bits_ctrl_isXSTrap = data_ctrl_isXSTrap; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_0_bits_ctrl_noSpecExec = data_ctrl_noSpecExec; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_0_bits_ctrl_blockBackward = data_ctrl_blockBackward; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_0_bits_ctrl_flushPipe = data_ctrl_flushPipe; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_0_bits_ctrl_selImm = data_ctrl_selImm; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_0_bits_ctrl_imm = data_ctrl_imm; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_0_bits_ctrl_commitType = data_ctrl_commitType; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_0_bits_ctrl_fpu_isAddSub = data_ctrl_fpu_isAddSub; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_0_bits_ctrl_fpu_typeTagIn = data_ctrl_fpu_typeTagIn; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_0_bits_ctrl_fpu_typeTagOut = data_ctrl_fpu_typeTagOut; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_0_bits_ctrl_fpu_fromInt = data_ctrl_fpu_fromInt; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_0_bits_ctrl_fpu_wflags = data_ctrl_fpu_wflags; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_0_bits_ctrl_fpu_fpWen = data_ctrl_fpu_fpWen; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_0_bits_ctrl_fpu_fmaCmd = data_ctrl_fpu_fmaCmd; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_0_bits_ctrl_fpu_div = data_ctrl_fpu_div; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_0_bits_ctrl_fpu_sqrt = data_ctrl_fpu_sqrt; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_0_bits_ctrl_fpu_fcvt = data_ctrl_fpu_fcvt; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_0_bits_ctrl_fpu_typ = data_ctrl_fpu_typ; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_0_bits_ctrl_fpu_fmt = data_ctrl_fpu_fmt; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_0_bits_ctrl_fpu_ren3 = data_ctrl_fpu_ren3; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_0_bits_ctrl_fpu_rm = data_ctrl_fpu_rm; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_0_bits_ctrl_isMove = data_ctrl_isMove; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_0_bits_psrc_0 = data_psrc_0; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_0_bits_psrc_1 = data_psrc_1; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_0_bits_psrc_2 = data_psrc_2; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_0_bits_pdest = data_pdest; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_0_bits_old_pdest = data_old_pdest; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_0_bits_robIdx_flag = data_robIdx_flag; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_0_bits_robIdx_value = data_robIdx_value; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_0_bits_eliminatedMove = data_eliminatedMove; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_1_valid = valid_1; // @[PipelineConnect.scala 117:17]
  assign dispatch_io_fromRename_1_bits_cf_foldpc = data_1_cf_foldpc; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_1_bits_cf_exceptionVec_1 = data_1_cf_exceptionVec_1; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_1_bits_cf_exceptionVec_2 = data_1_cf_exceptionVec_2; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_1_bits_cf_exceptionVec_12 = data_1_cf_exceptionVec_12; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_1_bits_cf_trigger_frontendHit_0 = data_1_cf_trigger_frontendHit_0; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_1_bits_cf_trigger_frontendHit_1 = data_1_cf_trigger_frontendHit_1; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_1_bits_cf_trigger_frontendHit_2 = data_1_cf_trigger_frontendHit_2; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_1_bits_cf_trigger_frontendHit_3 = data_1_cf_trigger_frontendHit_3; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_1_bits_cf_trigger_backendEn_0 = data_1_cf_trigger_backendEn_0; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_1_bits_cf_trigger_backendEn_1 = data_1_cf_trigger_backendEn_1; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_1_bits_cf_pd_isRVC = data_1_cf_pd_isRVC; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_1_bits_cf_pd_brType = data_1_cf_pd_brType; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_1_bits_cf_pd_isCall = data_1_cf_pd_isCall; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_1_bits_cf_pd_isRet = data_1_cf_pd_isRet; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_1_bits_cf_pred_taken = data_1_cf_pred_taken; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_1_bits_cf_crossPageIPFFix = data_1_cf_crossPageIPFFix; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_1_bits_cf_storeSetHit = data_1_cf_storeSetHit; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_1_bits_cf_loadWaitStrict = data_1_cf_loadWaitStrict; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_1_bits_cf_ssid = data_1_cf_ssid; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_1_bits_cf_ftqPtr_flag = data_1_cf_ftqPtr_flag; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_1_bits_cf_ftqPtr_value = data_1_cf_ftqPtr_value; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_1_bits_cf_ftqOffset = data_1_cf_ftqOffset; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_1_bits_ctrl_srcType_0 = data_1_ctrl_srcType_0; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_1_bits_ctrl_srcType_1 = data_1_ctrl_srcType_1; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_1_bits_ctrl_srcType_2 = data_1_ctrl_srcType_2; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_1_bits_ctrl_ldest = data_1_ctrl_ldest; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_1_bits_ctrl_fuType = data_1_ctrl_fuType; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_1_bits_ctrl_fuOpType = data_1_ctrl_fuOpType; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_1_bits_ctrl_rfWen = data_1_ctrl_rfWen; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_1_bits_ctrl_fpWen = data_1_ctrl_fpWen; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_1_bits_ctrl_isXSTrap = data_1_ctrl_isXSTrap; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_1_bits_ctrl_noSpecExec = data_1_ctrl_noSpecExec; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_1_bits_ctrl_blockBackward = data_1_ctrl_blockBackward; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_1_bits_ctrl_flushPipe = data_1_ctrl_flushPipe; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_1_bits_ctrl_selImm = data_1_ctrl_selImm; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_1_bits_ctrl_imm = data_1_ctrl_imm; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_1_bits_ctrl_fpu_isAddSub = data_1_ctrl_fpu_isAddSub; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_1_bits_ctrl_fpu_typeTagIn = data_1_ctrl_fpu_typeTagIn; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_1_bits_ctrl_fpu_typeTagOut = data_1_ctrl_fpu_typeTagOut; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_1_bits_ctrl_fpu_fromInt = data_1_ctrl_fpu_fromInt; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_1_bits_ctrl_fpu_wflags = data_1_ctrl_fpu_wflags; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_1_bits_ctrl_fpu_fpWen = data_1_ctrl_fpu_fpWen; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_1_bits_ctrl_fpu_fmaCmd = data_1_ctrl_fpu_fmaCmd; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_1_bits_ctrl_fpu_div = data_1_ctrl_fpu_div; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_1_bits_ctrl_fpu_sqrt = data_1_ctrl_fpu_sqrt; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_1_bits_ctrl_fpu_fcvt = data_1_ctrl_fpu_fcvt; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_1_bits_ctrl_fpu_typ = data_1_ctrl_fpu_typ; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_1_bits_ctrl_fpu_fmt = data_1_ctrl_fpu_fmt; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_1_bits_ctrl_fpu_ren3 = data_1_ctrl_fpu_ren3; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_1_bits_ctrl_fpu_rm = data_1_ctrl_fpu_rm; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_1_bits_ctrl_isMove = data_1_ctrl_isMove; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_1_bits_psrc_0 = data_1_psrc_0; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_1_bits_psrc_1 = data_1_psrc_1; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_1_bits_psrc_2 = data_1_psrc_2; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_1_bits_pdest = data_1_pdest; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_1_bits_old_pdest = data_1_old_pdest; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_1_bits_robIdx_flag = data_1_robIdx_flag; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_1_bits_robIdx_value = data_1_robIdx_value; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_fromRename_1_bits_eliminatedMove = data_1_eliminatedMove; // @[PipelineConnect.scala 116:16]
  assign dispatch_io_enqRob_canAccept = rob_io_enq_canAccept; // @[CtrlBlock.scala 496:22]
  assign dispatch_io_enqRob_isEmpty = rob_io_enq_isEmpty; // @[CtrlBlock.scala 496:22]
  assign dispatch_io_toIntDq_canAccept = intDq_io_enq_canAccept; // @[CtrlBlock.scala 497:23]
  assign dispatch_io_toFpDq_canAccept = fpDq_io_enq_canAccept; // @[CtrlBlock.scala 498:22]
  assign dispatch_io_toLsDq_canAccept = lsDq_io_enq_canAccept; // @[CtrlBlock.scala 499:22]
  assign dispatch_io_redirect_valid = flushRedirect_valid_REG ? flushRedirect_valid_REG :
    redirectGen_io_stage2Redirect_valid; // @[CtrlBlock.scala 302:27]
  assign dispatch_io_singleStep = dispatch_io_singleStep_REG; // @[CtrlBlock.scala 501:26]
  assign dispatch_io_lfst_resp_0_bits_shouldWait = lfst_io_dispatch_resp_0_bits_shouldWait; // @[CtrlBlock.scala 429:20]
  assign dispatch_io_lfst_resp_0_bits_robIdx_flag = lfst_io_dispatch_resp_0_bits_robIdx_flag; // @[CtrlBlock.scala 429:20]
  assign dispatch_io_lfst_resp_0_bits_robIdx_value = lfst_io_dispatch_resp_0_bits_robIdx_value; // @[CtrlBlock.scala 429:20]
  assign dispatch_io_lfst_resp_1_bits_shouldWait = lfst_io_dispatch_resp_1_bits_shouldWait; // @[CtrlBlock.scala 429:20]
  assign dispatch_io_lfst_resp_1_bits_robIdx_flag = lfst_io_dispatch_resp_1_bits_robIdx_flag; // @[CtrlBlock.scala 429:20]
  assign dispatch_io_lfst_resp_1_bits_robIdx_value = lfst_io_dispatch_resp_1_bits_robIdx_value; // @[CtrlBlock.scala 429:20]
  assign intDq_clock = clock;
  assign intDq_reset = reset;
  assign intDq_io_enq_needAlloc_0 = dispatch_io_toIntDq_needAlloc_0; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_needAlloc_1 = dispatch_io_toIntDq_needAlloc_1; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_0_valid = dispatch_io_toIntDq_req_0_valid; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_0_bits_cf_foldpc = dispatch_io_toIntDq_req_0_bits_cf_foldpc; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_0_bits_cf_trigger_backendEn_0 = dispatch_io_toIntDq_req_0_bits_cf_trigger_backendEn_0; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_0_bits_cf_trigger_backendEn_1 = dispatch_io_toIntDq_req_0_bits_cf_trigger_backendEn_1; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_0_bits_cf_pd_isRVC = dispatch_io_toIntDq_req_0_bits_cf_pd_isRVC; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_0_bits_cf_pd_brType = dispatch_io_toIntDq_req_0_bits_cf_pd_brType; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_0_bits_cf_pd_isCall = dispatch_io_toIntDq_req_0_bits_cf_pd_isCall; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_0_bits_cf_pd_isRet = dispatch_io_toIntDq_req_0_bits_cf_pd_isRet; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_0_bits_cf_pred_taken = dispatch_io_toIntDq_req_0_bits_cf_pred_taken; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_0_bits_cf_storeSetHit = dispatch_io_toIntDq_req_0_bits_cf_storeSetHit; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_0_bits_cf_waitForRobIdx_flag = dispatch_io_toIntDq_req_0_bits_cf_waitForRobIdx_flag; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_0_bits_cf_waitForRobIdx_value = dispatch_io_toIntDq_req_0_bits_cf_waitForRobIdx_value; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_0_bits_cf_loadWaitBit = dispatch_io_toIntDq_req_0_bits_cf_loadWaitBit; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_0_bits_cf_loadWaitStrict = dispatch_io_toIntDq_req_0_bits_cf_loadWaitStrict; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_0_bits_cf_ssid = dispatch_io_toIntDq_req_0_bits_cf_ssid; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_0_bits_cf_ftqPtr_flag = dispatch_io_toIntDq_req_0_bits_cf_ftqPtr_flag; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_0_bits_cf_ftqPtr_value = dispatch_io_toIntDq_req_0_bits_cf_ftqPtr_value; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_0_bits_cf_ftqOffset = dispatch_io_toIntDq_req_0_bits_cf_ftqOffset; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_0_bits_ctrl_srcType_0 = dispatch_io_toIntDq_req_0_bits_ctrl_srcType_0; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_0_bits_ctrl_srcType_1 = dispatch_io_toIntDq_req_0_bits_ctrl_srcType_1; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_0_bits_ctrl_srcType_2 = dispatch_io_toIntDq_req_0_bits_ctrl_srcType_2; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_0_bits_ctrl_fuType = dispatch_io_toIntDq_req_0_bits_ctrl_fuType; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_0_bits_ctrl_fuOpType = dispatch_io_toIntDq_req_0_bits_ctrl_fuOpType; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_0_bits_ctrl_rfWen = dispatch_io_toIntDq_req_0_bits_ctrl_rfWen; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_0_bits_ctrl_fpWen = dispatch_io_toIntDq_req_0_bits_ctrl_fpWen; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_0_bits_ctrl_flushPipe = dispatch_io_toIntDq_req_0_bits_ctrl_flushPipe; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_0_bits_ctrl_selImm = dispatch_io_toIntDq_req_0_bits_ctrl_selImm; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_0_bits_ctrl_imm = dispatch_io_toIntDq_req_0_bits_ctrl_imm; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_0_bits_ctrl_fpu_isAddSub = dispatch_io_toIntDq_req_0_bits_ctrl_fpu_isAddSub; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_0_bits_ctrl_fpu_typeTagIn = dispatch_io_toIntDq_req_0_bits_ctrl_fpu_typeTagIn; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_0_bits_ctrl_fpu_typeTagOut = dispatch_io_toIntDq_req_0_bits_ctrl_fpu_typeTagOut; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_0_bits_ctrl_fpu_fromInt = dispatch_io_toIntDq_req_0_bits_ctrl_fpu_fromInt; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_0_bits_ctrl_fpu_wflags = dispatch_io_toIntDq_req_0_bits_ctrl_fpu_wflags; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_0_bits_ctrl_fpu_fpWen = dispatch_io_toIntDq_req_0_bits_ctrl_fpu_fpWen; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_0_bits_ctrl_fpu_fmaCmd = dispatch_io_toIntDq_req_0_bits_ctrl_fpu_fmaCmd; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_0_bits_ctrl_fpu_div = dispatch_io_toIntDq_req_0_bits_ctrl_fpu_div; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_0_bits_ctrl_fpu_sqrt = dispatch_io_toIntDq_req_0_bits_ctrl_fpu_sqrt; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_0_bits_ctrl_fpu_fcvt = dispatch_io_toIntDq_req_0_bits_ctrl_fpu_fcvt; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_0_bits_ctrl_fpu_typ = dispatch_io_toIntDq_req_0_bits_ctrl_fpu_typ; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_0_bits_ctrl_fpu_fmt = dispatch_io_toIntDq_req_0_bits_ctrl_fpu_fmt; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_0_bits_ctrl_fpu_ren3 = dispatch_io_toIntDq_req_0_bits_ctrl_fpu_ren3; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_0_bits_ctrl_fpu_rm = dispatch_io_toIntDq_req_0_bits_ctrl_fpu_rm; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_0_bits_psrc_0 = dispatch_io_toIntDq_req_0_bits_psrc_0; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_0_bits_psrc_1 = dispatch_io_toIntDq_req_0_bits_psrc_1; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_0_bits_psrc_2 = dispatch_io_toIntDq_req_0_bits_psrc_2; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_0_bits_pdest = dispatch_io_toIntDq_req_0_bits_pdest; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_0_bits_robIdx_flag = dispatch_io_toIntDq_req_0_bits_robIdx_flag; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_0_bits_robIdx_value = dispatch_io_toIntDq_req_0_bits_robIdx_value; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_1_valid = dispatch_io_toIntDq_req_1_valid; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_1_bits_cf_foldpc = dispatch_io_toIntDq_req_1_bits_cf_foldpc; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_1_bits_cf_trigger_backendEn_0 = dispatch_io_toIntDq_req_1_bits_cf_trigger_backendEn_0; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_1_bits_cf_trigger_backendEn_1 = dispatch_io_toIntDq_req_1_bits_cf_trigger_backendEn_1; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_1_bits_cf_pd_isRVC = dispatch_io_toIntDq_req_1_bits_cf_pd_isRVC; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_1_bits_cf_pd_brType = dispatch_io_toIntDq_req_1_bits_cf_pd_brType; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_1_bits_cf_pd_isCall = dispatch_io_toIntDq_req_1_bits_cf_pd_isCall; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_1_bits_cf_pd_isRet = dispatch_io_toIntDq_req_1_bits_cf_pd_isRet; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_1_bits_cf_pred_taken = dispatch_io_toIntDq_req_1_bits_cf_pred_taken; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_1_bits_cf_storeSetHit = dispatch_io_toIntDq_req_1_bits_cf_storeSetHit; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_1_bits_cf_waitForRobIdx_flag = dispatch_io_toIntDq_req_1_bits_cf_waitForRobIdx_flag; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_1_bits_cf_waitForRobIdx_value = dispatch_io_toIntDq_req_1_bits_cf_waitForRobIdx_value; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_1_bits_cf_loadWaitBit = dispatch_io_toIntDq_req_1_bits_cf_loadWaitBit; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_1_bits_cf_loadWaitStrict = dispatch_io_toIntDq_req_1_bits_cf_loadWaitStrict; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_1_bits_cf_ssid = dispatch_io_toIntDq_req_1_bits_cf_ssid; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_1_bits_cf_ftqPtr_flag = dispatch_io_toIntDq_req_1_bits_cf_ftqPtr_flag; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_1_bits_cf_ftqPtr_value = dispatch_io_toIntDq_req_1_bits_cf_ftqPtr_value; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_1_bits_cf_ftqOffset = dispatch_io_toIntDq_req_1_bits_cf_ftqOffset; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_1_bits_ctrl_srcType_0 = dispatch_io_toIntDq_req_1_bits_ctrl_srcType_0; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_1_bits_ctrl_srcType_1 = dispatch_io_toIntDq_req_1_bits_ctrl_srcType_1; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_1_bits_ctrl_srcType_2 = dispatch_io_toIntDq_req_1_bits_ctrl_srcType_2; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_1_bits_ctrl_fuType = dispatch_io_toIntDq_req_1_bits_ctrl_fuType; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_1_bits_ctrl_fuOpType = dispatch_io_toIntDq_req_1_bits_ctrl_fuOpType; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_1_bits_ctrl_rfWen = dispatch_io_toIntDq_req_1_bits_ctrl_rfWen; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_1_bits_ctrl_fpWen = dispatch_io_toIntDq_req_1_bits_ctrl_fpWen; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_1_bits_ctrl_flushPipe = dispatch_io_toIntDq_req_1_bits_ctrl_flushPipe; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_1_bits_ctrl_selImm = dispatch_io_toIntDq_req_1_bits_ctrl_selImm; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_1_bits_ctrl_imm = dispatch_io_toIntDq_req_1_bits_ctrl_imm; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_1_bits_ctrl_fpu_isAddSub = dispatch_io_toIntDq_req_1_bits_ctrl_fpu_isAddSub; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_1_bits_ctrl_fpu_typeTagIn = dispatch_io_toIntDq_req_1_bits_ctrl_fpu_typeTagIn; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_1_bits_ctrl_fpu_typeTagOut = dispatch_io_toIntDq_req_1_bits_ctrl_fpu_typeTagOut; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_1_bits_ctrl_fpu_fromInt = dispatch_io_toIntDq_req_1_bits_ctrl_fpu_fromInt; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_1_bits_ctrl_fpu_wflags = dispatch_io_toIntDq_req_1_bits_ctrl_fpu_wflags; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_1_bits_ctrl_fpu_fpWen = dispatch_io_toIntDq_req_1_bits_ctrl_fpu_fpWen; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_1_bits_ctrl_fpu_fmaCmd = dispatch_io_toIntDq_req_1_bits_ctrl_fpu_fmaCmd; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_1_bits_ctrl_fpu_div = dispatch_io_toIntDq_req_1_bits_ctrl_fpu_div; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_1_bits_ctrl_fpu_sqrt = dispatch_io_toIntDq_req_1_bits_ctrl_fpu_sqrt; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_1_bits_ctrl_fpu_fcvt = dispatch_io_toIntDq_req_1_bits_ctrl_fpu_fcvt; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_1_bits_ctrl_fpu_typ = dispatch_io_toIntDq_req_1_bits_ctrl_fpu_typ; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_1_bits_ctrl_fpu_fmt = dispatch_io_toIntDq_req_1_bits_ctrl_fpu_fmt; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_1_bits_ctrl_fpu_ren3 = dispatch_io_toIntDq_req_1_bits_ctrl_fpu_ren3; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_1_bits_ctrl_fpu_rm = dispatch_io_toIntDq_req_1_bits_ctrl_fpu_rm; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_1_bits_psrc_0 = dispatch_io_toIntDq_req_1_bits_psrc_0; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_1_bits_psrc_1 = dispatch_io_toIntDq_req_1_bits_psrc_1; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_1_bits_psrc_2 = dispatch_io_toIntDq_req_1_bits_psrc_2; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_1_bits_pdest = dispatch_io_toIntDq_req_1_bits_pdest; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_1_bits_robIdx_flag = dispatch_io_toIntDq_req_1_bits_robIdx_flag; // @[CtrlBlock.scala 497:23]
  assign intDq_io_enq_req_1_bits_robIdx_value = dispatch_io_toIntDq_req_1_bits_robIdx_value; // @[CtrlBlock.scala 497:23]
  assign intDq_io_deq_0_ready = dispatch2_io_in_0_ready; // @[CtrlBlock.scala 533:21]
  assign intDq_io_deq_1_ready = dispatch2_io_in_1_ready; // @[CtrlBlock.scala 533:21]
  assign intDq_io_deq_2_ready = 1'h0; // @[CtrlBlock.scala 533:21]
  assign intDq_io_deq_3_ready = 1'h0; // @[CtrlBlock.scala 533:21]
  assign intDq_io_redirect_valid = redirectForExu_next_valid_REG; // @[BitUtils.scala 26:20 28:18]
  assign intDq_io_redirect_bits_robIdx_flag = redirectForExu_next_bits_rrobIdx_flag; // @[BitUtils.scala 26:20 33:15]
  assign intDq_io_redirect_bits_robIdx_value = redirectForExu_next_bits_rrobIdx_value; // @[BitUtils.scala 26:20 33:15]
  assign intDq_io_redirect_bits_level = redirectForExu_next_bits_rlevel; // @[BitUtils.scala 26:20 33:15]
  assign fpDq_clock = clock;
  assign fpDq_reset = reset;
  assign fpDq_io_enq_needAlloc_0 = dispatch_io_toFpDq_needAlloc_0; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_needAlloc_1 = dispatch_io_toFpDq_needAlloc_1; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_0_valid = dispatch_io_toFpDq_req_0_valid; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_0_bits_cf_foldpc = dispatch_io_toFpDq_req_0_bits_cf_foldpc; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_0_bits_cf_trigger_backendEn_0 = dispatch_io_toFpDq_req_0_bits_cf_trigger_backendEn_0; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_0_bits_cf_trigger_backendEn_1 = dispatch_io_toFpDq_req_0_bits_cf_trigger_backendEn_1; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_0_bits_cf_pd_isRVC = dispatch_io_toFpDq_req_0_bits_cf_pd_isRVC; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_0_bits_cf_pd_brType = dispatch_io_toFpDq_req_0_bits_cf_pd_brType; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_0_bits_cf_pd_isCall = dispatch_io_toFpDq_req_0_bits_cf_pd_isCall; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_0_bits_cf_pd_isRet = dispatch_io_toFpDq_req_0_bits_cf_pd_isRet; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_0_bits_cf_pred_taken = dispatch_io_toFpDq_req_0_bits_cf_pred_taken; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_0_bits_cf_storeSetHit = dispatch_io_toFpDq_req_0_bits_cf_storeSetHit; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_0_bits_cf_waitForRobIdx_flag = dispatch_io_toFpDq_req_0_bits_cf_waitForRobIdx_flag; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_0_bits_cf_waitForRobIdx_value = dispatch_io_toFpDq_req_0_bits_cf_waitForRobIdx_value; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_0_bits_cf_loadWaitBit = dispatch_io_toFpDq_req_0_bits_cf_loadWaitBit; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_0_bits_cf_loadWaitStrict = dispatch_io_toFpDq_req_0_bits_cf_loadWaitStrict; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_0_bits_cf_ssid = dispatch_io_toFpDq_req_0_bits_cf_ssid; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_0_bits_cf_ftqPtr_flag = dispatch_io_toFpDq_req_0_bits_cf_ftqPtr_flag; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_0_bits_cf_ftqPtr_value = dispatch_io_toFpDq_req_0_bits_cf_ftqPtr_value; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_0_bits_cf_ftqOffset = dispatch_io_toFpDq_req_0_bits_cf_ftqOffset; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_0_bits_ctrl_srcType_0 = dispatch_io_toFpDq_req_0_bits_ctrl_srcType_0; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_0_bits_ctrl_srcType_1 = dispatch_io_toFpDq_req_0_bits_ctrl_srcType_1; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_0_bits_ctrl_srcType_2 = dispatch_io_toFpDq_req_0_bits_ctrl_srcType_2; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_0_bits_ctrl_fuType = dispatch_io_toFpDq_req_0_bits_ctrl_fuType; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_0_bits_ctrl_fuOpType = dispatch_io_toFpDq_req_0_bits_ctrl_fuOpType; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_0_bits_ctrl_rfWen = dispatch_io_toFpDq_req_0_bits_ctrl_rfWen; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_0_bits_ctrl_fpWen = dispatch_io_toFpDq_req_0_bits_ctrl_fpWen; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_0_bits_ctrl_flushPipe = dispatch_io_toFpDq_req_0_bits_ctrl_flushPipe; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_0_bits_ctrl_selImm = dispatch_io_toFpDq_req_0_bits_ctrl_selImm; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_0_bits_ctrl_imm = dispatch_io_toFpDq_req_0_bits_ctrl_imm; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_0_bits_ctrl_fpu_isAddSub = dispatch_io_toFpDq_req_0_bits_ctrl_fpu_isAddSub; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_0_bits_ctrl_fpu_typeTagIn = dispatch_io_toFpDq_req_0_bits_ctrl_fpu_typeTagIn; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_0_bits_ctrl_fpu_typeTagOut = dispatch_io_toFpDq_req_0_bits_ctrl_fpu_typeTagOut; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_0_bits_ctrl_fpu_fromInt = dispatch_io_toFpDq_req_0_bits_ctrl_fpu_fromInt; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_0_bits_ctrl_fpu_wflags = dispatch_io_toFpDq_req_0_bits_ctrl_fpu_wflags; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_0_bits_ctrl_fpu_fpWen = dispatch_io_toFpDq_req_0_bits_ctrl_fpu_fpWen; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_0_bits_ctrl_fpu_fmaCmd = dispatch_io_toFpDq_req_0_bits_ctrl_fpu_fmaCmd; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_0_bits_ctrl_fpu_div = dispatch_io_toFpDq_req_0_bits_ctrl_fpu_div; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_0_bits_ctrl_fpu_sqrt = dispatch_io_toFpDq_req_0_bits_ctrl_fpu_sqrt; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_0_bits_ctrl_fpu_fcvt = dispatch_io_toFpDq_req_0_bits_ctrl_fpu_fcvt; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_0_bits_ctrl_fpu_typ = dispatch_io_toFpDq_req_0_bits_ctrl_fpu_typ; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_0_bits_ctrl_fpu_fmt = dispatch_io_toFpDq_req_0_bits_ctrl_fpu_fmt; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_0_bits_ctrl_fpu_ren3 = dispatch_io_toFpDq_req_0_bits_ctrl_fpu_ren3; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_0_bits_ctrl_fpu_rm = dispatch_io_toFpDq_req_0_bits_ctrl_fpu_rm; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_0_bits_psrc_0 = dispatch_io_toFpDq_req_0_bits_psrc_0; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_0_bits_psrc_1 = dispatch_io_toFpDq_req_0_bits_psrc_1; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_0_bits_psrc_2 = dispatch_io_toFpDq_req_0_bits_psrc_2; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_0_bits_pdest = dispatch_io_toFpDq_req_0_bits_pdest; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_0_bits_robIdx_flag = dispatch_io_toFpDq_req_0_bits_robIdx_flag; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_0_bits_robIdx_value = dispatch_io_toFpDq_req_0_bits_robIdx_value; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_1_valid = dispatch_io_toFpDq_req_1_valid; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_1_bits_cf_foldpc = dispatch_io_toFpDq_req_1_bits_cf_foldpc; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_1_bits_cf_trigger_backendEn_0 = dispatch_io_toFpDq_req_1_bits_cf_trigger_backendEn_0; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_1_bits_cf_trigger_backendEn_1 = dispatch_io_toFpDq_req_1_bits_cf_trigger_backendEn_1; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_1_bits_cf_pd_isRVC = dispatch_io_toFpDq_req_1_bits_cf_pd_isRVC; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_1_bits_cf_pd_brType = dispatch_io_toFpDq_req_1_bits_cf_pd_brType; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_1_bits_cf_pd_isCall = dispatch_io_toFpDq_req_1_bits_cf_pd_isCall; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_1_bits_cf_pd_isRet = dispatch_io_toFpDq_req_1_bits_cf_pd_isRet; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_1_bits_cf_pred_taken = dispatch_io_toFpDq_req_1_bits_cf_pred_taken; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_1_bits_cf_storeSetHit = dispatch_io_toFpDq_req_1_bits_cf_storeSetHit; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_1_bits_cf_waitForRobIdx_flag = dispatch_io_toFpDq_req_1_bits_cf_waitForRobIdx_flag; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_1_bits_cf_waitForRobIdx_value = dispatch_io_toFpDq_req_1_bits_cf_waitForRobIdx_value; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_1_bits_cf_loadWaitBit = dispatch_io_toFpDq_req_1_bits_cf_loadWaitBit; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_1_bits_cf_loadWaitStrict = dispatch_io_toFpDq_req_1_bits_cf_loadWaitStrict; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_1_bits_cf_ssid = dispatch_io_toFpDq_req_1_bits_cf_ssid; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_1_bits_cf_ftqPtr_flag = dispatch_io_toFpDq_req_1_bits_cf_ftqPtr_flag; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_1_bits_cf_ftqPtr_value = dispatch_io_toFpDq_req_1_bits_cf_ftqPtr_value; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_1_bits_cf_ftqOffset = dispatch_io_toFpDq_req_1_bits_cf_ftqOffset; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_1_bits_ctrl_srcType_0 = dispatch_io_toFpDq_req_1_bits_ctrl_srcType_0; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_1_bits_ctrl_srcType_1 = dispatch_io_toFpDq_req_1_bits_ctrl_srcType_1; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_1_bits_ctrl_srcType_2 = dispatch_io_toFpDq_req_1_bits_ctrl_srcType_2; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_1_bits_ctrl_fuType = dispatch_io_toFpDq_req_1_bits_ctrl_fuType; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_1_bits_ctrl_fuOpType = dispatch_io_toFpDq_req_1_bits_ctrl_fuOpType; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_1_bits_ctrl_rfWen = dispatch_io_toFpDq_req_1_bits_ctrl_rfWen; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_1_bits_ctrl_fpWen = dispatch_io_toFpDq_req_1_bits_ctrl_fpWen; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_1_bits_ctrl_flushPipe = dispatch_io_toFpDq_req_1_bits_ctrl_flushPipe; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_1_bits_ctrl_selImm = dispatch_io_toFpDq_req_1_bits_ctrl_selImm; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_1_bits_ctrl_imm = dispatch_io_toFpDq_req_1_bits_ctrl_imm; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_1_bits_ctrl_fpu_isAddSub = dispatch_io_toFpDq_req_1_bits_ctrl_fpu_isAddSub; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_1_bits_ctrl_fpu_typeTagIn = dispatch_io_toFpDq_req_1_bits_ctrl_fpu_typeTagIn; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_1_bits_ctrl_fpu_typeTagOut = dispatch_io_toFpDq_req_1_bits_ctrl_fpu_typeTagOut; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_1_bits_ctrl_fpu_fromInt = dispatch_io_toFpDq_req_1_bits_ctrl_fpu_fromInt; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_1_bits_ctrl_fpu_wflags = dispatch_io_toFpDq_req_1_bits_ctrl_fpu_wflags; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_1_bits_ctrl_fpu_fpWen = dispatch_io_toFpDq_req_1_bits_ctrl_fpu_fpWen; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_1_bits_ctrl_fpu_fmaCmd = dispatch_io_toFpDq_req_1_bits_ctrl_fpu_fmaCmd; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_1_bits_ctrl_fpu_div = dispatch_io_toFpDq_req_1_bits_ctrl_fpu_div; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_1_bits_ctrl_fpu_sqrt = dispatch_io_toFpDq_req_1_bits_ctrl_fpu_sqrt; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_1_bits_ctrl_fpu_fcvt = dispatch_io_toFpDq_req_1_bits_ctrl_fpu_fcvt; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_1_bits_ctrl_fpu_typ = dispatch_io_toFpDq_req_1_bits_ctrl_fpu_typ; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_1_bits_ctrl_fpu_fmt = dispatch_io_toFpDq_req_1_bits_ctrl_fpu_fmt; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_1_bits_ctrl_fpu_ren3 = dispatch_io_toFpDq_req_1_bits_ctrl_fpu_ren3; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_1_bits_ctrl_fpu_rm = dispatch_io_toFpDq_req_1_bits_ctrl_fpu_rm; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_1_bits_psrc_0 = dispatch_io_toFpDq_req_1_bits_psrc_0; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_1_bits_psrc_1 = dispatch_io_toFpDq_req_1_bits_psrc_1; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_1_bits_psrc_2 = dispatch_io_toFpDq_req_1_bits_psrc_2; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_1_bits_pdest = dispatch_io_toFpDq_req_1_bits_pdest; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_1_bits_robIdx_flag = dispatch_io_toFpDq_req_1_bits_robIdx_flag; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_enq_req_1_bits_robIdx_value = dispatch_io_toFpDq_req_1_bits_robIdx_value; // @[CtrlBlock.scala 498:22]
  assign fpDq_io_deq_0_ready = dispatch2_2_io_in_0_ready; // @[CtrlBlock.scala 533:21]
  assign fpDq_io_deq_1_ready = 1'h0; // @[CtrlBlock.scala 533:21]
  assign fpDq_io_deq_2_ready = 1'h0; // @[CtrlBlock.scala 533:21]
  assign fpDq_io_deq_3_ready = 1'h0; // @[CtrlBlock.scala 533:21]
  assign fpDq_io_redirect_valid = redirectForExu_next_valid_REG; // @[BitUtils.scala 26:20 28:18]
  assign fpDq_io_redirect_bits_robIdx_flag = redirectForExu_next_bits_rrobIdx_flag; // @[BitUtils.scala 26:20 33:15]
  assign fpDq_io_redirect_bits_robIdx_value = redirectForExu_next_bits_rrobIdx_value; // @[BitUtils.scala 26:20 33:15]
  assign fpDq_io_redirect_bits_level = redirectForExu_next_bits_rlevel; // @[BitUtils.scala 26:20 33:15]
  assign lsDq_clock = clock;
  assign lsDq_reset = reset;
  assign lsDq_io_enq_needAlloc_0 = dispatch_io_toLsDq_needAlloc_0; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_needAlloc_1 = dispatch_io_toLsDq_needAlloc_1; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_0_valid = dispatch_io_toLsDq_req_0_valid; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_0_bits_cf_foldpc = dispatch_io_toLsDq_req_0_bits_cf_foldpc; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_0_bits_cf_trigger_backendEn_0 = dispatch_io_toLsDq_req_0_bits_cf_trigger_backendEn_0; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_0_bits_cf_trigger_backendEn_1 = dispatch_io_toLsDq_req_0_bits_cf_trigger_backendEn_1; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_0_bits_cf_pd_isRVC = dispatch_io_toLsDq_req_0_bits_cf_pd_isRVC; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_0_bits_cf_pd_brType = dispatch_io_toLsDq_req_0_bits_cf_pd_brType; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_0_bits_cf_pd_isCall = dispatch_io_toLsDq_req_0_bits_cf_pd_isCall; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_0_bits_cf_pd_isRet = dispatch_io_toLsDq_req_0_bits_cf_pd_isRet; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_0_bits_cf_pred_taken = dispatch_io_toLsDq_req_0_bits_cf_pred_taken; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_0_bits_cf_storeSetHit = dispatch_io_toLsDq_req_0_bits_cf_storeSetHit; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_0_bits_cf_waitForRobIdx_flag = dispatch_io_toLsDq_req_0_bits_cf_waitForRobIdx_flag; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_0_bits_cf_waitForRobIdx_value = dispatch_io_toLsDq_req_0_bits_cf_waitForRobIdx_value; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_0_bits_cf_loadWaitBit = dispatch_io_toLsDq_req_0_bits_cf_loadWaitBit; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_0_bits_cf_loadWaitStrict = dispatch_io_toLsDq_req_0_bits_cf_loadWaitStrict; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_0_bits_cf_ssid = dispatch_io_toLsDq_req_0_bits_cf_ssid; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_0_bits_cf_ftqPtr_flag = dispatch_io_toLsDq_req_0_bits_cf_ftqPtr_flag; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_0_bits_cf_ftqPtr_value = dispatch_io_toLsDq_req_0_bits_cf_ftqPtr_value; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_0_bits_cf_ftqOffset = dispatch_io_toLsDq_req_0_bits_cf_ftqOffset; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_0_bits_ctrl_srcType_0 = dispatch_io_toLsDq_req_0_bits_ctrl_srcType_0; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_0_bits_ctrl_srcType_1 = dispatch_io_toLsDq_req_0_bits_ctrl_srcType_1; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_0_bits_ctrl_srcType_2 = dispatch_io_toLsDq_req_0_bits_ctrl_srcType_2; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_0_bits_ctrl_fuType = dispatch_io_toLsDq_req_0_bits_ctrl_fuType; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_0_bits_ctrl_fuOpType = dispatch_io_toLsDq_req_0_bits_ctrl_fuOpType; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_0_bits_ctrl_rfWen = dispatch_io_toLsDq_req_0_bits_ctrl_rfWen; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_0_bits_ctrl_fpWen = dispatch_io_toLsDq_req_0_bits_ctrl_fpWen; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_0_bits_ctrl_flushPipe = dispatch_io_toLsDq_req_0_bits_ctrl_flushPipe; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_0_bits_ctrl_selImm = dispatch_io_toLsDq_req_0_bits_ctrl_selImm; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_0_bits_ctrl_imm = dispatch_io_toLsDq_req_0_bits_ctrl_imm; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_0_bits_ctrl_fpu_isAddSub = dispatch_io_toLsDq_req_0_bits_ctrl_fpu_isAddSub; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_0_bits_ctrl_fpu_typeTagIn = dispatch_io_toLsDq_req_0_bits_ctrl_fpu_typeTagIn; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_0_bits_ctrl_fpu_typeTagOut = dispatch_io_toLsDq_req_0_bits_ctrl_fpu_typeTagOut; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_0_bits_ctrl_fpu_fromInt = dispatch_io_toLsDq_req_0_bits_ctrl_fpu_fromInt; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_0_bits_ctrl_fpu_wflags = dispatch_io_toLsDq_req_0_bits_ctrl_fpu_wflags; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_0_bits_ctrl_fpu_fpWen = dispatch_io_toLsDq_req_0_bits_ctrl_fpu_fpWen; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_0_bits_ctrl_fpu_fmaCmd = dispatch_io_toLsDq_req_0_bits_ctrl_fpu_fmaCmd; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_0_bits_ctrl_fpu_div = dispatch_io_toLsDq_req_0_bits_ctrl_fpu_div; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_0_bits_ctrl_fpu_sqrt = dispatch_io_toLsDq_req_0_bits_ctrl_fpu_sqrt; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_0_bits_ctrl_fpu_fcvt = dispatch_io_toLsDq_req_0_bits_ctrl_fpu_fcvt; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_0_bits_ctrl_fpu_typ = dispatch_io_toLsDq_req_0_bits_ctrl_fpu_typ; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_0_bits_ctrl_fpu_fmt = dispatch_io_toLsDq_req_0_bits_ctrl_fpu_fmt; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_0_bits_ctrl_fpu_ren3 = dispatch_io_toLsDq_req_0_bits_ctrl_fpu_ren3; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_0_bits_ctrl_fpu_rm = dispatch_io_toLsDq_req_0_bits_ctrl_fpu_rm; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_0_bits_psrc_0 = dispatch_io_toLsDq_req_0_bits_psrc_0; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_0_bits_psrc_1 = dispatch_io_toLsDq_req_0_bits_psrc_1; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_0_bits_psrc_2 = dispatch_io_toLsDq_req_0_bits_psrc_2; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_0_bits_pdest = dispatch_io_toLsDq_req_0_bits_pdest; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_0_bits_robIdx_flag = dispatch_io_toLsDq_req_0_bits_robIdx_flag; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_0_bits_robIdx_value = dispatch_io_toLsDq_req_0_bits_robIdx_value; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_1_valid = dispatch_io_toLsDq_req_1_valid; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_1_bits_cf_foldpc = dispatch_io_toLsDq_req_1_bits_cf_foldpc; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_1_bits_cf_trigger_backendEn_0 = dispatch_io_toLsDq_req_1_bits_cf_trigger_backendEn_0; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_1_bits_cf_trigger_backendEn_1 = dispatch_io_toLsDq_req_1_bits_cf_trigger_backendEn_1; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_1_bits_cf_pd_isRVC = dispatch_io_toLsDq_req_1_bits_cf_pd_isRVC; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_1_bits_cf_pd_brType = dispatch_io_toLsDq_req_1_bits_cf_pd_brType; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_1_bits_cf_pd_isCall = dispatch_io_toLsDq_req_1_bits_cf_pd_isCall; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_1_bits_cf_pd_isRet = dispatch_io_toLsDq_req_1_bits_cf_pd_isRet; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_1_bits_cf_pred_taken = dispatch_io_toLsDq_req_1_bits_cf_pred_taken; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_1_bits_cf_storeSetHit = dispatch_io_toLsDq_req_1_bits_cf_storeSetHit; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_1_bits_cf_waitForRobIdx_flag = dispatch_io_toLsDq_req_1_bits_cf_waitForRobIdx_flag; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_1_bits_cf_waitForRobIdx_value = dispatch_io_toLsDq_req_1_bits_cf_waitForRobIdx_value; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_1_bits_cf_loadWaitBit = dispatch_io_toLsDq_req_1_bits_cf_loadWaitBit; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_1_bits_cf_loadWaitStrict = dispatch_io_toLsDq_req_1_bits_cf_loadWaitStrict; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_1_bits_cf_ssid = dispatch_io_toLsDq_req_1_bits_cf_ssid; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_1_bits_cf_ftqPtr_flag = dispatch_io_toLsDq_req_1_bits_cf_ftqPtr_flag; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_1_bits_cf_ftqPtr_value = dispatch_io_toLsDq_req_1_bits_cf_ftqPtr_value; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_1_bits_cf_ftqOffset = dispatch_io_toLsDq_req_1_bits_cf_ftqOffset; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_1_bits_ctrl_srcType_0 = dispatch_io_toLsDq_req_1_bits_ctrl_srcType_0; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_1_bits_ctrl_srcType_1 = dispatch_io_toLsDq_req_1_bits_ctrl_srcType_1; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_1_bits_ctrl_srcType_2 = dispatch_io_toLsDq_req_1_bits_ctrl_srcType_2; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_1_bits_ctrl_fuType = dispatch_io_toLsDq_req_1_bits_ctrl_fuType; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_1_bits_ctrl_fuOpType = dispatch_io_toLsDq_req_1_bits_ctrl_fuOpType; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_1_bits_ctrl_rfWen = dispatch_io_toLsDq_req_1_bits_ctrl_rfWen; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_1_bits_ctrl_fpWen = dispatch_io_toLsDq_req_1_bits_ctrl_fpWen; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_1_bits_ctrl_flushPipe = dispatch_io_toLsDq_req_1_bits_ctrl_flushPipe; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_1_bits_ctrl_selImm = dispatch_io_toLsDq_req_1_bits_ctrl_selImm; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_1_bits_ctrl_imm = dispatch_io_toLsDq_req_1_bits_ctrl_imm; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_1_bits_ctrl_fpu_isAddSub = dispatch_io_toLsDq_req_1_bits_ctrl_fpu_isAddSub; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_1_bits_ctrl_fpu_typeTagIn = dispatch_io_toLsDq_req_1_bits_ctrl_fpu_typeTagIn; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_1_bits_ctrl_fpu_typeTagOut = dispatch_io_toLsDq_req_1_bits_ctrl_fpu_typeTagOut; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_1_bits_ctrl_fpu_fromInt = dispatch_io_toLsDq_req_1_bits_ctrl_fpu_fromInt; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_1_bits_ctrl_fpu_wflags = dispatch_io_toLsDq_req_1_bits_ctrl_fpu_wflags; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_1_bits_ctrl_fpu_fpWen = dispatch_io_toLsDq_req_1_bits_ctrl_fpu_fpWen; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_1_bits_ctrl_fpu_fmaCmd = dispatch_io_toLsDq_req_1_bits_ctrl_fpu_fmaCmd; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_1_bits_ctrl_fpu_div = dispatch_io_toLsDq_req_1_bits_ctrl_fpu_div; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_1_bits_ctrl_fpu_sqrt = dispatch_io_toLsDq_req_1_bits_ctrl_fpu_sqrt; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_1_bits_ctrl_fpu_fcvt = dispatch_io_toLsDq_req_1_bits_ctrl_fpu_fcvt; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_1_bits_ctrl_fpu_typ = dispatch_io_toLsDq_req_1_bits_ctrl_fpu_typ; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_1_bits_ctrl_fpu_fmt = dispatch_io_toLsDq_req_1_bits_ctrl_fpu_fmt; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_1_bits_ctrl_fpu_ren3 = dispatch_io_toLsDq_req_1_bits_ctrl_fpu_ren3; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_1_bits_ctrl_fpu_rm = dispatch_io_toLsDq_req_1_bits_ctrl_fpu_rm; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_1_bits_psrc_0 = dispatch_io_toLsDq_req_1_bits_psrc_0; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_1_bits_psrc_1 = dispatch_io_toLsDq_req_1_bits_psrc_1; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_1_bits_psrc_2 = dispatch_io_toLsDq_req_1_bits_psrc_2; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_1_bits_pdest = dispatch_io_toLsDq_req_1_bits_pdest; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_1_bits_robIdx_flag = dispatch_io_toLsDq_req_1_bits_robIdx_flag; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_enq_req_1_bits_robIdx_value = dispatch_io_toLsDq_req_1_bits_robIdx_value; // @[CtrlBlock.scala 499:22]
  assign lsDq_io_deq_0_ready = dispatch2_1_io_in_0_ready; // @[CtrlBlock.scala 533:21]
  assign lsDq_io_deq_1_ready = dispatch2_1_io_in_1_ready; // @[CtrlBlock.scala 533:21]
  assign lsDq_io_deq_2_ready = dispatch2_1_io_in_2_ready; // @[CtrlBlock.scala 533:21]
  assign lsDq_io_deq_3_ready = dispatch2_1_io_in_3_ready; // @[CtrlBlock.scala 533:21]
  assign lsDq_io_redirect_valid = redirectForExu_next_valid_REG; // @[BitUtils.scala 26:20 28:18]
  assign lsDq_io_redirect_bits_robIdx_flag = redirectForExu_next_bits_rrobIdx_flag; // @[BitUtils.scala 26:20 33:15]
  assign lsDq_io_redirect_bits_robIdx_value = redirectForExu_next_bits_rrobIdx_value; // @[BitUtils.scala 26:20 33:15]
  assign lsDq_io_redirect_bits_level = redirectForExu_next_bits_rlevel; // @[BitUtils.scala 26:20 33:15]
  assign redirectGen_clock = clock;
  assign redirectGen_reset = reset;
  assign redirectGen_io_exuMispredict_0_valid = exuRedirect_delayed_valid_REG; // @[CtrlBlock.scala 309:23 310:19]
  assign redirectGen_io_exuMispredict_0_bits_uop_cf_pd_isRVC = exuRedirect_delayed_bits_ruop_cf_pd_isRVC; // @[CtrlBlock.scala 309:23 311:18]
  assign redirectGen_io_exuMispredict_0_bits_uop_cf_pd_brType = exuRedirect_delayed_bits_ruop_cf_pd_brType; // @[CtrlBlock.scala 309:23 311:18]
  assign redirectGen_io_exuMispredict_0_bits_uop_cf_pd_isCall = exuRedirect_delayed_bits_ruop_cf_pd_isCall; // @[CtrlBlock.scala 309:23 311:18]
  assign redirectGen_io_exuMispredict_0_bits_uop_cf_pd_isRet = exuRedirect_delayed_bits_ruop_cf_pd_isRet; // @[CtrlBlock.scala 309:23 311:18]
  assign redirectGen_io_exuMispredict_0_bits_uop_ctrl_imm = exuRedirect_delayed_bits_ruop_ctrl_imm; // @[CtrlBlock.scala 309:23 311:18]
  assign redirectGen_io_exuMispredict_0_bits_redirect_robIdx_flag = exuRedirect_delayed_bits_rredirect_robIdx_flag; // @[CtrlBlock.scala 309:23 311:18]
  assign redirectGen_io_exuMispredict_0_bits_redirect_robIdx_value = exuRedirect_delayed_bits_rredirect_robIdx_value; // @[CtrlBlock.scala 309:23 311:18]
  assign redirectGen_io_exuMispredict_0_bits_redirect_ftqIdx_flag = exuRedirect_delayed_bits_rredirect_ftqIdx_flag; // @[CtrlBlock.scala 309:23 311:18]
  assign redirectGen_io_exuMispredict_0_bits_redirect_ftqIdx_value = exuRedirect_delayed_bits_rredirect_ftqIdx_value; // @[CtrlBlock.scala 309:23 311:18]
  assign redirectGen_io_exuMispredict_0_bits_redirect_ftqOffset = exuRedirect_delayed_bits_rredirect_ftqOffset; // @[CtrlBlock.scala 309:23 311:18]
  assign redirectGen_io_exuMispredict_0_bits_redirect_cfiUpdate_target =
    exuRedirect_delayed_bits_rredirect_cfiUpdate_target; // @[CtrlBlock.scala 309:23 311:18]
  assign redirectGen_io_exuMispredict_0_bits_redirect_cfiUpdate_isMisPred =
    exuRedirect_delayed_bits_rredirect_cfiUpdate_isMisPred; // @[CtrlBlock.scala 309:23 311:18]
  assign redirectGen_io_exuMispredict_1_valid = exuRedirect_delayed_valid_REG_1; // @[CtrlBlock.scala 309:23 310:19]
  assign redirectGen_io_exuMispredict_1_bits_uop_cf_pd_isRVC = exuRedirect_delayed_bits_r1_uop_cf_pd_isRVC; // @[CtrlBlock.scala 309:23 311:18]
  assign redirectGen_io_exuMispredict_1_bits_uop_cf_pd_brType = exuRedirect_delayed_bits_r1_uop_cf_pd_brType; // @[CtrlBlock.scala 309:23 311:18]
  assign redirectGen_io_exuMispredict_1_bits_uop_cf_pd_isCall = exuRedirect_delayed_bits_r1_uop_cf_pd_isCall; // @[CtrlBlock.scala 309:23 311:18]
  assign redirectGen_io_exuMispredict_1_bits_uop_cf_pd_isRet = exuRedirect_delayed_bits_r1_uop_cf_pd_isRet; // @[CtrlBlock.scala 309:23 311:18]
  assign redirectGen_io_exuMispredict_1_bits_uop_ctrl_imm = exuRedirect_delayed_bits_r1_uop_ctrl_imm; // @[CtrlBlock.scala 309:23 311:18]
  assign redirectGen_io_exuMispredict_1_bits_redirect_robIdx_flag = exuRedirect_delayed_bits_r1_redirect_robIdx_flag; // @[CtrlBlock.scala 309:23 311:18]
  assign redirectGen_io_exuMispredict_1_bits_redirect_robIdx_value = exuRedirect_delayed_bits_r1_redirect_robIdx_value; // @[CtrlBlock.scala 309:23 311:18]
  assign redirectGen_io_exuMispredict_1_bits_redirect_ftqIdx_flag = exuRedirect_delayed_bits_r1_redirect_ftqIdx_flag; // @[CtrlBlock.scala 309:23 311:18]
  assign redirectGen_io_exuMispredict_1_bits_redirect_ftqIdx_value = exuRedirect_delayed_bits_r1_redirect_ftqIdx_value; // @[CtrlBlock.scala 309:23 311:18]
  assign redirectGen_io_exuMispredict_1_bits_redirect_ftqOffset = exuRedirect_delayed_bits_r1_redirect_ftqOffset; // @[CtrlBlock.scala 309:23 311:18]
  assign redirectGen_io_exuMispredict_1_bits_redirect_cfiUpdate_taken =
    exuRedirect_delayed_bits_r1_redirect_cfiUpdate_taken; // @[CtrlBlock.scala 309:23 311:18]
  assign redirectGen_io_exuMispredict_1_bits_redirect_cfiUpdate_isMisPred =
    exuRedirect_delayed_bits_r1_redirect_cfiUpdate_isMisPred; // @[CtrlBlock.scala 309:23 311:18]
  assign redirectGen_io_exuMispredict_2_valid = exuRedirect_delayed_valid_REG_2; // @[CtrlBlock.scala 309:23 310:19]
  assign redirectGen_io_exuMispredict_2_bits_uop_cf_pd_isRVC = exuRedirect_delayed_bits_r2_uop_cf_pd_isRVC; // @[CtrlBlock.scala 309:23 311:18]
  assign redirectGen_io_exuMispredict_2_bits_uop_cf_pd_brType = exuRedirect_delayed_bits_r2_uop_cf_pd_brType; // @[CtrlBlock.scala 309:23 311:18]
  assign redirectGen_io_exuMispredict_2_bits_uop_cf_pd_isCall = exuRedirect_delayed_bits_r2_uop_cf_pd_isCall; // @[CtrlBlock.scala 309:23 311:18]
  assign redirectGen_io_exuMispredict_2_bits_uop_cf_pd_isRet = exuRedirect_delayed_bits_r2_uop_cf_pd_isRet; // @[CtrlBlock.scala 309:23 311:18]
  assign redirectGen_io_exuMispredict_2_bits_uop_ctrl_imm = exuRedirect_delayed_bits_r2_uop_ctrl_imm; // @[CtrlBlock.scala 309:23 311:18]
  assign redirectGen_io_exuMispredict_2_bits_redirect_robIdx_flag = exuRedirect_delayed_bits_r2_redirect_robIdx_flag; // @[CtrlBlock.scala 309:23 311:18]
  assign redirectGen_io_exuMispredict_2_bits_redirect_robIdx_value = exuRedirect_delayed_bits_r2_redirect_robIdx_value; // @[CtrlBlock.scala 309:23 311:18]
  assign redirectGen_io_exuMispredict_2_bits_redirect_ftqIdx_flag = exuRedirect_delayed_bits_r2_redirect_ftqIdx_flag; // @[CtrlBlock.scala 309:23 311:18]
  assign redirectGen_io_exuMispredict_2_bits_redirect_ftqIdx_value = exuRedirect_delayed_bits_r2_redirect_ftqIdx_value; // @[CtrlBlock.scala 309:23 311:18]
  assign redirectGen_io_exuMispredict_2_bits_redirect_ftqOffset = exuRedirect_delayed_bits_r2_redirect_ftqOffset; // @[CtrlBlock.scala 309:23 311:18]
  assign redirectGen_io_exuMispredict_2_bits_redirect_cfiUpdate_taken =
    exuRedirect_delayed_bits_r2_redirect_cfiUpdate_taken; // @[CtrlBlock.scala 309:23 311:18]
  assign redirectGen_io_exuMispredict_2_bits_redirect_cfiUpdate_isMisPred =
    exuRedirect_delayed_bits_r2_redirect_cfiUpdate_isMisPred; // @[CtrlBlock.scala 309:23 311:18]
  assign redirectGen_io_loadReplay_valid = loadReplay_valid_REG; // @[CtrlBlock.scala 314:24 315:20]
  assign redirectGen_io_loadReplay_bits_robIdx_flag = loadReplay_bits_rrobIdx_flag; // @[CtrlBlock.scala 314:24 319:19]
  assign redirectGen_io_loadReplay_bits_robIdx_value = loadReplay_bits_rrobIdx_value; // @[CtrlBlock.scala 314:24 319:19]
  assign redirectGen_io_loadReplay_bits_ftqIdx_flag = loadReplay_bits_rftqIdx_flag; // @[CtrlBlock.scala 314:24 319:19]
  assign redirectGen_io_loadReplay_bits_ftqIdx_value = loadReplay_bits_rftqIdx_value; // @[CtrlBlock.scala 314:24 319:19]
  assign redirectGen_io_loadReplay_bits_ftqOffset = loadReplay_bits_rftqOffset; // @[CtrlBlock.scala 314:24 319:19]
  assign redirectGen_io_loadReplay_bits_stFtqIdx_value = loadReplay_bits_rstFtqIdx_value; // @[CtrlBlock.scala 314:24 319:19]
  assign redirectGen_io_loadReplay_bits_stFtqOffset = loadReplay_bits_rstFtqOffset; // @[CtrlBlock.scala 314:24 319:19]
  assign redirectGen_io_flush = flushRedirect_valid_REG; // @[CtrlBlock.scala 294:27 295:23]
  assign redirectGen_io_redirectPcRead_data = {redirectGen_io_redirectPcRead_data_hi,1'h0}; // @[Cat.scala 31:58]
  assign redirectGen_io_memPredPcRead_data = {redirectGen_io_memPredPcRead_data_hi,1'h0}; // @[Cat.scala 31:58]
  assign pcMem_clock = clock;
  assign pcMem_io_raddr_0 = intDq_io_deqNext_0_cf_ftqPtr_value; // @[CtrlBlock.scala 541:21]
  assign pcMem_io_raddr_2 = redirectGen_io_redirectPcRead_ptr_value; // @[CtrlBlock.scala 320:21]
  assign pcMem_io_raddr_3 = redirectGen_io_memPredPcRead_ptr_value; // @[CtrlBlock.scala 322:21]
  assign pcMem_io_raddr_4 = _pcMem_io_raddr_4_new_ptr_T_2[2:0]; // @[CircularQueuePtr.scala 39:59]
  assign pcMem_io_raddr_7 = rob_io_flushOut_bits_ftqIdx_value; // @[CtrlBlock.scala 291:23]
  assign pcMem_io_wen_0 = pcMem_io_wen_0_REG; // @[CtrlBlock.scala 287:23]
  assign pcMem_io_waddr_0 = pcMem_io_waddr_0_REG; // @[CtrlBlock.scala 288:23]
  assign pcMem_io_wdata_0_startAddr = pcMem_io_wdata_0_REG_startAddr; // @[CtrlBlock.scala 289:23]
  assign pcMem_io_wdata_0_nextLineAddr = pcMem_io_wdata_0_REG_nextLineAddr; // @[CtrlBlock.scala 289:23]
  assign pcMem_io_wdata_0_isNextMask_0 = pcMem_io_wdata_0_REG_isNextMask_0; // @[CtrlBlock.scala 289:23]
  assign pcMem_io_wdata_0_isNextMask_1 = pcMem_io_wdata_0_REG_isNextMask_1; // @[CtrlBlock.scala 289:23]
  assign pcMem_io_wdata_0_isNextMask_2 = pcMem_io_wdata_0_REG_isNextMask_2; // @[CtrlBlock.scala 289:23]
  assign pcMem_io_wdata_0_isNextMask_3 = pcMem_io_wdata_0_REG_isNextMask_3; // @[CtrlBlock.scala 289:23]
  assign pcMem_io_wdata_0_isNextMask_4 = pcMem_io_wdata_0_REG_isNextMask_4; // @[CtrlBlock.scala 289:23]
  assign pcMem_io_wdata_0_isNextMask_5 = pcMem_io_wdata_0_REG_isNextMask_5; // @[CtrlBlock.scala 289:23]
  assign pcMem_io_wdata_0_isNextMask_6 = pcMem_io_wdata_0_REG_isNextMask_6; // @[CtrlBlock.scala 289:23]
  assign pcMem_io_wdata_0_isNextMask_7 = pcMem_io_wdata_0_REG_isNextMask_7; // @[CtrlBlock.scala 289:23]
  assign frontendFlushValid_delay_clock = clock;
  assign frontendFlushValid_delay_io_in = flushRedirect_valid_REG; // @[CtrlBlock.scala 294:27 295:23]
  assign pc_from_csr_delay_clock = clock;
  assign pc_from_csr_delay_io_in = rob_io_exception_valid; // @[Hold.scala 98:17]
  assign lfst_clock = clock;
  assign lfst_reset = reset;
  assign lfst_io_redirect_valid = lfst_io_redirect_REG_valid; // @[CtrlBlock.scala 426:20]
  assign lfst_io_redirect_bits_robIdx_flag = lfst_io_redirect_REG_bits_robIdx_flag; // @[CtrlBlock.scala 426:20]
  assign lfst_io_redirect_bits_robIdx_value = lfst_io_redirect_REG_bits_robIdx_value; // @[CtrlBlock.scala 426:20]
  assign lfst_io_redirect_bits_level = lfst_io_redirect_REG_bits_level; // @[CtrlBlock.scala 426:20]
  assign lfst_io_dispatch_req_0_valid = dispatch_io_lfst_req_0_valid; // @[CtrlBlock.scala 429:20]
  assign lfst_io_dispatch_req_0_bits_isstore = dispatch_io_lfst_req_0_bits_isstore; // @[CtrlBlock.scala 429:20]
  assign lfst_io_dispatch_req_0_bits_ssid = dispatch_io_lfst_req_0_bits_ssid; // @[CtrlBlock.scala 429:20]
  assign lfst_io_dispatch_req_0_bits_robIdx_flag = dispatch_io_lfst_req_0_bits_robIdx_flag; // @[CtrlBlock.scala 429:20]
  assign lfst_io_dispatch_req_0_bits_robIdx_value = dispatch_io_lfst_req_0_bits_robIdx_value; // @[CtrlBlock.scala 429:20]
  assign lfst_io_dispatch_req_1_valid = dispatch_io_lfst_req_1_valid; // @[CtrlBlock.scala 429:20]
  assign lfst_io_dispatch_req_1_bits_isstore = dispatch_io_lfst_req_1_bits_isstore; // @[CtrlBlock.scala 429:20]
  assign lfst_io_dispatch_req_1_bits_ssid = dispatch_io_lfst_req_1_bits_ssid; // @[CtrlBlock.scala 429:20]
  assign lfst_io_dispatch_req_1_bits_robIdx_flag = dispatch_io_lfst_req_1_bits_robIdx_flag; // @[CtrlBlock.scala 429:20]
  assign lfst_io_dispatch_req_1_bits_robIdx_value = dispatch_io_lfst_req_1_bits_robIdx_value; // @[CtrlBlock.scala 429:20]
  assign lfst_io_storeIssue_0_valid = REG_1_0_valid; // @[CtrlBlock.scala 427:22]
  assign lfst_io_storeIssue_0_bits_uop_cf_storeSetHit = REG_1_0_bits_uop_cf_storeSetHit; // @[CtrlBlock.scala 427:22]
  assign lfst_io_storeIssue_0_bits_uop_cf_ssid = REG_1_0_bits_uop_cf_ssid; // @[CtrlBlock.scala 427:22]
  assign lfst_io_storeIssue_0_bits_uop_robIdx_value = REG_1_0_bits_uop_robIdx_value; // @[CtrlBlock.scala 427:22]
  assign lfst_io_storeIssue_1_valid = REG_1_1_valid; // @[CtrlBlock.scala 427:22]
  assign lfst_io_storeIssue_1_bits_uop_cf_storeSetHit = REG_1_1_bits_uop_cf_storeSetHit; // @[CtrlBlock.scala 427:22]
  assign lfst_io_storeIssue_1_bits_uop_cf_ssid = REG_1_1_bits_uop_cf_ssid; // @[CtrlBlock.scala 427:22]
  assign lfst_io_storeIssue_1_bits_uop_robIdx_value = REG_1_1_bits_uop_robIdx_value; // @[CtrlBlock.scala 427:22]
  assign lfst_io_csrCtrl_lvpred_disable = lfst_io_csrCtrl_REG_lvpred_disable; // @[CtrlBlock.scala 428:19]
  assign lfst_io_csrCtrl_no_spec_load = lfst_io_csrCtrl_REG_no_spec_load; // @[CtrlBlock.scala 428:19]
  assign lfst_io_csrCtrl_storeset_wait_store = lfst_io_csrCtrl_REG_storeset_wait_store; // @[CtrlBlock.scala 428:19]
  assign lsqCtrl_clock = clock;
  assign lsqCtrl_reset = reset;
  assign lsqCtrl_io_redirect_valid = redirectForExu_next_valid_REG; // @[BitUtils.scala 26:20 28:18]
  assign lsqCtrl_io_enq_needAlloc_0 = dispatch2_1_io_enqLsq_needAlloc_0; // @[CtrlBlock.scala 521:22]
  assign lsqCtrl_io_enq_needAlloc_1 = dispatch2_1_io_enqLsq_needAlloc_1; // @[CtrlBlock.scala 521:22]
  assign lsqCtrl_io_enq_needAlloc_2 = dispatch2_1_io_enqLsq_needAlloc_2; // @[CtrlBlock.scala 521:22]
  assign lsqCtrl_io_enq_needAlloc_3 = dispatch2_1_io_enqLsq_needAlloc_3; // @[CtrlBlock.scala 521:22]
  assign lsqCtrl_io_enq_req_0_valid = dispatch2_1_io_enqLsq_req_0_valid; // @[CtrlBlock.scala 521:22]
  assign lsqCtrl_io_enq_req_0_bits_cf_trigger_backendEn_0 = dispatch2_1_io_enqLsq_req_0_bits_cf_trigger_backendEn_0; // @[CtrlBlock.scala 521:22]
  assign lsqCtrl_io_enq_req_0_bits_cf_trigger_backendEn_1 = dispatch2_1_io_enqLsq_req_0_bits_cf_trigger_backendEn_1; // @[CtrlBlock.scala 521:22]
  assign lsqCtrl_io_enq_req_0_bits_ctrl_fuOpType = dispatch2_1_io_enqLsq_req_0_bits_ctrl_fuOpType; // @[CtrlBlock.scala 521:22]
  assign lsqCtrl_io_enq_req_0_bits_ctrl_rfWen = dispatch2_1_io_enqLsq_req_0_bits_ctrl_rfWen; // @[CtrlBlock.scala 521:22]
  assign lsqCtrl_io_enq_req_0_bits_ctrl_fpWen = dispatch2_1_io_enqLsq_req_0_bits_ctrl_fpWen; // @[CtrlBlock.scala 521:22]
  assign lsqCtrl_io_enq_req_0_bits_ctrl_flushPipe = dispatch2_1_io_enqLsq_req_0_bits_ctrl_flushPipe; // @[CtrlBlock.scala 521:22]
  assign lsqCtrl_io_enq_req_0_bits_ctrl_replayInst = dispatch2_1_io_enqLsq_req_0_bits_ctrl_replayInst; // @[CtrlBlock.scala 521:22]
  assign lsqCtrl_io_enq_req_0_bits_pdest = dispatch2_1_io_enqLsq_req_0_bits_pdest; // @[CtrlBlock.scala 521:22]
  assign lsqCtrl_io_enq_req_0_bits_robIdx_flag = dispatch2_1_io_enqLsq_req_0_bits_robIdx_flag; // @[CtrlBlock.scala 521:22]
  assign lsqCtrl_io_enq_req_0_bits_robIdx_value = dispatch2_1_io_enqLsq_req_0_bits_robIdx_value; // @[CtrlBlock.scala 521:22]
  assign lsqCtrl_io_enq_req_1_valid = dispatch2_1_io_enqLsq_req_1_valid; // @[CtrlBlock.scala 521:22]
  assign lsqCtrl_io_enq_req_1_bits_cf_trigger_backendEn_0 = dispatch2_1_io_enqLsq_req_1_bits_cf_trigger_backendEn_0; // @[CtrlBlock.scala 521:22]
  assign lsqCtrl_io_enq_req_1_bits_cf_trigger_backendEn_1 = dispatch2_1_io_enqLsq_req_1_bits_cf_trigger_backendEn_1; // @[CtrlBlock.scala 521:22]
  assign lsqCtrl_io_enq_req_1_bits_ctrl_fuOpType = dispatch2_1_io_enqLsq_req_1_bits_ctrl_fuOpType; // @[CtrlBlock.scala 521:22]
  assign lsqCtrl_io_enq_req_1_bits_ctrl_rfWen = dispatch2_1_io_enqLsq_req_1_bits_ctrl_rfWen; // @[CtrlBlock.scala 521:22]
  assign lsqCtrl_io_enq_req_1_bits_ctrl_fpWen = dispatch2_1_io_enqLsq_req_1_bits_ctrl_fpWen; // @[CtrlBlock.scala 521:22]
  assign lsqCtrl_io_enq_req_1_bits_ctrl_flushPipe = dispatch2_1_io_enqLsq_req_1_bits_ctrl_flushPipe; // @[CtrlBlock.scala 521:22]
  assign lsqCtrl_io_enq_req_1_bits_ctrl_replayInst = dispatch2_1_io_enqLsq_req_1_bits_ctrl_replayInst; // @[CtrlBlock.scala 521:22]
  assign lsqCtrl_io_enq_req_1_bits_pdest = dispatch2_1_io_enqLsq_req_1_bits_pdest; // @[CtrlBlock.scala 521:22]
  assign lsqCtrl_io_enq_req_1_bits_robIdx_flag = dispatch2_1_io_enqLsq_req_1_bits_robIdx_flag; // @[CtrlBlock.scala 521:22]
  assign lsqCtrl_io_enq_req_1_bits_robIdx_value = dispatch2_1_io_enqLsq_req_1_bits_robIdx_value; // @[CtrlBlock.scala 521:22]
  assign lsqCtrl_io_enq_req_2_valid = dispatch2_1_io_enqLsq_req_2_valid; // @[CtrlBlock.scala 521:22]
  assign lsqCtrl_io_enq_req_2_bits_cf_trigger_backendEn_0 = dispatch2_1_io_enqLsq_req_2_bits_cf_trigger_backendEn_0; // @[CtrlBlock.scala 521:22]
  assign lsqCtrl_io_enq_req_2_bits_cf_trigger_backendEn_1 = dispatch2_1_io_enqLsq_req_2_bits_cf_trigger_backendEn_1; // @[CtrlBlock.scala 521:22]
  assign lsqCtrl_io_enq_req_2_bits_ctrl_fuOpType = dispatch2_1_io_enqLsq_req_2_bits_ctrl_fuOpType; // @[CtrlBlock.scala 521:22]
  assign lsqCtrl_io_enq_req_2_bits_ctrl_rfWen = dispatch2_1_io_enqLsq_req_2_bits_ctrl_rfWen; // @[CtrlBlock.scala 521:22]
  assign lsqCtrl_io_enq_req_2_bits_ctrl_fpWen = dispatch2_1_io_enqLsq_req_2_bits_ctrl_fpWen; // @[CtrlBlock.scala 521:22]
  assign lsqCtrl_io_enq_req_2_bits_ctrl_flushPipe = dispatch2_1_io_enqLsq_req_2_bits_ctrl_flushPipe; // @[CtrlBlock.scala 521:22]
  assign lsqCtrl_io_enq_req_2_bits_ctrl_replayInst = dispatch2_1_io_enqLsq_req_2_bits_ctrl_replayInst; // @[CtrlBlock.scala 521:22]
  assign lsqCtrl_io_enq_req_2_bits_pdest = dispatch2_1_io_enqLsq_req_2_bits_pdest; // @[CtrlBlock.scala 521:22]
  assign lsqCtrl_io_enq_req_2_bits_robIdx_flag = dispatch2_1_io_enqLsq_req_2_bits_robIdx_flag; // @[CtrlBlock.scala 521:22]
  assign lsqCtrl_io_enq_req_2_bits_robIdx_value = dispatch2_1_io_enqLsq_req_2_bits_robIdx_value; // @[CtrlBlock.scala 521:22]
  assign lsqCtrl_io_enq_req_3_valid = dispatch2_1_io_enqLsq_req_3_valid; // @[CtrlBlock.scala 521:22]
  assign lsqCtrl_io_enq_req_3_bits_cf_trigger_backendEn_0 = dispatch2_1_io_enqLsq_req_3_bits_cf_trigger_backendEn_0; // @[CtrlBlock.scala 521:22]
  assign lsqCtrl_io_enq_req_3_bits_cf_trigger_backendEn_1 = dispatch2_1_io_enqLsq_req_3_bits_cf_trigger_backendEn_1; // @[CtrlBlock.scala 521:22]
  assign lsqCtrl_io_enq_req_3_bits_ctrl_fuOpType = dispatch2_1_io_enqLsq_req_3_bits_ctrl_fuOpType; // @[CtrlBlock.scala 521:22]
  assign lsqCtrl_io_enq_req_3_bits_ctrl_rfWen = dispatch2_1_io_enqLsq_req_3_bits_ctrl_rfWen; // @[CtrlBlock.scala 521:22]
  assign lsqCtrl_io_enq_req_3_bits_ctrl_fpWen = dispatch2_1_io_enqLsq_req_3_bits_ctrl_fpWen; // @[CtrlBlock.scala 521:22]
  assign lsqCtrl_io_enq_req_3_bits_ctrl_flushPipe = dispatch2_1_io_enqLsq_req_3_bits_ctrl_flushPipe; // @[CtrlBlock.scala 521:22]
  assign lsqCtrl_io_enq_req_3_bits_ctrl_replayInst = dispatch2_1_io_enqLsq_req_3_bits_ctrl_replayInst; // @[CtrlBlock.scala 521:22]
  assign lsqCtrl_io_enq_req_3_bits_pdest = dispatch2_1_io_enqLsq_req_3_bits_pdest; // @[CtrlBlock.scala 521:22]
  assign lsqCtrl_io_enq_req_3_bits_robIdx_flag = dispatch2_1_io_enqLsq_req_3_bits_robIdx_flag; // @[CtrlBlock.scala 521:22]
  assign lsqCtrl_io_enq_req_3_bits_robIdx_value = dispatch2_1_io_enqLsq_req_3_bits_robIdx_value; // @[CtrlBlock.scala 521:22]
  assign lsqCtrl_io_lcommit = io_lqDeq; // @[CtrlBlock.scala 522:26]
  assign lsqCtrl_io_scommit = io_sqDeq; // @[CtrlBlock.scala 523:26]
  assign lsqCtrl_io_lqCancelCnt = io_lqCancelCnt; // @[CtrlBlock.scala 524:30]
  assign lsqCtrl_io_sqCancelCnt = io_sqCancelCnt; // @[CtrlBlock.scala 525:30]
  assign io_cpu_halt_delay_clock = clock;
  assign io_cpu_halt_delay_io_in = rob_io_cpu_halt; // @[Hold.scala 98:17]
  assign pfevent_clock = clock;
  assign pfevent_reset = reset;
  assign pfevent_io_distribute_csr_wvalid = pfevent_io_distribute_csr_REG_wvalid; // @[CtrlBlock.scala 586:29]
  assign pfevent_io_distribute_csr_waddr = pfevent_io_distribute_csr_REG_waddr; // @[CtrlBlock.scala 586:29]
  assign pfevent_io_distribute_csr_wdata = pfevent_io_distribute_csr_REG_wdata; // @[CtrlBlock.scala 586:29]
  assign hpm_clock = clock;
  assign hpm_io_hpm_event_0 = pfevent_io_hpmevent_8; // @[PerfCounterUtils.scala 256:22]
  assign hpm_io_hpm_event_1 = pfevent_io_hpmevent_9; // @[PerfCounterUtils.scala 256:22]
  assign hpm_io_hpm_event_2 = pfevent_io_hpmevent_10; // @[PerfCounterUtils.scala 256:22]
  assign hpm_io_hpm_event_3 = pfevent_io_hpmevent_11; // @[PerfCounterUtils.scala 256:22]
  assign hpm_io_hpm_event_4 = pfevent_io_hpmevent_12; // @[PerfCounterUtils.scala 256:22]
  assign hpm_io_hpm_event_5 = pfevent_io_hpmevent_13; // @[PerfCounterUtils.scala 256:22]
  assign hpm_io_hpm_event_6 = pfevent_io_hpmevent_14; // @[PerfCounterUtils.scala 256:22]
  assign hpm_io_hpm_event_7 = pfevent_io_hpmevent_15; // @[PerfCounterUtils.scala 256:22]
  assign hpm_io_events_sets_0_value = decode_io_perf_0_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_1_value = decode_io_perf_1_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_2_value = decode_io_perf_2_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_3_value = decode_io_perf_3_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_4_value = rename_io_perf_0_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_5_value = rename_io_perf_1_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_6_value = rename_io_perf_2_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_7_value = rename_io_perf_3_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_8_value = rename_io_perf_4_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_9_value = rename_io_perf_5_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_10_value = rename_io_perf_6_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_11_value = rename_io_perf_7_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_12_value = rename_io_perf_8_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_13_value = rename_io_perf_9_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_14_value = rename_io_perf_10_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_15_value = rename_io_perf_11_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_16_value = rename_io_perf_12_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_17_value = rename_io_perf_13_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_18_value = dispatch_io_perf_0_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_19_value = dispatch_io_perf_1_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_20_value = dispatch_io_perf_2_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_21_value = dispatch_io_perf_3_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_23_value = dispatch_io_perf_5_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_24_value = dispatch_io_perf_6_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_25_value = dispatch_io_perf_7_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_26_value = dispatch_io_perf_8_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_27_value = intDq_io_perf_0_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_28_value = intDq_io_perf_1_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_29_value = intDq_io_perf_2_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_30_value = intDq_io_perf_3_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_31_value = intDq_io_perf_4_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_32_value = intDq_io_perf_5_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_33_value = intDq_io_perf_6_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_34_value = intDq_io_perf_7_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_35_value = fpDq_io_perf_0_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_36_value = fpDq_io_perf_1_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_37_value = fpDq_io_perf_2_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_38_value = fpDq_io_perf_3_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_39_value = fpDq_io_perf_4_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_40_value = fpDq_io_perf_5_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_41_value = fpDq_io_perf_6_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_42_value = fpDq_io_perf_7_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_43_value = lsDq_io_perf_0_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_44_value = lsDq_io_perf_1_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_45_value = lsDq_io_perf_2_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_46_value = lsDq_io_perf_3_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_47_value = lsDq_io_perf_4_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_48_value = lsDq_io_perf_5_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_49_value = lsDq_io_perf_6_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_50_value = lsDq_io_perf_7_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_51_value = rob_io_perf_0_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_52_value = rob_io_perf_1_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_53_value = rob_io_perf_2_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_54_value = rob_io_perf_3_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_55_value = rob_io_perf_4_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_56_value = rob_io_perf_5_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_57_value = rob_io_perf_6_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_58_value = rob_io_perf_7_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_59_value = rob_io_perf_8_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_60_value = rob_io_perf_9_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_61_value = rob_io_perf_10_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_62_value = rob_io_perf_11_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_63_value = rob_io_perf_12_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_64_value = rob_io_perf_13_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_65_value = rob_io_perf_14_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_66_value = rob_io_perf_15_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_67_value = rob_io_perf_16_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_68_value = rob_io_perf_17_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_69_value = perfinfo_perfEventsEu0_0_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_70_value = perfinfo_perfEventsEu0_1_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_71_value = perfinfo_perfEventsEu0_2_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_72_value = perfinfo_perfEventsEu0_3_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_73_value = perfinfo_perfEventsEu0_4_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_74_value = perfinfo_perfEventsEu0_5_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_75_value = perfinfo_perfEventsEu1_0_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_76_value = perfinfo_perfEventsEu1_1_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_77_value = perfinfo_perfEventsEu1_2_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_78_value = perfinfo_perfEventsEu1_3_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_79_value = perfinfo_perfEventsEu1_4_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_80_value = perfinfo_perfEventsEu1_5_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_81_value = perfinfo_perfEventsRs_0_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_82_value = perfinfo_perfEventsRs_1_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_83_value = perfinfo_perfEventsRs_2_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_84_value = perfinfo_perfEventsRs_3_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_85_value = perfinfo_perfEventsRs_4_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_86_value = perfinfo_perfEventsRs_5_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_87_value = perfinfo_perfEventsRs_6_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_88_value = perfinfo_perfEventsRs_7_value; // @[PerfCounterUtils.scala 257:24]
  always @(posedge clock) begin
    pcMem_io_wen_0_REG <= io_frontend_fromFtq_pc_mem_wen; // @[CtrlBlock.scala 287:33]
    pcMem_io_waddr_0_REG <= io_frontend_fromFtq_pc_mem_waddr; // @[CtrlBlock.scala 288:33]
    pcMem_io_wdata_0_REG_startAddr <= io_frontend_fromFtq_pc_mem_wdata_startAddr; // @[CtrlBlock.scala 289:33]
    pcMem_io_wdata_0_REG_nextLineAddr <= io_frontend_fromFtq_pc_mem_wdata_nextLineAddr; // @[CtrlBlock.scala 289:33]
    pcMem_io_wdata_0_REG_isNextMask_0 <= io_frontend_fromFtq_pc_mem_wdata_isNextMask_0; // @[CtrlBlock.scala 289:33]
    pcMem_io_wdata_0_REG_isNextMask_1 <= io_frontend_fromFtq_pc_mem_wdata_isNextMask_1; // @[CtrlBlock.scala 289:33]
    pcMem_io_wdata_0_REG_isNextMask_2 <= io_frontend_fromFtq_pc_mem_wdata_isNextMask_2; // @[CtrlBlock.scala 289:33]
    pcMem_io_wdata_0_REG_isNextMask_3 <= io_frontend_fromFtq_pc_mem_wdata_isNextMask_3; // @[CtrlBlock.scala 289:33]
    pcMem_io_wdata_0_REG_isNextMask_4 <= io_frontend_fromFtq_pc_mem_wdata_isNextMask_4; // @[CtrlBlock.scala 289:33]
    pcMem_io_wdata_0_REG_isNextMask_5 <= io_frontend_fromFtq_pc_mem_wdata_isNextMask_5; // @[CtrlBlock.scala 289:33]
    pcMem_io_wdata_0_REG_isNextMask_6 <= io_frontend_fromFtq_pc_mem_wdata_isNextMask_6; // @[CtrlBlock.scala 289:33]
    pcMem_io_wdata_0_REG_isNextMask_7 <= io_frontend_fromFtq_pc_mem_wdata_isNextMask_7; // @[CtrlBlock.scala 289:33]
    flushPC_REG <= rob_io_flushOut_bits_ftqOffset; // @[CtrlBlock.scala 292:50]
    flushRedirect_valid_REG <= rob_io_flushOut_valid; // @[CtrlBlock.scala 295:33]
    if (rob_io_flushOut_valid) begin // @[Reg.scala 17:18]
      flushRedirect_bits_rrobIdx_flag <= rob_io_flushOut_bits_robIdx_flag; // @[Reg.scala 17:22]
    end
    if (rob_io_flushOut_valid) begin // @[Reg.scala 17:18]
      flushRedirect_bits_rrobIdx_value <= rob_io_flushOut_bits_robIdx_value; // @[Reg.scala 17:22]
    end
    if (rob_io_flushOut_valid) begin // @[Reg.scala 17:18]
      flushRedirect_bits_rftqIdx_flag <= rob_io_flushOut_bits_ftqIdx_flag; // @[Reg.scala 17:22]
    end
    if (rob_io_flushOut_valid) begin // @[Reg.scala 17:18]
      flushRedirect_bits_rftqIdx_value <= rob_io_flushOut_bits_ftqIdx_value; // @[Reg.scala 17:22]
    end
    if (rob_io_flushOut_valid) begin // @[Reg.scala 17:18]
      flushRedirect_bits_rftqOffset <= rob_io_flushOut_bits_ftqOffset; // @[Reg.scala 17:22]
    end
    if (rob_io_flushOut_valid) begin // @[Reg.scala 17:18]
      flushRedirect_bits_rlevel <= rob_io_flushOut_bits_level; // @[Reg.scala 17:22]
    end
    if (stage2Redirect_valid) begin // @[Reg.scala 17:18]
      if (flushRedirect_valid_REG) begin // @[CtrlBlock.scala 302:27]
        redirectForExu_next_bits_rrobIdx_flag <= flushRedirect_bits_rrobIdx_flag;
      end else begin
        redirectForExu_next_bits_rrobIdx_flag <= redirectGen_io_stage2Redirect_bits_robIdx_flag;
      end
    end
    if (stage2Redirect_valid) begin // @[Reg.scala 17:18]
      if (flushRedirect_valid_REG) begin // @[CtrlBlock.scala 302:27]
        redirectForExu_next_bits_rrobIdx_value <= flushRedirect_bits_rrobIdx_value;
      end else begin
        redirectForExu_next_bits_rrobIdx_value <= redirectGen_io_stage2Redirect_bits_robIdx_value;
      end
    end
    if (stage2Redirect_valid) begin // @[Reg.scala 17:18]
      if (flushRedirect_valid_REG) begin // @[CtrlBlock.scala 302:27]
        redirectForExu_next_bits_rlevel <= flushRedirect_bits_rlevel;
      end else begin
        redirectForExu_next_bits_rlevel <= redirectGen_io_stage2Redirect_bits_level;
      end
    end
    if (io_exuRedirect_0_valid) begin // @[Reg.scala 17:18]
      exuRedirect_delayed_bits_ruop_cf_pd_isRVC <= io_exuRedirect_0_bits_uop_cf_pd_isRVC; // @[Reg.scala 17:22]
    end
    if (io_exuRedirect_0_valid) begin // @[Reg.scala 17:18]
      exuRedirect_delayed_bits_ruop_cf_pd_brType <= io_exuRedirect_0_bits_uop_cf_pd_brType; // @[Reg.scala 17:22]
    end
    if (io_exuRedirect_0_valid) begin // @[Reg.scala 17:18]
      exuRedirect_delayed_bits_ruop_cf_pd_isCall <= io_exuRedirect_0_bits_uop_cf_pd_isCall; // @[Reg.scala 17:22]
    end
    if (io_exuRedirect_0_valid) begin // @[Reg.scala 17:18]
      exuRedirect_delayed_bits_ruop_cf_pd_isRet <= io_exuRedirect_0_bits_uop_cf_pd_isRet; // @[Reg.scala 17:22]
    end
    if (io_exuRedirect_0_valid) begin // @[Reg.scala 17:18]
      exuRedirect_delayed_bits_ruop_ctrl_imm <= io_exuRedirect_0_bits_uop_ctrl_imm; // @[Reg.scala 17:22]
    end
    if (io_exuRedirect_0_valid) begin // @[Reg.scala 17:18]
      exuRedirect_delayed_bits_rredirect_robIdx_flag <= io_exuRedirect_0_bits_redirect_robIdx_flag; // @[Reg.scala 17:22]
    end
    if (io_exuRedirect_0_valid) begin // @[Reg.scala 17:18]
      exuRedirect_delayed_bits_rredirect_robIdx_value <= io_exuRedirect_0_bits_redirect_robIdx_value; // @[Reg.scala 17:22]
    end
    if (io_exuRedirect_0_valid) begin // @[Reg.scala 17:18]
      exuRedirect_delayed_bits_rredirect_ftqIdx_flag <= io_exuRedirect_0_bits_redirect_ftqIdx_flag; // @[Reg.scala 17:22]
    end
    if (io_exuRedirect_0_valid) begin // @[Reg.scala 17:18]
      exuRedirect_delayed_bits_rredirect_ftqIdx_value <= io_exuRedirect_0_bits_redirect_ftqIdx_value; // @[Reg.scala 17:22]
    end
    if (io_exuRedirect_0_valid) begin // @[Reg.scala 17:18]
      exuRedirect_delayed_bits_rredirect_ftqOffset <= io_exuRedirect_0_bits_redirect_ftqOffset; // @[Reg.scala 17:22]
    end
    if (io_exuRedirect_0_valid) begin // @[Reg.scala 17:18]
      exuRedirect_delayed_bits_rredirect_cfiUpdate_target <= io_exuRedirect_0_bits_redirect_cfiUpdate_target; // @[Reg.scala 17:22]
    end
    if (io_exuRedirect_0_valid) begin // @[Reg.scala 17:18]
      exuRedirect_delayed_bits_rredirect_cfiUpdate_isMisPred <= io_exuRedirect_0_bits_redirect_cfiUpdate_isMisPred; // @[Reg.scala 17:22]
    end
    if (io_exuRedirect_1_valid) begin // @[Reg.scala 17:18]
      exuRedirect_delayed_bits_r1_uop_cf_pd_isRVC <= io_exuRedirect_1_bits_uop_cf_pd_isRVC; // @[Reg.scala 17:22]
    end
    if (io_exuRedirect_1_valid) begin // @[Reg.scala 17:18]
      exuRedirect_delayed_bits_r1_uop_cf_pd_brType <= io_exuRedirect_1_bits_uop_cf_pd_brType; // @[Reg.scala 17:22]
    end
    if (io_exuRedirect_1_valid) begin // @[Reg.scala 17:18]
      exuRedirect_delayed_bits_r1_uop_cf_pd_isCall <= io_exuRedirect_1_bits_uop_cf_pd_isCall; // @[Reg.scala 17:22]
    end
    if (io_exuRedirect_1_valid) begin // @[Reg.scala 17:18]
      exuRedirect_delayed_bits_r1_uop_cf_pd_isRet <= io_exuRedirect_1_bits_uop_cf_pd_isRet; // @[Reg.scala 17:22]
    end
    if (io_exuRedirect_1_valid) begin // @[Reg.scala 17:18]
      exuRedirect_delayed_bits_r1_uop_ctrl_imm <= io_exuRedirect_1_bits_uop_ctrl_imm; // @[Reg.scala 17:22]
    end
    if (io_exuRedirect_1_valid) begin // @[Reg.scala 17:18]
      exuRedirect_delayed_bits_r1_redirect_robIdx_flag <= io_exuRedirect_1_bits_redirect_robIdx_flag; // @[Reg.scala 17:22]
    end
    if (io_exuRedirect_1_valid) begin // @[Reg.scala 17:18]
      exuRedirect_delayed_bits_r1_redirect_robIdx_value <= io_exuRedirect_1_bits_redirect_robIdx_value; // @[Reg.scala 17:22]
    end
    if (io_exuRedirect_1_valid) begin // @[Reg.scala 17:18]
      exuRedirect_delayed_bits_r1_redirect_ftqIdx_flag <= io_exuRedirect_1_bits_redirect_ftqIdx_flag; // @[Reg.scala 17:22]
    end
    if (io_exuRedirect_1_valid) begin // @[Reg.scala 17:18]
      exuRedirect_delayed_bits_r1_redirect_ftqIdx_value <= io_exuRedirect_1_bits_redirect_ftqIdx_value; // @[Reg.scala 17:22]
    end
    if (io_exuRedirect_1_valid) begin // @[Reg.scala 17:18]
      exuRedirect_delayed_bits_r1_redirect_ftqOffset <= io_exuRedirect_1_bits_redirect_ftqOffset; // @[Reg.scala 17:22]
    end
    if (io_exuRedirect_1_valid) begin // @[Reg.scala 17:18]
      exuRedirect_delayed_bits_r1_redirect_cfiUpdate_taken <= io_exuRedirect_1_bits_redirect_cfiUpdate_taken; // @[Reg.scala 17:22]
    end
    if (io_exuRedirect_1_valid) begin // @[Reg.scala 17:18]
      exuRedirect_delayed_bits_r1_redirect_cfiUpdate_isMisPred <= io_exuRedirect_1_bits_redirect_cfiUpdate_isMisPred; // @[Reg.scala 17:22]
    end
    if (io_exuRedirect_2_valid) begin // @[Reg.scala 17:18]
      exuRedirect_delayed_bits_r2_uop_cf_pd_isRVC <= io_exuRedirect_2_bits_uop_cf_pd_isRVC; // @[Reg.scala 17:22]
    end
    if (io_exuRedirect_2_valid) begin // @[Reg.scala 17:18]
      exuRedirect_delayed_bits_r2_uop_cf_pd_brType <= io_exuRedirect_2_bits_uop_cf_pd_brType; // @[Reg.scala 17:22]
    end
    if (io_exuRedirect_2_valid) begin // @[Reg.scala 17:18]
      exuRedirect_delayed_bits_r2_uop_cf_pd_isCall <= io_exuRedirect_2_bits_uop_cf_pd_isCall; // @[Reg.scala 17:22]
    end
    if (io_exuRedirect_2_valid) begin // @[Reg.scala 17:18]
      exuRedirect_delayed_bits_r2_uop_cf_pd_isRet <= io_exuRedirect_2_bits_uop_cf_pd_isRet; // @[Reg.scala 17:22]
    end
    if (io_exuRedirect_2_valid) begin // @[Reg.scala 17:18]
      exuRedirect_delayed_bits_r2_uop_ctrl_imm <= io_exuRedirect_2_bits_uop_ctrl_imm; // @[Reg.scala 17:22]
    end
    if (io_exuRedirect_2_valid) begin // @[Reg.scala 17:18]
      exuRedirect_delayed_bits_r2_redirect_robIdx_flag <= io_exuRedirect_2_bits_redirect_robIdx_flag; // @[Reg.scala 17:22]
    end
    if (io_exuRedirect_2_valid) begin // @[Reg.scala 17:18]
      exuRedirect_delayed_bits_r2_redirect_robIdx_value <= io_exuRedirect_2_bits_redirect_robIdx_value; // @[Reg.scala 17:22]
    end
    if (io_exuRedirect_2_valid) begin // @[Reg.scala 17:18]
      exuRedirect_delayed_bits_r2_redirect_ftqIdx_flag <= io_exuRedirect_2_bits_redirect_ftqIdx_flag; // @[Reg.scala 17:22]
    end
    if (io_exuRedirect_2_valid) begin // @[Reg.scala 17:18]
      exuRedirect_delayed_bits_r2_redirect_ftqIdx_value <= io_exuRedirect_2_bits_redirect_ftqIdx_value; // @[Reg.scala 17:22]
    end
    if (io_exuRedirect_2_valid) begin // @[Reg.scala 17:18]
      exuRedirect_delayed_bits_r2_redirect_ftqOffset <= io_exuRedirect_2_bits_redirect_ftqOffset; // @[Reg.scala 17:22]
    end
    if (io_exuRedirect_2_valid) begin // @[Reg.scala 17:18]
      exuRedirect_delayed_bits_r2_redirect_cfiUpdate_taken <= io_exuRedirect_2_bits_redirect_cfiUpdate_taken; // @[Reg.scala 17:22]
    end
    if (io_exuRedirect_2_valid) begin // @[Reg.scala 17:18]
      exuRedirect_delayed_bits_r2_redirect_cfiUpdate_isMisPred <= io_exuRedirect_2_bits_redirect_cfiUpdate_isMisPred; // @[Reg.scala 17:22]
    end
    if (io_memoryViolation_valid) begin // @[Reg.scala 17:18]
      loadReplay_bits_rrobIdx_flag <= io_memoryViolation_bits_robIdx_flag; // @[Reg.scala 17:22]
    end
    if (io_memoryViolation_valid) begin // @[Reg.scala 17:18]
      loadReplay_bits_rrobIdx_value <= io_memoryViolation_bits_robIdx_value; // @[Reg.scala 17:22]
    end
    if (io_memoryViolation_valid) begin // @[Reg.scala 17:18]
      loadReplay_bits_rftqIdx_flag <= io_memoryViolation_bits_ftqIdx_flag; // @[Reg.scala 17:22]
    end
    if (io_memoryViolation_valid) begin // @[Reg.scala 17:18]
      loadReplay_bits_rftqIdx_value <= io_memoryViolation_bits_ftqIdx_value; // @[Reg.scala 17:22]
    end
    if (io_memoryViolation_valid) begin // @[Reg.scala 17:18]
      loadReplay_bits_rftqOffset <= io_memoryViolation_bits_ftqOffset; // @[Reg.scala 17:22]
    end
    if (io_memoryViolation_valid) begin // @[Reg.scala 17:18]
      loadReplay_bits_rstFtqIdx_value <= io_memoryViolation_bits_stFtqIdx_value; // @[Reg.scala 17:22]
    end
    if (io_memoryViolation_valid) begin // @[Reg.scala 17:18]
      loadReplay_bits_rstFtqOffset <= io_memoryViolation_bits_stFtqOffset; // @[Reg.scala 17:22]
    end
    redirectGen_io_redirectPcRead_data_REG <= redirectGen_io_redirectPcRead_offset; // @[CtrlBlock.scala 321:72]
    redirectGen_io_memPredPcRead_data_REG <= redirectGen_io_memPredPcRead_offset; // @[CtrlBlock.scala 323:71]
    if (flushRedirect_valid_REG) begin // @[Reg.scala 17:18]
      frontendFlushBits_ftqIdx_flag <= flushRedirect_bits_rftqIdx_flag; // @[Reg.scala 17:22]
    end
    if (flushRedirect_valid_REG) begin // @[Reg.scala 17:18]
      frontendFlushBits_ftqIdx_value <= flushRedirect_bits_rftqIdx_value; // @[Reg.scala 17:22]
    end
    if (flushRedirect_valid_REG) begin // @[Reg.scala 17:18]
      frontendFlushBits_ftqOffset <= flushRedirect_bits_rftqOffset; // @[Reg.scala 17:22]
    end
    if (flushRedirect_valid_REG) begin // @[Reg.scala 17:18]
      frontendFlushBits_level <= flushRedirect_bits_rlevel; // @[Reg.scala 17:22]
    end
    io_frontend_toFtq_rob_commits_0_valid_REG <= rob_io_commits_commitValid_0 & rob_io_commits_isCommit & ~
      rob_io_flushOut_valid; // @[CtrlBlock.scala 337:78]
    if (is_commit) begin // @[Reg.scala 17:18]
      io_frontend_toFtq_rob_commits_0_bits_rcommitType <= rob_io_commits_info_0_commitType; // @[Reg.scala 17:22]
    end
    if (is_commit) begin // @[Reg.scala 17:18]
      io_frontend_toFtq_rob_commits_0_bits_rftqIdx_flag <= rob_io_commits_info_0_ftqIdx_flag; // @[Reg.scala 17:22]
    end
    if (is_commit) begin // @[Reg.scala 17:18]
      io_frontend_toFtq_rob_commits_0_bits_rftqIdx_value <= rob_io_commits_info_0_ftqIdx_value; // @[Reg.scala 17:22]
    end
    if (is_commit) begin // @[Reg.scala 17:18]
      io_frontend_toFtq_rob_commits_0_bits_rftqOffset <= rob_io_commits_info_0_ftqOffset; // @[Reg.scala 17:22]
    end
    io_frontend_toFtq_rob_commits_1_valid_REG <= rob_io_commits_commitValid_1 & rob_io_commits_isCommit & ~
      rob_io_flushOut_valid; // @[CtrlBlock.scala 337:78]
    if (is_commit_1) begin // @[Reg.scala 17:18]
      io_frontend_toFtq_rob_commits_1_bits_rcommitType <= rob_io_commits_info_1_commitType; // @[Reg.scala 17:22]
    end
    if (is_commit_1) begin // @[Reg.scala 17:18]
      io_frontend_toFtq_rob_commits_1_bits_rftqIdx_flag <= rob_io_commits_info_1_ftqIdx_flag; // @[Reg.scala 17:22]
    end
    if (is_commit_1) begin // @[Reg.scala 17:18]
      io_frontend_toFtq_rob_commits_1_bits_rftqIdx_value <= rob_io_commits_info_1_ftqIdx_value; // @[Reg.scala 17:22]
    end
    if (is_commit_1) begin // @[Reg.scala 17:18]
      io_frontend_toFtq_rob_commits_1_bits_rftqOffset <= rob_io_commits_info_1_ftqOffset; // @[Reg.scala 17:22]
    end
    if (flushRedirect_valid_REG) begin // @[Reg.scala 17:18]
      if (flushRedirect_bits_rlevel) begin // @[CtrlBlock.scala 351:35]
        rob_flush_pc <= flushPC;
      end else begin
        rob_flush_pc <= _rob_flush_pc_T_2;
      end
    end
    if (pc_from_csr) begin // @[CtrlBlock.scala 355:24]
      io_frontend_toFtq_redirect_bits_cfiUpdate_target_REG <= io_robio_toCSR_trapTarget;
    end else begin
      io_frontend_toFtq_redirect_bits_cfiUpdate_target_REG <= rob_flush_pc;
    end
    REG <= io_frontend_toFtq_redirect_valid; // @[CtrlBlock.scala 365:22]
    decode_io_csrCtrl_REG_fusion_enable <= io_csrCtrl_fusion_enable; // @[CtrlBlock.scala 403:31]
    decode_io_csrCtrl_REG_wfi_enable <= io_csrCtrl_wfi_enable; // @[CtrlBlock.scala 403:31]
    decode_io_csrCtrl_REG_svinval_enable <= io_csrCtrl_svinval_enable; // @[CtrlBlock.scala 403:31]
    decode_io_csrCtrl_REG_singlestep <= io_csrCtrl_singlestep; // @[CtrlBlock.scala 403:31]
    ssit_io_update_REG_valid <= redirectGen_io_memPredUpdate_valid; // @[CtrlBlock.scala 419:28]
    ssit_io_update_REG_ldpc <= redirectGen_io_memPredUpdate_ldpc; // @[CtrlBlock.scala 419:28]
    ssit_io_update_REG_stpc <= redirectGen_io_memPredUpdate_stpc; // @[CtrlBlock.scala 419:28]
    ssit_io_csrCtrl_REG_lvpred_timeout <= io_csrCtrl_lvpred_timeout; // @[CtrlBlock.scala 420:29]
    lfst_io_redirect_REG_valid <= io_redirect_valid; // @[CtrlBlock.scala 426:30]
    lfst_io_redirect_REG_bits_robIdx_flag <= io_redirect_bits_robIdx_flag; // @[CtrlBlock.scala 426:30]
    lfst_io_redirect_REG_bits_robIdx_value <= io_redirect_bits_robIdx_value; // @[CtrlBlock.scala 426:30]
    lfst_io_redirect_REG_bits_level <= io_redirect_bits_level; // @[CtrlBlock.scala 426:30]
    REG_1_0_valid <= io_stIn_0_valid; // @[CtrlBlock.scala 427:32]
    REG_1_0_bits_uop_cf_storeSetHit <= io_stIn_0_bits_uop_cf_storeSetHit; // @[CtrlBlock.scala 427:32]
    REG_1_0_bits_uop_cf_ssid <= io_stIn_0_bits_uop_cf_ssid; // @[CtrlBlock.scala 427:32]
    REG_1_0_bits_uop_robIdx_value <= io_stIn_0_bits_uop_robIdx_value; // @[CtrlBlock.scala 427:32]
    REG_1_1_valid <= io_stIn_1_valid; // @[CtrlBlock.scala 427:32]
    REG_1_1_bits_uop_cf_storeSetHit <= io_stIn_1_bits_uop_cf_storeSetHit; // @[CtrlBlock.scala 427:32]
    REG_1_1_bits_uop_cf_ssid <= io_stIn_1_bits_uop_cf_ssid; // @[CtrlBlock.scala 427:32]
    REG_1_1_bits_uop_robIdx_value <= io_stIn_1_bits_uop_robIdx_value; // @[CtrlBlock.scala 427:32]
    lfst_io_csrCtrl_REG_lvpred_disable <= io_csrCtrl_lvpred_disable; // @[CtrlBlock.scala 428:29]
    lfst_io_csrCtrl_REG_no_spec_load <= io_csrCtrl_no_spec_load; // @[CtrlBlock.scala 428:29]
    lfst_io_csrCtrl_REG_storeset_wait_store <= io_csrCtrl_storeset_wait_store; // @[CtrlBlock.scala 428:29]
    if (renamePipe_leftFire) begin // @[Reg.scala 17:18]
      renamePipe_data_cf_foldpc <= decode_io_out_0_bits_cf_foldpc; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire) begin // @[Reg.scala 17:18]
      renamePipe_data_cf_exceptionVec_1 <= decode_io_out_0_bits_cf_exceptionVec_1; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire) begin // @[Reg.scala 17:18]
      renamePipe_data_cf_exceptionVec_2 <= decode_io_out_0_bits_cf_exceptionVec_2; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire) begin // @[Reg.scala 17:18]
      renamePipe_data_cf_exceptionVec_12 <= decode_io_out_0_bits_cf_exceptionVec_12; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire) begin // @[Reg.scala 17:18]
      renamePipe_data_cf_trigger_frontendHit_0 <= decode_io_out_0_bits_cf_trigger_frontendHit_0; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire) begin // @[Reg.scala 17:18]
      renamePipe_data_cf_trigger_frontendHit_1 <= decode_io_out_0_bits_cf_trigger_frontendHit_1; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire) begin // @[Reg.scala 17:18]
      renamePipe_data_cf_trigger_frontendHit_2 <= decode_io_out_0_bits_cf_trigger_frontendHit_2; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire) begin // @[Reg.scala 17:18]
      renamePipe_data_cf_trigger_frontendHit_3 <= decode_io_out_0_bits_cf_trigger_frontendHit_3; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire) begin // @[Reg.scala 17:18]
      renamePipe_data_cf_trigger_backendEn_0 <= decode_io_out_0_bits_cf_trigger_backendEn_0; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire) begin // @[Reg.scala 17:18]
      renamePipe_data_cf_trigger_backendEn_1 <= decode_io_out_0_bits_cf_trigger_backendEn_1; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire) begin // @[Reg.scala 17:18]
      renamePipe_data_cf_pd_isRVC <= decode_io_out_0_bits_cf_pd_isRVC; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire) begin // @[Reg.scala 17:18]
      renamePipe_data_cf_pd_brType <= decode_io_out_0_bits_cf_pd_brType; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire) begin // @[Reg.scala 17:18]
      renamePipe_data_cf_pd_isCall <= decode_io_out_0_bits_cf_pd_isCall; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire) begin // @[Reg.scala 17:18]
      renamePipe_data_cf_pd_isRet <= decode_io_out_0_bits_cf_pd_isRet; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire) begin // @[Reg.scala 17:18]
      renamePipe_data_cf_pred_taken <= decode_io_out_0_bits_cf_pred_taken; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire) begin // @[Reg.scala 17:18]
      renamePipe_data_cf_crossPageIPFFix <= decode_io_out_0_bits_cf_crossPageIPFFix; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire) begin // @[Reg.scala 17:18]
      renamePipe_data_cf_ftqPtr_flag <= decode_io_out_0_bits_cf_ftqPtr_flag; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire) begin // @[Reg.scala 17:18]
      renamePipe_data_cf_ftqPtr_value <= decode_io_out_0_bits_cf_ftqPtr_value; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire) begin // @[Reg.scala 17:18]
      renamePipe_data_cf_ftqOffset <= decode_io_out_0_bits_cf_ftqOffset; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire) begin // @[Reg.scala 17:18]
      renamePipe_data_ctrl_srcType_0 <= decode_io_out_0_bits_ctrl_srcType_0; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire) begin // @[Reg.scala 17:18]
      renamePipe_data_ctrl_srcType_1 <= decode_io_out_0_bits_ctrl_srcType_1; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire) begin // @[Reg.scala 17:18]
      renamePipe_data_ctrl_srcType_2 <= decode_io_out_0_bits_ctrl_srcType_2; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire) begin // @[Reg.scala 17:18]
      renamePipe_data_ctrl_lsrc_0 <= decode_io_out_0_bits_ctrl_lsrc_0; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire) begin // @[Reg.scala 17:18]
      renamePipe_data_ctrl_lsrc_1 <= decode_io_out_0_bits_ctrl_lsrc_1; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire) begin // @[Reg.scala 17:18]
      renamePipe_data_ctrl_ldest <= decode_io_out_0_bits_ctrl_ldest; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire) begin // @[Reg.scala 17:18]
      renamePipe_data_ctrl_fuType <= decode_io_out_0_bits_ctrl_fuType; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire) begin // @[Reg.scala 17:18]
      renamePipe_data_ctrl_fuOpType <= decode_io_out_0_bits_ctrl_fuOpType; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire) begin // @[Reg.scala 17:18]
      renamePipe_data_ctrl_rfWen <= decode_io_out_0_bits_ctrl_rfWen; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire) begin // @[Reg.scala 17:18]
      renamePipe_data_ctrl_fpWen <= decode_io_out_0_bits_ctrl_fpWen; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire) begin // @[Reg.scala 17:18]
      renamePipe_data_ctrl_isXSTrap <= decode_io_out_0_bits_ctrl_isXSTrap; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire) begin // @[Reg.scala 17:18]
      renamePipe_data_ctrl_noSpecExec <= decode_io_out_0_bits_ctrl_noSpecExec; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire) begin // @[Reg.scala 17:18]
      renamePipe_data_ctrl_blockBackward <= decode_io_out_0_bits_ctrl_blockBackward; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire) begin // @[Reg.scala 17:18]
      renamePipe_data_ctrl_flushPipe <= decode_io_out_0_bits_ctrl_flushPipe; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire) begin // @[Reg.scala 17:18]
      renamePipe_data_ctrl_selImm <= decode_io_out_0_bits_ctrl_selImm; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire) begin // @[Reg.scala 17:18]
      renamePipe_data_ctrl_imm <= decode_io_out_0_bits_ctrl_imm; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire) begin // @[Reg.scala 17:18]
      renamePipe_data_ctrl_fpu_isAddSub <= decode_io_out_0_bits_ctrl_fpu_isAddSub; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire) begin // @[Reg.scala 17:18]
      renamePipe_data_ctrl_fpu_typeTagIn <= decode_io_out_0_bits_ctrl_fpu_typeTagIn; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire) begin // @[Reg.scala 17:18]
      renamePipe_data_ctrl_fpu_typeTagOut <= decode_io_out_0_bits_ctrl_fpu_typeTagOut; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire) begin // @[Reg.scala 17:18]
      renamePipe_data_ctrl_fpu_fromInt <= decode_io_out_0_bits_ctrl_fpu_fromInt; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire) begin // @[Reg.scala 17:18]
      renamePipe_data_ctrl_fpu_wflags <= decode_io_out_0_bits_ctrl_fpu_wflags; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire) begin // @[Reg.scala 17:18]
      renamePipe_data_ctrl_fpu_fpWen <= decode_io_out_0_bits_ctrl_fpu_fpWen; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire) begin // @[Reg.scala 17:18]
      renamePipe_data_ctrl_fpu_fmaCmd <= decode_io_out_0_bits_ctrl_fpu_fmaCmd; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire) begin // @[Reg.scala 17:18]
      renamePipe_data_ctrl_fpu_div <= decode_io_out_0_bits_ctrl_fpu_div; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire) begin // @[Reg.scala 17:18]
      renamePipe_data_ctrl_fpu_sqrt <= decode_io_out_0_bits_ctrl_fpu_sqrt; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire) begin // @[Reg.scala 17:18]
      renamePipe_data_ctrl_fpu_fcvt <= decode_io_out_0_bits_ctrl_fpu_fcvt; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire) begin // @[Reg.scala 17:18]
      renamePipe_data_ctrl_fpu_typ <= decode_io_out_0_bits_ctrl_fpu_typ; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire) begin // @[Reg.scala 17:18]
      renamePipe_data_ctrl_fpu_fmt <= decode_io_out_0_bits_ctrl_fpu_fmt; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire) begin // @[Reg.scala 17:18]
      renamePipe_data_ctrl_fpu_ren3 <= decode_io_out_0_bits_ctrl_fpu_ren3; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire) begin // @[Reg.scala 17:18]
      renamePipe_data_ctrl_fpu_rm <= decode_io_out_0_bits_ctrl_fpu_rm; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire) begin // @[Reg.scala 17:18]
      renamePipe_data_ctrl_isMove <= decode_io_out_0_bits_ctrl_isMove; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire_1) begin // @[Reg.scala 17:18]
      renamePipe_data_1_cf_foldpc <= decode_io_out_1_bits_cf_foldpc; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire_1) begin // @[Reg.scala 17:18]
      renamePipe_data_1_cf_exceptionVec_1 <= decode_io_out_1_bits_cf_exceptionVec_1; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire_1) begin // @[Reg.scala 17:18]
      renamePipe_data_1_cf_exceptionVec_2 <= decode_io_out_1_bits_cf_exceptionVec_2; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire_1) begin // @[Reg.scala 17:18]
      renamePipe_data_1_cf_exceptionVec_12 <= decode_io_out_1_bits_cf_exceptionVec_12; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire_1) begin // @[Reg.scala 17:18]
      renamePipe_data_1_cf_trigger_frontendHit_0 <= decode_io_out_1_bits_cf_trigger_frontendHit_0; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire_1) begin // @[Reg.scala 17:18]
      renamePipe_data_1_cf_trigger_frontendHit_1 <= decode_io_out_1_bits_cf_trigger_frontendHit_1; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire_1) begin // @[Reg.scala 17:18]
      renamePipe_data_1_cf_trigger_frontendHit_2 <= decode_io_out_1_bits_cf_trigger_frontendHit_2; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire_1) begin // @[Reg.scala 17:18]
      renamePipe_data_1_cf_trigger_frontendHit_3 <= decode_io_out_1_bits_cf_trigger_frontendHit_3; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire_1) begin // @[Reg.scala 17:18]
      renamePipe_data_1_cf_trigger_backendEn_0 <= decode_io_out_1_bits_cf_trigger_backendEn_0; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire_1) begin // @[Reg.scala 17:18]
      renamePipe_data_1_cf_trigger_backendEn_1 <= decode_io_out_1_bits_cf_trigger_backendEn_1; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire_1) begin // @[Reg.scala 17:18]
      renamePipe_data_1_cf_pd_isRVC <= decode_io_out_1_bits_cf_pd_isRVC; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire_1) begin // @[Reg.scala 17:18]
      renamePipe_data_1_cf_pd_brType <= decode_io_out_1_bits_cf_pd_brType; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire_1) begin // @[Reg.scala 17:18]
      renamePipe_data_1_cf_pd_isCall <= decode_io_out_1_bits_cf_pd_isCall; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire_1) begin // @[Reg.scala 17:18]
      renamePipe_data_1_cf_pd_isRet <= decode_io_out_1_bits_cf_pd_isRet; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire_1) begin // @[Reg.scala 17:18]
      renamePipe_data_1_cf_pred_taken <= decode_io_out_1_bits_cf_pred_taken; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire_1) begin // @[Reg.scala 17:18]
      renamePipe_data_1_cf_crossPageIPFFix <= decode_io_out_1_bits_cf_crossPageIPFFix; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire_1) begin // @[Reg.scala 17:18]
      renamePipe_data_1_cf_ftqPtr_flag <= decode_io_out_1_bits_cf_ftqPtr_flag; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire_1) begin // @[Reg.scala 17:18]
      renamePipe_data_1_cf_ftqPtr_value <= decode_io_out_1_bits_cf_ftqPtr_value; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire_1) begin // @[Reg.scala 17:18]
      renamePipe_data_1_cf_ftqOffset <= decode_io_out_1_bits_cf_ftqOffset; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire_1) begin // @[Reg.scala 17:18]
      renamePipe_data_1_ctrl_srcType_0 <= decode_io_out_1_bits_ctrl_srcType_0; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire_1) begin // @[Reg.scala 17:18]
      renamePipe_data_1_ctrl_srcType_1 <= decode_io_out_1_bits_ctrl_srcType_1; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire_1) begin // @[Reg.scala 17:18]
      renamePipe_data_1_ctrl_srcType_2 <= decode_io_out_1_bits_ctrl_srcType_2; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire_1) begin // @[Reg.scala 17:18]
      renamePipe_data_1_ctrl_lsrc_0 <= decode_io_out_1_bits_ctrl_lsrc_0; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire_1) begin // @[Reg.scala 17:18]
      renamePipe_data_1_ctrl_lsrc_1 <= decode_io_out_1_bits_ctrl_lsrc_1; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire_1) begin // @[Reg.scala 17:18]
      renamePipe_data_1_ctrl_lsrc_2 <= decode_io_out_1_bits_ctrl_lsrc_2; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire_1) begin // @[Reg.scala 17:18]
      renamePipe_data_1_ctrl_ldest <= decode_io_out_1_bits_ctrl_ldest; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire_1) begin // @[Reg.scala 17:18]
      renamePipe_data_1_ctrl_fuType <= decode_io_out_1_bits_ctrl_fuType; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire_1) begin // @[Reg.scala 17:18]
      renamePipe_data_1_ctrl_fuOpType <= decode_io_out_1_bits_ctrl_fuOpType; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire_1) begin // @[Reg.scala 17:18]
      renamePipe_data_1_ctrl_rfWen <= decode_io_out_1_bits_ctrl_rfWen; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire_1) begin // @[Reg.scala 17:18]
      renamePipe_data_1_ctrl_fpWen <= decode_io_out_1_bits_ctrl_fpWen; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire_1) begin // @[Reg.scala 17:18]
      renamePipe_data_1_ctrl_isXSTrap <= decode_io_out_1_bits_ctrl_isXSTrap; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire_1) begin // @[Reg.scala 17:18]
      renamePipe_data_1_ctrl_noSpecExec <= decode_io_out_1_bits_ctrl_noSpecExec; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire_1) begin // @[Reg.scala 17:18]
      renamePipe_data_1_ctrl_blockBackward <= decode_io_out_1_bits_ctrl_blockBackward; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire_1) begin // @[Reg.scala 17:18]
      renamePipe_data_1_ctrl_flushPipe <= decode_io_out_1_bits_ctrl_flushPipe; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire_1) begin // @[Reg.scala 17:18]
      renamePipe_data_1_ctrl_selImm <= decode_io_out_1_bits_ctrl_selImm; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire_1) begin // @[Reg.scala 17:18]
      renamePipe_data_1_ctrl_imm <= decode_io_out_1_bits_ctrl_imm; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire_1) begin // @[Reg.scala 17:18]
      renamePipe_data_1_ctrl_fpu_isAddSub <= decode_io_out_1_bits_ctrl_fpu_isAddSub; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire_1) begin // @[Reg.scala 17:18]
      renamePipe_data_1_ctrl_fpu_typeTagIn <= decode_io_out_1_bits_ctrl_fpu_typeTagIn; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire_1) begin // @[Reg.scala 17:18]
      renamePipe_data_1_ctrl_fpu_typeTagOut <= decode_io_out_1_bits_ctrl_fpu_typeTagOut; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire_1) begin // @[Reg.scala 17:18]
      renamePipe_data_1_ctrl_fpu_fromInt <= decode_io_out_1_bits_ctrl_fpu_fromInt; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire_1) begin // @[Reg.scala 17:18]
      renamePipe_data_1_ctrl_fpu_wflags <= decode_io_out_1_bits_ctrl_fpu_wflags; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire_1) begin // @[Reg.scala 17:18]
      renamePipe_data_1_ctrl_fpu_fpWen <= decode_io_out_1_bits_ctrl_fpu_fpWen; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire_1) begin // @[Reg.scala 17:18]
      renamePipe_data_1_ctrl_fpu_fmaCmd <= decode_io_out_1_bits_ctrl_fpu_fmaCmd; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire_1) begin // @[Reg.scala 17:18]
      renamePipe_data_1_ctrl_fpu_div <= decode_io_out_1_bits_ctrl_fpu_div; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire_1) begin // @[Reg.scala 17:18]
      renamePipe_data_1_ctrl_fpu_sqrt <= decode_io_out_1_bits_ctrl_fpu_sqrt; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire_1) begin // @[Reg.scala 17:18]
      renamePipe_data_1_ctrl_fpu_fcvt <= decode_io_out_1_bits_ctrl_fpu_fcvt; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire_1) begin // @[Reg.scala 17:18]
      renamePipe_data_1_ctrl_fpu_typ <= decode_io_out_1_bits_ctrl_fpu_typ; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire_1) begin // @[Reg.scala 17:18]
      renamePipe_data_1_ctrl_fpu_fmt <= decode_io_out_1_bits_ctrl_fpu_fmt; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire_1) begin // @[Reg.scala 17:18]
      renamePipe_data_1_ctrl_fpu_ren3 <= decode_io_out_1_bits_ctrl_fpu_ren3; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire_1) begin // @[Reg.scala 17:18]
      renamePipe_data_1_ctrl_fpu_rm <= decode_io_out_1_bits_ctrl_fpu_rm; // @[Reg.scala 17:22]
    end
    if (renamePipe_leftFire_1) begin // @[Reg.scala 17:18]
      renamePipe_data_1_ctrl_isMove <= decode_io_out_1_bits_ctrl_isMove; // @[Reg.scala 17:22]
    end
    if (leftFire) begin // @[Reg.scala 17:18]
      data_cf_foldpc <= rename_io_out_0_bits_cf_foldpc; // @[Reg.scala 17:22]
    end
    if (leftFire) begin // @[Reg.scala 17:18]
      data_cf_exceptionVec_1 <= rename_io_out_0_bits_cf_exceptionVec_1; // @[Reg.scala 17:22]
    end
    if (leftFire) begin // @[Reg.scala 17:18]
      data_cf_exceptionVec_2 <= rename_io_out_0_bits_cf_exceptionVec_2; // @[Reg.scala 17:22]
    end
    if (leftFire) begin // @[Reg.scala 17:18]
      data_cf_exceptionVec_12 <= rename_io_out_0_bits_cf_exceptionVec_12; // @[Reg.scala 17:22]
    end
    if (leftFire) begin // @[Reg.scala 17:18]
      data_cf_trigger_frontendHit_0 <= rename_io_out_0_bits_cf_trigger_frontendHit_0; // @[Reg.scala 17:22]
    end
    if (leftFire) begin // @[Reg.scala 17:18]
      data_cf_trigger_frontendHit_1 <= rename_io_out_0_bits_cf_trigger_frontendHit_1; // @[Reg.scala 17:22]
    end
    if (leftFire) begin // @[Reg.scala 17:18]
      data_cf_trigger_frontendHit_2 <= rename_io_out_0_bits_cf_trigger_frontendHit_2; // @[Reg.scala 17:22]
    end
    if (leftFire) begin // @[Reg.scala 17:18]
      data_cf_trigger_frontendHit_3 <= rename_io_out_0_bits_cf_trigger_frontendHit_3; // @[Reg.scala 17:22]
    end
    if (leftFire) begin // @[Reg.scala 17:18]
      data_cf_trigger_backendEn_0 <= rename_io_out_0_bits_cf_trigger_backendEn_0; // @[Reg.scala 17:22]
    end
    if (leftFire) begin // @[Reg.scala 17:18]
      data_cf_trigger_backendEn_1 <= rename_io_out_0_bits_cf_trigger_backendEn_1; // @[Reg.scala 17:22]
    end
    if (leftFire) begin // @[Reg.scala 17:18]
      data_cf_pd_isRVC <= rename_io_out_0_bits_cf_pd_isRVC; // @[Reg.scala 17:22]
    end
    if (leftFire) begin // @[Reg.scala 17:18]
      data_cf_pd_brType <= rename_io_out_0_bits_cf_pd_brType; // @[Reg.scala 17:22]
    end
    if (leftFire) begin // @[Reg.scala 17:18]
      data_cf_pd_isCall <= rename_io_out_0_bits_cf_pd_isCall; // @[Reg.scala 17:22]
    end
    if (leftFire) begin // @[Reg.scala 17:18]
      data_cf_pd_isRet <= rename_io_out_0_bits_cf_pd_isRet; // @[Reg.scala 17:22]
    end
    if (leftFire) begin // @[Reg.scala 17:18]
      data_cf_pred_taken <= rename_io_out_0_bits_cf_pred_taken; // @[Reg.scala 17:22]
    end
    if (leftFire) begin // @[Reg.scala 17:18]
      data_cf_crossPageIPFFix <= rename_io_out_0_bits_cf_crossPageIPFFix; // @[Reg.scala 17:22]
    end
    if (leftFire) begin // @[Reg.scala 17:18]
      data_cf_storeSetHit <= rename_io_out_0_bits_cf_storeSetHit; // @[Reg.scala 17:22]
    end
    if (leftFire) begin // @[Reg.scala 17:18]
      data_cf_loadWaitStrict <= rename_io_out_0_bits_cf_loadWaitStrict; // @[Reg.scala 17:22]
    end
    if (leftFire) begin // @[Reg.scala 17:18]
      data_cf_ssid <= rename_io_out_0_bits_cf_ssid; // @[Reg.scala 17:22]
    end
    if (leftFire) begin // @[Reg.scala 17:18]
      data_cf_ftqPtr_flag <= rename_io_out_0_bits_cf_ftqPtr_flag; // @[Reg.scala 17:22]
    end
    if (leftFire) begin // @[Reg.scala 17:18]
      data_cf_ftqPtr_value <= rename_io_out_0_bits_cf_ftqPtr_value; // @[Reg.scala 17:22]
    end
    if (leftFire) begin // @[Reg.scala 17:18]
      data_cf_ftqOffset <= rename_io_out_0_bits_cf_ftqOffset; // @[Reg.scala 17:22]
    end
    if (leftFire) begin // @[Reg.scala 17:18]
      data_ctrl_srcType_0 <= rename_io_out_0_bits_ctrl_srcType_0; // @[Reg.scala 17:22]
    end
    if (leftFire) begin // @[Reg.scala 17:18]
      data_ctrl_srcType_1 <= rename_io_out_0_bits_ctrl_srcType_1; // @[Reg.scala 17:22]
    end
    if (leftFire) begin // @[Reg.scala 17:18]
      data_ctrl_srcType_2 <= rename_io_out_0_bits_ctrl_srcType_2; // @[Reg.scala 17:22]
    end
    if (leftFire) begin // @[Reg.scala 17:18]
      data_ctrl_ldest <= rename_io_out_0_bits_ctrl_ldest; // @[Reg.scala 17:22]
    end
    if (leftFire) begin // @[Reg.scala 17:18]
      data_ctrl_fuType <= rename_io_out_0_bits_ctrl_fuType; // @[Reg.scala 17:22]
    end
    if (leftFire) begin // @[Reg.scala 17:18]
      data_ctrl_fuOpType <= rename_io_out_0_bits_ctrl_fuOpType; // @[Reg.scala 17:22]
    end
    if (leftFire) begin // @[Reg.scala 17:18]
      data_ctrl_rfWen <= rename_io_out_0_bits_ctrl_rfWen; // @[Reg.scala 17:22]
    end
    if (leftFire) begin // @[Reg.scala 17:18]
      data_ctrl_fpWen <= rename_io_out_0_bits_ctrl_fpWen; // @[Reg.scala 17:22]
    end
    if (leftFire) begin // @[Reg.scala 17:18]
      data_ctrl_isXSTrap <= rename_io_out_0_bits_ctrl_isXSTrap; // @[Reg.scala 17:22]
    end
    if (leftFire) begin // @[Reg.scala 17:18]
      data_ctrl_noSpecExec <= rename_io_out_0_bits_ctrl_noSpecExec; // @[Reg.scala 17:22]
    end
    if (leftFire) begin // @[Reg.scala 17:18]
      data_ctrl_blockBackward <= rename_io_out_0_bits_ctrl_blockBackward; // @[Reg.scala 17:22]
    end
    if (leftFire) begin // @[Reg.scala 17:18]
      data_ctrl_flushPipe <= rename_io_out_0_bits_ctrl_flushPipe; // @[Reg.scala 17:22]
    end
    if (leftFire) begin // @[Reg.scala 17:18]
      data_ctrl_selImm <= rename_io_out_0_bits_ctrl_selImm; // @[Reg.scala 17:22]
    end
    if (leftFire) begin // @[Reg.scala 17:18]
      data_ctrl_imm <= rename_io_out_0_bits_ctrl_imm; // @[Reg.scala 17:22]
    end
    if (leftFire) begin // @[Reg.scala 17:18]
      data_ctrl_commitType <= rename_io_out_0_bits_ctrl_commitType; // @[Reg.scala 17:22]
    end
    if (leftFire) begin // @[Reg.scala 17:18]
      data_ctrl_fpu_isAddSub <= rename_io_out_0_bits_ctrl_fpu_isAddSub; // @[Reg.scala 17:22]
    end
    if (leftFire) begin // @[Reg.scala 17:18]
      data_ctrl_fpu_typeTagIn <= rename_io_out_0_bits_ctrl_fpu_typeTagIn; // @[Reg.scala 17:22]
    end
    if (leftFire) begin // @[Reg.scala 17:18]
      data_ctrl_fpu_typeTagOut <= rename_io_out_0_bits_ctrl_fpu_typeTagOut; // @[Reg.scala 17:22]
    end
    if (leftFire) begin // @[Reg.scala 17:18]
      data_ctrl_fpu_fromInt <= rename_io_out_0_bits_ctrl_fpu_fromInt; // @[Reg.scala 17:22]
    end
    if (leftFire) begin // @[Reg.scala 17:18]
      data_ctrl_fpu_wflags <= rename_io_out_0_bits_ctrl_fpu_wflags; // @[Reg.scala 17:22]
    end
    if (leftFire) begin // @[Reg.scala 17:18]
      data_ctrl_fpu_fpWen <= rename_io_out_0_bits_ctrl_fpu_fpWen; // @[Reg.scala 17:22]
    end
    if (leftFire) begin // @[Reg.scala 17:18]
      data_ctrl_fpu_fmaCmd <= rename_io_out_0_bits_ctrl_fpu_fmaCmd; // @[Reg.scala 17:22]
    end
    if (leftFire) begin // @[Reg.scala 17:18]
      data_ctrl_fpu_div <= rename_io_out_0_bits_ctrl_fpu_div; // @[Reg.scala 17:22]
    end
    if (leftFire) begin // @[Reg.scala 17:18]
      data_ctrl_fpu_sqrt <= rename_io_out_0_bits_ctrl_fpu_sqrt; // @[Reg.scala 17:22]
    end
    if (leftFire) begin // @[Reg.scala 17:18]
      data_ctrl_fpu_fcvt <= rename_io_out_0_bits_ctrl_fpu_fcvt; // @[Reg.scala 17:22]
    end
    if (leftFire) begin // @[Reg.scala 17:18]
      data_ctrl_fpu_typ <= rename_io_out_0_bits_ctrl_fpu_typ; // @[Reg.scala 17:22]
    end
    if (leftFire) begin // @[Reg.scala 17:18]
      data_ctrl_fpu_fmt <= rename_io_out_0_bits_ctrl_fpu_fmt; // @[Reg.scala 17:22]
    end
    if (leftFire) begin // @[Reg.scala 17:18]
      data_ctrl_fpu_ren3 <= rename_io_out_0_bits_ctrl_fpu_ren3; // @[Reg.scala 17:22]
    end
    if (leftFire) begin // @[Reg.scala 17:18]
      data_ctrl_fpu_rm <= rename_io_out_0_bits_ctrl_fpu_rm; // @[Reg.scala 17:22]
    end
    if (leftFire) begin // @[Reg.scala 17:18]
      data_ctrl_isMove <= rename_io_out_0_bits_ctrl_isMove; // @[Reg.scala 17:22]
    end
    if (leftFire) begin // @[Reg.scala 17:18]
      data_psrc_0 <= rename_io_out_0_bits_psrc_0; // @[Reg.scala 17:22]
    end
    if (leftFire) begin // @[Reg.scala 17:18]
      data_psrc_1 <= rename_io_out_0_bits_psrc_1; // @[Reg.scala 17:22]
    end
    if (leftFire) begin // @[Reg.scala 17:18]
      data_psrc_2 <= rename_io_out_0_bits_psrc_2; // @[Reg.scala 17:22]
    end
    if (leftFire) begin // @[Reg.scala 17:18]
      data_pdest <= rename_io_out_0_bits_pdest; // @[Reg.scala 17:22]
    end
    if (leftFire) begin // @[Reg.scala 17:18]
      data_old_pdest <= rename_io_out_0_bits_old_pdest; // @[Reg.scala 17:22]
    end
    if (leftFire) begin // @[Reg.scala 17:18]
      data_robIdx_flag <= rename_io_out_0_bits_robIdx_flag; // @[Reg.scala 17:22]
    end
    if (leftFire) begin // @[Reg.scala 17:18]
      data_robIdx_value <= rename_io_out_0_bits_robIdx_value; // @[Reg.scala 17:22]
    end
    if (leftFire) begin // @[Reg.scala 17:18]
      data_eliminatedMove <= rename_io_out_0_bits_eliminatedMove; // @[Reg.scala 17:22]
    end
    if (leftFire_1) begin // @[Reg.scala 17:18]
      data_1_cf_foldpc <= rename_io_out_1_bits_cf_foldpc; // @[Reg.scala 17:22]
    end
    if (leftFire_1) begin // @[Reg.scala 17:18]
      data_1_cf_exceptionVec_1 <= rename_io_out_1_bits_cf_exceptionVec_1; // @[Reg.scala 17:22]
    end
    if (leftFire_1) begin // @[Reg.scala 17:18]
      data_1_cf_exceptionVec_2 <= rename_io_out_1_bits_cf_exceptionVec_2; // @[Reg.scala 17:22]
    end
    if (leftFire_1) begin // @[Reg.scala 17:18]
      data_1_cf_exceptionVec_12 <= rename_io_out_1_bits_cf_exceptionVec_12; // @[Reg.scala 17:22]
    end
    if (leftFire_1) begin // @[Reg.scala 17:18]
      data_1_cf_trigger_frontendHit_0 <= rename_io_out_1_bits_cf_trigger_frontendHit_0; // @[Reg.scala 17:22]
    end
    if (leftFire_1) begin // @[Reg.scala 17:18]
      data_1_cf_trigger_frontendHit_1 <= rename_io_out_1_bits_cf_trigger_frontendHit_1; // @[Reg.scala 17:22]
    end
    if (leftFire_1) begin // @[Reg.scala 17:18]
      data_1_cf_trigger_frontendHit_2 <= rename_io_out_1_bits_cf_trigger_frontendHit_2; // @[Reg.scala 17:22]
    end
    if (leftFire_1) begin // @[Reg.scala 17:18]
      data_1_cf_trigger_frontendHit_3 <= rename_io_out_1_bits_cf_trigger_frontendHit_3; // @[Reg.scala 17:22]
    end
    if (leftFire_1) begin // @[Reg.scala 17:18]
      data_1_cf_trigger_backendEn_0 <= rename_io_out_1_bits_cf_trigger_backendEn_0; // @[Reg.scala 17:22]
    end
    if (leftFire_1) begin // @[Reg.scala 17:18]
      data_1_cf_trigger_backendEn_1 <= rename_io_out_1_bits_cf_trigger_backendEn_1; // @[Reg.scala 17:22]
    end
    if (leftFire_1) begin // @[Reg.scala 17:18]
      data_1_cf_pd_isRVC <= rename_io_out_1_bits_cf_pd_isRVC; // @[Reg.scala 17:22]
    end
    if (leftFire_1) begin // @[Reg.scala 17:18]
      data_1_cf_pd_brType <= rename_io_out_1_bits_cf_pd_brType; // @[Reg.scala 17:22]
    end
    if (leftFire_1) begin // @[Reg.scala 17:18]
      data_1_cf_pd_isCall <= rename_io_out_1_bits_cf_pd_isCall; // @[Reg.scala 17:22]
    end
    if (leftFire_1) begin // @[Reg.scala 17:18]
      data_1_cf_pd_isRet <= rename_io_out_1_bits_cf_pd_isRet; // @[Reg.scala 17:22]
    end
    if (leftFire_1) begin // @[Reg.scala 17:18]
      data_1_cf_pred_taken <= rename_io_out_1_bits_cf_pred_taken; // @[Reg.scala 17:22]
    end
    if (leftFire_1) begin // @[Reg.scala 17:18]
      data_1_cf_crossPageIPFFix <= rename_io_out_1_bits_cf_crossPageIPFFix; // @[Reg.scala 17:22]
    end
    if (leftFire_1) begin // @[Reg.scala 17:18]
      data_1_cf_storeSetHit <= rename_io_out_1_bits_cf_storeSetHit; // @[Reg.scala 17:22]
    end
    if (leftFire_1) begin // @[Reg.scala 17:18]
      data_1_cf_loadWaitStrict <= rename_io_out_1_bits_cf_loadWaitStrict; // @[Reg.scala 17:22]
    end
    if (leftFire_1) begin // @[Reg.scala 17:18]
      data_1_cf_ssid <= rename_io_out_1_bits_cf_ssid; // @[Reg.scala 17:22]
    end
    if (leftFire_1) begin // @[Reg.scala 17:18]
      data_1_cf_ftqPtr_flag <= rename_io_out_1_bits_cf_ftqPtr_flag; // @[Reg.scala 17:22]
    end
    if (leftFire_1) begin // @[Reg.scala 17:18]
      data_1_cf_ftqPtr_value <= rename_io_out_1_bits_cf_ftqPtr_value; // @[Reg.scala 17:22]
    end
    if (leftFire_1) begin // @[Reg.scala 17:18]
      data_1_cf_ftqOffset <= rename_io_out_1_bits_cf_ftqOffset; // @[Reg.scala 17:22]
    end
    if (leftFire_1) begin // @[Reg.scala 17:18]
      data_1_ctrl_srcType_0 <= rename_io_out_1_bits_ctrl_srcType_0; // @[Reg.scala 17:22]
    end
    if (leftFire_1) begin // @[Reg.scala 17:18]
      data_1_ctrl_srcType_1 <= rename_io_out_1_bits_ctrl_srcType_1; // @[Reg.scala 17:22]
    end
    if (leftFire_1) begin // @[Reg.scala 17:18]
      data_1_ctrl_srcType_2 <= rename_io_out_1_bits_ctrl_srcType_2; // @[Reg.scala 17:22]
    end
    if (leftFire_1) begin // @[Reg.scala 17:18]
      data_1_ctrl_ldest <= rename_io_out_1_bits_ctrl_ldest; // @[Reg.scala 17:22]
    end
    if (leftFire_1) begin // @[Reg.scala 17:18]
      data_1_ctrl_fuType <= rename_io_out_1_bits_ctrl_fuType; // @[Reg.scala 17:22]
    end
    if (leftFire_1) begin // @[Reg.scala 17:18]
      data_1_ctrl_fuOpType <= rename_io_out_1_bits_ctrl_fuOpType; // @[Reg.scala 17:22]
    end
    if (leftFire_1) begin // @[Reg.scala 17:18]
      data_1_ctrl_rfWen <= rename_io_out_1_bits_ctrl_rfWen; // @[Reg.scala 17:22]
    end
    if (leftFire_1) begin // @[Reg.scala 17:18]
      data_1_ctrl_fpWen <= rename_io_out_1_bits_ctrl_fpWen; // @[Reg.scala 17:22]
    end
    if (leftFire_1) begin // @[Reg.scala 17:18]
      data_1_ctrl_isXSTrap <= rename_io_out_1_bits_ctrl_isXSTrap; // @[Reg.scala 17:22]
    end
    if (leftFire_1) begin // @[Reg.scala 17:18]
      data_1_ctrl_noSpecExec <= rename_io_out_1_bits_ctrl_noSpecExec; // @[Reg.scala 17:22]
    end
    if (leftFire_1) begin // @[Reg.scala 17:18]
      data_1_ctrl_blockBackward <= rename_io_out_1_bits_ctrl_blockBackward; // @[Reg.scala 17:22]
    end
    if (leftFire_1) begin // @[Reg.scala 17:18]
      data_1_ctrl_flushPipe <= rename_io_out_1_bits_ctrl_flushPipe; // @[Reg.scala 17:22]
    end
    if (leftFire_1) begin // @[Reg.scala 17:18]
      data_1_ctrl_selImm <= rename_io_out_1_bits_ctrl_selImm; // @[Reg.scala 17:22]
    end
    if (leftFire_1) begin // @[Reg.scala 17:18]
      data_1_ctrl_imm <= rename_io_out_1_bits_ctrl_imm; // @[Reg.scala 17:22]
    end
    if (leftFire_1) begin // @[Reg.scala 17:18]
      data_1_ctrl_fpu_isAddSub <= rename_io_out_1_bits_ctrl_fpu_isAddSub; // @[Reg.scala 17:22]
    end
    if (leftFire_1) begin // @[Reg.scala 17:18]
      data_1_ctrl_fpu_typeTagIn <= rename_io_out_1_bits_ctrl_fpu_typeTagIn; // @[Reg.scala 17:22]
    end
    if (leftFire_1) begin // @[Reg.scala 17:18]
      data_1_ctrl_fpu_typeTagOut <= rename_io_out_1_bits_ctrl_fpu_typeTagOut; // @[Reg.scala 17:22]
    end
    if (leftFire_1) begin // @[Reg.scala 17:18]
      data_1_ctrl_fpu_fromInt <= rename_io_out_1_bits_ctrl_fpu_fromInt; // @[Reg.scala 17:22]
    end
    if (leftFire_1) begin // @[Reg.scala 17:18]
      data_1_ctrl_fpu_wflags <= rename_io_out_1_bits_ctrl_fpu_wflags; // @[Reg.scala 17:22]
    end
    if (leftFire_1) begin // @[Reg.scala 17:18]
      data_1_ctrl_fpu_fpWen <= rename_io_out_1_bits_ctrl_fpu_fpWen; // @[Reg.scala 17:22]
    end
    if (leftFire_1) begin // @[Reg.scala 17:18]
      data_1_ctrl_fpu_fmaCmd <= rename_io_out_1_bits_ctrl_fpu_fmaCmd; // @[Reg.scala 17:22]
    end
    if (leftFire_1) begin // @[Reg.scala 17:18]
      data_1_ctrl_fpu_div <= rename_io_out_1_bits_ctrl_fpu_div; // @[Reg.scala 17:22]
    end
    if (leftFire_1) begin // @[Reg.scala 17:18]
      data_1_ctrl_fpu_sqrt <= rename_io_out_1_bits_ctrl_fpu_sqrt; // @[Reg.scala 17:22]
    end
    if (leftFire_1) begin // @[Reg.scala 17:18]
      data_1_ctrl_fpu_fcvt <= rename_io_out_1_bits_ctrl_fpu_fcvt; // @[Reg.scala 17:22]
    end
    if (leftFire_1) begin // @[Reg.scala 17:18]
      data_1_ctrl_fpu_typ <= rename_io_out_1_bits_ctrl_fpu_typ; // @[Reg.scala 17:22]
    end
    if (leftFire_1) begin // @[Reg.scala 17:18]
      data_1_ctrl_fpu_fmt <= rename_io_out_1_bits_ctrl_fpu_fmt; // @[Reg.scala 17:22]
    end
    if (leftFire_1) begin // @[Reg.scala 17:18]
      data_1_ctrl_fpu_ren3 <= rename_io_out_1_bits_ctrl_fpu_ren3; // @[Reg.scala 17:22]
    end
    if (leftFire_1) begin // @[Reg.scala 17:18]
      data_1_ctrl_fpu_rm <= rename_io_out_1_bits_ctrl_fpu_rm; // @[Reg.scala 17:22]
    end
    if (leftFire_1) begin // @[Reg.scala 17:18]
      data_1_ctrl_isMove <= rename_io_out_1_bits_ctrl_isMove; // @[Reg.scala 17:22]
    end
    if (leftFire_1) begin // @[Reg.scala 17:18]
      data_1_psrc_0 <= rename_io_out_1_bits_psrc_0; // @[Reg.scala 17:22]
    end
    if (leftFire_1) begin // @[Reg.scala 17:18]
      data_1_psrc_1 <= rename_io_out_1_bits_psrc_1; // @[Reg.scala 17:22]
    end
    if (leftFire_1) begin // @[Reg.scala 17:18]
      data_1_psrc_2 <= rename_io_out_1_bits_psrc_2; // @[Reg.scala 17:22]
    end
    if (leftFire_1) begin // @[Reg.scala 17:18]
      data_1_pdest <= rename_io_out_1_bits_pdest; // @[Reg.scala 17:22]
    end
    if (leftFire_1) begin // @[Reg.scala 17:18]
      data_1_old_pdest <= rename_io_out_1_bits_old_pdest; // @[Reg.scala 17:22]
    end
    if (leftFire_1) begin // @[Reg.scala 17:18]
      data_1_robIdx_flag <= rename_io_out_1_bits_robIdx_flag; // @[Reg.scala 17:22]
    end
    if (leftFire_1) begin // @[Reg.scala 17:18]
      data_1_robIdx_value <= rename_io_out_1_bits_robIdx_value; // @[Reg.scala 17:22]
    end
    if (leftFire_1) begin // @[Reg.scala 17:18]
      data_1_eliminatedMove <= rename_io_out_1_bits_eliminatedMove; // @[Reg.scala 17:22]
    end
    dispatch_io_singleStep_REG <= io_csrCtrl_singlestep; // @[CtrlBlock.scala 501:36]
    jumpPcRead0_REG <= intDq_io_deqNext_0_cf_ftqOffset; // @[CtrlBlock.scala 543:52]
    read_from_newest_entry_REG_flag <= io_dispatch_0_bits_cf_ftqPtr_flag; // @[CtrlBlock.scala 546:30]
    read_from_newest_entry_REG_value <= io_dispatch_0_bits_cf_ftqPtr_value; // @[CtrlBlock.scala 546:30]
    read_from_newest_entry_REG_1_flag <= io_frontend_fromFtq_newest_entry_ptr_flag; // @[CtrlBlock.scala 551:70]
    read_from_newest_entry_REG_1_value <= io_frontend_fromFtq_newest_entry_ptr_value; // @[CtrlBlock.scala 551:70]
    io_jalr_target_REG <= io_frontend_fromFtq_newest_entry_target; // @[CtrlBlock.scala 552:56]
    sources_source_exuOutput_3_valid_REG <= io_writeback_0_3_valid & ~_sources_exuOutput_3_valid_T_7; // @[CtrlBlock.scala 255:43]
    sources_source_exuOutput_3_bits_REG_uop_cf_exceptionVec_2 <= io_writeback_0_3_bits_uop_cf_exceptionVec_2; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_3_bits_REG_uop_cf_exceptionVec_3 <= io_writeback_0_3_bits_uop_cf_exceptionVec_3; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_3_bits_REG_uop_cf_exceptionVec_8 <= io_writeback_0_3_bits_uop_cf_exceptionVec_8; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_3_bits_REG_uop_cf_exceptionVec_9 <= io_writeback_0_3_bits_uop_cf_exceptionVec_9; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_3_bits_REG_uop_cf_exceptionVec_11 <= io_writeback_0_3_bits_uop_cf_exceptionVec_11; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_3_bits_REG_uop_ctrl_flushPipe <= io_writeback_0_3_bits_uop_ctrl_flushPipe; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_3_bits_REG_uop_robIdx_flag <= io_writeback_0_3_bits_uop_robIdx_flag; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_3_bits_REG_uop_robIdx_value <= io_writeback_0_3_bits_uop_robIdx_value; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_3_bits_REG_fflags <= io_writeback_0_3_bits_fflags; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_4_valid_REG <= io_writeback_0_4_valid & ~_sources_exuOutput_4_valid_T_7; // @[CtrlBlock.scala 255:43]
    sources_source_exuOutput_4_bits_REG_uop_robIdx_value <= io_writeback_0_4_bits_uop_robIdx_value; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_4_bits_REG_fflags <= io_writeback_0_4_bits_fflags; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_5_valid_REG <= io_writeback_0_5_valid & ~_sources_exuOutput_5_valid_T_7; // @[CtrlBlock.scala 255:43]
    sources_source_exuOutput_5_bits_REG_uop_robIdx_value <= io_writeback_0_5_bits_uop_robIdx_value; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_5_bits_REG_fflags <= io_writeback_0_5_bits_fflags; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_6_valid_REG <= io_writeback_0_6_valid & ~_sources_exuOutput_6_valid_T_7; // @[CtrlBlock.scala 255:43]
    sources_source_exuOutput_6_bits_REG_uop_cf_exceptionVec_4 <= io_writeback_0_6_bits_uop_cf_exceptionVec_4; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_6_bits_REG_uop_cf_exceptionVec_5 <= io_writeback_0_6_bits_uop_cf_exceptionVec_5; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_6_bits_REG_uop_cf_exceptionVec_13 <= io_writeback_0_6_bits_uop_cf_exceptionVec_13; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_6_bits_REG_uop_cf_trigger_backendHit_0 <= io_writeback_0_6_bits_uop_cf_trigger_backendHit_0
      ; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_6_bits_REG_uop_cf_trigger_backendHit_1 <= io_writeback_0_6_bits_uop_cf_trigger_backendHit_1
      ; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_6_bits_REG_uop_cf_trigger_backendHit_2 <= io_writeback_0_6_bits_uop_cf_trigger_backendHit_2
      ; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_6_bits_REG_uop_cf_trigger_backendHit_3 <= io_writeback_0_6_bits_uop_cf_trigger_backendHit_3
      ; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_6_bits_REG_uop_cf_trigger_backendHit_4 <= io_writeback_0_6_bits_uop_cf_trigger_backendHit_4
      ; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_6_bits_REG_uop_cf_trigger_backendHit_5 <= io_writeback_0_6_bits_uop_cf_trigger_backendHit_5
      ; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_6_bits_REG_uop_ctrl_flushPipe <= io_writeback_0_6_bits_uop_ctrl_flushPipe; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_6_bits_REG_uop_ctrl_replayInst <= io_writeback_0_6_bits_uop_ctrl_replayInst; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_6_bits_REG_uop_robIdx_flag <= io_writeback_0_6_bits_uop_robIdx_flag; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_6_bits_REG_uop_robIdx_value <= io_writeback_0_6_bits_uop_robIdx_value; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_7_valid_REG <= io_writeback_0_7_valid & ~_sources_exuOutput_7_valid_T_7; // @[CtrlBlock.scala 255:43]
    sources_source_exuOutput_7_bits_REG_uop_cf_exceptionVec_4 <= io_writeback_0_7_bits_uop_cf_exceptionVec_4; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_7_bits_REG_uop_cf_exceptionVec_5 <= io_writeback_0_7_bits_uop_cf_exceptionVec_5; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_7_bits_REG_uop_cf_exceptionVec_13 <= io_writeback_0_7_bits_uop_cf_exceptionVec_13; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_7_bits_REG_uop_cf_trigger_backendHit_0 <= io_writeback_0_7_bits_uop_cf_trigger_backendHit_0
      ; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_7_bits_REG_uop_cf_trigger_backendHit_1 <= io_writeback_0_7_bits_uop_cf_trigger_backendHit_1
      ; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_7_bits_REG_uop_cf_trigger_backendHit_2 <= io_writeback_0_7_bits_uop_cf_trigger_backendHit_2
      ; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_7_bits_REG_uop_cf_trigger_backendHit_3 <= io_writeback_0_7_bits_uop_cf_trigger_backendHit_3
      ; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_7_bits_REG_uop_cf_trigger_backendHit_4 <= io_writeback_0_7_bits_uop_cf_trigger_backendHit_4
      ; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_7_bits_REG_uop_cf_trigger_backendHit_5 <= io_writeback_0_7_bits_uop_cf_trigger_backendHit_5
      ; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_7_bits_REG_uop_ctrl_flushPipe <= io_writeback_0_7_bits_uop_ctrl_flushPipe; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_7_bits_REG_uop_ctrl_replayInst <= io_writeback_0_7_bits_uop_ctrl_replayInst; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_7_bits_REG_uop_robIdx_flag <= io_writeback_0_7_bits_uop_robIdx_flag; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_7_bits_REG_uop_robIdx_value <= io_writeback_0_7_bits_uop_robIdx_value; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_8_valid_REG <= io_writeback_0_8_valid & ~_sources_exuOutput_8_valid_T_7; // @[CtrlBlock.scala 255:43]
    sources_source_exuOutput_8_bits_REG_uop_cf_exceptionVec_4 <= io_writeback_0_8_bits_uop_cf_exceptionVec_4; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_8_bits_REG_uop_cf_exceptionVec_5 <= io_writeback_0_8_bits_uop_cf_exceptionVec_5; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_8_bits_REG_uop_cf_exceptionVec_6 <= io_writeback_0_8_bits_uop_cf_exceptionVec_6; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_8_bits_REG_uop_cf_exceptionVec_7 <= io_writeback_0_8_bits_uop_cf_exceptionVec_7; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_8_bits_REG_uop_cf_exceptionVec_13 <= io_writeback_0_8_bits_uop_cf_exceptionVec_13; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_8_bits_REG_uop_cf_exceptionVec_15 <= io_writeback_0_8_bits_uop_cf_exceptionVec_15; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_8_bits_REG_uop_cf_trigger_backendHit_0 <= io_writeback_0_8_bits_uop_cf_trigger_backendHit_0
      ; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_8_bits_REG_uop_cf_trigger_backendHit_1 <= io_writeback_0_8_bits_uop_cf_trigger_backendHit_1
      ; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_8_bits_REG_uop_cf_trigger_backendHit_2 <= io_writeback_0_8_bits_uop_cf_trigger_backendHit_2
      ; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_8_bits_REG_uop_cf_trigger_backendHit_3 <= io_writeback_0_8_bits_uop_cf_trigger_backendHit_3
      ; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_8_bits_REG_uop_cf_trigger_backendHit_4 <= io_writeback_0_8_bits_uop_cf_trigger_backendHit_4
      ; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_8_bits_REG_uop_cf_trigger_backendHit_5 <= io_writeback_0_8_bits_uop_cf_trigger_backendHit_5
      ; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_8_bits_REG_uop_robIdx_flag <= io_writeback_0_8_bits_uop_robIdx_flag; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_8_bits_REG_uop_robIdx_value <= io_writeback_0_8_bits_uop_robIdx_value; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_9_valid_REG <= io_writeback_0_9_valid & ~_sources_exuOutput_9_valid_T_7; // @[CtrlBlock.scala 255:43]
    sources_source_exuOutput_9_bits_REG_uop_cf_exceptionVec_6 <= io_writeback_0_9_bits_uop_cf_exceptionVec_6; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_9_bits_REG_uop_cf_exceptionVec_7 <= io_writeback_0_9_bits_uop_cf_exceptionVec_7; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_9_bits_REG_uop_cf_exceptionVec_15 <= io_writeback_0_9_bits_uop_cf_exceptionVec_15; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_9_bits_REG_uop_cf_trigger_backendHit_0 <= io_writeback_0_9_bits_uop_cf_trigger_backendHit_0
      ; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_9_bits_REG_uop_cf_trigger_backendHit_1 <= io_writeback_0_9_bits_uop_cf_trigger_backendHit_1
      ; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_9_bits_REG_uop_cf_trigger_backendHit_4 <= io_writeback_0_9_bits_uop_cf_trigger_backendHit_4
      ; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_9_bits_REG_uop_robIdx_flag <= io_writeback_0_9_bits_uop_robIdx_flag; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_9_bits_REG_uop_robIdx_value <= io_writeback_0_9_bits_uop_robIdx_value; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_0_valid_REG_3 <= io_writeback_1_0_valid & ~_sources_exuOutput_0_valid_T_17; // @[CtrlBlock.scala 255:43]
    sources_source_exuOutput_0_bits_REG_3_uop_robIdx_value <= io_writeback_1_0_bits_uop_robIdx_value; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_0_bits_REG_3_redirectValid <= io_writeback_1_0_bits_redirectValid; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_0_bits_REG_3_redirect_cfiUpdate_isMisPred <=
      io_writeback_1_0_bits_redirect_cfiUpdate_isMisPred; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_1_valid_REG_3 <= io_writeback_1_1_valid & ~_sources_exuOutput_1_valid_T_17; // @[CtrlBlock.scala 255:43]
    sources_source_exuOutput_1_bits_REG_3_uop_robIdx_value <= io_writeback_1_1_bits_uop_robIdx_value; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_1_bits_REG_3_redirectValid <= io_writeback_1_1_bits_redirectValid; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_1_bits_REG_3_redirect_cfiUpdate_isMisPred <=
      io_writeback_1_1_bits_redirect_cfiUpdate_isMisPred; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_2_valid_REG_3 <= io_writeback_1_2_valid & ~_sources_exuOutput_2_valid_T_17; // @[CtrlBlock.scala 255:43]
    sources_source_exuOutput_2_bits_REG_3_uop_cf_exceptionVec_4 <= io_writeback_1_2_bits_uop_cf_exceptionVec_4; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_2_bits_REG_3_uop_cf_exceptionVec_5 <= io_writeback_1_2_bits_uop_cf_exceptionVec_5; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_2_bits_REG_3_uop_cf_exceptionVec_13 <= io_writeback_1_2_bits_uop_cf_exceptionVec_13; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_2_bits_REG_3_uop_cf_trigger_backendHit_0 <=
      io_writeback_1_2_bits_uop_cf_trigger_backendHit_0; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_2_bits_REG_3_uop_cf_trigger_backendHit_1 <=
      io_writeback_1_2_bits_uop_cf_trigger_backendHit_1; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_2_bits_REG_3_uop_cf_trigger_backendHit_2 <=
      io_writeback_1_2_bits_uop_cf_trigger_backendHit_2; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_2_bits_REG_3_uop_cf_trigger_backendHit_3 <=
      io_writeback_1_2_bits_uop_cf_trigger_backendHit_3; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_2_bits_REG_3_uop_cf_trigger_backendHit_4 <=
      io_writeback_1_2_bits_uop_cf_trigger_backendHit_4; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_2_bits_REG_3_uop_cf_trigger_backendHit_5 <=
      io_writeback_1_2_bits_uop_cf_trigger_backendHit_5; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_2_bits_REG_3_uop_ctrl_flushPipe <= io_writeback_1_2_bits_uop_ctrl_flushPipe; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_2_bits_REG_3_uop_ctrl_replayInst <= io_writeback_1_2_bits_uop_ctrl_replayInst; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_2_bits_REG_3_uop_robIdx_value <= io_writeback_1_2_bits_uop_robIdx_value; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_2_bits_REG_3_debug_isMMIO <= io_writeback_1_2_bits_debug_isMMIO; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_3_valid_REG_3 <= io_writeback_1_3_valid & ~_sources_exuOutput_3_valid_T_17; // @[CtrlBlock.scala 255:43]
    sources_source_exuOutput_3_bits_REG_3_uop_cf_exceptionVec_4 <= io_writeback_1_3_bits_uop_cf_exceptionVec_4; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_3_bits_REG_3_uop_cf_exceptionVec_5 <= io_writeback_1_3_bits_uop_cf_exceptionVec_5; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_3_bits_REG_3_uop_cf_exceptionVec_13 <= io_writeback_1_3_bits_uop_cf_exceptionVec_13; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_3_bits_REG_3_uop_cf_trigger_backendHit_0 <=
      io_writeback_1_3_bits_uop_cf_trigger_backendHit_0; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_3_bits_REG_3_uop_cf_trigger_backendHit_1 <=
      io_writeback_1_3_bits_uop_cf_trigger_backendHit_1; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_3_bits_REG_3_uop_cf_trigger_backendHit_2 <=
      io_writeback_1_3_bits_uop_cf_trigger_backendHit_2; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_3_bits_REG_3_uop_cf_trigger_backendHit_3 <=
      io_writeback_1_3_bits_uop_cf_trigger_backendHit_3; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_3_bits_REG_3_uop_cf_trigger_backendHit_4 <=
      io_writeback_1_3_bits_uop_cf_trigger_backendHit_4; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_3_bits_REG_3_uop_cf_trigger_backendHit_5 <=
      io_writeback_1_3_bits_uop_cf_trigger_backendHit_5; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_3_bits_REG_3_uop_ctrl_flushPipe <= io_writeback_1_3_bits_uop_ctrl_flushPipe; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_3_bits_REG_3_uop_ctrl_replayInst <= io_writeback_1_3_bits_uop_ctrl_replayInst; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_3_bits_REG_3_uop_robIdx_value <= io_writeback_1_3_bits_uop_robIdx_value; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_3_bits_REG_3_debug_isMMIO <= io_writeback_1_3_bits_debug_isMMIO; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_4_valid_REG_3 <= io_writeback_1_4_valid & ~_sources_exuOutput_4_valid_T_17; // @[CtrlBlock.scala 255:43]
    sources_source_exuOutput_4_bits_REG_3_uop_cf_exceptionVec_2 <= io_writeback_1_4_bits_uop_cf_exceptionVec_2; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_4_bits_REG_3_uop_cf_exceptionVec_3 <= io_writeback_1_4_bits_uop_cf_exceptionVec_3; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_4_bits_REG_3_uop_cf_exceptionVec_8 <= io_writeback_1_4_bits_uop_cf_exceptionVec_8; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_4_bits_REG_3_uop_cf_exceptionVec_9 <= io_writeback_1_4_bits_uop_cf_exceptionVec_9; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_4_bits_REG_3_uop_cf_exceptionVec_11 <= io_writeback_1_4_bits_uop_cf_exceptionVec_11; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_4_bits_REG_3_uop_ctrl_flushPipe <= io_writeback_1_4_bits_uop_ctrl_flushPipe; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_4_bits_REG_3_uop_robIdx_value <= io_writeback_1_4_bits_uop_robIdx_value; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_4_bits_REG_3_redirectValid <= io_writeback_1_4_bits_redirectValid; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_4_bits_REG_3_redirect_cfiUpdate_isMisPred <=
      io_writeback_1_4_bits_redirect_cfiUpdate_isMisPred; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_4_bits_REG_3_debug_isPerfCnt <= io_writeback_1_4_bits_debug_isPerfCnt; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_5_valid_REG_3 <= io_writeback_1_5_valid & ~_sources_exuOutput_5_valid_T_17; // @[CtrlBlock.scala 255:43]
    sources_source_exuOutput_5_bits_REG_3_uop_cf_trigger_backendHit_0 <=
      io_writeback_1_5_bits_uop_cf_trigger_backendHit_0; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_5_bits_REG_3_uop_cf_trigger_backendHit_1 <=
      io_writeback_1_5_bits_uop_cf_trigger_backendHit_1; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_5_bits_REG_3_uop_cf_trigger_backendHit_2 <=
      io_writeback_1_5_bits_uop_cf_trigger_backendHit_2; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_5_bits_REG_3_uop_cf_trigger_backendHit_3 <=
      io_writeback_1_5_bits_uop_cf_trigger_backendHit_3; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_5_bits_REG_3_uop_cf_trigger_backendHit_4 <=
      io_writeback_1_5_bits_uop_cf_trigger_backendHit_4; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_5_bits_REG_3_uop_cf_trigger_backendHit_5 <=
      io_writeback_1_5_bits_uop_cf_trigger_backendHit_5; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_5_bits_REG_3_uop_robIdx_value <= io_writeback_1_5_bits_uop_robIdx_value; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_6_valid_REG_3 <= io_writeback_1_6_valid & ~_sources_exuOutput_6_valid_T_17; // @[CtrlBlock.scala 255:43]
    sources_source_exuOutput_6_bits_REG_3_uop_cf_exceptionVec_2 <= io_writeback_1_6_bits_uop_cf_exceptionVec_2; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_6_bits_REG_3_uop_cf_exceptionVec_3 <= io_writeback_1_6_bits_uop_cf_exceptionVec_3; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_6_bits_REG_3_uop_cf_exceptionVec_8 <= io_writeback_1_6_bits_uop_cf_exceptionVec_8; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_6_bits_REG_3_uop_cf_exceptionVec_9 <= io_writeback_1_6_bits_uop_cf_exceptionVec_9; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_6_bits_REG_3_uop_cf_exceptionVec_11 <= io_writeback_1_6_bits_uop_cf_exceptionVec_11; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_6_bits_REG_3_uop_ctrl_flushPipe <= io_writeback_1_6_bits_uop_ctrl_flushPipe; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_6_bits_REG_3_uop_robIdx_value <= io_writeback_1_6_bits_uop_robIdx_value; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_6_bits_REG_3_redirectValid <= io_writeback_1_6_bits_redirectValid; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_6_bits_REG_3_redirect_cfiUpdate_isMisPred <=
      io_writeback_1_6_bits_redirect_cfiUpdate_isMisPred; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_6_bits_REG_3_debug_isPerfCnt <= io_writeback_1_6_bits_debug_isPerfCnt; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_7_valid_REG_3 <= io_writeback_1_7_valid & ~_sources_exuOutput_7_valid_T_17; // @[CtrlBlock.scala 255:43]
    sources_source_exuOutput_7_bits_REG_3_uop_cf_exceptionVec_4 <= io_writeback_1_7_bits_uop_cf_exceptionVec_4; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_7_bits_REG_3_uop_cf_exceptionVec_5 <= io_writeback_1_7_bits_uop_cf_exceptionVec_5; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_7_bits_REG_3_uop_cf_exceptionVec_6 <= io_writeback_1_7_bits_uop_cf_exceptionVec_6; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_7_bits_REG_3_uop_cf_exceptionVec_7 <= io_writeback_1_7_bits_uop_cf_exceptionVec_7; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_7_bits_REG_3_uop_cf_exceptionVec_13 <= io_writeback_1_7_bits_uop_cf_exceptionVec_13; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_7_bits_REG_3_uop_cf_exceptionVec_15 <= io_writeback_1_7_bits_uop_cf_exceptionVec_15; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_7_bits_REG_3_uop_cf_trigger_backendHit_0 <=
      io_writeback_1_7_bits_uop_cf_trigger_backendHit_0; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_7_bits_REG_3_uop_cf_trigger_backendHit_1 <=
      io_writeback_1_7_bits_uop_cf_trigger_backendHit_1; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_7_bits_REG_3_uop_cf_trigger_backendHit_2 <=
      io_writeback_1_7_bits_uop_cf_trigger_backendHit_2; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_7_bits_REG_3_uop_cf_trigger_backendHit_3 <=
      io_writeback_1_7_bits_uop_cf_trigger_backendHit_3; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_7_bits_REG_3_uop_cf_trigger_backendHit_4 <=
      io_writeback_1_7_bits_uop_cf_trigger_backendHit_4; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_7_bits_REG_3_uop_cf_trigger_backendHit_5 <=
      io_writeback_1_7_bits_uop_cf_trigger_backendHit_5; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_7_bits_REG_3_uop_robIdx_value <= io_writeback_1_7_bits_uop_robIdx_value; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_7_bits_REG_3_redirectValid <= io_writeback_1_7_bits_redirectValid; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_7_bits_REG_3_redirect_cfiUpdate_isMisPred <=
      io_writeback_1_7_bits_redirect_cfiUpdate_isMisPred; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_7_bits_REG_3_debug_isMMIO <= io_writeback_1_7_bits_debug_isMMIO; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_7_bits_REG_3_debug_isPerfCnt <= io_writeback_1_7_bits_debug_isPerfCnt; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_8_valid_REG_3 <= io_writeback_1_8_valid & ~_sources_exuOutput_8_valid_T_17; // @[CtrlBlock.scala 255:43]
    sources_source_exuOutput_8_bits_REG_3_uop_cf_exceptionVec_4 <= io_writeback_1_8_bits_uop_cf_exceptionVec_4; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_8_bits_REG_3_uop_cf_exceptionVec_5 <= io_writeback_1_8_bits_uop_cf_exceptionVec_5; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_8_bits_REG_3_uop_cf_exceptionVec_6 <= io_writeback_1_8_bits_uop_cf_exceptionVec_6; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_8_bits_REG_3_uop_cf_exceptionVec_7 <= io_writeback_1_8_bits_uop_cf_exceptionVec_7; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_8_bits_REG_3_uop_cf_exceptionVec_13 <= io_writeback_1_8_bits_uop_cf_exceptionVec_13; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_8_bits_REG_3_uop_cf_exceptionVec_15 <= io_writeback_1_8_bits_uop_cf_exceptionVec_15; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_8_bits_REG_3_uop_cf_trigger_backendHit_0 <=
      io_writeback_1_8_bits_uop_cf_trigger_backendHit_0; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_8_bits_REG_3_uop_cf_trigger_backendHit_1 <=
      io_writeback_1_8_bits_uop_cf_trigger_backendHit_1; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_8_bits_REG_3_uop_cf_trigger_backendHit_2 <=
      io_writeback_1_8_bits_uop_cf_trigger_backendHit_2; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_8_bits_REG_3_uop_cf_trigger_backendHit_3 <=
      io_writeback_1_8_bits_uop_cf_trigger_backendHit_3; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_8_bits_REG_3_uop_cf_trigger_backendHit_4 <=
      io_writeback_1_8_bits_uop_cf_trigger_backendHit_4; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_8_bits_REG_3_uop_cf_trigger_backendHit_5 <=
      io_writeback_1_8_bits_uop_cf_trigger_backendHit_5; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_8_bits_REG_3_uop_robIdx_value <= io_writeback_1_8_bits_uop_robIdx_value; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_8_bits_REG_3_redirectValid <= io_writeback_1_8_bits_redirectValid; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_8_bits_REG_3_redirect_cfiUpdate_isMisPred <=
      io_writeback_1_8_bits_redirect_cfiUpdate_isMisPred; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_8_bits_REG_3_debug_isMMIO <= io_writeback_1_8_bits_debug_isMMIO; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_8_bits_REG_3_debug_isPerfCnt <= io_writeback_1_8_bits_debug_isPerfCnt; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_9_valid_REG_3 <= io_writeback_1_9_valid & ~_sources_exuOutput_9_valid_T_17; // @[CtrlBlock.scala 255:43]
    sources_source_exuOutput_9_bits_REG_3_uop_robIdx_value <= io_writeback_1_9_bits_uop_robIdx_value; // @[CtrlBlock.scala 256:32]
    sources_source_exuOutput_10_valid_REG_3 <= io_writeback_1_10_valid & ~_sources_exuOutput_10_valid_T_17; // @[CtrlBlock.scala 255:43]
    sources_source_exuOutput_10_bits_REG_3_uop_robIdx_value <= io_writeback_1_10_bits_uop_robIdx_value; // @[CtrlBlock.scala 256:32]
    io_robio_toCSR_perfinfo_retiredInstr_REG <= rob_io_csr_perfinfo_retiredInstr; // @[CtrlBlock.scala 571:50]
    pfevent_io_distribute_csr_REG_wvalid <= io_csrCtrl_distribute_csr_wvalid; // @[CtrlBlock.scala 586:39]
    pfevent_io_distribute_csr_REG_waddr <= io_csrCtrl_distribute_csr_waddr; // @[CtrlBlock.scala 586:39]
    pfevent_io_distribute_csr_REG_wdata <= io_csrCtrl_distribute_csr_wdata; // @[CtrlBlock.scala 586:39]
    io_perf_0_value_REG <= hpm_io_perf_0_value; // @[PerfCounterUtils.scala 188:35]
    io_perf_0_value_REG_1 <= io_perf_0_value_REG; // @[PerfCounterUtils.scala 188:27]
    io_perf_1_value_REG <= hpm_io_perf_1_value; // @[PerfCounterUtils.scala 188:35]
    io_perf_1_value_REG_1 <= io_perf_1_value_REG; // @[PerfCounterUtils.scala 188:27]
    io_perf_2_value_REG <= hpm_io_perf_2_value; // @[PerfCounterUtils.scala 188:35]
    io_perf_2_value_REG_1 <= io_perf_2_value_REG; // @[PerfCounterUtils.scala 188:27]
    io_perf_3_value_REG <= hpm_io_perf_3_value; // @[PerfCounterUtils.scala 188:35]
    io_perf_3_value_REG_1 <= io_perf_3_value_REG; // @[PerfCounterUtils.scala 188:27]
    io_perf_4_value_REG <= hpm_io_perf_4_value; // @[PerfCounterUtils.scala 188:35]
    io_perf_4_value_REG_1 <= io_perf_4_value_REG; // @[PerfCounterUtils.scala 188:27]
    io_perf_5_value_REG <= hpm_io_perf_5_value; // @[PerfCounterUtils.scala 188:35]
    io_perf_5_value_REG_1 <= io_perf_5_value_REG; // @[PerfCounterUtils.scala 188:27]
    io_perf_6_value_REG <= hpm_io_perf_6_value; // @[PerfCounterUtils.scala 188:35]
    io_perf_6_value_REG_1 <= io_perf_6_value_REG; // @[PerfCounterUtils.scala 188:27]
    io_perf_7_value_REG <= hpm_io_perf_7_value; // @[PerfCounterUtils.scala 188:35]
    io_perf_7_value_REG_1 <= io_perf_7_value_REG; // @[PerfCounterUtils.scala 188:27]
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[CtrlBlock.scala 302:27]
      redirectForExu_next_valid_REG <= 1'h0;
    end else if (flushRedirect_valid_REG) begin
      redirectForExu_next_valid_REG <= flushRedirect_valid_REG;
    end else begin
      redirectForExu_next_valid_REG <= redirectGen_io_stage2Redirect_valid;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[CtrlBlock.scala 310:36]
      exuRedirect_delayed_valid_REG <= 1'h0;
    end else begin
      exuRedirect_delayed_valid_REG <= exuRedirect_valid & ~exuRedirect_killedByOlder;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[CtrlBlock.scala 310:36]
      exuRedirect_delayed_valid_REG_1 <= 1'h0;
    end else begin
      exuRedirect_delayed_valid_REG_1 <= exuRedirect_valid_1 & ~exuRedirect_killedByOlder_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[CtrlBlock.scala 310:36]
      exuRedirect_delayed_valid_REG_2 <= 1'h0;
    end else begin
      exuRedirect_delayed_valid_REG_2 <= exuRedirect_valid_2 & ~exuRedirect_killedByOlder_2;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[CtrlBlock.scala 315:56]
      loadReplay_valid_REG <= 1'h0;
    end else begin
      loadReplay_valid_REG <= io_memoryViolation_valid & _loadReplay_valid_T_8;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[CtrlBlock.scala 363:31]
      pendingRedirect <= 1'h0; // @[CtrlBlock.scala 364:21]
    end else begin
      pendingRedirect <= stage2Redirect_valid | _GEN_996;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PipelineConnect.scala 112:20]
      renamePipe_valid <= 1'h0; // @[PipelineConnect.scala 112:28]
    end else if (_renamePipe_T) begin
      renamePipe_valid <= 1'h0;
    end else begin
      renamePipe_valid <= _GEN_999;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PipelineConnect.scala 112:20]
      renamePipe_valid_1 <= 1'h0; // @[PipelineConnect.scala 112:28]
    end else if (_renamePipe_T) begin
      renamePipe_valid_1 <= 1'h0;
    end else begin
      renamePipe_valid_1 <= _GEN_1095;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PipelineConnect.scala 112:20]
      valid <= 1'h0; // @[PipelineConnect.scala 112:28]
    end else if (stage2Redirect_valid) begin
      valid <= 1'h0;
    end else begin
      valid <= _GEN_1182;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PipelineConnect.scala 112:20]
      valid_1 <= 1'h0; // @[PipelineConnect.scala 112:28]
    end else if (stage2Redirect_valid) begin
      valid_1 <= 1'h0;
    end else begin
      valid_1 <= _GEN_1293;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  pcMem_io_wen_0_REG = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  pcMem_io_waddr_0_REG = _RAND_1[2:0];
  _RAND_2 = {2{`RANDOM}};
  pcMem_io_wdata_0_REG_startAddr = _RAND_2[38:0];
  _RAND_3 = {2{`RANDOM}};
  pcMem_io_wdata_0_REG_nextLineAddr = _RAND_3[38:0];
  _RAND_4 = {1{`RANDOM}};
  pcMem_io_wdata_0_REG_isNextMask_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  pcMem_io_wdata_0_REG_isNextMask_1 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  pcMem_io_wdata_0_REG_isNextMask_2 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  pcMem_io_wdata_0_REG_isNextMask_3 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  pcMem_io_wdata_0_REG_isNextMask_4 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  pcMem_io_wdata_0_REG_isNextMask_5 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  pcMem_io_wdata_0_REG_isNextMask_6 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  pcMem_io_wdata_0_REG_isNextMask_7 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  flushPC_REG = _RAND_12[2:0];
  _RAND_13 = {1{`RANDOM}};
  flushRedirect_valid_REG = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  flushRedirect_bits_rrobIdx_flag = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  flushRedirect_bits_rrobIdx_value = _RAND_15[4:0];
  _RAND_16 = {1{`RANDOM}};
  flushRedirect_bits_rftqIdx_flag = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  flushRedirect_bits_rftqIdx_value = _RAND_17[2:0];
  _RAND_18 = {1{`RANDOM}};
  flushRedirect_bits_rftqOffset = _RAND_18[2:0];
  _RAND_19 = {1{`RANDOM}};
  flushRedirect_bits_rlevel = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  redirectForExu_next_valid_REG = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  redirectForExu_next_bits_rrobIdx_flag = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  redirectForExu_next_bits_rrobIdx_value = _RAND_22[4:0];
  _RAND_23 = {1{`RANDOM}};
  redirectForExu_next_bits_rlevel = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  exuRedirect_delayed_valid_REG = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  exuRedirect_delayed_bits_ruop_cf_pd_isRVC = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  exuRedirect_delayed_bits_ruop_cf_pd_brType = _RAND_26[1:0];
  _RAND_27 = {1{`RANDOM}};
  exuRedirect_delayed_bits_ruop_cf_pd_isCall = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  exuRedirect_delayed_bits_ruop_cf_pd_isRet = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  exuRedirect_delayed_bits_ruop_ctrl_imm = _RAND_29[19:0];
  _RAND_30 = {1{`RANDOM}};
  exuRedirect_delayed_bits_rredirect_robIdx_flag = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  exuRedirect_delayed_bits_rredirect_robIdx_value = _RAND_31[4:0];
  _RAND_32 = {1{`RANDOM}};
  exuRedirect_delayed_bits_rredirect_ftqIdx_flag = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  exuRedirect_delayed_bits_rredirect_ftqIdx_value = _RAND_33[2:0];
  _RAND_34 = {1{`RANDOM}};
  exuRedirect_delayed_bits_rredirect_ftqOffset = _RAND_34[2:0];
  _RAND_35 = {2{`RANDOM}};
  exuRedirect_delayed_bits_rredirect_cfiUpdate_target = _RAND_35[38:0];
  _RAND_36 = {1{`RANDOM}};
  exuRedirect_delayed_bits_rredirect_cfiUpdate_isMisPred = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  exuRedirect_delayed_valid_REG_1 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  exuRedirect_delayed_bits_r1_uop_cf_pd_isRVC = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  exuRedirect_delayed_bits_r1_uop_cf_pd_brType = _RAND_39[1:0];
  _RAND_40 = {1{`RANDOM}};
  exuRedirect_delayed_bits_r1_uop_cf_pd_isCall = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  exuRedirect_delayed_bits_r1_uop_cf_pd_isRet = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  exuRedirect_delayed_bits_r1_uop_ctrl_imm = _RAND_42[19:0];
  _RAND_43 = {1{`RANDOM}};
  exuRedirect_delayed_bits_r1_redirect_robIdx_flag = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  exuRedirect_delayed_bits_r1_redirect_robIdx_value = _RAND_44[4:0];
  _RAND_45 = {1{`RANDOM}};
  exuRedirect_delayed_bits_r1_redirect_ftqIdx_flag = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  exuRedirect_delayed_bits_r1_redirect_ftqIdx_value = _RAND_46[2:0];
  _RAND_47 = {1{`RANDOM}};
  exuRedirect_delayed_bits_r1_redirect_ftqOffset = _RAND_47[2:0];
  _RAND_48 = {1{`RANDOM}};
  exuRedirect_delayed_bits_r1_redirect_cfiUpdate_taken = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  exuRedirect_delayed_bits_r1_redirect_cfiUpdate_isMisPred = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  exuRedirect_delayed_valid_REG_2 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  exuRedirect_delayed_bits_r2_uop_cf_pd_isRVC = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  exuRedirect_delayed_bits_r2_uop_cf_pd_brType = _RAND_52[1:0];
  _RAND_53 = {1{`RANDOM}};
  exuRedirect_delayed_bits_r2_uop_cf_pd_isCall = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  exuRedirect_delayed_bits_r2_uop_cf_pd_isRet = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  exuRedirect_delayed_bits_r2_uop_ctrl_imm = _RAND_55[19:0];
  _RAND_56 = {1{`RANDOM}};
  exuRedirect_delayed_bits_r2_redirect_robIdx_flag = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  exuRedirect_delayed_bits_r2_redirect_robIdx_value = _RAND_57[4:0];
  _RAND_58 = {1{`RANDOM}};
  exuRedirect_delayed_bits_r2_redirect_ftqIdx_flag = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  exuRedirect_delayed_bits_r2_redirect_ftqIdx_value = _RAND_59[2:0];
  _RAND_60 = {1{`RANDOM}};
  exuRedirect_delayed_bits_r2_redirect_ftqOffset = _RAND_60[2:0];
  _RAND_61 = {1{`RANDOM}};
  exuRedirect_delayed_bits_r2_redirect_cfiUpdate_taken = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  exuRedirect_delayed_bits_r2_redirect_cfiUpdate_isMisPred = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  loadReplay_valid_REG = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  loadReplay_bits_rrobIdx_flag = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  loadReplay_bits_rrobIdx_value = _RAND_65[4:0];
  _RAND_66 = {1{`RANDOM}};
  loadReplay_bits_rftqIdx_flag = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  loadReplay_bits_rftqIdx_value = _RAND_67[2:0];
  _RAND_68 = {1{`RANDOM}};
  loadReplay_bits_rftqOffset = _RAND_68[2:0];
  _RAND_69 = {1{`RANDOM}};
  loadReplay_bits_rstFtqIdx_value = _RAND_69[2:0];
  _RAND_70 = {1{`RANDOM}};
  loadReplay_bits_rstFtqOffset = _RAND_70[2:0];
  _RAND_71 = {1{`RANDOM}};
  redirectGen_io_redirectPcRead_data_REG = _RAND_71[2:0];
  _RAND_72 = {1{`RANDOM}};
  redirectGen_io_memPredPcRead_data_REG = _RAND_72[2:0];
  _RAND_73 = {1{`RANDOM}};
  frontendFlushBits_ftqIdx_flag = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  frontendFlushBits_ftqIdx_value = _RAND_74[2:0];
  _RAND_75 = {1{`RANDOM}};
  frontendFlushBits_ftqOffset = _RAND_75[2:0];
  _RAND_76 = {1{`RANDOM}};
  frontendFlushBits_level = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  io_frontend_toFtq_rob_commits_0_valid_REG = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  io_frontend_toFtq_rob_commits_0_bits_rcommitType = _RAND_78[2:0];
  _RAND_79 = {1{`RANDOM}};
  io_frontend_toFtq_rob_commits_0_bits_rftqIdx_flag = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  io_frontend_toFtq_rob_commits_0_bits_rftqIdx_value = _RAND_80[2:0];
  _RAND_81 = {1{`RANDOM}};
  io_frontend_toFtq_rob_commits_0_bits_rftqOffset = _RAND_81[2:0];
  _RAND_82 = {1{`RANDOM}};
  io_frontend_toFtq_rob_commits_1_valid_REG = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  io_frontend_toFtq_rob_commits_1_bits_rcommitType = _RAND_83[2:0];
  _RAND_84 = {1{`RANDOM}};
  io_frontend_toFtq_rob_commits_1_bits_rftqIdx_flag = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  io_frontend_toFtq_rob_commits_1_bits_rftqIdx_value = _RAND_85[2:0];
  _RAND_86 = {1{`RANDOM}};
  io_frontend_toFtq_rob_commits_1_bits_rftqOffset = _RAND_86[2:0];
  _RAND_87 = {2{`RANDOM}};
  rob_flush_pc = _RAND_87[38:0];
  _RAND_88 = {2{`RANDOM}};
  io_frontend_toFtq_redirect_bits_cfiUpdate_target_REG = _RAND_88[38:0];
  _RAND_89 = {1{`RANDOM}};
  pendingRedirect = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  REG = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  decode_io_csrCtrl_REG_fusion_enable = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  decode_io_csrCtrl_REG_wfi_enable = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  decode_io_csrCtrl_REG_svinval_enable = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  decode_io_csrCtrl_REG_singlestep = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  ssit_io_update_REG_valid = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  ssit_io_update_REG_ldpc = _RAND_96[9:0];
  _RAND_97 = {1{`RANDOM}};
  ssit_io_update_REG_stpc = _RAND_97[9:0];
  _RAND_98 = {1{`RANDOM}};
  ssit_io_csrCtrl_REG_lvpred_timeout = _RAND_98[4:0];
  _RAND_99 = {1{`RANDOM}};
  lfst_io_redirect_REG_valid = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  lfst_io_redirect_REG_bits_robIdx_flag = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  lfst_io_redirect_REG_bits_robIdx_value = _RAND_101[4:0];
  _RAND_102 = {1{`RANDOM}};
  lfst_io_redirect_REG_bits_level = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  REG_1_0_valid = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  REG_1_0_bits_uop_cf_storeSetHit = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  REG_1_0_bits_uop_cf_ssid = _RAND_105[4:0];
  _RAND_106 = {1{`RANDOM}};
  REG_1_0_bits_uop_robIdx_value = _RAND_106[4:0];
  _RAND_107 = {1{`RANDOM}};
  REG_1_1_valid = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  REG_1_1_bits_uop_cf_storeSetHit = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  REG_1_1_bits_uop_cf_ssid = _RAND_109[4:0];
  _RAND_110 = {1{`RANDOM}};
  REG_1_1_bits_uop_robIdx_value = _RAND_110[4:0];
  _RAND_111 = {1{`RANDOM}};
  lfst_io_csrCtrl_REG_lvpred_disable = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  lfst_io_csrCtrl_REG_no_spec_load = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  lfst_io_csrCtrl_REG_storeset_wait_store = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  renamePipe_valid = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  renamePipe_data_cf_foldpc = _RAND_115[9:0];
  _RAND_116 = {1{`RANDOM}};
  renamePipe_data_cf_exceptionVec_1 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  renamePipe_data_cf_exceptionVec_2 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  renamePipe_data_cf_exceptionVec_12 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  renamePipe_data_cf_trigger_frontendHit_0 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  renamePipe_data_cf_trigger_frontendHit_1 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  renamePipe_data_cf_trigger_frontendHit_2 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  renamePipe_data_cf_trigger_frontendHit_3 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  renamePipe_data_cf_trigger_backendEn_0 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  renamePipe_data_cf_trigger_backendEn_1 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  renamePipe_data_cf_pd_isRVC = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  renamePipe_data_cf_pd_brType = _RAND_126[1:0];
  _RAND_127 = {1{`RANDOM}};
  renamePipe_data_cf_pd_isCall = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  renamePipe_data_cf_pd_isRet = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  renamePipe_data_cf_pred_taken = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  renamePipe_data_cf_crossPageIPFFix = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  renamePipe_data_cf_ftqPtr_flag = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  renamePipe_data_cf_ftqPtr_value = _RAND_132[2:0];
  _RAND_133 = {1{`RANDOM}};
  renamePipe_data_cf_ftqOffset = _RAND_133[2:0];
  _RAND_134 = {1{`RANDOM}};
  renamePipe_data_ctrl_srcType_0 = _RAND_134[1:0];
  _RAND_135 = {1{`RANDOM}};
  renamePipe_data_ctrl_srcType_1 = _RAND_135[1:0];
  _RAND_136 = {1{`RANDOM}};
  renamePipe_data_ctrl_srcType_2 = _RAND_136[1:0];
  _RAND_137 = {1{`RANDOM}};
  renamePipe_data_ctrl_lsrc_0 = _RAND_137[4:0];
  _RAND_138 = {1{`RANDOM}};
  renamePipe_data_ctrl_lsrc_1 = _RAND_138[4:0];
  _RAND_139 = {1{`RANDOM}};
  renamePipe_data_ctrl_ldest = _RAND_139[4:0];
  _RAND_140 = {1{`RANDOM}};
  renamePipe_data_ctrl_fuType = _RAND_140[3:0];
  _RAND_141 = {1{`RANDOM}};
  renamePipe_data_ctrl_fuOpType = _RAND_141[6:0];
  _RAND_142 = {1{`RANDOM}};
  renamePipe_data_ctrl_rfWen = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  renamePipe_data_ctrl_fpWen = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  renamePipe_data_ctrl_isXSTrap = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  renamePipe_data_ctrl_noSpecExec = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  renamePipe_data_ctrl_blockBackward = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  renamePipe_data_ctrl_flushPipe = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  renamePipe_data_ctrl_selImm = _RAND_148[3:0];
  _RAND_149 = {1{`RANDOM}};
  renamePipe_data_ctrl_imm = _RAND_149[19:0];
  _RAND_150 = {1{`RANDOM}};
  renamePipe_data_ctrl_fpu_isAddSub = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  renamePipe_data_ctrl_fpu_typeTagIn = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  renamePipe_data_ctrl_fpu_typeTagOut = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  renamePipe_data_ctrl_fpu_fromInt = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  renamePipe_data_ctrl_fpu_wflags = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  renamePipe_data_ctrl_fpu_fpWen = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  renamePipe_data_ctrl_fpu_fmaCmd = _RAND_156[1:0];
  _RAND_157 = {1{`RANDOM}};
  renamePipe_data_ctrl_fpu_div = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  renamePipe_data_ctrl_fpu_sqrt = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  renamePipe_data_ctrl_fpu_fcvt = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  renamePipe_data_ctrl_fpu_typ = _RAND_160[1:0];
  _RAND_161 = {1{`RANDOM}};
  renamePipe_data_ctrl_fpu_fmt = _RAND_161[1:0];
  _RAND_162 = {1{`RANDOM}};
  renamePipe_data_ctrl_fpu_ren3 = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  renamePipe_data_ctrl_fpu_rm = _RAND_163[2:0];
  _RAND_164 = {1{`RANDOM}};
  renamePipe_data_ctrl_isMove = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  renamePipe_valid_1 = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  renamePipe_data_1_cf_foldpc = _RAND_166[9:0];
  _RAND_167 = {1{`RANDOM}};
  renamePipe_data_1_cf_exceptionVec_1 = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  renamePipe_data_1_cf_exceptionVec_2 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  renamePipe_data_1_cf_exceptionVec_12 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  renamePipe_data_1_cf_trigger_frontendHit_0 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  renamePipe_data_1_cf_trigger_frontendHit_1 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  renamePipe_data_1_cf_trigger_frontendHit_2 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  renamePipe_data_1_cf_trigger_frontendHit_3 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  renamePipe_data_1_cf_trigger_backendEn_0 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  renamePipe_data_1_cf_trigger_backendEn_1 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  renamePipe_data_1_cf_pd_isRVC = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  renamePipe_data_1_cf_pd_brType = _RAND_177[1:0];
  _RAND_178 = {1{`RANDOM}};
  renamePipe_data_1_cf_pd_isCall = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  renamePipe_data_1_cf_pd_isRet = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  renamePipe_data_1_cf_pred_taken = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  renamePipe_data_1_cf_crossPageIPFFix = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  renamePipe_data_1_cf_ftqPtr_flag = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  renamePipe_data_1_cf_ftqPtr_value = _RAND_183[2:0];
  _RAND_184 = {1{`RANDOM}};
  renamePipe_data_1_cf_ftqOffset = _RAND_184[2:0];
  _RAND_185 = {1{`RANDOM}};
  renamePipe_data_1_ctrl_srcType_0 = _RAND_185[1:0];
  _RAND_186 = {1{`RANDOM}};
  renamePipe_data_1_ctrl_srcType_1 = _RAND_186[1:0];
  _RAND_187 = {1{`RANDOM}};
  renamePipe_data_1_ctrl_srcType_2 = _RAND_187[1:0];
  _RAND_188 = {1{`RANDOM}};
  renamePipe_data_1_ctrl_lsrc_0 = _RAND_188[4:0];
  _RAND_189 = {1{`RANDOM}};
  renamePipe_data_1_ctrl_lsrc_1 = _RAND_189[4:0];
  _RAND_190 = {1{`RANDOM}};
  renamePipe_data_1_ctrl_lsrc_2 = _RAND_190[4:0];
  _RAND_191 = {1{`RANDOM}};
  renamePipe_data_1_ctrl_ldest = _RAND_191[4:0];
  _RAND_192 = {1{`RANDOM}};
  renamePipe_data_1_ctrl_fuType = _RAND_192[3:0];
  _RAND_193 = {1{`RANDOM}};
  renamePipe_data_1_ctrl_fuOpType = _RAND_193[6:0];
  _RAND_194 = {1{`RANDOM}};
  renamePipe_data_1_ctrl_rfWen = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  renamePipe_data_1_ctrl_fpWen = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  renamePipe_data_1_ctrl_isXSTrap = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  renamePipe_data_1_ctrl_noSpecExec = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  renamePipe_data_1_ctrl_blockBackward = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  renamePipe_data_1_ctrl_flushPipe = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  renamePipe_data_1_ctrl_selImm = _RAND_200[3:0];
  _RAND_201 = {1{`RANDOM}};
  renamePipe_data_1_ctrl_imm = _RAND_201[19:0];
  _RAND_202 = {1{`RANDOM}};
  renamePipe_data_1_ctrl_fpu_isAddSub = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  renamePipe_data_1_ctrl_fpu_typeTagIn = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  renamePipe_data_1_ctrl_fpu_typeTagOut = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  renamePipe_data_1_ctrl_fpu_fromInt = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  renamePipe_data_1_ctrl_fpu_wflags = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  renamePipe_data_1_ctrl_fpu_fpWen = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  renamePipe_data_1_ctrl_fpu_fmaCmd = _RAND_208[1:0];
  _RAND_209 = {1{`RANDOM}};
  renamePipe_data_1_ctrl_fpu_div = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  renamePipe_data_1_ctrl_fpu_sqrt = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  renamePipe_data_1_ctrl_fpu_fcvt = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  renamePipe_data_1_ctrl_fpu_typ = _RAND_212[1:0];
  _RAND_213 = {1{`RANDOM}};
  renamePipe_data_1_ctrl_fpu_fmt = _RAND_213[1:0];
  _RAND_214 = {1{`RANDOM}};
  renamePipe_data_1_ctrl_fpu_ren3 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  renamePipe_data_1_ctrl_fpu_rm = _RAND_215[2:0];
  _RAND_216 = {1{`RANDOM}};
  renamePipe_data_1_ctrl_isMove = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  valid = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  data_cf_foldpc = _RAND_218[9:0];
  _RAND_219 = {1{`RANDOM}};
  data_cf_exceptionVec_1 = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  data_cf_exceptionVec_2 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  data_cf_exceptionVec_12 = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  data_cf_trigger_frontendHit_0 = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  data_cf_trigger_frontendHit_1 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  data_cf_trigger_frontendHit_2 = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  data_cf_trigger_frontendHit_3 = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  data_cf_trigger_backendEn_0 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  data_cf_trigger_backendEn_1 = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  data_cf_pd_isRVC = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  data_cf_pd_brType = _RAND_229[1:0];
  _RAND_230 = {1{`RANDOM}};
  data_cf_pd_isCall = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  data_cf_pd_isRet = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  data_cf_pred_taken = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  data_cf_crossPageIPFFix = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  data_cf_storeSetHit = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  data_cf_loadWaitStrict = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  data_cf_ssid = _RAND_236[4:0];
  _RAND_237 = {1{`RANDOM}};
  data_cf_ftqPtr_flag = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  data_cf_ftqPtr_value = _RAND_238[2:0];
  _RAND_239 = {1{`RANDOM}};
  data_cf_ftqOffset = _RAND_239[2:0];
  _RAND_240 = {1{`RANDOM}};
  data_ctrl_srcType_0 = _RAND_240[1:0];
  _RAND_241 = {1{`RANDOM}};
  data_ctrl_srcType_1 = _RAND_241[1:0];
  _RAND_242 = {1{`RANDOM}};
  data_ctrl_srcType_2 = _RAND_242[1:0];
  _RAND_243 = {1{`RANDOM}};
  data_ctrl_ldest = _RAND_243[4:0];
  _RAND_244 = {1{`RANDOM}};
  data_ctrl_fuType = _RAND_244[3:0];
  _RAND_245 = {1{`RANDOM}};
  data_ctrl_fuOpType = _RAND_245[6:0];
  _RAND_246 = {1{`RANDOM}};
  data_ctrl_rfWen = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  data_ctrl_fpWen = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  data_ctrl_isXSTrap = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  data_ctrl_noSpecExec = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  data_ctrl_blockBackward = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  data_ctrl_flushPipe = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  data_ctrl_selImm = _RAND_252[3:0];
  _RAND_253 = {1{`RANDOM}};
  data_ctrl_imm = _RAND_253[19:0];
  _RAND_254 = {1{`RANDOM}};
  data_ctrl_commitType = _RAND_254[2:0];
  _RAND_255 = {1{`RANDOM}};
  data_ctrl_fpu_isAddSub = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  data_ctrl_fpu_typeTagIn = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  data_ctrl_fpu_typeTagOut = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  data_ctrl_fpu_fromInt = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  data_ctrl_fpu_wflags = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  data_ctrl_fpu_fpWen = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  data_ctrl_fpu_fmaCmd = _RAND_261[1:0];
  _RAND_262 = {1{`RANDOM}};
  data_ctrl_fpu_div = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  data_ctrl_fpu_sqrt = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  data_ctrl_fpu_fcvt = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  data_ctrl_fpu_typ = _RAND_265[1:0];
  _RAND_266 = {1{`RANDOM}};
  data_ctrl_fpu_fmt = _RAND_266[1:0];
  _RAND_267 = {1{`RANDOM}};
  data_ctrl_fpu_ren3 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  data_ctrl_fpu_rm = _RAND_268[2:0];
  _RAND_269 = {1{`RANDOM}};
  data_ctrl_isMove = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  data_psrc_0 = _RAND_270[5:0];
  _RAND_271 = {1{`RANDOM}};
  data_psrc_1 = _RAND_271[5:0];
  _RAND_272 = {1{`RANDOM}};
  data_psrc_2 = _RAND_272[5:0];
  _RAND_273 = {1{`RANDOM}};
  data_pdest = _RAND_273[5:0];
  _RAND_274 = {1{`RANDOM}};
  data_old_pdest = _RAND_274[5:0];
  _RAND_275 = {1{`RANDOM}};
  data_robIdx_flag = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  data_robIdx_value = _RAND_276[4:0];
  _RAND_277 = {1{`RANDOM}};
  data_eliminatedMove = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  valid_1 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  data_1_cf_foldpc = _RAND_279[9:0];
  _RAND_280 = {1{`RANDOM}};
  data_1_cf_exceptionVec_1 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  data_1_cf_exceptionVec_2 = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  data_1_cf_exceptionVec_12 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  data_1_cf_trigger_frontendHit_0 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  data_1_cf_trigger_frontendHit_1 = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  data_1_cf_trigger_frontendHit_2 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  data_1_cf_trigger_frontendHit_3 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  data_1_cf_trigger_backendEn_0 = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  data_1_cf_trigger_backendEn_1 = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  data_1_cf_pd_isRVC = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  data_1_cf_pd_brType = _RAND_290[1:0];
  _RAND_291 = {1{`RANDOM}};
  data_1_cf_pd_isCall = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  data_1_cf_pd_isRet = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  data_1_cf_pred_taken = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  data_1_cf_crossPageIPFFix = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  data_1_cf_storeSetHit = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  data_1_cf_loadWaitStrict = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  data_1_cf_ssid = _RAND_297[4:0];
  _RAND_298 = {1{`RANDOM}};
  data_1_cf_ftqPtr_flag = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  data_1_cf_ftqPtr_value = _RAND_299[2:0];
  _RAND_300 = {1{`RANDOM}};
  data_1_cf_ftqOffset = _RAND_300[2:0];
  _RAND_301 = {1{`RANDOM}};
  data_1_ctrl_srcType_0 = _RAND_301[1:0];
  _RAND_302 = {1{`RANDOM}};
  data_1_ctrl_srcType_1 = _RAND_302[1:0];
  _RAND_303 = {1{`RANDOM}};
  data_1_ctrl_srcType_2 = _RAND_303[1:0];
  _RAND_304 = {1{`RANDOM}};
  data_1_ctrl_ldest = _RAND_304[4:0];
  _RAND_305 = {1{`RANDOM}};
  data_1_ctrl_fuType = _RAND_305[3:0];
  _RAND_306 = {1{`RANDOM}};
  data_1_ctrl_fuOpType = _RAND_306[6:0];
  _RAND_307 = {1{`RANDOM}};
  data_1_ctrl_rfWen = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  data_1_ctrl_fpWen = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  data_1_ctrl_isXSTrap = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  data_1_ctrl_noSpecExec = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  data_1_ctrl_blockBackward = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  data_1_ctrl_flushPipe = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  data_1_ctrl_selImm = _RAND_313[3:0];
  _RAND_314 = {1{`RANDOM}};
  data_1_ctrl_imm = _RAND_314[19:0];
  _RAND_315 = {1{`RANDOM}};
  data_1_ctrl_fpu_isAddSub = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  data_1_ctrl_fpu_typeTagIn = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  data_1_ctrl_fpu_typeTagOut = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  data_1_ctrl_fpu_fromInt = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  data_1_ctrl_fpu_wflags = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  data_1_ctrl_fpu_fpWen = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  data_1_ctrl_fpu_fmaCmd = _RAND_321[1:0];
  _RAND_322 = {1{`RANDOM}};
  data_1_ctrl_fpu_div = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  data_1_ctrl_fpu_sqrt = _RAND_323[0:0];
  _RAND_324 = {1{`RANDOM}};
  data_1_ctrl_fpu_fcvt = _RAND_324[0:0];
  _RAND_325 = {1{`RANDOM}};
  data_1_ctrl_fpu_typ = _RAND_325[1:0];
  _RAND_326 = {1{`RANDOM}};
  data_1_ctrl_fpu_fmt = _RAND_326[1:0];
  _RAND_327 = {1{`RANDOM}};
  data_1_ctrl_fpu_ren3 = _RAND_327[0:0];
  _RAND_328 = {1{`RANDOM}};
  data_1_ctrl_fpu_rm = _RAND_328[2:0];
  _RAND_329 = {1{`RANDOM}};
  data_1_ctrl_isMove = _RAND_329[0:0];
  _RAND_330 = {1{`RANDOM}};
  data_1_psrc_0 = _RAND_330[5:0];
  _RAND_331 = {1{`RANDOM}};
  data_1_psrc_1 = _RAND_331[5:0];
  _RAND_332 = {1{`RANDOM}};
  data_1_psrc_2 = _RAND_332[5:0];
  _RAND_333 = {1{`RANDOM}};
  data_1_pdest = _RAND_333[5:0];
  _RAND_334 = {1{`RANDOM}};
  data_1_old_pdest = _RAND_334[5:0];
  _RAND_335 = {1{`RANDOM}};
  data_1_robIdx_flag = _RAND_335[0:0];
  _RAND_336 = {1{`RANDOM}};
  data_1_robIdx_value = _RAND_336[4:0];
  _RAND_337 = {1{`RANDOM}};
  data_1_eliminatedMove = _RAND_337[0:0];
  _RAND_338 = {1{`RANDOM}};
  dispatch_io_singleStep_REG = _RAND_338[0:0];
  _RAND_339 = {1{`RANDOM}};
  jumpPcRead0_REG = _RAND_339[2:0];
  _RAND_340 = {1{`RANDOM}};
  read_from_newest_entry_REG_flag = _RAND_340[0:0];
  _RAND_341 = {1{`RANDOM}};
  read_from_newest_entry_REG_value = _RAND_341[2:0];
  _RAND_342 = {1{`RANDOM}};
  read_from_newest_entry_REG_1_flag = _RAND_342[0:0];
  _RAND_343 = {1{`RANDOM}};
  read_from_newest_entry_REG_1_value = _RAND_343[2:0];
  _RAND_344 = {2{`RANDOM}};
  io_jalr_target_REG = _RAND_344[38:0];
  _RAND_345 = {1{`RANDOM}};
  sources_source_exuOutput_3_valid_REG = _RAND_345[0:0];
  _RAND_346 = {1{`RANDOM}};
  sources_source_exuOutput_3_bits_REG_uop_cf_exceptionVec_2 = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  sources_source_exuOutput_3_bits_REG_uop_cf_exceptionVec_3 = _RAND_347[0:0];
  _RAND_348 = {1{`RANDOM}};
  sources_source_exuOutput_3_bits_REG_uop_cf_exceptionVec_8 = _RAND_348[0:0];
  _RAND_349 = {1{`RANDOM}};
  sources_source_exuOutput_3_bits_REG_uop_cf_exceptionVec_9 = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  sources_source_exuOutput_3_bits_REG_uop_cf_exceptionVec_11 = _RAND_350[0:0];
  _RAND_351 = {1{`RANDOM}};
  sources_source_exuOutput_3_bits_REG_uop_ctrl_flushPipe = _RAND_351[0:0];
  _RAND_352 = {1{`RANDOM}};
  sources_source_exuOutput_3_bits_REG_uop_robIdx_flag = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  sources_source_exuOutput_3_bits_REG_uop_robIdx_value = _RAND_353[4:0];
  _RAND_354 = {1{`RANDOM}};
  sources_source_exuOutput_3_bits_REG_fflags = _RAND_354[4:0];
  _RAND_355 = {1{`RANDOM}};
  sources_source_exuOutput_4_valid_REG = _RAND_355[0:0];
  _RAND_356 = {1{`RANDOM}};
  sources_source_exuOutput_4_bits_REG_uop_robIdx_value = _RAND_356[4:0];
  _RAND_357 = {1{`RANDOM}};
  sources_source_exuOutput_4_bits_REG_fflags = _RAND_357[4:0];
  _RAND_358 = {1{`RANDOM}};
  sources_source_exuOutput_5_valid_REG = _RAND_358[0:0];
  _RAND_359 = {1{`RANDOM}};
  sources_source_exuOutput_5_bits_REG_uop_robIdx_value = _RAND_359[4:0];
  _RAND_360 = {1{`RANDOM}};
  sources_source_exuOutput_5_bits_REG_fflags = _RAND_360[4:0];
  _RAND_361 = {1{`RANDOM}};
  sources_source_exuOutput_6_valid_REG = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  sources_source_exuOutput_6_bits_REG_uop_cf_exceptionVec_4 = _RAND_362[0:0];
  _RAND_363 = {1{`RANDOM}};
  sources_source_exuOutput_6_bits_REG_uop_cf_exceptionVec_5 = _RAND_363[0:0];
  _RAND_364 = {1{`RANDOM}};
  sources_source_exuOutput_6_bits_REG_uop_cf_exceptionVec_13 = _RAND_364[0:0];
  _RAND_365 = {1{`RANDOM}};
  sources_source_exuOutput_6_bits_REG_uop_cf_trigger_backendHit_0 = _RAND_365[0:0];
  _RAND_366 = {1{`RANDOM}};
  sources_source_exuOutput_6_bits_REG_uop_cf_trigger_backendHit_1 = _RAND_366[0:0];
  _RAND_367 = {1{`RANDOM}};
  sources_source_exuOutput_6_bits_REG_uop_cf_trigger_backendHit_2 = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  sources_source_exuOutput_6_bits_REG_uop_cf_trigger_backendHit_3 = _RAND_368[0:0];
  _RAND_369 = {1{`RANDOM}};
  sources_source_exuOutput_6_bits_REG_uop_cf_trigger_backendHit_4 = _RAND_369[0:0];
  _RAND_370 = {1{`RANDOM}};
  sources_source_exuOutput_6_bits_REG_uop_cf_trigger_backendHit_5 = _RAND_370[0:0];
  _RAND_371 = {1{`RANDOM}};
  sources_source_exuOutput_6_bits_REG_uop_ctrl_flushPipe = _RAND_371[0:0];
  _RAND_372 = {1{`RANDOM}};
  sources_source_exuOutput_6_bits_REG_uop_ctrl_replayInst = _RAND_372[0:0];
  _RAND_373 = {1{`RANDOM}};
  sources_source_exuOutput_6_bits_REG_uop_robIdx_flag = _RAND_373[0:0];
  _RAND_374 = {1{`RANDOM}};
  sources_source_exuOutput_6_bits_REG_uop_robIdx_value = _RAND_374[4:0];
  _RAND_375 = {1{`RANDOM}};
  sources_source_exuOutput_7_valid_REG = _RAND_375[0:0];
  _RAND_376 = {1{`RANDOM}};
  sources_source_exuOutput_7_bits_REG_uop_cf_exceptionVec_4 = _RAND_376[0:0];
  _RAND_377 = {1{`RANDOM}};
  sources_source_exuOutput_7_bits_REG_uop_cf_exceptionVec_5 = _RAND_377[0:0];
  _RAND_378 = {1{`RANDOM}};
  sources_source_exuOutput_7_bits_REG_uop_cf_exceptionVec_13 = _RAND_378[0:0];
  _RAND_379 = {1{`RANDOM}};
  sources_source_exuOutput_7_bits_REG_uop_cf_trigger_backendHit_0 = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  sources_source_exuOutput_7_bits_REG_uop_cf_trigger_backendHit_1 = _RAND_380[0:0];
  _RAND_381 = {1{`RANDOM}};
  sources_source_exuOutput_7_bits_REG_uop_cf_trigger_backendHit_2 = _RAND_381[0:0];
  _RAND_382 = {1{`RANDOM}};
  sources_source_exuOutput_7_bits_REG_uop_cf_trigger_backendHit_3 = _RAND_382[0:0];
  _RAND_383 = {1{`RANDOM}};
  sources_source_exuOutput_7_bits_REG_uop_cf_trigger_backendHit_4 = _RAND_383[0:0];
  _RAND_384 = {1{`RANDOM}};
  sources_source_exuOutput_7_bits_REG_uop_cf_trigger_backendHit_5 = _RAND_384[0:0];
  _RAND_385 = {1{`RANDOM}};
  sources_source_exuOutput_7_bits_REG_uop_ctrl_flushPipe = _RAND_385[0:0];
  _RAND_386 = {1{`RANDOM}};
  sources_source_exuOutput_7_bits_REG_uop_ctrl_replayInst = _RAND_386[0:0];
  _RAND_387 = {1{`RANDOM}};
  sources_source_exuOutput_7_bits_REG_uop_robIdx_flag = _RAND_387[0:0];
  _RAND_388 = {1{`RANDOM}};
  sources_source_exuOutput_7_bits_REG_uop_robIdx_value = _RAND_388[4:0];
  _RAND_389 = {1{`RANDOM}};
  sources_source_exuOutput_8_valid_REG = _RAND_389[0:0];
  _RAND_390 = {1{`RANDOM}};
  sources_source_exuOutput_8_bits_REG_uop_cf_exceptionVec_4 = _RAND_390[0:0];
  _RAND_391 = {1{`RANDOM}};
  sources_source_exuOutput_8_bits_REG_uop_cf_exceptionVec_5 = _RAND_391[0:0];
  _RAND_392 = {1{`RANDOM}};
  sources_source_exuOutput_8_bits_REG_uop_cf_exceptionVec_6 = _RAND_392[0:0];
  _RAND_393 = {1{`RANDOM}};
  sources_source_exuOutput_8_bits_REG_uop_cf_exceptionVec_7 = _RAND_393[0:0];
  _RAND_394 = {1{`RANDOM}};
  sources_source_exuOutput_8_bits_REG_uop_cf_exceptionVec_13 = _RAND_394[0:0];
  _RAND_395 = {1{`RANDOM}};
  sources_source_exuOutput_8_bits_REG_uop_cf_exceptionVec_15 = _RAND_395[0:0];
  _RAND_396 = {1{`RANDOM}};
  sources_source_exuOutput_8_bits_REG_uop_cf_trigger_backendHit_0 = _RAND_396[0:0];
  _RAND_397 = {1{`RANDOM}};
  sources_source_exuOutput_8_bits_REG_uop_cf_trigger_backendHit_1 = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  sources_source_exuOutput_8_bits_REG_uop_cf_trigger_backendHit_2 = _RAND_398[0:0];
  _RAND_399 = {1{`RANDOM}};
  sources_source_exuOutput_8_bits_REG_uop_cf_trigger_backendHit_3 = _RAND_399[0:0];
  _RAND_400 = {1{`RANDOM}};
  sources_source_exuOutput_8_bits_REG_uop_cf_trigger_backendHit_4 = _RAND_400[0:0];
  _RAND_401 = {1{`RANDOM}};
  sources_source_exuOutput_8_bits_REG_uop_cf_trigger_backendHit_5 = _RAND_401[0:0];
  _RAND_402 = {1{`RANDOM}};
  sources_source_exuOutput_8_bits_REG_uop_robIdx_flag = _RAND_402[0:0];
  _RAND_403 = {1{`RANDOM}};
  sources_source_exuOutput_8_bits_REG_uop_robIdx_value = _RAND_403[4:0];
  _RAND_404 = {1{`RANDOM}};
  sources_source_exuOutput_9_valid_REG = _RAND_404[0:0];
  _RAND_405 = {1{`RANDOM}};
  sources_source_exuOutput_9_bits_REG_uop_cf_exceptionVec_6 = _RAND_405[0:0];
  _RAND_406 = {1{`RANDOM}};
  sources_source_exuOutput_9_bits_REG_uop_cf_exceptionVec_7 = _RAND_406[0:0];
  _RAND_407 = {1{`RANDOM}};
  sources_source_exuOutput_9_bits_REG_uop_cf_exceptionVec_15 = _RAND_407[0:0];
  _RAND_408 = {1{`RANDOM}};
  sources_source_exuOutput_9_bits_REG_uop_cf_trigger_backendHit_0 = _RAND_408[0:0];
  _RAND_409 = {1{`RANDOM}};
  sources_source_exuOutput_9_bits_REG_uop_cf_trigger_backendHit_1 = _RAND_409[0:0];
  _RAND_410 = {1{`RANDOM}};
  sources_source_exuOutput_9_bits_REG_uop_cf_trigger_backendHit_4 = _RAND_410[0:0];
  _RAND_411 = {1{`RANDOM}};
  sources_source_exuOutput_9_bits_REG_uop_robIdx_flag = _RAND_411[0:0];
  _RAND_412 = {1{`RANDOM}};
  sources_source_exuOutput_9_bits_REG_uop_robIdx_value = _RAND_412[4:0];
  _RAND_413 = {1{`RANDOM}};
  sources_source_exuOutput_0_valid_REG_3 = _RAND_413[0:0];
  _RAND_414 = {1{`RANDOM}};
  sources_source_exuOutput_0_bits_REG_3_uop_robIdx_value = _RAND_414[4:0];
  _RAND_415 = {1{`RANDOM}};
  sources_source_exuOutput_0_bits_REG_3_redirectValid = _RAND_415[0:0];
  _RAND_416 = {1{`RANDOM}};
  sources_source_exuOutput_0_bits_REG_3_redirect_cfiUpdate_isMisPred = _RAND_416[0:0];
  _RAND_417 = {1{`RANDOM}};
  sources_source_exuOutput_1_valid_REG_3 = _RAND_417[0:0];
  _RAND_418 = {1{`RANDOM}};
  sources_source_exuOutput_1_bits_REG_3_uop_robIdx_value = _RAND_418[4:0];
  _RAND_419 = {1{`RANDOM}};
  sources_source_exuOutput_1_bits_REG_3_redirectValid = _RAND_419[0:0];
  _RAND_420 = {1{`RANDOM}};
  sources_source_exuOutput_1_bits_REG_3_redirect_cfiUpdate_isMisPred = _RAND_420[0:0];
  _RAND_421 = {1{`RANDOM}};
  sources_source_exuOutput_2_valid_REG_3 = _RAND_421[0:0];
  _RAND_422 = {1{`RANDOM}};
  sources_source_exuOutput_2_bits_REG_3_uop_cf_exceptionVec_4 = _RAND_422[0:0];
  _RAND_423 = {1{`RANDOM}};
  sources_source_exuOutput_2_bits_REG_3_uop_cf_exceptionVec_5 = _RAND_423[0:0];
  _RAND_424 = {1{`RANDOM}};
  sources_source_exuOutput_2_bits_REG_3_uop_cf_exceptionVec_13 = _RAND_424[0:0];
  _RAND_425 = {1{`RANDOM}};
  sources_source_exuOutput_2_bits_REG_3_uop_cf_trigger_backendHit_0 = _RAND_425[0:0];
  _RAND_426 = {1{`RANDOM}};
  sources_source_exuOutput_2_bits_REG_3_uop_cf_trigger_backendHit_1 = _RAND_426[0:0];
  _RAND_427 = {1{`RANDOM}};
  sources_source_exuOutput_2_bits_REG_3_uop_cf_trigger_backendHit_2 = _RAND_427[0:0];
  _RAND_428 = {1{`RANDOM}};
  sources_source_exuOutput_2_bits_REG_3_uop_cf_trigger_backendHit_3 = _RAND_428[0:0];
  _RAND_429 = {1{`RANDOM}};
  sources_source_exuOutput_2_bits_REG_3_uop_cf_trigger_backendHit_4 = _RAND_429[0:0];
  _RAND_430 = {1{`RANDOM}};
  sources_source_exuOutput_2_bits_REG_3_uop_cf_trigger_backendHit_5 = _RAND_430[0:0];
  _RAND_431 = {1{`RANDOM}};
  sources_source_exuOutput_2_bits_REG_3_uop_ctrl_flushPipe = _RAND_431[0:0];
  _RAND_432 = {1{`RANDOM}};
  sources_source_exuOutput_2_bits_REG_3_uop_ctrl_replayInst = _RAND_432[0:0];
  _RAND_433 = {1{`RANDOM}};
  sources_source_exuOutput_2_bits_REG_3_uop_robIdx_value = _RAND_433[4:0];
  _RAND_434 = {1{`RANDOM}};
  sources_source_exuOutput_2_bits_REG_3_debug_isMMIO = _RAND_434[0:0];
  _RAND_435 = {1{`RANDOM}};
  sources_source_exuOutput_3_valid_REG_3 = _RAND_435[0:0];
  _RAND_436 = {1{`RANDOM}};
  sources_source_exuOutput_3_bits_REG_3_uop_cf_exceptionVec_4 = _RAND_436[0:0];
  _RAND_437 = {1{`RANDOM}};
  sources_source_exuOutput_3_bits_REG_3_uop_cf_exceptionVec_5 = _RAND_437[0:0];
  _RAND_438 = {1{`RANDOM}};
  sources_source_exuOutput_3_bits_REG_3_uop_cf_exceptionVec_13 = _RAND_438[0:0];
  _RAND_439 = {1{`RANDOM}};
  sources_source_exuOutput_3_bits_REG_3_uop_cf_trigger_backendHit_0 = _RAND_439[0:0];
  _RAND_440 = {1{`RANDOM}};
  sources_source_exuOutput_3_bits_REG_3_uop_cf_trigger_backendHit_1 = _RAND_440[0:0];
  _RAND_441 = {1{`RANDOM}};
  sources_source_exuOutput_3_bits_REG_3_uop_cf_trigger_backendHit_2 = _RAND_441[0:0];
  _RAND_442 = {1{`RANDOM}};
  sources_source_exuOutput_3_bits_REG_3_uop_cf_trigger_backendHit_3 = _RAND_442[0:0];
  _RAND_443 = {1{`RANDOM}};
  sources_source_exuOutput_3_bits_REG_3_uop_cf_trigger_backendHit_4 = _RAND_443[0:0];
  _RAND_444 = {1{`RANDOM}};
  sources_source_exuOutput_3_bits_REG_3_uop_cf_trigger_backendHit_5 = _RAND_444[0:0];
  _RAND_445 = {1{`RANDOM}};
  sources_source_exuOutput_3_bits_REG_3_uop_ctrl_flushPipe = _RAND_445[0:0];
  _RAND_446 = {1{`RANDOM}};
  sources_source_exuOutput_3_bits_REG_3_uop_ctrl_replayInst = _RAND_446[0:0];
  _RAND_447 = {1{`RANDOM}};
  sources_source_exuOutput_3_bits_REG_3_uop_robIdx_value = _RAND_447[4:0];
  _RAND_448 = {1{`RANDOM}};
  sources_source_exuOutput_3_bits_REG_3_debug_isMMIO = _RAND_448[0:0];
  _RAND_449 = {1{`RANDOM}};
  sources_source_exuOutput_4_valid_REG_3 = _RAND_449[0:0];
  _RAND_450 = {1{`RANDOM}};
  sources_source_exuOutput_4_bits_REG_3_uop_cf_exceptionVec_2 = _RAND_450[0:0];
  _RAND_451 = {1{`RANDOM}};
  sources_source_exuOutput_4_bits_REG_3_uop_cf_exceptionVec_3 = _RAND_451[0:0];
  _RAND_452 = {1{`RANDOM}};
  sources_source_exuOutput_4_bits_REG_3_uop_cf_exceptionVec_8 = _RAND_452[0:0];
  _RAND_453 = {1{`RANDOM}};
  sources_source_exuOutput_4_bits_REG_3_uop_cf_exceptionVec_9 = _RAND_453[0:0];
  _RAND_454 = {1{`RANDOM}};
  sources_source_exuOutput_4_bits_REG_3_uop_cf_exceptionVec_11 = _RAND_454[0:0];
  _RAND_455 = {1{`RANDOM}};
  sources_source_exuOutput_4_bits_REG_3_uop_ctrl_flushPipe = _RAND_455[0:0];
  _RAND_456 = {1{`RANDOM}};
  sources_source_exuOutput_4_bits_REG_3_uop_robIdx_value = _RAND_456[4:0];
  _RAND_457 = {1{`RANDOM}};
  sources_source_exuOutput_4_bits_REG_3_redirectValid = _RAND_457[0:0];
  _RAND_458 = {1{`RANDOM}};
  sources_source_exuOutput_4_bits_REG_3_redirect_cfiUpdate_isMisPred = _RAND_458[0:0];
  _RAND_459 = {1{`RANDOM}};
  sources_source_exuOutput_4_bits_REG_3_debug_isPerfCnt = _RAND_459[0:0];
  _RAND_460 = {1{`RANDOM}};
  sources_source_exuOutput_5_valid_REG_3 = _RAND_460[0:0];
  _RAND_461 = {1{`RANDOM}};
  sources_source_exuOutput_5_bits_REG_3_uop_cf_trigger_backendHit_0 = _RAND_461[0:0];
  _RAND_462 = {1{`RANDOM}};
  sources_source_exuOutput_5_bits_REG_3_uop_cf_trigger_backendHit_1 = _RAND_462[0:0];
  _RAND_463 = {1{`RANDOM}};
  sources_source_exuOutput_5_bits_REG_3_uop_cf_trigger_backendHit_2 = _RAND_463[0:0];
  _RAND_464 = {1{`RANDOM}};
  sources_source_exuOutput_5_bits_REG_3_uop_cf_trigger_backendHit_3 = _RAND_464[0:0];
  _RAND_465 = {1{`RANDOM}};
  sources_source_exuOutput_5_bits_REG_3_uop_cf_trigger_backendHit_4 = _RAND_465[0:0];
  _RAND_466 = {1{`RANDOM}};
  sources_source_exuOutput_5_bits_REG_3_uop_cf_trigger_backendHit_5 = _RAND_466[0:0];
  _RAND_467 = {1{`RANDOM}};
  sources_source_exuOutput_5_bits_REG_3_uop_robIdx_value = _RAND_467[4:0];
  _RAND_468 = {1{`RANDOM}};
  sources_source_exuOutput_6_valid_REG_3 = _RAND_468[0:0];
  _RAND_469 = {1{`RANDOM}};
  sources_source_exuOutput_6_bits_REG_3_uop_cf_exceptionVec_2 = _RAND_469[0:0];
  _RAND_470 = {1{`RANDOM}};
  sources_source_exuOutput_6_bits_REG_3_uop_cf_exceptionVec_3 = _RAND_470[0:0];
  _RAND_471 = {1{`RANDOM}};
  sources_source_exuOutput_6_bits_REG_3_uop_cf_exceptionVec_8 = _RAND_471[0:0];
  _RAND_472 = {1{`RANDOM}};
  sources_source_exuOutput_6_bits_REG_3_uop_cf_exceptionVec_9 = _RAND_472[0:0];
  _RAND_473 = {1{`RANDOM}};
  sources_source_exuOutput_6_bits_REG_3_uop_cf_exceptionVec_11 = _RAND_473[0:0];
  _RAND_474 = {1{`RANDOM}};
  sources_source_exuOutput_6_bits_REG_3_uop_ctrl_flushPipe = _RAND_474[0:0];
  _RAND_475 = {1{`RANDOM}};
  sources_source_exuOutput_6_bits_REG_3_uop_robIdx_value = _RAND_475[4:0];
  _RAND_476 = {1{`RANDOM}};
  sources_source_exuOutput_6_bits_REG_3_redirectValid = _RAND_476[0:0];
  _RAND_477 = {1{`RANDOM}};
  sources_source_exuOutput_6_bits_REG_3_redirect_cfiUpdate_isMisPred = _RAND_477[0:0];
  _RAND_478 = {1{`RANDOM}};
  sources_source_exuOutput_6_bits_REG_3_debug_isPerfCnt = _RAND_478[0:0];
  _RAND_479 = {1{`RANDOM}};
  sources_source_exuOutput_7_valid_REG_3 = _RAND_479[0:0];
  _RAND_480 = {1{`RANDOM}};
  sources_source_exuOutput_7_bits_REG_3_uop_cf_exceptionVec_4 = _RAND_480[0:0];
  _RAND_481 = {1{`RANDOM}};
  sources_source_exuOutput_7_bits_REG_3_uop_cf_exceptionVec_5 = _RAND_481[0:0];
  _RAND_482 = {1{`RANDOM}};
  sources_source_exuOutput_7_bits_REG_3_uop_cf_exceptionVec_6 = _RAND_482[0:0];
  _RAND_483 = {1{`RANDOM}};
  sources_source_exuOutput_7_bits_REG_3_uop_cf_exceptionVec_7 = _RAND_483[0:0];
  _RAND_484 = {1{`RANDOM}};
  sources_source_exuOutput_7_bits_REG_3_uop_cf_exceptionVec_13 = _RAND_484[0:0];
  _RAND_485 = {1{`RANDOM}};
  sources_source_exuOutput_7_bits_REG_3_uop_cf_exceptionVec_15 = _RAND_485[0:0];
  _RAND_486 = {1{`RANDOM}};
  sources_source_exuOutput_7_bits_REG_3_uop_cf_trigger_backendHit_0 = _RAND_486[0:0];
  _RAND_487 = {1{`RANDOM}};
  sources_source_exuOutput_7_bits_REG_3_uop_cf_trigger_backendHit_1 = _RAND_487[0:0];
  _RAND_488 = {1{`RANDOM}};
  sources_source_exuOutput_7_bits_REG_3_uop_cf_trigger_backendHit_2 = _RAND_488[0:0];
  _RAND_489 = {1{`RANDOM}};
  sources_source_exuOutput_7_bits_REG_3_uop_cf_trigger_backendHit_3 = _RAND_489[0:0];
  _RAND_490 = {1{`RANDOM}};
  sources_source_exuOutput_7_bits_REG_3_uop_cf_trigger_backendHit_4 = _RAND_490[0:0];
  _RAND_491 = {1{`RANDOM}};
  sources_source_exuOutput_7_bits_REG_3_uop_cf_trigger_backendHit_5 = _RAND_491[0:0];
  _RAND_492 = {1{`RANDOM}};
  sources_source_exuOutput_7_bits_REG_3_uop_robIdx_value = _RAND_492[4:0];
  _RAND_493 = {1{`RANDOM}};
  sources_source_exuOutput_7_bits_REG_3_redirectValid = _RAND_493[0:0];
  _RAND_494 = {1{`RANDOM}};
  sources_source_exuOutput_7_bits_REG_3_redirect_cfiUpdate_isMisPred = _RAND_494[0:0];
  _RAND_495 = {1{`RANDOM}};
  sources_source_exuOutput_7_bits_REG_3_debug_isMMIO = _RAND_495[0:0];
  _RAND_496 = {1{`RANDOM}};
  sources_source_exuOutput_7_bits_REG_3_debug_isPerfCnt = _RAND_496[0:0];
  _RAND_497 = {1{`RANDOM}};
  sources_source_exuOutput_8_valid_REG_3 = _RAND_497[0:0];
  _RAND_498 = {1{`RANDOM}};
  sources_source_exuOutput_8_bits_REG_3_uop_cf_exceptionVec_4 = _RAND_498[0:0];
  _RAND_499 = {1{`RANDOM}};
  sources_source_exuOutput_8_bits_REG_3_uop_cf_exceptionVec_5 = _RAND_499[0:0];
  _RAND_500 = {1{`RANDOM}};
  sources_source_exuOutput_8_bits_REG_3_uop_cf_exceptionVec_6 = _RAND_500[0:0];
  _RAND_501 = {1{`RANDOM}};
  sources_source_exuOutput_8_bits_REG_3_uop_cf_exceptionVec_7 = _RAND_501[0:0];
  _RAND_502 = {1{`RANDOM}};
  sources_source_exuOutput_8_bits_REG_3_uop_cf_exceptionVec_13 = _RAND_502[0:0];
  _RAND_503 = {1{`RANDOM}};
  sources_source_exuOutput_8_bits_REG_3_uop_cf_exceptionVec_15 = _RAND_503[0:0];
  _RAND_504 = {1{`RANDOM}};
  sources_source_exuOutput_8_bits_REG_3_uop_cf_trigger_backendHit_0 = _RAND_504[0:0];
  _RAND_505 = {1{`RANDOM}};
  sources_source_exuOutput_8_bits_REG_3_uop_cf_trigger_backendHit_1 = _RAND_505[0:0];
  _RAND_506 = {1{`RANDOM}};
  sources_source_exuOutput_8_bits_REG_3_uop_cf_trigger_backendHit_2 = _RAND_506[0:0];
  _RAND_507 = {1{`RANDOM}};
  sources_source_exuOutput_8_bits_REG_3_uop_cf_trigger_backendHit_3 = _RAND_507[0:0];
  _RAND_508 = {1{`RANDOM}};
  sources_source_exuOutput_8_bits_REG_3_uop_cf_trigger_backendHit_4 = _RAND_508[0:0];
  _RAND_509 = {1{`RANDOM}};
  sources_source_exuOutput_8_bits_REG_3_uop_cf_trigger_backendHit_5 = _RAND_509[0:0];
  _RAND_510 = {1{`RANDOM}};
  sources_source_exuOutput_8_bits_REG_3_uop_robIdx_value = _RAND_510[4:0];
  _RAND_511 = {1{`RANDOM}};
  sources_source_exuOutput_8_bits_REG_3_redirectValid = _RAND_511[0:0];
  _RAND_512 = {1{`RANDOM}};
  sources_source_exuOutput_8_bits_REG_3_redirect_cfiUpdate_isMisPred = _RAND_512[0:0];
  _RAND_513 = {1{`RANDOM}};
  sources_source_exuOutput_8_bits_REG_3_debug_isMMIO = _RAND_513[0:0];
  _RAND_514 = {1{`RANDOM}};
  sources_source_exuOutput_8_bits_REG_3_debug_isPerfCnt = _RAND_514[0:0];
  _RAND_515 = {1{`RANDOM}};
  sources_source_exuOutput_9_valid_REG_3 = _RAND_515[0:0];
  _RAND_516 = {1{`RANDOM}};
  sources_source_exuOutput_9_bits_REG_3_uop_robIdx_value = _RAND_516[4:0];
  _RAND_517 = {1{`RANDOM}};
  sources_source_exuOutput_10_valid_REG_3 = _RAND_517[0:0];
  _RAND_518 = {1{`RANDOM}};
  sources_source_exuOutput_10_bits_REG_3_uop_robIdx_value = _RAND_518[4:0];
  _RAND_519 = {1{`RANDOM}};
  io_robio_toCSR_perfinfo_retiredInstr_REG = _RAND_519[2:0];
  _RAND_520 = {1{`RANDOM}};
  pfevent_io_distribute_csr_REG_wvalid = _RAND_520[0:0];
  _RAND_521 = {1{`RANDOM}};
  pfevent_io_distribute_csr_REG_waddr = _RAND_521[11:0];
  _RAND_522 = {2{`RANDOM}};
  pfevent_io_distribute_csr_REG_wdata = _RAND_522[63:0];
  _RAND_523 = {1{`RANDOM}};
  io_perf_0_value_REG = _RAND_523[5:0];
  _RAND_524 = {1{`RANDOM}};
  io_perf_0_value_REG_1 = _RAND_524[5:0];
  _RAND_525 = {1{`RANDOM}};
  io_perf_1_value_REG = _RAND_525[5:0];
  _RAND_526 = {1{`RANDOM}};
  io_perf_1_value_REG_1 = _RAND_526[5:0];
  _RAND_527 = {1{`RANDOM}};
  io_perf_2_value_REG = _RAND_527[5:0];
  _RAND_528 = {1{`RANDOM}};
  io_perf_2_value_REG_1 = _RAND_528[5:0];
  _RAND_529 = {1{`RANDOM}};
  io_perf_3_value_REG = _RAND_529[5:0];
  _RAND_530 = {1{`RANDOM}};
  io_perf_3_value_REG_1 = _RAND_530[5:0];
  _RAND_531 = {1{`RANDOM}};
  io_perf_4_value_REG = _RAND_531[5:0];
  _RAND_532 = {1{`RANDOM}};
  io_perf_4_value_REG_1 = _RAND_532[5:0];
  _RAND_533 = {1{`RANDOM}};
  io_perf_5_value_REG = _RAND_533[5:0];
  _RAND_534 = {1{`RANDOM}};
  io_perf_5_value_REG_1 = _RAND_534[5:0];
  _RAND_535 = {1{`RANDOM}};
  io_perf_6_value_REG = _RAND_535[5:0];
  _RAND_536 = {1{`RANDOM}};
  io_perf_6_value_REG_1 = _RAND_536[5:0];
  _RAND_537 = {1{`RANDOM}};
  io_perf_7_value_REG = _RAND_537[5:0];
  _RAND_538 = {1{`RANDOM}};
  io_perf_7_value_REG_1 = _RAND_538[5:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    redirectForExu_next_valid_REG = 1'h0;
  end
  if (reset) begin
    exuRedirect_delayed_valid_REG = 1'h0;
  end
  if (reset) begin
    exuRedirect_delayed_valid_REG_1 = 1'h0;
  end
  if (reset) begin
    exuRedirect_delayed_valid_REG_2 = 1'h0;
  end
  if (reset) begin
    loadReplay_valid_REG = 1'h0;
  end
  if (reset) begin
    pendingRedirect = 1'h0;
  end
  if (reset) begin
    renamePipe_valid = 1'h0;
  end
  if (reset) begin
    renamePipe_valid_1 = 1'h0;
  end
  if (reset) begin
    valid = 1'h0;
  end
  if (reset) begin
    valid_1 = 1'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule

