module L1FlagMetaArray(
  input        clock,
  input        reset,
  input        io_read_0_valid,
  input  [5:0] io_read_0_bits_idx,
  input        io_read_1_valid,
  input  [5:0] io_read_1_bits_idx,
  input        io_read_2_valid,
  input  [5:0] io_read_2_bits_idx,
  output       io_resp_0_0,
  output       io_resp_0_1,
  output       io_resp_0_2,
  output       io_resp_0_3,
  output       io_resp_0_4,
  output       io_resp_0_5,
  output       io_resp_0_6,
  output       io_resp_0_7,
  output       io_resp_1_0,
  output       io_resp_1_1,
  output       io_resp_1_2,
  output       io_resp_1_3,
  output       io_resp_1_4,
  output       io_resp_1_5,
  output       io_resp_1_6,
  output       io_resp_1_7,
  output       io_resp_2_0,
  output       io_resp_2_1,
  output       io_resp_2_2,
  output       io_resp_2_3,
  output       io_resp_2_4,
  output       io_resp_2_5,
  output       io_resp_2_6,
  output       io_resp_2_7,
  input        io_write_0_valid,
  input  [5:0] io_write_0_bits_idx,
  input  [7:0] io_write_0_bits_way_en,
  input        io_write_0_bits_flag,
  input        io_write_1_valid,
  input  [5:0] io_write_1_bits_idx,
  input  [7:0] io_write_1_bits_way_en,
  input        io_write_1_bits_flag
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
`endif // RANDOMIZE_REG_INIT
  reg  meta_array_0_0; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_0_1; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_0_2; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_0_3; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_0_4; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_0_5; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_0_6; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_0_7; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_1_0; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_1_1; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_1_2; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_1_3; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_1_4; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_1_5; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_1_6; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_1_7; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_2_0; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_2_1; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_2_2; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_2_3; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_2_4; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_2_5; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_2_6; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_2_7; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_3_0; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_3_1; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_3_2; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_3_3; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_3_4; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_3_5; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_3_6; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_3_7; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_4_0; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_4_1; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_4_2; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_4_3; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_4_4; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_4_5; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_4_6; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_4_7; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_5_0; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_5_1; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_5_2; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_5_3; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_5_4; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_5_5; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_5_6; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_5_7; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_6_0; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_6_1; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_6_2; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_6_3; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_6_4; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_6_5; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_6_6; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_6_7; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_7_0; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_7_1; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_7_2; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_7_3; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_7_4; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_7_5; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_7_6; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_7_7; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_8_0; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_8_1; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_8_2; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_8_3; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_8_4; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_8_5; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_8_6; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_8_7; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_9_0; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_9_1; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_9_2; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_9_3; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_9_4; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_9_5; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_9_6; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_9_7; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_10_0; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_10_1; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_10_2; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_10_3; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_10_4; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_10_5; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_10_6; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_10_7; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_11_0; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_11_1; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_11_2; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_11_3; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_11_4; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_11_5; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_11_6; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_11_7; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_12_0; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_12_1; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_12_2; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_12_3; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_12_4; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_12_5; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_12_6; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_12_7; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_13_0; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_13_1; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_13_2; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_13_3; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_13_4; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_13_5; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_13_6; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_13_7; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_14_0; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_14_1; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_14_2; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_14_3; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_14_4; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_14_5; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_14_6; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_14_7; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_15_0; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_15_1; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_15_2; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_15_3; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_15_4; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_15_5; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_15_6; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_15_7; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_16_0; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_16_1; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_16_2; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_16_3; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_16_4; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_16_5; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_16_6; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_16_7; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_17_0; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_17_1; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_17_2; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_17_3; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_17_4; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_17_5; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_17_6; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_17_7; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_18_0; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_18_1; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_18_2; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_18_3; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_18_4; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_18_5; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_18_6; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_18_7; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_19_0; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_19_1; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_19_2; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_19_3; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_19_4; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_19_5; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_19_6; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_19_7; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_20_0; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_20_1; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_20_2; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_20_3; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_20_4; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_20_5; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_20_6; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_20_7; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_21_0; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_21_1; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_21_2; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_21_3; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_21_4; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_21_5; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_21_6; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_21_7; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_22_0; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_22_1; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_22_2; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_22_3; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_22_4; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_22_5; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_22_6; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_22_7; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_23_0; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_23_1; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_23_2; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_23_3; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_23_4; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_23_5; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_23_6; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_23_7; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_24_0; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_24_1; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_24_2; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_24_3; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_24_4; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_24_5; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_24_6; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_24_7; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_25_0; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_25_1; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_25_2; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_25_3; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_25_4; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_25_5; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_25_6; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_25_7; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_26_0; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_26_1; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_26_2; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_26_3; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_26_4; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_26_5; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_26_6; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_26_7; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_27_0; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_27_1; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_27_2; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_27_3; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_27_4; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_27_5; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_27_6; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_27_7; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_28_0; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_28_1; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_28_2; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_28_3; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_28_4; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_28_5; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_28_6; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_28_7; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_29_0; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_29_1; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_29_2; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_29_3; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_29_4; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_29_5; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_29_6; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_29_7; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_30_0; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_30_1; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_30_2; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_30_3; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_30_4; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_30_5; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_30_6; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_30_7; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_31_0; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_31_1; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_31_2; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_31_3; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_31_4; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_31_5; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_31_6; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_31_7; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_32_0; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_32_1; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_32_2; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_32_3; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_32_4; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_32_5; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_32_6; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_32_7; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_33_0; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_33_1; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_33_2; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_33_3; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_33_4; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_33_5; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_33_6; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_33_7; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_34_0; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_34_1; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_34_2; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_34_3; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_34_4; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_34_5; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_34_6; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_34_7; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_35_0; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_35_1; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_35_2; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_35_3; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_35_4; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_35_5; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_35_6; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_35_7; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_36_0; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_36_1; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_36_2; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_36_3; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_36_4; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_36_5; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_36_6; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_36_7; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_37_0; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_37_1; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_37_2; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_37_3; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_37_4; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_37_5; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_37_6; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_37_7; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_38_0; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_38_1; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_38_2; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_38_3; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_38_4; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_38_5; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_38_6; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_38_7; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_39_0; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_39_1; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_39_2; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_39_3; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_39_4; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_39_5; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_39_6; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_39_7; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_40_0; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_40_1; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_40_2; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_40_3; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_40_4; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_40_5; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_40_6; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_40_7; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_41_0; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_41_1; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_41_2; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_41_3; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_41_4; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_41_5; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_41_6; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_41_7; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_42_0; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_42_1; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_42_2; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_42_3; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_42_4; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_42_5; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_42_6; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_42_7; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_43_0; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_43_1; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_43_2; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_43_3; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_43_4; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_43_5; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_43_6; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_43_7; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_44_0; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_44_1; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_44_2; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_44_3; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_44_4; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_44_5; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_44_6; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_44_7; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_45_0; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_45_1; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_45_2; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_45_3; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_45_4; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_45_5; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_45_6; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_45_7; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_46_0; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_46_1; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_46_2; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_46_3; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_46_4; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_46_5; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_46_6; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_46_7; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_47_0; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_47_1; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_47_2; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_47_3; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_47_4; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_47_5; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_47_6; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_47_7; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_48_0; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_48_1; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_48_2; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_48_3; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_48_4; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_48_5; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_48_6; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_48_7; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_49_0; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_49_1; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_49_2; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_49_3; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_49_4; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_49_5; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_49_6; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_49_7; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_50_0; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_50_1; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_50_2; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_50_3; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_50_4; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_50_5; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_50_6; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_50_7; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_51_0; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_51_1; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_51_2; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_51_3; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_51_4; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_51_5; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_51_6; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_51_7; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_52_0; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_52_1; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_52_2; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_52_3; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_52_4; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_52_5; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_52_6; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_52_7; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_53_0; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_53_1; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_53_2; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_53_3; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_53_4; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_53_5; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_53_6; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_53_7; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_54_0; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_54_1; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_54_2; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_54_3; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_54_4; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_54_5; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_54_6; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_54_7; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_55_0; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_55_1; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_55_2; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_55_3; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_55_4; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_55_5; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_55_6; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_55_7; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_56_0; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_56_1; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_56_2; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_56_3; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_56_4; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_56_5; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_56_6; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_56_7; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_57_0; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_57_1; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_57_2; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_57_3; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_57_4; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_57_5; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_57_6; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_57_7; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_58_0; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_58_1; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_58_2; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_58_3; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_58_4; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_58_5; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_58_6; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_58_7; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_59_0; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_59_1; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_59_2; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_59_3; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_59_4; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_59_5; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_59_6; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_59_7; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_60_0; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_60_1; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_60_2; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_60_3; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_60_4; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_60_5; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_60_6; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_60_7; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_61_0; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_61_1; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_61_2; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_61_3; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_61_4; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_61_5; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_61_6; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_61_7; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_62_0; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_62_1; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_62_2; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_62_3; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_62_4; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_62_5; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_62_6; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_62_7; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_63_0; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_63_1; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_63_2; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_63_3; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_63_4; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_63_5; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_63_6; // @[AsynchronousMetaArray.scala 115:27]
  reg  meta_array_63_7; // @[AsynchronousMetaArray.scala 115:27]
  reg [5:0] s1_way_waddr_0_0_r; // @[Reg.scala 16:16]
  reg  s1_way_wen_0_0_REG; // @[AsynchronousMetaArray.scala 153:44]
  reg  s1_way_wdata_0_0_r; // @[Reg.scala 16:16]
  reg [5:0] s1_way_waddr_0_1_r; // @[Reg.scala 16:16]
  reg  s1_way_wen_0_1_REG; // @[AsynchronousMetaArray.scala 153:44]
  wire  read_way_bypass = s1_way_wen_0_1_REG & s1_way_waddr_0_1_r == io_read_0_bits_idx | s1_way_wen_0_0_REG &
    s1_way_waddr_0_0_r == io_read_0_bits_idx; // @[AsynchronousMetaArray.scala 134:85 135:29]
  reg  s1_way_wdata_0_1_r; // @[Reg.scala 16:16]
  reg  io_resp_0_0_r; // @[Reg.scala 16:16]
  reg  io_resp_0_0_r1; // @[Reg.scala 16:16]
  reg [5:0] io_resp_0_0_r2; // @[Reg.scala 16:16]
  wire  _GEN_8 = 6'h1 == io_resp_0_0_r2 ? meta_array_1_0 : meta_array_0_0; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_9 = 6'h2 == io_resp_0_0_r2 ? meta_array_2_0 : _GEN_8; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_10 = 6'h3 == io_resp_0_0_r2 ? meta_array_3_0 : _GEN_9; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_11 = 6'h4 == io_resp_0_0_r2 ? meta_array_4_0 : _GEN_10; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_12 = 6'h5 == io_resp_0_0_r2 ? meta_array_5_0 : _GEN_11; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_13 = 6'h6 == io_resp_0_0_r2 ? meta_array_6_0 : _GEN_12; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_14 = 6'h7 == io_resp_0_0_r2 ? meta_array_7_0 : _GEN_13; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_15 = 6'h8 == io_resp_0_0_r2 ? meta_array_8_0 : _GEN_14; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_16 = 6'h9 == io_resp_0_0_r2 ? meta_array_9_0 : _GEN_15; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_17 = 6'ha == io_resp_0_0_r2 ? meta_array_10_0 : _GEN_16; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_18 = 6'hb == io_resp_0_0_r2 ? meta_array_11_0 : _GEN_17; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_19 = 6'hc == io_resp_0_0_r2 ? meta_array_12_0 : _GEN_18; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_20 = 6'hd == io_resp_0_0_r2 ? meta_array_13_0 : _GEN_19; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_21 = 6'he == io_resp_0_0_r2 ? meta_array_14_0 : _GEN_20; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_22 = 6'hf == io_resp_0_0_r2 ? meta_array_15_0 : _GEN_21; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_23 = 6'h10 == io_resp_0_0_r2 ? meta_array_16_0 : _GEN_22; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_24 = 6'h11 == io_resp_0_0_r2 ? meta_array_17_0 : _GEN_23; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_25 = 6'h12 == io_resp_0_0_r2 ? meta_array_18_0 : _GEN_24; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_26 = 6'h13 == io_resp_0_0_r2 ? meta_array_19_0 : _GEN_25; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_27 = 6'h14 == io_resp_0_0_r2 ? meta_array_20_0 : _GEN_26; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_28 = 6'h15 == io_resp_0_0_r2 ? meta_array_21_0 : _GEN_27; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_29 = 6'h16 == io_resp_0_0_r2 ? meta_array_22_0 : _GEN_28; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_30 = 6'h17 == io_resp_0_0_r2 ? meta_array_23_0 : _GEN_29; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_31 = 6'h18 == io_resp_0_0_r2 ? meta_array_24_0 : _GEN_30; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_32 = 6'h19 == io_resp_0_0_r2 ? meta_array_25_0 : _GEN_31; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_33 = 6'h1a == io_resp_0_0_r2 ? meta_array_26_0 : _GEN_32; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_34 = 6'h1b == io_resp_0_0_r2 ? meta_array_27_0 : _GEN_33; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_35 = 6'h1c == io_resp_0_0_r2 ? meta_array_28_0 : _GEN_34; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_36 = 6'h1d == io_resp_0_0_r2 ? meta_array_29_0 : _GEN_35; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_37 = 6'h1e == io_resp_0_0_r2 ? meta_array_30_0 : _GEN_36; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_38 = 6'h1f == io_resp_0_0_r2 ? meta_array_31_0 : _GEN_37; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_39 = 6'h20 == io_resp_0_0_r2 ? meta_array_32_0 : _GEN_38; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_40 = 6'h21 == io_resp_0_0_r2 ? meta_array_33_0 : _GEN_39; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_41 = 6'h22 == io_resp_0_0_r2 ? meta_array_34_0 : _GEN_40; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_42 = 6'h23 == io_resp_0_0_r2 ? meta_array_35_0 : _GEN_41; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_43 = 6'h24 == io_resp_0_0_r2 ? meta_array_36_0 : _GEN_42; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_44 = 6'h25 == io_resp_0_0_r2 ? meta_array_37_0 : _GEN_43; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_45 = 6'h26 == io_resp_0_0_r2 ? meta_array_38_0 : _GEN_44; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_46 = 6'h27 == io_resp_0_0_r2 ? meta_array_39_0 : _GEN_45; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_47 = 6'h28 == io_resp_0_0_r2 ? meta_array_40_0 : _GEN_46; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_48 = 6'h29 == io_resp_0_0_r2 ? meta_array_41_0 : _GEN_47; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_49 = 6'h2a == io_resp_0_0_r2 ? meta_array_42_0 : _GEN_48; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_50 = 6'h2b == io_resp_0_0_r2 ? meta_array_43_0 : _GEN_49; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_51 = 6'h2c == io_resp_0_0_r2 ? meta_array_44_0 : _GEN_50; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_52 = 6'h2d == io_resp_0_0_r2 ? meta_array_45_0 : _GEN_51; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_53 = 6'h2e == io_resp_0_0_r2 ? meta_array_46_0 : _GEN_52; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_54 = 6'h2f == io_resp_0_0_r2 ? meta_array_47_0 : _GEN_53; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_55 = 6'h30 == io_resp_0_0_r2 ? meta_array_48_0 : _GEN_54; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_56 = 6'h31 == io_resp_0_0_r2 ? meta_array_49_0 : _GEN_55; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_57 = 6'h32 == io_resp_0_0_r2 ? meta_array_50_0 : _GEN_56; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_58 = 6'h33 == io_resp_0_0_r2 ? meta_array_51_0 : _GEN_57; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_59 = 6'h34 == io_resp_0_0_r2 ? meta_array_52_0 : _GEN_58; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_60 = 6'h35 == io_resp_0_0_r2 ? meta_array_53_0 : _GEN_59; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_61 = 6'h36 == io_resp_0_0_r2 ? meta_array_54_0 : _GEN_60; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_62 = 6'h37 == io_resp_0_0_r2 ? meta_array_55_0 : _GEN_61; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_63 = 6'h38 == io_resp_0_0_r2 ? meta_array_56_0 : _GEN_62; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_64 = 6'h39 == io_resp_0_0_r2 ? meta_array_57_0 : _GEN_63; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_65 = 6'h3a == io_resp_0_0_r2 ? meta_array_58_0 : _GEN_64; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_66 = 6'h3b == io_resp_0_0_r2 ? meta_array_59_0 : _GEN_65; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_67 = 6'h3c == io_resp_0_0_r2 ? meta_array_60_0 : _GEN_66; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_68 = 6'h3d == io_resp_0_0_r2 ? meta_array_61_0 : _GEN_67; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_69 = 6'h3e == io_resp_0_0_r2 ? meta_array_62_0 : _GEN_68; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_70 = 6'h3f == io_resp_0_0_r2 ? meta_array_63_0 : _GEN_69; // @[AsynchronousMetaArray.scala 139:{25,25}]
  reg [5:0] s1_way_waddr_1_0_r; // @[Reg.scala 16:16]
  reg  s1_way_wen_1_0_REG; // @[AsynchronousMetaArray.scala 153:44]
  reg  s1_way_wdata_1_0_r; // @[Reg.scala 16:16]
  reg [5:0] s1_way_waddr_1_1_r; // @[Reg.scala 16:16]
  reg  s1_way_wen_1_1_REG; // @[AsynchronousMetaArray.scala 153:44]
  wire  read_way_bypass_1 = s1_way_wen_1_1_REG & s1_way_waddr_1_1_r == io_read_0_bits_idx | s1_way_wen_1_0_REG &
    s1_way_waddr_1_0_r == io_read_0_bits_idx; // @[AsynchronousMetaArray.scala 134:85 135:29]
  reg  s1_way_wdata_1_1_r; // @[Reg.scala 16:16]
  reg  io_resp_0_1_r; // @[Reg.scala 16:16]
  reg  io_resp_0_1_r1; // @[Reg.scala 16:16]
  reg [5:0] io_resp_0_1_r2; // @[Reg.scala 16:16]
  wire  _GEN_79 = 6'h1 == io_resp_0_1_r2 ? meta_array_1_1 : meta_array_0_1; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_80 = 6'h2 == io_resp_0_1_r2 ? meta_array_2_1 : _GEN_79; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_81 = 6'h3 == io_resp_0_1_r2 ? meta_array_3_1 : _GEN_80; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_82 = 6'h4 == io_resp_0_1_r2 ? meta_array_4_1 : _GEN_81; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_83 = 6'h5 == io_resp_0_1_r2 ? meta_array_5_1 : _GEN_82; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_84 = 6'h6 == io_resp_0_1_r2 ? meta_array_6_1 : _GEN_83; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_85 = 6'h7 == io_resp_0_1_r2 ? meta_array_7_1 : _GEN_84; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_86 = 6'h8 == io_resp_0_1_r2 ? meta_array_8_1 : _GEN_85; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_87 = 6'h9 == io_resp_0_1_r2 ? meta_array_9_1 : _GEN_86; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_88 = 6'ha == io_resp_0_1_r2 ? meta_array_10_1 : _GEN_87; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_89 = 6'hb == io_resp_0_1_r2 ? meta_array_11_1 : _GEN_88; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_90 = 6'hc == io_resp_0_1_r2 ? meta_array_12_1 : _GEN_89; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_91 = 6'hd == io_resp_0_1_r2 ? meta_array_13_1 : _GEN_90; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_92 = 6'he == io_resp_0_1_r2 ? meta_array_14_1 : _GEN_91; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_93 = 6'hf == io_resp_0_1_r2 ? meta_array_15_1 : _GEN_92; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_94 = 6'h10 == io_resp_0_1_r2 ? meta_array_16_1 : _GEN_93; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_95 = 6'h11 == io_resp_0_1_r2 ? meta_array_17_1 : _GEN_94; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_96 = 6'h12 == io_resp_0_1_r2 ? meta_array_18_1 : _GEN_95; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_97 = 6'h13 == io_resp_0_1_r2 ? meta_array_19_1 : _GEN_96; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_98 = 6'h14 == io_resp_0_1_r2 ? meta_array_20_1 : _GEN_97; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_99 = 6'h15 == io_resp_0_1_r2 ? meta_array_21_1 : _GEN_98; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_100 = 6'h16 == io_resp_0_1_r2 ? meta_array_22_1 : _GEN_99; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_101 = 6'h17 == io_resp_0_1_r2 ? meta_array_23_1 : _GEN_100; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_102 = 6'h18 == io_resp_0_1_r2 ? meta_array_24_1 : _GEN_101; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_103 = 6'h19 == io_resp_0_1_r2 ? meta_array_25_1 : _GEN_102; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_104 = 6'h1a == io_resp_0_1_r2 ? meta_array_26_1 : _GEN_103; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_105 = 6'h1b == io_resp_0_1_r2 ? meta_array_27_1 : _GEN_104; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_106 = 6'h1c == io_resp_0_1_r2 ? meta_array_28_1 : _GEN_105; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_107 = 6'h1d == io_resp_0_1_r2 ? meta_array_29_1 : _GEN_106; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_108 = 6'h1e == io_resp_0_1_r2 ? meta_array_30_1 : _GEN_107; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_109 = 6'h1f == io_resp_0_1_r2 ? meta_array_31_1 : _GEN_108; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_110 = 6'h20 == io_resp_0_1_r2 ? meta_array_32_1 : _GEN_109; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_111 = 6'h21 == io_resp_0_1_r2 ? meta_array_33_1 : _GEN_110; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_112 = 6'h22 == io_resp_0_1_r2 ? meta_array_34_1 : _GEN_111; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_113 = 6'h23 == io_resp_0_1_r2 ? meta_array_35_1 : _GEN_112; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_114 = 6'h24 == io_resp_0_1_r2 ? meta_array_36_1 : _GEN_113; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_115 = 6'h25 == io_resp_0_1_r2 ? meta_array_37_1 : _GEN_114; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_116 = 6'h26 == io_resp_0_1_r2 ? meta_array_38_1 : _GEN_115; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_117 = 6'h27 == io_resp_0_1_r2 ? meta_array_39_1 : _GEN_116; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_118 = 6'h28 == io_resp_0_1_r2 ? meta_array_40_1 : _GEN_117; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_119 = 6'h29 == io_resp_0_1_r2 ? meta_array_41_1 : _GEN_118; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_120 = 6'h2a == io_resp_0_1_r2 ? meta_array_42_1 : _GEN_119; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_121 = 6'h2b == io_resp_0_1_r2 ? meta_array_43_1 : _GEN_120; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_122 = 6'h2c == io_resp_0_1_r2 ? meta_array_44_1 : _GEN_121; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_123 = 6'h2d == io_resp_0_1_r2 ? meta_array_45_1 : _GEN_122; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_124 = 6'h2e == io_resp_0_1_r2 ? meta_array_46_1 : _GEN_123; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_125 = 6'h2f == io_resp_0_1_r2 ? meta_array_47_1 : _GEN_124; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_126 = 6'h30 == io_resp_0_1_r2 ? meta_array_48_1 : _GEN_125; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_127 = 6'h31 == io_resp_0_1_r2 ? meta_array_49_1 : _GEN_126; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_128 = 6'h32 == io_resp_0_1_r2 ? meta_array_50_1 : _GEN_127; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_129 = 6'h33 == io_resp_0_1_r2 ? meta_array_51_1 : _GEN_128; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_130 = 6'h34 == io_resp_0_1_r2 ? meta_array_52_1 : _GEN_129; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_131 = 6'h35 == io_resp_0_1_r2 ? meta_array_53_1 : _GEN_130; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_132 = 6'h36 == io_resp_0_1_r2 ? meta_array_54_1 : _GEN_131; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_133 = 6'h37 == io_resp_0_1_r2 ? meta_array_55_1 : _GEN_132; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_134 = 6'h38 == io_resp_0_1_r2 ? meta_array_56_1 : _GEN_133; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_135 = 6'h39 == io_resp_0_1_r2 ? meta_array_57_1 : _GEN_134; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_136 = 6'h3a == io_resp_0_1_r2 ? meta_array_58_1 : _GEN_135; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_137 = 6'h3b == io_resp_0_1_r2 ? meta_array_59_1 : _GEN_136; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_138 = 6'h3c == io_resp_0_1_r2 ? meta_array_60_1 : _GEN_137; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_139 = 6'h3d == io_resp_0_1_r2 ? meta_array_61_1 : _GEN_138; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_140 = 6'h3e == io_resp_0_1_r2 ? meta_array_62_1 : _GEN_139; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_141 = 6'h3f == io_resp_0_1_r2 ? meta_array_63_1 : _GEN_140; // @[AsynchronousMetaArray.scala 139:{25,25}]
  reg [5:0] s1_way_waddr_2_0_r; // @[Reg.scala 16:16]
  reg  s1_way_wen_2_0_REG; // @[AsynchronousMetaArray.scala 153:44]
  reg  s1_way_wdata_2_0_r; // @[Reg.scala 16:16]
  reg [5:0] s1_way_waddr_2_1_r; // @[Reg.scala 16:16]
  reg  s1_way_wen_2_1_REG; // @[AsynchronousMetaArray.scala 153:44]
  wire  read_way_bypass_2 = s1_way_wen_2_1_REG & s1_way_waddr_2_1_r == io_read_0_bits_idx | s1_way_wen_2_0_REG &
    s1_way_waddr_2_0_r == io_read_0_bits_idx; // @[AsynchronousMetaArray.scala 134:85 135:29]
  reg  s1_way_wdata_2_1_r; // @[Reg.scala 16:16]
  reg  io_resp_0_2_r; // @[Reg.scala 16:16]
  reg  io_resp_0_2_r1; // @[Reg.scala 16:16]
  reg [5:0] io_resp_0_2_r2; // @[Reg.scala 16:16]
  wire  _GEN_150 = 6'h1 == io_resp_0_2_r2 ? meta_array_1_2 : meta_array_0_2; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_151 = 6'h2 == io_resp_0_2_r2 ? meta_array_2_2 : _GEN_150; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_152 = 6'h3 == io_resp_0_2_r2 ? meta_array_3_2 : _GEN_151; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_153 = 6'h4 == io_resp_0_2_r2 ? meta_array_4_2 : _GEN_152; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_154 = 6'h5 == io_resp_0_2_r2 ? meta_array_5_2 : _GEN_153; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_155 = 6'h6 == io_resp_0_2_r2 ? meta_array_6_2 : _GEN_154; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_156 = 6'h7 == io_resp_0_2_r2 ? meta_array_7_2 : _GEN_155; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_157 = 6'h8 == io_resp_0_2_r2 ? meta_array_8_2 : _GEN_156; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_158 = 6'h9 == io_resp_0_2_r2 ? meta_array_9_2 : _GEN_157; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_159 = 6'ha == io_resp_0_2_r2 ? meta_array_10_2 : _GEN_158; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_160 = 6'hb == io_resp_0_2_r2 ? meta_array_11_2 : _GEN_159; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_161 = 6'hc == io_resp_0_2_r2 ? meta_array_12_2 : _GEN_160; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_162 = 6'hd == io_resp_0_2_r2 ? meta_array_13_2 : _GEN_161; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_163 = 6'he == io_resp_0_2_r2 ? meta_array_14_2 : _GEN_162; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_164 = 6'hf == io_resp_0_2_r2 ? meta_array_15_2 : _GEN_163; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_165 = 6'h10 == io_resp_0_2_r2 ? meta_array_16_2 : _GEN_164; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_166 = 6'h11 == io_resp_0_2_r2 ? meta_array_17_2 : _GEN_165; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_167 = 6'h12 == io_resp_0_2_r2 ? meta_array_18_2 : _GEN_166; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_168 = 6'h13 == io_resp_0_2_r2 ? meta_array_19_2 : _GEN_167; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_169 = 6'h14 == io_resp_0_2_r2 ? meta_array_20_2 : _GEN_168; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_170 = 6'h15 == io_resp_0_2_r2 ? meta_array_21_2 : _GEN_169; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_171 = 6'h16 == io_resp_0_2_r2 ? meta_array_22_2 : _GEN_170; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_172 = 6'h17 == io_resp_0_2_r2 ? meta_array_23_2 : _GEN_171; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_173 = 6'h18 == io_resp_0_2_r2 ? meta_array_24_2 : _GEN_172; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_174 = 6'h19 == io_resp_0_2_r2 ? meta_array_25_2 : _GEN_173; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_175 = 6'h1a == io_resp_0_2_r2 ? meta_array_26_2 : _GEN_174; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_176 = 6'h1b == io_resp_0_2_r2 ? meta_array_27_2 : _GEN_175; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_177 = 6'h1c == io_resp_0_2_r2 ? meta_array_28_2 : _GEN_176; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_178 = 6'h1d == io_resp_0_2_r2 ? meta_array_29_2 : _GEN_177; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_179 = 6'h1e == io_resp_0_2_r2 ? meta_array_30_2 : _GEN_178; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_180 = 6'h1f == io_resp_0_2_r2 ? meta_array_31_2 : _GEN_179; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_181 = 6'h20 == io_resp_0_2_r2 ? meta_array_32_2 : _GEN_180; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_182 = 6'h21 == io_resp_0_2_r2 ? meta_array_33_2 : _GEN_181; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_183 = 6'h22 == io_resp_0_2_r2 ? meta_array_34_2 : _GEN_182; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_184 = 6'h23 == io_resp_0_2_r2 ? meta_array_35_2 : _GEN_183; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_185 = 6'h24 == io_resp_0_2_r2 ? meta_array_36_2 : _GEN_184; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_186 = 6'h25 == io_resp_0_2_r2 ? meta_array_37_2 : _GEN_185; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_187 = 6'h26 == io_resp_0_2_r2 ? meta_array_38_2 : _GEN_186; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_188 = 6'h27 == io_resp_0_2_r2 ? meta_array_39_2 : _GEN_187; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_189 = 6'h28 == io_resp_0_2_r2 ? meta_array_40_2 : _GEN_188; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_190 = 6'h29 == io_resp_0_2_r2 ? meta_array_41_2 : _GEN_189; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_191 = 6'h2a == io_resp_0_2_r2 ? meta_array_42_2 : _GEN_190; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_192 = 6'h2b == io_resp_0_2_r2 ? meta_array_43_2 : _GEN_191; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_193 = 6'h2c == io_resp_0_2_r2 ? meta_array_44_2 : _GEN_192; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_194 = 6'h2d == io_resp_0_2_r2 ? meta_array_45_2 : _GEN_193; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_195 = 6'h2e == io_resp_0_2_r2 ? meta_array_46_2 : _GEN_194; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_196 = 6'h2f == io_resp_0_2_r2 ? meta_array_47_2 : _GEN_195; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_197 = 6'h30 == io_resp_0_2_r2 ? meta_array_48_2 : _GEN_196; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_198 = 6'h31 == io_resp_0_2_r2 ? meta_array_49_2 : _GEN_197; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_199 = 6'h32 == io_resp_0_2_r2 ? meta_array_50_2 : _GEN_198; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_200 = 6'h33 == io_resp_0_2_r2 ? meta_array_51_2 : _GEN_199; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_201 = 6'h34 == io_resp_0_2_r2 ? meta_array_52_2 : _GEN_200; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_202 = 6'h35 == io_resp_0_2_r2 ? meta_array_53_2 : _GEN_201; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_203 = 6'h36 == io_resp_0_2_r2 ? meta_array_54_2 : _GEN_202; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_204 = 6'h37 == io_resp_0_2_r2 ? meta_array_55_2 : _GEN_203; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_205 = 6'h38 == io_resp_0_2_r2 ? meta_array_56_2 : _GEN_204; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_206 = 6'h39 == io_resp_0_2_r2 ? meta_array_57_2 : _GEN_205; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_207 = 6'h3a == io_resp_0_2_r2 ? meta_array_58_2 : _GEN_206; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_208 = 6'h3b == io_resp_0_2_r2 ? meta_array_59_2 : _GEN_207; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_209 = 6'h3c == io_resp_0_2_r2 ? meta_array_60_2 : _GEN_208; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_210 = 6'h3d == io_resp_0_2_r2 ? meta_array_61_2 : _GEN_209; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_211 = 6'h3e == io_resp_0_2_r2 ? meta_array_62_2 : _GEN_210; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_212 = 6'h3f == io_resp_0_2_r2 ? meta_array_63_2 : _GEN_211; // @[AsynchronousMetaArray.scala 139:{25,25}]
  reg [5:0] s1_way_waddr_3_0_r; // @[Reg.scala 16:16]
  reg  s1_way_wen_3_0_REG; // @[AsynchronousMetaArray.scala 153:44]
  reg  s1_way_wdata_3_0_r; // @[Reg.scala 16:16]
  reg [5:0] s1_way_waddr_3_1_r; // @[Reg.scala 16:16]
  reg  s1_way_wen_3_1_REG; // @[AsynchronousMetaArray.scala 153:44]
  wire  read_way_bypass_3 = s1_way_wen_3_1_REG & s1_way_waddr_3_1_r == io_read_0_bits_idx | s1_way_wen_3_0_REG &
    s1_way_waddr_3_0_r == io_read_0_bits_idx; // @[AsynchronousMetaArray.scala 134:85 135:29]
  reg  s1_way_wdata_3_1_r; // @[Reg.scala 16:16]
  reg  io_resp_0_3_r; // @[Reg.scala 16:16]
  reg  io_resp_0_3_r1; // @[Reg.scala 16:16]
  reg [5:0] io_resp_0_3_r2; // @[Reg.scala 16:16]
  wire  _GEN_221 = 6'h1 == io_resp_0_3_r2 ? meta_array_1_3 : meta_array_0_3; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_222 = 6'h2 == io_resp_0_3_r2 ? meta_array_2_3 : _GEN_221; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_223 = 6'h3 == io_resp_0_3_r2 ? meta_array_3_3 : _GEN_222; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_224 = 6'h4 == io_resp_0_3_r2 ? meta_array_4_3 : _GEN_223; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_225 = 6'h5 == io_resp_0_3_r2 ? meta_array_5_3 : _GEN_224; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_226 = 6'h6 == io_resp_0_3_r2 ? meta_array_6_3 : _GEN_225; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_227 = 6'h7 == io_resp_0_3_r2 ? meta_array_7_3 : _GEN_226; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_228 = 6'h8 == io_resp_0_3_r2 ? meta_array_8_3 : _GEN_227; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_229 = 6'h9 == io_resp_0_3_r2 ? meta_array_9_3 : _GEN_228; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_230 = 6'ha == io_resp_0_3_r2 ? meta_array_10_3 : _GEN_229; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_231 = 6'hb == io_resp_0_3_r2 ? meta_array_11_3 : _GEN_230; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_232 = 6'hc == io_resp_0_3_r2 ? meta_array_12_3 : _GEN_231; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_233 = 6'hd == io_resp_0_3_r2 ? meta_array_13_3 : _GEN_232; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_234 = 6'he == io_resp_0_3_r2 ? meta_array_14_3 : _GEN_233; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_235 = 6'hf == io_resp_0_3_r2 ? meta_array_15_3 : _GEN_234; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_236 = 6'h10 == io_resp_0_3_r2 ? meta_array_16_3 : _GEN_235; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_237 = 6'h11 == io_resp_0_3_r2 ? meta_array_17_3 : _GEN_236; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_238 = 6'h12 == io_resp_0_3_r2 ? meta_array_18_3 : _GEN_237; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_239 = 6'h13 == io_resp_0_3_r2 ? meta_array_19_3 : _GEN_238; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_240 = 6'h14 == io_resp_0_3_r2 ? meta_array_20_3 : _GEN_239; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_241 = 6'h15 == io_resp_0_3_r2 ? meta_array_21_3 : _GEN_240; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_242 = 6'h16 == io_resp_0_3_r2 ? meta_array_22_3 : _GEN_241; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_243 = 6'h17 == io_resp_0_3_r2 ? meta_array_23_3 : _GEN_242; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_244 = 6'h18 == io_resp_0_3_r2 ? meta_array_24_3 : _GEN_243; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_245 = 6'h19 == io_resp_0_3_r2 ? meta_array_25_3 : _GEN_244; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_246 = 6'h1a == io_resp_0_3_r2 ? meta_array_26_3 : _GEN_245; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_247 = 6'h1b == io_resp_0_3_r2 ? meta_array_27_3 : _GEN_246; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_248 = 6'h1c == io_resp_0_3_r2 ? meta_array_28_3 : _GEN_247; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_249 = 6'h1d == io_resp_0_3_r2 ? meta_array_29_3 : _GEN_248; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_250 = 6'h1e == io_resp_0_3_r2 ? meta_array_30_3 : _GEN_249; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_251 = 6'h1f == io_resp_0_3_r2 ? meta_array_31_3 : _GEN_250; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_252 = 6'h20 == io_resp_0_3_r2 ? meta_array_32_3 : _GEN_251; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_253 = 6'h21 == io_resp_0_3_r2 ? meta_array_33_3 : _GEN_252; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_254 = 6'h22 == io_resp_0_3_r2 ? meta_array_34_3 : _GEN_253; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_255 = 6'h23 == io_resp_0_3_r2 ? meta_array_35_3 : _GEN_254; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_256 = 6'h24 == io_resp_0_3_r2 ? meta_array_36_3 : _GEN_255; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_257 = 6'h25 == io_resp_0_3_r2 ? meta_array_37_3 : _GEN_256; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_258 = 6'h26 == io_resp_0_3_r2 ? meta_array_38_3 : _GEN_257; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_259 = 6'h27 == io_resp_0_3_r2 ? meta_array_39_3 : _GEN_258; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_260 = 6'h28 == io_resp_0_3_r2 ? meta_array_40_3 : _GEN_259; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_261 = 6'h29 == io_resp_0_3_r2 ? meta_array_41_3 : _GEN_260; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_262 = 6'h2a == io_resp_0_3_r2 ? meta_array_42_3 : _GEN_261; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_263 = 6'h2b == io_resp_0_3_r2 ? meta_array_43_3 : _GEN_262; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_264 = 6'h2c == io_resp_0_3_r2 ? meta_array_44_3 : _GEN_263; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_265 = 6'h2d == io_resp_0_3_r2 ? meta_array_45_3 : _GEN_264; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_266 = 6'h2e == io_resp_0_3_r2 ? meta_array_46_3 : _GEN_265; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_267 = 6'h2f == io_resp_0_3_r2 ? meta_array_47_3 : _GEN_266; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_268 = 6'h30 == io_resp_0_3_r2 ? meta_array_48_3 : _GEN_267; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_269 = 6'h31 == io_resp_0_3_r2 ? meta_array_49_3 : _GEN_268; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_270 = 6'h32 == io_resp_0_3_r2 ? meta_array_50_3 : _GEN_269; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_271 = 6'h33 == io_resp_0_3_r2 ? meta_array_51_3 : _GEN_270; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_272 = 6'h34 == io_resp_0_3_r2 ? meta_array_52_3 : _GEN_271; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_273 = 6'h35 == io_resp_0_3_r2 ? meta_array_53_3 : _GEN_272; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_274 = 6'h36 == io_resp_0_3_r2 ? meta_array_54_3 : _GEN_273; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_275 = 6'h37 == io_resp_0_3_r2 ? meta_array_55_3 : _GEN_274; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_276 = 6'h38 == io_resp_0_3_r2 ? meta_array_56_3 : _GEN_275; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_277 = 6'h39 == io_resp_0_3_r2 ? meta_array_57_3 : _GEN_276; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_278 = 6'h3a == io_resp_0_3_r2 ? meta_array_58_3 : _GEN_277; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_279 = 6'h3b == io_resp_0_3_r2 ? meta_array_59_3 : _GEN_278; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_280 = 6'h3c == io_resp_0_3_r2 ? meta_array_60_3 : _GEN_279; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_281 = 6'h3d == io_resp_0_3_r2 ? meta_array_61_3 : _GEN_280; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_282 = 6'h3e == io_resp_0_3_r2 ? meta_array_62_3 : _GEN_281; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_283 = 6'h3f == io_resp_0_3_r2 ? meta_array_63_3 : _GEN_282; // @[AsynchronousMetaArray.scala 139:{25,25}]
  reg [5:0] s1_way_waddr_4_0_r; // @[Reg.scala 16:16]
  reg  s1_way_wen_4_0_REG; // @[AsynchronousMetaArray.scala 153:44]
  reg  s1_way_wdata_4_0_r; // @[Reg.scala 16:16]
  reg [5:0] s1_way_waddr_4_1_r; // @[Reg.scala 16:16]
  reg  s1_way_wen_4_1_REG; // @[AsynchronousMetaArray.scala 153:44]
  wire  read_way_bypass_4 = s1_way_wen_4_1_REG & s1_way_waddr_4_1_r == io_read_0_bits_idx | s1_way_wen_4_0_REG &
    s1_way_waddr_4_0_r == io_read_0_bits_idx; // @[AsynchronousMetaArray.scala 134:85 135:29]
  reg  s1_way_wdata_4_1_r; // @[Reg.scala 16:16]
  reg  io_resp_0_4_r; // @[Reg.scala 16:16]
  reg  io_resp_0_4_r1; // @[Reg.scala 16:16]
  reg [5:0] io_resp_0_4_r2; // @[Reg.scala 16:16]
  wire  _GEN_292 = 6'h1 == io_resp_0_4_r2 ? meta_array_1_4 : meta_array_0_4; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_293 = 6'h2 == io_resp_0_4_r2 ? meta_array_2_4 : _GEN_292; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_294 = 6'h3 == io_resp_0_4_r2 ? meta_array_3_4 : _GEN_293; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_295 = 6'h4 == io_resp_0_4_r2 ? meta_array_4_4 : _GEN_294; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_296 = 6'h5 == io_resp_0_4_r2 ? meta_array_5_4 : _GEN_295; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_297 = 6'h6 == io_resp_0_4_r2 ? meta_array_6_4 : _GEN_296; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_298 = 6'h7 == io_resp_0_4_r2 ? meta_array_7_4 : _GEN_297; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_299 = 6'h8 == io_resp_0_4_r2 ? meta_array_8_4 : _GEN_298; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_300 = 6'h9 == io_resp_0_4_r2 ? meta_array_9_4 : _GEN_299; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_301 = 6'ha == io_resp_0_4_r2 ? meta_array_10_4 : _GEN_300; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_302 = 6'hb == io_resp_0_4_r2 ? meta_array_11_4 : _GEN_301; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_303 = 6'hc == io_resp_0_4_r2 ? meta_array_12_4 : _GEN_302; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_304 = 6'hd == io_resp_0_4_r2 ? meta_array_13_4 : _GEN_303; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_305 = 6'he == io_resp_0_4_r2 ? meta_array_14_4 : _GEN_304; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_306 = 6'hf == io_resp_0_4_r2 ? meta_array_15_4 : _GEN_305; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_307 = 6'h10 == io_resp_0_4_r2 ? meta_array_16_4 : _GEN_306; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_308 = 6'h11 == io_resp_0_4_r2 ? meta_array_17_4 : _GEN_307; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_309 = 6'h12 == io_resp_0_4_r2 ? meta_array_18_4 : _GEN_308; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_310 = 6'h13 == io_resp_0_4_r2 ? meta_array_19_4 : _GEN_309; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_311 = 6'h14 == io_resp_0_4_r2 ? meta_array_20_4 : _GEN_310; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_312 = 6'h15 == io_resp_0_4_r2 ? meta_array_21_4 : _GEN_311; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_313 = 6'h16 == io_resp_0_4_r2 ? meta_array_22_4 : _GEN_312; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_314 = 6'h17 == io_resp_0_4_r2 ? meta_array_23_4 : _GEN_313; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_315 = 6'h18 == io_resp_0_4_r2 ? meta_array_24_4 : _GEN_314; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_316 = 6'h19 == io_resp_0_4_r2 ? meta_array_25_4 : _GEN_315; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_317 = 6'h1a == io_resp_0_4_r2 ? meta_array_26_4 : _GEN_316; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_318 = 6'h1b == io_resp_0_4_r2 ? meta_array_27_4 : _GEN_317; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_319 = 6'h1c == io_resp_0_4_r2 ? meta_array_28_4 : _GEN_318; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_320 = 6'h1d == io_resp_0_4_r2 ? meta_array_29_4 : _GEN_319; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_321 = 6'h1e == io_resp_0_4_r2 ? meta_array_30_4 : _GEN_320; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_322 = 6'h1f == io_resp_0_4_r2 ? meta_array_31_4 : _GEN_321; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_323 = 6'h20 == io_resp_0_4_r2 ? meta_array_32_4 : _GEN_322; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_324 = 6'h21 == io_resp_0_4_r2 ? meta_array_33_4 : _GEN_323; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_325 = 6'h22 == io_resp_0_4_r2 ? meta_array_34_4 : _GEN_324; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_326 = 6'h23 == io_resp_0_4_r2 ? meta_array_35_4 : _GEN_325; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_327 = 6'h24 == io_resp_0_4_r2 ? meta_array_36_4 : _GEN_326; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_328 = 6'h25 == io_resp_0_4_r2 ? meta_array_37_4 : _GEN_327; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_329 = 6'h26 == io_resp_0_4_r2 ? meta_array_38_4 : _GEN_328; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_330 = 6'h27 == io_resp_0_4_r2 ? meta_array_39_4 : _GEN_329; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_331 = 6'h28 == io_resp_0_4_r2 ? meta_array_40_4 : _GEN_330; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_332 = 6'h29 == io_resp_0_4_r2 ? meta_array_41_4 : _GEN_331; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_333 = 6'h2a == io_resp_0_4_r2 ? meta_array_42_4 : _GEN_332; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_334 = 6'h2b == io_resp_0_4_r2 ? meta_array_43_4 : _GEN_333; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_335 = 6'h2c == io_resp_0_4_r2 ? meta_array_44_4 : _GEN_334; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_336 = 6'h2d == io_resp_0_4_r2 ? meta_array_45_4 : _GEN_335; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_337 = 6'h2e == io_resp_0_4_r2 ? meta_array_46_4 : _GEN_336; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_338 = 6'h2f == io_resp_0_4_r2 ? meta_array_47_4 : _GEN_337; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_339 = 6'h30 == io_resp_0_4_r2 ? meta_array_48_4 : _GEN_338; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_340 = 6'h31 == io_resp_0_4_r2 ? meta_array_49_4 : _GEN_339; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_341 = 6'h32 == io_resp_0_4_r2 ? meta_array_50_4 : _GEN_340; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_342 = 6'h33 == io_resp_0_4_r2 ? meta_array_51_4 : _GEN_341; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_343 = 6'h34 == io_resp_0_4_r2 ? meta_array_52_4 : _GEN_342; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_344 = 6'h35 == io_resp_0_4_r2 ? meta_array_53_4 : _GEN_343; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_345 = 6'h36 == io_resp_0_4_r2 ? meta_array_54_4 : _GEN_344; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_346 = 6'h37 == io_resp_0_4_r2 ? meta_array_55_4 : _GEN_345; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_347 = 6'h38 == io_resp_0_4_r2 ? meta_array_56_4 : _GEN_346; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_348 = 6'h39 == io_resp_0_4_r2 ? meta_array_57_4 : _GEN_347; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_349 = 6'h3a == io_resp_0_4_r2 ? meta_array_58_4 : _GEN_348; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_350 = 6'h3b == io_resp_0_4_r2 ? meta_array_59_4 : _GEN_349; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_351 = 6'h3c == io_resp_0_4_r2 ? meta_array_60_4 : _GEN_350; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_352 = 6'h3d == io_resp_0_4_r2 ? meta_array_61_4 : _GEN_351; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_353 = 6'h3e == io_resp_0_4_r2 ? meta_array_62_4 : _GEN_352; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_354 = 6'h3f == io_resp_0_4_r2 ? meta_array_63_4 : _GEN_353; // @[AsynchronousMetaArray.scala 139:{25,25}]
  reg [5:0] s1_way_waddr_5_0_r; // @[Reg.scala 16:16]
  reg  s1_way_wen_5_0_REG; // @[AsynchronousMetaArray.scala 153:44]
  reg  s1_way_wdata_5_0_r; // @[Reg.scala 16:16]
  reg [5:0] s1_way_waddr_5_1_r; // @[Reg.scala 16:16]
  reg  s1_way_wen_5_1_REG; // @[AsynchronousMetaArray.scala 153:44]
  wire  read_way_bypass_5 = s1_way_wen_5_1_REG & s1_way_waddr_5_1_r == io_read_0_bits_idx | s1_way_wen_5_0_REG &
    s1_way_waddr_5_0_r == io_read_0_bits_idx; // @[AsynchronousMetaArray.scala 134:85 135:29]
  reg  s1_way_wdata_5_1_r; // @[Reg.scala 16:16]
  reg  io_resp_0_5_r; // @[Reg.scala 16:16]
  reg  io_resp_0_5_r1; // @[Reg.scala 16:16]
  reg [5:0] io_resp_0_5_r2; // @[Reg.scala 16:16]
  wire  _GEN_363 = 6'h1 == io_resp_0_5_r2 ? meta_array_1_5 : meta_array_0_5; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_364 = 6'h2 == io_resp_0_5_r2 ? meta_array_2_5 : _GEN_363; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_365 = 6'h3 == io_resp_0_5_r2 ? meta_array_3_5 : _GEN_364; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_366 = 6'h4 == io_resp_0_5_r2 ? meta_array_4_5 : _GEN_365; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_367 = 6'h5 == io_resp_0_5_r2 ? meta_array_5_5 : _GEN_366; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_368 = 6'h6 == io_resp_0_5_r2 ? meta_array_6_5 : _GEN_367; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_369 = 6'h7 == io_resp_0_5_r2 ? meta_array_7_5 : _GEN_368; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_370 = 6'h8 == io_resp_0_5_r2 ? meta_array_8_5 : _GEN_369; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_371 = 6'h9 == io_resp_0_5_r2 ? meta_array_9_5 : _GEN_370; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_372 = 6'ha == io_resp_0_5_r2 ? meta_array_10_5 : _GEN_371; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_373 = 6'hb == io_resp_0_5_r2 ? meta_array_11_5 : _GEN_372; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_374 = 6'hc == io_resp_0_5_r2 ? meta_array_12_5 : _GEN_373; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_375 = 6'hd == io_resp_0_5_r2 ? meta_array_13_5 : _GEN_374; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_376 = 6'he == io_resp_0_5_r2 ? meta_array_14_5 : _GEN_375; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_377 = 6'hf == io_resp_0_5_r2 ? meta_array_15_5 : _GEN_376; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_378 = 6'h10 == io_resp_0_5_r2 ? meta_array_16_5 : _GEN_377; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_379 = 6'h11 == io_resp_0_5_r2 ? meta_array_17_5 : _GEN_378; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_380 = 6'h12 == io_resp_0_5_r2 ? meta_array_18_5 : _GEN_379; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_381 = 6'h13 == io_resp_0_5_r2 ? meta_array_19_5 : _GEN_380; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_382 = 6'h14 == io_resp_0_5_r2 ? meta_array_20_5 : _GEN_381; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_383 = 6'h15 == io_resp_0_5_r2 ? meta_array_21_5 : _GEN_382; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_384 = 6'h16 == io_resp_0_5_r2 ? meta_array_22_5 : _GEN_383; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_385 = 6'h17 == io_resp_0_5_r2 ? meta_array_23_5 : _GEN_384; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_386 = 6'h18 == io_resp_0_5_r2 ? meta_array_24_5 : _GEN_385; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_387 = 6'h19 == io_resp_0_5_r2 ? meta_array_25_5 : _GEN_386; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_388 = 6'h1a == io_resp_0_5_r2 ? meta_array_26_5 : _GEN_387; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_389 = 6'h1b == io_resp_0_5_r2 ? meta_array_27_5 : _GEN_388; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_390 = 6'h1c == io_resp_0_5_r2 ? meta_array_28_5 : _GEN_389; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_391 = 6'h1d == io_resp_0_5_r2 ? meta_array_29_5 : _GEN_390; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_392 = 6'h1e == io_resp_0_5_r2 ? meta_array_30_5 : _GEN_391; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_393 = 6'h1f == io_resp_0_5_r2 ? meta_array_31_5 : _GEN_392; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_394 = 6'h20 == io_resp_0_5_r2 ? meta_array_32_5 : _GEN_393; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_395 = 6'h21 == io_resp_0_5_r2 ? meta_array_33_5 : _GEN_394; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_396 = 6'h22 == io_resp_0_5_r2 ? meta_array_34_5 : _GEN_395; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_397 = 6'h23 == io_resp_0_5_r2 ? meta_array_35_5 : _GEN_396; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_398 = 6'h24 == io_resp_0_5_r2 ? meta_array_36_5 : _GEN_397; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_399 = 6'h25 == io_resp_0_5_r2 ? meta_array_37_5 : _GEN_398; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_400 = 6'h26 == io_resp_0_5_r2 ? meta_array_38_5 : _GEN_399; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_401 = 6'h27 == io_resp_0_5_r2 ? meta_array_39_5 : _GEN_400; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_402 = 6'h28 == io_resp_0_5_r2 ? meta_array_40_5 : _GEN_401; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_403 = 6'h29 == io_resp_0_5_r2 ? meta_array_41_5 : _GEN_402; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_404 = 6'h2a == io_resp_0_5_r2 ? meta_array_42_5 : _GEN_403; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_405 = 6'h2b == io_resp_0_5_r2 ? meta_array_43_5 : _GEN_404; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_406 = 6'h2c == io_resp_0_5_r2 ? meta_array_44_5 : _GEN_405; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_407 = 6'h2d == io_resp_0_5_r2 ? meta_array_45_5 : _GEN_406; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_408 = 6'h2e == io_resp_0_5_r2 ? meta_array_46_5 : _GEN_407; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_409 = 6'h2f == io_resp_0_5_r2 ? meta_array_47_5 : _GEN_408; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_410 = 6'h30 == io_resp_0_5_r2 ? meta_array_48_5 : _GEN_409; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_411 = 6'h31 == io_resp_0_5_r2 ? meta_array_49_5 : _GEN_410; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_412 = 6'h32 == io_resp_0_5_r2 ? meta_array_50_5 : _GEN_411; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_413 = 6'h33 == io_resp_0_5_r2 ? meta_array_51_5 : _GEN_412; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_414 = 6'h34 == io_resp_0_5_r2 ? meta_array_52_5 : _GEN_413; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_415 = 6'h35 == io_resp_0_5_r2 ? meta_array_53_5 : _GEN_414; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_416 = 6'h36 == io_resp_0_5_r2 ? meta_array_54_5 : _GEN_415; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_417 = 6'h37 == io_resp_0_5_r2 ? meta_array_55_5 : _GEN_416; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_418 = 6'h38 == io_resp_0_5_r2 ? meta_array_56_5 : _GEN_417; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_419 = 6'h39 == io_resp_0_5_r2 ? meta_array_57_5 : _GEN_418; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_420 = 6'h3a == io_resp_0_5_r2 ? meta_array_58_5 : _GEN_419; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_421 = 6'h3b == io_resp_0_5_r2 ? meta_array_59_5 : _GEN_420; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_422 = 6'h3c == io_resp_0_5_r2 ? meta_array_60_5 : _GEN_421; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_423 = 6'h3d == io_resp_0_5_r2 ? meta_array_61_5 : _GEN_422; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_424 = 6'h3e == io_resp_0_5_r2 ? meta_array_62_5 : _GEN_423; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_425 = 6'h3f == io_resp_0_5_r2 ? meta_array_63_5 : _GEN_424; // @[AsynchronousMetaArray.scala 139:{25,25}]
  reg [5:0] s1_way_waddr_6_0_r; // @[Reg.scala 16:16]
  reg  s1_way_wen_6_0_REG; // @[AsynchronousMetaArray.scala 153:44]
  reg  s1_way_wdata_6_0_r; // @[Reg.scala 16:16]
  reg [5:0] s1_way_waddr_6_1_r; // @[Reg.scala 16:16]
  reg  s1_way_wen_6_1_REG; // @[AsynchronousMetaArray.scala 153:44]
  wire  read_way_bypass_6 = s1_way_wen_6_1_REG & s1_way_waddr_6_1_r == io_read_0_bits_idx | s1_way_wen_6_0_REG &
    s1_way_waddr_6_0_r == io_read_0_bits_idx; // @[AsynchronousMetaArray.scala 134:85 135:29]
  reg  s1_way_wdata_6_1_r; // @[Reg.scala 16:16]
  reg  io_resp_0_6_r; // @[Reg.scala 16:16]
  reg  io_resp_0_6_r1; // @[Reg.scala 16:16]
  reg [5:0] io_resp_0_6_r2; // @[Reg.scala 16:16]
  wire  _GEN_434 = 6'h1 == io_resp_0_6_r2 ? meta_array_1_6 : meta_array_0_6; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_435 = 6'h2 == io_resp_0_6_r2 ? meta_array_2_6 : _GEN_434; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_436 = 6'h3 == io_resp_0_6_r2 ? meta_array_3_6 : _GEN_435; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_437 = 6'h4 == io_resp_0_6_r2 ? meta_array_4_6 : _GEN_436; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_438 = 6'h5 == io_resp_0_6_r2 ? meta_array_5_6 : _GEN_437; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_439 = 6'h6 == io_resp_0_6_r2 ? meta_array_6_6 : _GEN_438; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_440 = 6'h7 == io_resp_0_6_r2 ? meta_array_7_6 : _GEN_439; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_441 = 6'h8 == io_resp_0_6_r2 ? meta_array_8_6 : _GEN_440; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_442 = 6'h9 == io_resp_0_6_r2 ? meta_array_9_6 : _GEN_441; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_443 = 6'ha == io_resp_0_6_r2 ? meta_array_10_6 : _GEN_442; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_444 = 6'hb == io_resp_0_6_r2 ? meta_array_11_6 : _GEN_443; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_445 = 6'hc == io_resp_0_6_r2 ? meta_array_12_6 : _GEN_444; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_446 = 6'hd == io_resp_0_6_r2 ? meta_array_13_6 : _GEN_445; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_447 = 6'he == io_resp_0_6_r2 ? meta_array_14_6 : _GEN_446; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_448 = 6'hf == io_resp_0_6_r2 ? meta_array_15_6 : _GEN_447; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_449 = 6'h10 == io_resp_0_6_r2 ? meta_array_16_6 : _GEN_448; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_450 = 6'h11 == io_resp_0_6_r2 ? meta_array_17_6 : _GEN_449; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_451 = 6'h12 == io_resp_0_6_r2 ? meta_array_18_6 : _GEN_450; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_452 = 6'h13 == io_resp_0_6_r2 ? meta_array_19_6 : _GEN_451; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_453 = 6'h14 == io_resp_0_6_r2 ? meta_array_20_6 : _GEN_452; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_454 = 6'h15 == io_resp_0_6_r2 ? meta_array_21_6 : _GEN_453; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_455 = 6'h16 == io_resp_0_6_r2 ? meta_array_22_6 : _GEN_454; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_456 = 6'h17 == io_resp_0_6_r2 ? meta_array_23_6 : _GEN_455; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_457 = 6'h18 == io_resp_0_6_r2 ? meta_array_24_6 : _GEN_456; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_458 = 6'h19 == io_resp_0_6_r2 ? meta_array_25_6 : _GEN_457; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_459 = 6'h1a == io_resp_0_6_r2 ? meta_array_26_6 : _GEN_458; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_460 = 6'h1b == io_resp_0_6_r2 ? meta_array_27_6 : _GEN_459; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_461 = 6'h1c == io_resp_0_6_r2 ? meta_array_28_6 : _GEN_460; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_462 = 6'h1d == io_resp_0_6_r2 ? meta_array_29_6 : _GEN_461; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_463 = 6'h1e == io_resp_0_6_r2 ? meta_array_30_6 : _GEN_462; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_464 = 6'h1f == io_resp_0_6_r2 ? meta_array_31_6 : _GEN_463; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_465 = 6'h20 == io_resp_0_6_r2 ? meta_array_32_6 : _GEN_464; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_466 = 6'h21 == io_resp_0_6_r2 ? meta_array_33_6 : _GEN_465; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_467 = 6'h22 == io_resp_0_6_r2 ? meta_array_34_6 : _GEN_466; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_468 = 6'h23 == io_resp_0_6_r2 ? meta_array_35_6 : _GEN_467; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_469 = 6'h24 == io_resp_0_6_r2 ? meta_array_36_6 : _GEN_468; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_470 = 6'h25 == io_resp_0_6_r2 ? meta_array_37_6 : _GEN_469; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_471 = 6'h26 == io_resp_0_6_r2 ? meta_array_38_6 : _GEN_470; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_472 = 6'h27 == io_resp_0_6_r2 ? meta_array_39_6 : _GEN_471; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_473 = 6'h28 == io_resp_0_6_r2 ? meta_array_40_6 : _GEN_472; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_474 = 6'h29 == io_resp_0_6_r2 ? meta_array_41_6 : _GEN_473; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_475 = 6'h2a == io_resp_0_6_r2 ? meta_array_42_6 : _GEN_474; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_476 = 6'h2b == io_resp_0_6_r2 ? meta_array_43_6 : _GEN_475; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_477 = 6'h2c == io_resp_0_6_r2 ? meta_array_44_6 : _GEN_476; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_478 = 6'h2d == io_resp_0_6_r2 ? meta_array_45_6 : _GEN_477; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_479 = 6'h2e == io_resp_0_6_r2 ? meta_array_46_6 : _GEN_478; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_480 = 6'h2f == io_resp_0_6_r2 ? meta_array_47_6 : _GEN_479; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_481 = 6'h30 == io_resp_0_6_r2 ? meta_array_48_6 : _GEN_480; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_482 = 6'h31 == io_resp_0_6_r2 ? meta_array_49_6 : _GEN_481; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_483 = 6'h32 == io_resp_0_6_r2 ? meta_array_50_6 : _GEN_482; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_484 = 6'h33 == io_resp_0_6_r2 ? meta_array_51_6 : _GEN_483; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_485 = 6'h34 == io_resp_0_6_r2 ? meta_array_52_6 : _GEN_484; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_486 = 6'h35 == io_resp_0_6_r2 ? meta_array_53_6 : _GEN_485; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_487 = 6'h36 == io_resp_0_6_r2 ? meta_array_54_6 : _GEN_486; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_488 = 6'h37 == io_resp_0_6_r2 ? meta_array_55_6 : _GEN_487; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_489 = 6'h38 == io_resp_0_6_r2 ? meta_array_56_6 : _GEN_488; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_490 = 6'h39 == io_resp_0_6_r2 ? meta_array_57_6 : _GEN_489; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_491 = 6'h3a == io_resp_0_6_r2 ? meta_array_58_6 : _GEN_490; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_492 = 6'h3b == io_resp_0_6_r2 ? meta_array_59_6 : _GEN_491; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_493 = 6'h3c == io_resp_0_6_r2 ? meta_array_60_6 : _GEN_492; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_494 = 6'h3d == io_resp_0_6_r2 ? meta_array_61_6 : _GEN_493; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_495 = 6'h3e == io_resp_0_6_r2 ? meta_array_62_6 : _GEN_494; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_496 = 6'h3f == io_resp_0_6_r2 ? meta_array_63_6 : _GEN_495; // @[AsynchronousMetaArray.scala 139:{25,25}]
  reg [5:0] s1_way_waddr_7_0_r; // @[Reg.scala 16:16]
  reg  s1_way_wen_7_0_REG; // @[AsynchronousMetaArray.scala 153:44]
  reg  s1_way_wdata_7_0_r; // @[Reg.scala 16:16]
  reg [5:0] s1_way_waddr_7_1_r; // @[Reg.scala 16:16]
  reg  s1_way_wen_7_1_REG; // @[AsynchronousMetaArray.scala 153:44]
  wire  read_way_bypass_7 = s1_way_wen_7_1_REG & s1_way_waddr_7_1_r == io_read_0_bits_idx | s1_way_wen_7_0_REG &
    s1_way_waddr_7_0_r == io_read_0_bits_idx; // @[AsynchronousMetaArray.scala 134:85 135:29]
  reg  s1_way_wdata_7_1_r; // @[Reg.scala 16:16]
  reg  io_resp_0_7_r; // @[Reg.scala 16:16]
  reg  io_resp_0_7_r1; // @[Reg.scala 16:16]
  reg [5:0] io_resp_0_7_r2; // @[Reg.scala 16:16]
  wire  _GEN_505 = 6'h1 == io_resp_0_7_r2 ? meta_array_1_7 : meta_array_0_7; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_506 = 6'h2 == io_resp_0_7_r2 ? meta_array_2_7 : _GEN_505; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_507 = 6'h3 == io_resp_0_7_r2 ? meta_array_3_7 : _GEN_506; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_508 = 6'h4 == io_resp_0_7_r2 ? meta_array_4_7 : _GEN_507; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_509 = 6'h5 == io_resp_0_7_r2 ? meta_array_5_7 : _GEN_508; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_510 = 6'h6 == io_resp_0_7_r2 ? meta_array_6_7 : _GEN_509; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_511 = 6'h7 == io_resp_0_7_r2 ? meta_array_7_7 : _GEN_510; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_512 = 6'h8 == io_resp_0_7_r2 ? meta_array_8_7 : _GEN_511; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_513 = 6'h9 == io_resp_0_7_r2 ? meta_array_9_7 : _GEN_512; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_514 = 6'ha == io_resp_0_7_r2 ? meta_array_10_7 : _GEN_513; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_515 = 6'hb == io_resp_0_7_r2 ? meta_array_11_7 : _GEN_514; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_516 = 6'hc == io_resp_0_7_r2 ? meta_array_12_7 : _GEN_515; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_517 = 6'hd == io_resp_0_7_r2 ? meta_array_13_7 : _GEN_516; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_518 = 6'he == io_resp_0_7_r2 ? meta_array_14_7 : _GEN_517; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_519 = 6'hf == io_resp_0_7_r2 ? meta_array_15_7 : _GEN_518; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_520 = 6'h10 == io_resp_0_7_r2 ? meta_array_16_7 : _GEN_519; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_521 = 6'h11 == io_resp_0_7_r2 ? meta_array_17_7 : _GEN_520; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_522 = 6'h12 == io_resp_0_7_r2 ? meta_array_18_7 : _GEN_521; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_523 = 6'h13 == io_resp_0_7_r2 ? meta_array_19_7 : _GEN_522; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_524 = 6'h14 == io_resp_0_7_r2 ? meta_array_20_7 : _GEN_523; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_525 = 6'h15 == io_resp_0_7_r2 ? meta_array_21_7 : _GEN_524; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_526 = 6'h16 == io_resp_0_7_r2 ? meta_array_22_7 : _GEN_525; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_527 = 6'h17 == io_resp_0_7_r2 ? meta_array_23_7 : _GEN_526; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_528 = 6'h18 == io_resp_0_7_r2 ? meta_array_24_7 : _GEN_527; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_529 = 6'h19 == io_resp_0_7_r2 ? meta_array_25_7 : _GEN_528; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_530 = 6'h1a == io_resp_0_7_r2 ? meta_array_26_7 : _GEN_529; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_531 = 6'h1b == io_resp_0_7_r2 ? meta_array_27_7 : _GEN_530; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_532 = 6'h1c == io_resp_0_7_r2 ? meta_array_28_7 : _GEN_531; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_533 = 6'h1d == io_resp_0_7_r2 ? meta_array_29_7 : _GEN_532; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_534 = 6'h1e == io_resp_0_7_r2 ? meta_array_30_7 : _GEN_533; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_535 = 6'h1f == io_resp_0_7_r2 ? meta_array_31_7 : _GEN_534; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_536 = 6'h20 == io_resp_0_7_r2 ? meta_array_32_7 : _GEN_535; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_537 = 6'h21 == io_resp_0_7_r2 ? meta_array_33_7 : _GEN_536; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_538 = 6'h22 == io_resp_0_7_r2 ? meta_array_34_7 : _GEN_537; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_539 = 6'h23 == io_resp_0_7_r2 ? meta_array_35_7 : _GEN_538; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_540 = 6'h24 == io_resp_0_7_r2 ? meta_array_36_7 : _GEN_539; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_541 = 6'h25 == io_resp_0_7_r2 ? meta_array_37_7 : _GEN_540; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_542 = 6'h26 == io_resp_0_7_r2 ? meta_array_38_7 : _GEN_541; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_543 = 6'h27 == io_resp_0_7_r2 ? meta_array_39_7 : _GEN_542; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_544 = 6'h28 == io_resp_0_7_r2 ? meta_array_40_7 : _GEN_543; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_545 = 6'h29 == io_resp_0_7_r2 ? meta_array_41_7 : _GEN_544; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_546 = 6'h2a == io_resp_0_7_r2 ? meta_array_42_7 : _GEN_545; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_547 = 6'h2b == io_resp_0_7_r2 ? meta_array_43_7 : _GEN_546; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_548 = 6'h2c == io_resp_0_7_r2 ? meta_array_44_7 : _GEN_547; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_549 = 6'h2d == io_resp_0_7_r2 ? meta_array_45_7 : _GEN_548; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_550 = 6'h2e == io_resp_0_7_r2 ? meta_array_46_7 : _GEN_549; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_551 = 6'h2f == io_resp_0_7_r2 ? meta_array_47_7 : _GEN_550; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_552 = 6'h30 == io_resp_0_7_r2 ? meta_array_48_7 : _GEN_551; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_553 = 6'h31 == io_resp_0_7_r2 ? meta_array_49_7 : _GEN_552; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_554 = 6'h32 == io_resp_0_7_r2 ? meta_array_50_7 : _GEN_553; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_555 = 6'h33 == io_resp_0_7_r2 ? meta_array_51_7 : _GEN_554; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_556 = 6'h34 == io_resp_0_7_r2 ? meta_array_52_7 : _GEN_555; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_557 = 6'h35 == io_resp_0_7_r2 ? meta_array_53_7 : _GEN_556; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_558 = 6'h36 == io_resp_0_7_r2 ? meta_array_54_7 : _GEN_557; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_559 = 6'h37 == io_resp_0_7_r2 ? meta_array_55_7 : _GEN_558; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_560 = 6'h38 == io_resp_0_7_r2 ? meta_array_56_7 : _GEN_559; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_561 = 6'h39 == io_resp_0_7_r2 ? meta_array_57_7 : _GEN_560; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_562 = 6'h3a == io_resp_0_7_r2 ? meta_array_58_7 : _GEN_561; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_563 = 6'h3b == io_resp_0_7_r2 ? meta_array_59_7 : _GEN_562; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_564 = 6'h3c == io_resp_0_7_r2 ? meta_array_60_7 : _GEN_563; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_565 = 6'h3d == io_resp_0_7_r2 ? meta_array_61_7 : _GEN_564; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_566 = 6'h3e == io_resp_0_7_r2 ? meta_array_62_7 : _GEN_565; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_567 = 6'h3f == io_resp_0_7_r2 ? meta_array_63_7 : _GEN_566; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  read_way_bypass_8 = s1_way_wen_0_1_REG & s1_way_waddr_0_1_r == io_read_1_bits_idx | s1_way_wen_0_0_REG &
    s1_way_waddr_0_0_r == io_read_1_bits_idx; // @[AsynchronousMetaArray.scala 134:85 135:29]
  reg  io_resp_1_0_r; // @[Reg.scala 16:16]
  reg  io_resp_1_0_r1; // @[Reg.scala 16:16]
  reg [5:0] io_resp_1_0_r2; // @[Reg.scala 16:16]
  wire  _GEN_576 = 6'h1 == io_resp_1_0_r2 ? meta_array_1_0 : meta_array_0_0; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_577 = 6'h2 == io_resp_1_0_r2 ? meta_array_2_0 : _GEN_576; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_578 = 6'h3 == io_resp_1_0_r2 ? meta_array_3_0 : _GEN_577; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_579 = 6'h4 == io_resp_1_0_r2 ? meta_array_4_0 : _GEN_578; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_580 = 6'h5 == io_resp_1_0_r2 ? meta_array_5_0 : _GEN_579; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_581 = 6'h6 == io_resp_1_0_r2 ? meta_array_6_0 : _GEN_580; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_582 = 6'h7 == io_resp_1_0_r2 ? meta_array_7_0 : _GEN_581; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_583 = 6'h8 == io_resp_1_0_r2 ? meta_array_8_0 : _GEN_582; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_584 = 6'h9 == io_resp_1_0_r2 ? meta_array_9_0 : _GEN_583; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_585 = 6'ha == io_resp_1_0_r2 ? meta_array_10_0 : _GEN_584; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_586 = 6'hb == io_resp_1_0_r2 ? meta_array_11_0 : _GEN_585; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_587 = 6'hc == io_resp_1_0_r2 ? meta_array_12_0 : _GEN_586; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_588 = 6'hd == io_resp_1_0_r2 ? meta_array_13_0 : _GEN_587; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_589 = 6'he == io_resp_1_0_r2 ? meta_array_14_0 : _GEN_588; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_590 = 6'hf == io_resp_1_0_r2 ? meta_array_15_0 : _GEN_589; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_591 = 6'h10 == io_resp_1_0_r2 ? meta_array_16_0 : _GEN_590; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_592 = 6'h11 == io_resp_1_0_r2 ? meta_array_17_0 : _GEN_591; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_593 = 6'h12 == io_resp_1_0_r2 ? meta_array_18_0 : _GEN_592; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_594 = 6'h13 == io_resp_1_0_r2 ? meta_array_19_0 : _GEN_593; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_595 = 6'h14 == io_resp_1_0_r2 ? meta_array_20_0 : _GEN_594; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_596 = 6'h15 == io_resp_1_0_r2 ? meta_array_21_0 : _GEN_595; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_597 = 6'h16 == io_resp_1_0_r2 ? meta_array_22_0 : _GEN_596; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_598 = 6'h17 == io_resp_1_0_r2 ? meta_array_23_0 : _GEN_597; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_599 = 6'h18 == io_resp_1_0_r2 ? meta_array_24_0 : _GEN_598; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_600 = 6'h19 == io_resp_1_0_r2 ? meta_array_25_0 : _GEN_599; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_601 = 6'h1a == io_resp_1_0_r2 ? meta_array_26_0 : _GEN_600; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_602 = 6'h1b == io_resp_1_0_r2 ? meta_array_27_0 : _GEN_601; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_603 = 6'h1c == io_resp_1_0_r2 ? meta_array_28_0 : _GEN_602; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_604 = 6'h1d == io_resp_1_0_r2 ? meta_array_29_0 : _GEN_603; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_605 = 6'h1e == io_resp_1_0_r2 ? meta_array_30_0 : _GEN_604; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_606 = 6'h1f == io_resp_1_0_r2 ? meta_array_31_0 : _GEN_605; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_607 = 6'h20 == io_resp_1_0_r2 ? meta_array_32_0 : _GEN_606; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_608 = 6'h21 == io_resp_1_0_r2 ? meta_array_33_0 : _GEN_607; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_609 = 6'h22 == io_resp_1_0_r2 ? meta_array_34_0 : _GEN_608; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_610 = 6'h23 == io_resp_1_0_r2 ? meta_array_35_0 : _GEN_609; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_611 = 6'h24 == io_resp_1_0_r2 ? meta_array_36_0 : _GEN_610; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_612 = 6'h25 == io_resp_1_0_r2 ? meta_array_37_0 : _GEN_611; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_613 = 6'h26 == io_resp_1_0_r2 ? meta_array_38_0 : _GEN_612; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_614 = 6'h27 == io_resp_1_0_r2 ? meta_array_39_0 : _GEN_613; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_615 = 6'h28 == io_resp_1_0_r2 ? meta_array_40_0 : _GEN_614; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_616 = 6'h29 == io_resp_1_0_r2 ? meta_array_41_0 : _GEN_615; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_617 = 6'h2a == io_resp_1_0_r2 ? meta_array_42_0 : _GEN_616; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_618 = 6'h2b == io_resp_1_0_r2 ? meta_array_43_0 : _GEN_617; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_619 = 6'h2c == io_resp_1_0_r2 ? meta_array_44_0 : _GEN_618; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_620 = 6'h2d == io_resp_1_0_r2 ? meta_array_45_0 : _GEN_619; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_621 = 6'h2e == io_resp_1_0_r2 ? meta_array_46_0 : _GEN_620; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_622 = 6'h2f == io_resp_1_0_r2 ? meta_array_47_0 : _GEN_621; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_623 = 6'h30 == io_resp_1_0_r2 ? meta_array_48_0 : _GEN_622; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_624 = 6'h31 == io_resp_1_0_r2 ? meta_array_49_0 : _GEN_623; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_625 = 6'h32 == io_resp_1_0_r2 ? meta_array_50_0 : _GEN_624; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_626 = 6'h33 == io_resp_1_0_r2 ? meta_array_51_0 : _GEN_625; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_627 = 6'h34 == io_resp_1_0_r2 ? meta_array_52_0 : _GEN_626; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_628 = 6'h35 == io_resp_1_0_r2 ? meta_array_53_0 : _GEN_627; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_629 = 6'h36 == io_resp_1_0_r2 ? meta_array_54_0 : _GEN_628; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_630 = 6'h37 == io_resp_1_0_r2 ? meta_array_55_0 : _GEN_629; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_631 = 6'h38 == io_resp_1_0_r2 ? meta_array_56_0 : _GEN_630; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_632 = 6'h39 == io_resp_1_0_r2 ? meta_array_57_0 : _GEN_631; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_633 = 6'h3a == io_resp_1_0_r2 ? meta_array_58_0 : _GEN_632; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_634 = 6'h3b == io_resp_1_0_r2 ? meta_array_59_0 : _GEN_633; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_635 = 6'h3c == io_resp_1_0_r2 ? meta_array_60_0 : _GEN_634; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_636 = 6'h3d == io_resp_1_0_r2 ? meta_array_61_0 : _GEN_635; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_637 = 6'h3e == io_resp_1_0_r2 ? meta_array_62_0 : _GEN_636; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_638 = 6'h3f == io_resp_1_0_r2 ? meta_array_63_0 : _GEN_637; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  read_way_bypass_9 = s1_way_wen_1_1_REG & s1_way_waddr_1_1_r == io_read_1_bits_idx | s1_way_wen_1_0_REG &
    s1_way_waddr_1_0_r == io_read_1_bits_idx; // @[AsynchronousMetaArray.scala 134:85 135:29]
  reg  io_resp_1_1_r; // @[Reg.scala 16:16]
  reg  io_resp_1_1_r1; // @[Reg.scala 16:16]
  reg [5:0] io_resp_1_1_r2; // @[Reg.scala 16:16]
  wire  _GEN_647 = 6'h1 == io_resp_1_1_r2 ? meta_array_1_1 : meta_array_0_1; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_648 = 6'h2 == io_resp_1_1_r2 ? meta_array_2_1 : _GEN_647; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_649 = 6'h3 == io_resp_1_1_r2 ? meta_array_3_1 : _GEN_648; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_650 = 6'h4 == io_resp_1_1_r2 ? meta_array_4_1 : _GEN_649; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_651 = 6'h5 == io_resp_1_1_r2 ? meta_array_5_1 : _GEN_650; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_652 = 6'h6 == io_resp_1_1_r2 ? meta_array_6_1 : _GEN_651; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_653 = 6'h7 == io_resp_1_1_r2 ? meta_array_7_1 : _GEN_652; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_654 = 6'h8 == io_resp_1_1_r2 ? meta_array_8_1 : _GEN_653; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_655 = 6'h9 == io_resp_1_1_r2 ? meta_array_9_1 : _GEN_654; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_656 = 6'ha == io_resp_1_1_r2 ? meta_array_10_1 : _GEN_655; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_657 = 6'hb == io_resp_1_1_r2 ? meta_array_11_1 : _GEN_656; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_658 = 6'hc == io_resp_1_1_r2 ? meta_array_12_1 : _GEN_657; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_659 = 6'hd == io_resp_1_1_r2 ? meta_array_13_1 : _GEN_658; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_660 = 6'he == io_resp_1_1_r2 ? meta_array_14_1 : _GEN_659; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_661 = 6'hf == io_resp_1_1_r2 ? meta_array_15_1 : _GEN_660; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_662 = 6'h10 == io_resp_1_1_r2 ? meta_array_16_1 : _GEN_661; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_663 = 6'h11 == io_resp_1_1_r2 ? meta_array_17_1 : _GEN_662; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_664 = 6'h12 == io_resp_1_1_r2 ? meta_array_18_1 : _GEN_663; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_665 = 6'h13 == io_resp_1_1_r2 ? meta_array_19_1 : _GEN_664; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_666 = 6'h14 == io_resp_1_1_r2 ? meta_array_20_1 : _GEN_665; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_667 = 6'h15 == io_resp_1_1_r2 ? meta_array_21_1 : _GEN_666; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_668 = 6'h16 == io_resp_1_1_r2 ? meta_array_22_1 : _GEN_667; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_669 = 6'h17 == io_resp_1_1_r2 ? meta_array_23_1 : _GEN_668; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_670 = 6'h18 == io_resp_1_1_r2 ? meta_array_24_1 : _GEN_669; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_671 = 6'h19 == io_resp_1_1_r2 ? meta_array_25_1 : _GEN_670; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_672 = 6'h1a == io_resp_1_1_r2 ? meta_array_26_1 : _GEN_671; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_673 = 6'h1b == io_resp_1_1_r2 ? meta_array_27_1 : _GEN_672; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_674 = 6'h1c == io_resp_1_1_r2 ? meta_array_28_1 : _GEN_673; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_675 = 6'h1d == io_resp_1_1_r2 ? meta_array_29_1 : _GEN_674; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_676 = 6'h1e == io_resp_1_1_r2 ? meta_array_30_1 : _GEN_675; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_677 = 6'h1f == io_resp_1_1_r2 ? meta_array_31_1 : _GEN_676; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_678 = 6'h20 == io_resp_1_1_r2 ? meta_array_32_1 : _GEN_677; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_679 = 6'h21 == io_resp_1_1_r2 ? meta_array_33_1 : _GEN_678; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_680 = 6'h22 == io_resp_1_1_r2 ? meta_array_34_1 : _GEN_679; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_681 = 6'h23 == io_resp_1_1_r2 ? meta_array_35_1 : _GEN_680; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_682 = 6'h24 == io_resp_1_1_r2 ? meta_array_36_1 : _GEN_681; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_683 = 6'h25 == io_resp_1_1_r2 ? meta_array_37_1 : _GEN_682; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_684 = 6'h26 == io_resp_1_1_r2 ? meta_array_38_1 : _GEN_683; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_685 = 6'h27 == io_resp_1_1_r2 ? meta_array_39_1 : _GEN_684; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_686 = 6'h28 == io_resp_1_1_r2 ? meta_array_40_1 : _GEN_685; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_687 = 6'h29 == io_resp_1_1_r2 ? meta_array_41_1 : _GEN_686; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_688 = 6'h2a == io_resp_1_1_r2 ? meta_array_42_1 : _GEN_687; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_689 = 6'h2b == io_resp_1_1_r2 ? meta_array_43_1 : _GEN_688; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_690 = 6'h2c == io_resp_1_1_r2 ? meta_array_44_1 : _GEN_689; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_691 = 6'h2d == io_resp_1_1_r2 ? meta_array_45_1 : _GEN_690; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_692 = 6'h2e == io_resp_1_1_r2 ? meta_array_46_1 : _GEN_691; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_693 = 6'h2f == io_resp_1_1_r2 ? meta_array_47_1 : _GEN_692; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_694 = 6'h30 == io_resp_1_1_r2 ? meta_array_48_1 : _GEN_693; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_695 = 6'h31 == io_resp_1_1_r2 ? meta_array_49_1 : _GEN_694; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_696 = 6'h32 == io_resp_1_1_r2 ? meta_array_50_1 : _GEN_695; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_697 = 6'h33 == io_resp_1_1_r2 ? meta_array_51_1 : _GEN_696; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_698 = 6'h34 == io_resp_1_1_r2 ? meta_array_52_1 : _GEN_697; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_699 = 6'h35 == io_resp_1_1_r2 ? meta_array_53_1 : _GEN_698; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_700 = 6'h36 == io_resp_1_1_r2 ? meta_array_54_1 : _GEN_699; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_701 = 6'h37 == io_resp_1_1_r2 ? meta_array_55_1 : _GEN_700; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_702 = 6'h38 == io_resp_1_1_r2 ? meta_array_56_1 : _GEN_701; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_703 = 6'h39 == io_resp_1_1_r2 ? meta_array_57_1 : _GEN_702; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_704 = 6'h3a == io_resp_1_1_r2 ? meta_array_58_1 : _GEN_703; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_705 = 6'h3b == io_resp_1_1_r2 ? meta_array_59_1 : _GEN_704; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_706 = 6'h3c == io_resp_1_1_r2 ? meta_array_60_1 : _GEN_705; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_707 = 6'h3d == io_resp_1_1_r2 ? meta_array_61_1 : _GEN_706; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_708 = 6'h3e == io_resp_1_1_r2 ? meta_array_62_1 : _GEN_707; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_709 = 6'h3f == io_resp_1_1_r2 ? meta_array_63_1 : _GEN_708; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  read_way_bypass_10 = s1_way_wen_2_1_REG & s1_way_waddr_2_1_r == io_read_1_bits_idx | s1_way_wen_2_0_REG &
    s1_way_waddr_2_0_r == io_read_1_bits_idx; // @[AsynchronousMetaArray.scala 134:85 135:29]
  reg  io_resp_1_2_r; // @[Reg.scala 16:16]
  reg  io_resp_1_2_r1; // @[Reg.scala 16:16]
  reg [5:0] io_resp_1_2_r2; // @[Reg.scala 16:16]
  wire  _GEN_718 = 6'h1 == io_resp_1_2_r2 ? meta_array_1_2 : meta_array_0_2; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_719 = 6'h2 == io_resp_1_2_r2 ? meta_array_2_2 : _GEN_718; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_720 = 6'h3 == io_resp_1_2_r2 ? meta_array_3_2 : _GEN_719; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_721 = 6'h4 == io_resp_1_2_r2 ? meta_array_4_2 : _GEN_720; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_722 = 6'h5 == io_resp_1_2_r2 ? meta_array_5_2 : _GEN_721; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_723 = 6'h6 == io_resp_1_2_r2 ? meta_array_6_2 : _GEN_722; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_724 = 6'h7 == io_resp_1_2_r2 ? meta_array_7_2 : _GEN_723; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_725 = 6'h8 == io_resp_1_2_r2 ? meta_array_8_2 : _GEN_724; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_726 = 6'h9 == io_resp_1_2_r2 ? meta_array_9_2 : _GEN_725; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_727 = 6'ha == io_resp_1_2_r2 ? meta_array_10_2 : _GEN_726; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_728 = 6'hb == io_resp_1_2_r2 ? meta_array_11_2 : _GEN_727; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_729 = 6'hc == io_resp_1_2_r2 ? meta_array_12_2 : _GEN_728; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_730 = 6'hd == io_resp_1_2_r2 ? meta_array_13_2 : _GEN_729; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_731 = 6'he == io_resp_1_2_r2 ? meta_array_14_2 : _GEN_730; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_732 = 6'hf == io_resp_1_2_r2 ? meta_array_15_2 : _GEN_731; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_733 = 6'h10 == io_resp_1_2_r2 ? meta_array_16_2 : _GEN_732; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_734 = 6'h11 == io_resp_1_2_r2 ? meta_array_17_2 : _GEN_733; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_735 = 6'h12 == io_resp_1_2_r2 ? meta_array_18_2 : _GEN_734; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_736 = 6'h13 == io_resp_1_2_r2 ? meta_array_19_2 : _GEN_735; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_737 = 6'h14 == io_resp_1_2_r2 ? meta_array_20_2 : _GEN_736; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_738 = 6'h15 == io_resp_1_2_r2 ? meta_array_21_2 : _GEN_737; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_739 = 6'h16 == io_resp_1_2_r2 ? meta_array_22_2 : _GEN_738; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_740 = 6'h17 == io_resp_1_2_r2 ? meta_array_23_2 : _GEN_739; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_741 = 6'h18 == io_resp_1_2_r2 ? meta_array_24_2 : _GEN_740; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_742 = 6'h19 == io_resp_1_2_r2 ? meta_array_25_2 : _GEN_741; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_743 = 6'h1a == io_resp_1_2_r2 ? meta_array_26_2 : _GEN_742; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_744 = 6'h1b == io_resp_1_2_r2 ? meta_array_27_2 : _GEN_743; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_745 = 6'h1c == io_resp_1_2_r2 ? meta_array_28_2 : _GEN_744; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_746 = 6'h1d == io_resp_1_2_r2 ? meta_array_29_2 : _GEN_745; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_747 = 6'h1e == io_resp_1_2_r2 ? meta_array_30_2 : _GEN_746; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_748 = 6'h1f == io_resp_1_2_r2 ? meta_array_31_2 : _GEN_747; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_749 = 6'h20 == io_resp_1_2_r2 ? meta_array_32_2 : _GEN_748; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_750 = 6'h21 == io_resp_1_2_r2 ? meta_array_33_2 : _GEN_749; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_751 = 6'h22 == io_resp_1_2_r2 ? meta_array_34_2 : _GEN_750; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_752 = 6'h23 == io_resp_1_2_r2 ? meta_array_35_2 : _GEN_751; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_753 = 6'h24 == io_resp_1_2_r2 ? meta_array_36_2 : _GEN_752; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_754 = 6'h25 == io_resp_1_2_r2 ? meta_array_37_2 : _GEN_753; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_755 = 6'h26 == io_resp_1_2_r2 ? meta_array_38_2 : _GEN_754; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_756 = 6'h27 == io_resp_1_2_r2 ? meta_array_39_2 : _GEN_755; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_757 = 6'h28 == io_resp_1_2_r2 ? meta_array_40_2 : _GEN_756; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_758 = 6'h29 == io_resp_1_2_r2 ? meta_array_41_2 : _GEN_757; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_759 = 6'h2a == io_resp_1_2_r2 ? meta_array_42_2 : _GEN_758; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_760 = 6'h2b == io_resp_1_2_r2 ? meta_array_43_2 : _GEN_759; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_761 = 6'h2c == io_resp_1_2_r2 ? meta_array_44_2 : _GEN_760; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_762 = 6'h2d == io_resp_1_2_r2 ? meta_array_45_2 : _GEN_761; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_763 = 6'h2e == io_resp_1_2_r2 ? meta_array_46_2 : _GEN_762; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_764 = 6'h2f == io_resp_1_2_r2 ? meta_array_47_2 : _GEN_763; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_765 = 6'h30 == io_resp_1_2_r2 ? meta_array_48_2 : _GEN_764; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_766 = 6'h31 == io_resp_1_2_r2 ? meta_array_49_2 : _GEN_765; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_767 = 6'h32 == io_resp_1_2_r2 ? meta_array_50_2 : _GEN_766; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_768 = 6'h33 == io_resp_1_2_r2 ? meta_array_51_2 : _GEN_767; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_769 = 6'h34 == io_resp_1_2_r2 ? meta_array_52_2 : _GEN_768; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_770 = 6'h35 == io_resp_1_2_r2 ? meta_array_53_2 : _GEN_769; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_771 = 6'h36 == io_resp_1_2_r2 ? meta_array_54_2 : _GEN_770; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_772 = 6'h37 == io_resp_1_2_r2 ? meta_array_55_2 : _GEN_771; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_773 = 6'h38 == io_resp_1_2_r2 ? meta_array_56_2 : _GEN_772; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_774 = 6'h39 == io_resp_1_2_r2 ? meta_array_57_2 : _GEN_773; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_775 = 6'h3a == io_resp_1_2_r2 ? meta_array_58_2 : _GEN_774; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_776 = 6'h3b == io_resp_1_2_r2 ? meta_array_59_2 : _GEN_775; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_777 = 6'h3c == io_resp_1_2_r2 ? meta_array_60_2 : _GEN_776; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_778 = 6'h3d == io_resp_1_2_r2 ? meta_array_61_2 : _GEN_777; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_779 = 6'h3e == io_resp_1_2_r2 ? meta_array_62_2 : _GEN_778; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_780 = 6'h3f == io_resp_1_2_r2 ? meta_array_63_2 : _GEN_779; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  read_way_bypass_11 = s1_way_wen_3_1_REG & s1_way_waddr_3_1_r == io_read_1_bits_idx | s1_way_wen_3_0_REG &
    s1_way_waddr_3_0_r == io_read_1_bits_idx; // @[AsynchronousMetaArray.scala 134:85 135:29]
  reg  io_resp_1_3_r; // @[Reg.scala 16:16]
  reg  io_resp_1_3_r1; // @[Reg.scala 16:16]
  reg [5:0] io_resp_1_3_r2; // @[Reg.scala 16:16]
  wire  _GEN_789 = 6'h1 == io_resp_1_3_r2 ? meta_array_1_3 : meta_array_0_3; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_790 = 6'h2 == io_resp_1_3_r2 ? meta_array_2_3 : _GEN_789; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_791 = 6'h3 == io_resp_1_3_r2 ? meta_array_3_3 : _GEN_790; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_792 = 6'h4 == io_resp_1_3_r2 ? meta_array_4_3 : _GEN_791; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_793 = 6'h5 == io_resp_1_3_r2 ? meta_array_5_3 : _GEN_792; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_794 = 6'h6 == io_resp_1_3_r2 ? meta_array_6_3 : _GEN_793; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_795 = 6'h7 == io_resp_1_3_r2 ? meta_array_7_3 : _GEN_794; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_796 = 6'h8 == io_resp_1_3_r2 ? meta_array_8_3 : _GEN_795; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_797 = 6'h9 == io_resp_1_3_r2 ? meta_array_9_3 : _GEN_796; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_798 = 6'ha == io_resp_1_3_r2 ? meta_array_10_3 : _GEN_797; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_799 = 6'hb == io_resp_1_3_r2 ? meta_array_11_3 : _GEN_798; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_800 = 6'hc == io_resp_1_3_r2 ? meta_array_12_3 : _GEN_799; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_801 = 6'hd == io_resp_1_3_r2 ? meta_array_13_3 : _GEN_800; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_802 = 6'he == io_resp_1_3_r2 ? meta_array_14_3 : _GEN_801; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_803 = 6'hf == io_resp_1_3_r2 ? meta_array_15_3 : _GEN_802; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_804 = 6'h10 == io_resp_1_3_r2 ? meta_array_16_3 : _GEN_803; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_805 = 6'h11 == io_resp_1_3_r2 ? meta_array_17_3 : _GEN_804; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_806 = 6'h12 == io_resp_1_3_r2 ? meta_array_18_3 : _GEN_805; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_807 = 6'h13 == io_resp_1_3_r2 ? meta_array_19_3 : _GEN_806; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_808 = 6'h14 == io_resp_1_3_r2 ? meta_array_20_3 : _GEN_807; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_809 = 6'h15 == io_resp_1_3_r2 ? meta_array_21_3 : _GEN_808; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_810 = 6'h16 == io_resp_1_3_r2 ? meta_array_22_3 : _GEN_809; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_811 = 6'h17 == io_resp_1_3_r2 ? meta_array_23_3 : _GEN_810; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_812 = 6'h18 == io_resp_1_3_r2 ? meta_array_24_3 : _GEN_811; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_813 = 6'h19 == io_resp_1_3_r2 ? meta_array_25_3 : _GEN_812; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_814 = 6'h1a == io_resp_1_3_r2 ? meta_array_26_3 : _GEN_813; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_815 = 6'h1b == io_resp_1_3_r2 ? meta_array_27_3 : _GEN_814; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_816 = 6'h1c == io_resp_1_3_r2 ? meta_array_28_3 : _GEN_815; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_817 = 6'h1d == io_resp_1_3_r2 ? meta_array_29_3 : _GEN_816; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_818 = 6'h1e == io_resp_1_3_r2 ? meta_array_30_3 : _GEN_817; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_819 = 6'h1f == io_resp_1_3_r2 ? meta_array_31_3 : _GEN_818; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_820 = 6'h20 == io_resp_1_3_r2 ? meta_array_32_3 : _GEN_819; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_821 = 6'h21 == io_resp_1_3_r2 ? meta_array_33_3 : _GEN_820; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_822 = 6'h22 == io_resp_1_3_r2 ? meta_array_34_3 : _GEN_821; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_823 = 6'h23 == io_resp_1_3_r2 ? meta_array_35_3 : _GEN_822; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_824 = 6'h24 == io_resp_1_3_r2 ? meta_array_36_3 : _GEN_823; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_825 = 6'h25 == io_resp_1_3_r2 ? meta_array_37_3 : _GEN_824; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_826 = 6'h26 == io_resp_1_3_r2 ? meta_array_38_3 : _GEN_825; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_827 = 6'h27 == io_resp_1_3_r2 ? meta_array_39_3 : _GEN_826; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_828 = 6'h28 == io_resp_1_3_r2 ? meta_array_40_3 : _GEN_827; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_829 = 6'h29 == io_resp_1_3_r2 ? meta_array_41_3 : _GEN_828; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_830 = 6'h2a == io_resp_1_3_r2 ? meta_array_42_3 : _GEN_829; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_831 = 6'h2b == io_resp_1_3_r2 ? meta_array_43_3 : _GEN_830; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_832 = 6'h2c == io_resp_1_3_r2 ? meta_array_44_3 : _GEN_831; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_833 = 6'h2d == io_resp_1_3_r2 ? meta_array_45_3 : _GEN_832; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_834 = 6'h2e == io_resp_1_3_r2 ? meta_array_46_3 : _GEN_833; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_835 = 6'h2f == io_resp_1_3_r2 ? meta_array_47_3 : _GEN_834; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_836 = 6'h30 == io_resp_1_3_r2 ? meta_array_48_3 : _GEN_835; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_837 = 6'h31 == io_resp_1_3_r2 ? meta_array_49_3 : _GEN_836; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_838 = 6'h32 == io_resp_1_3_r2 ? meta_array_50_3 : _GEN_837; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_839 = 6'h33 == io_resp_1_3_r2 ? meta_array_51_3 : _GEN_838; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_840 = 6'h34 == io_resp_1_3_r2 ? meta_array_52_3 : _GEN_839; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_841 = 6'h35 == io_resp_1_3_r2 ? meta_array_53_3 : _GEN_840; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_842 = 6'h36 == io_resp_1_3_r2 ? meta_array_54_3 : _GEN_841; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_843 = 6'h37 == io_resp_1_3_r2 ? meta_array_55_3 : _GEN_842; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_844 = 6'h38 == io_resp_1_3_r2 ? meta_array_56_3 : _GEN_843; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_845 = 6'h39 == io_resp_1_3_r2 ? meta_array_57_3 : _GEN_844; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_846 = 6'h3a == io_resp_1_3_r2 ? meta_array_58_3 : _GEN_845; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_847 = 6'h3b == io_resp_1_3_r2 ? meta_array_59_3 : _GEN_846; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_848 = 6'h3c == io_resp_1_3_r2 ? meta_array_60_3 : _GEN_847; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_849 = 6'h3d == io_resp_1_3_r2 ? meta_array_61_3 : _GEN_848; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_850 = 6'h3e == io_resp_1_3_r2 ? meta_array_62_3 : _GEN_849; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_851 = 6'h3f == io_resp_1_3_r2 ? meta_array_63_3 : _GEN_850; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  read_way_bypass_12 = s1_way_wen_4_1_REG & s1_way_waddr_4_1_r == io_read_1_bits_idx | s1_way_wen_4_0_REG &
    s1_way_waddr_4_0_r == io_read_1_bits_idx; // @[AsynchronousMetaArray.scala 134:85 135:29]
  reg  io_resp_1_4_r; // @[Reg.scala 16:16]
  reg  io_resp_1_4_r1; // @[Reg.scala 16:16]
  reg [5:0] io_resp_1_4_r2; // @[Reg.scala 16:16]
  wire  _GEN_860 = 6'h1 == io_resp_1_4_r2 ? meta_array_1_4 : meta_array_0_4; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_861 = 6'h2 == io_resp_1_4_r2 ? meta_array_2_4 : _GEN_860; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_862 = 6'h3 == io_resp_1_4_r2 ? meta_array_3_4 : _GEN_861; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_863 = 6'h4 == io_resp_1_4_r2 ? meta_array_4_4 : _GEN_862; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_864 = 6'h5 == io_resp_1_4_r2 ? meta_array_5_4 : _GEN_863; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_865 = 6'h6 == io_resp_1_4_r2 ? meta_array_6_4 : _GEN_864; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_866 = 6'h7 == io_resp_1_4_r2 ? meta_array_7_4 : _GEN_865; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_867 = 6'h8 == io_resp_1_4_r2 ? meta_array_8_4 : _GEN_866; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_868 = 6'h9 == io_resp_1_4_r2 ? meta_array_9_4 : _GEN_867; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_869 = 6'ha == io_resp_1_4_r2 ? meta_array_10_4 : _GEN_868; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_870 = 6'hb == io_resp_1_4_r2 ? meta_array_11_4 : _GEN_869; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_871 = 6'hc == io_resp_1_4_r2 ? meta_array_12_4 : _GEN_870; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_872 = 6'hd == io_resp_1_4_r2 ? meta_array_13_4 : _GEN_871; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_873 = 6'he == io_resp_1_4_r2 ? meta_array_14_4 : _GEN_872; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_874 = 6'hf == io_resp_1_4_r2 ? meta_array_15_4 : _GEN_873; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_875 = 6'h10 == io_resp_1_4_r2 ? meta_array_16_4 : _GEN_874; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_876 = 6'h11 == io_resp_1_4_r2 ? meta_array_17_4 : _GEN_875; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_877 = 6'h12 == io_resp_1_4_r2 ? meta_array_18_4 : _GEN_876; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_878 = 6'h13 == io_resp_1_4_r2 ? meta_array_19_4 : _GEN_877; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_879 = 6'h14 == io_resp_1_4_r2 ? meta_array_20_4 : _GEN_878; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_880 = 6'h15 == io_resp_1_4_r2 ? meta_array_21_4 : _GEN_879; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_881 = 6'h16 == io_resp_1_4_r2 ? meta_array_22_4 : _GEN_880; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_882 = 6'h17 == io_resp_1_4_r2 ? meta_array_23_4 : _GEN_881; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_883 = 6'h18 == io_resp_1_4_r2 ? meta_array_24_4 : _GEN_882; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_884 = 6'h19 == io_resp_1_4_r2 ? meta_array_25_4 : _GEN_883; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_885 = 6'h1a == io_resp_1_4_r2 ? meta_array_26_4 : _GEN_884; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_886 = 6'h1b == io_resp_1_4_r2 ? meta_array_27_4 : _GEN_885; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_887 = 6'h1c == io_resp_1_4_r2 ? meta_array_28_4 : _GEN_886; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_888 = 6'h1d == io_resp_1_4_r2 ? meta_array_29_4 : _GEN_887; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_889 = 6'h1e == io_resp_1_4_r2 ? meta_array_30_4 : _GEN_888; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_890 = 6'h1f == io_resp_1_4_r2 ? meta_array_31_4 : _GEN_889; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_891 = 6'h20 == io_resp_1_4_r2 ? meta_array_32_4 : _GEN_890; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_892 = 6'h21 == io_resp_1_4_r2 ? meta_array_33_4 : _GEN_891; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_893 = 6'h22 == io_resp_1_4_r2 ? meta_array_34_4 : _GEN_892; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_894 = 6'h23 == io_resp_1_4_r2 ? meta_array_35_4 : _GEN_893; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_895 = 6'h24 == io_resp_1_4_r2 ? meta_array_36_4 : _GEN_894; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_896 = 6'h25 == io_resp_1_4_r2 ? meta_array_37_4 : _GEN_895; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_897 = 6'h26 == io_resp_1_4_r2 ? meta_array_38_4 : _GEN_896; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_898 = 6'h27 == io_resp_1_4_r2 ? meta_array_39_4 : _GEN_897; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_899 = 6'h28 == io_resp_1_4_r2 ? meta_array_40_4 : _GEN_898; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_900 = 6'h29 == io_resp_1_4_r2 ? meta_array_41_4 : _GEN_899; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_901 = 6'h2a == io_resp_1_4_r2 ? meta_array_42_4 : _GEN_900; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_902 = 6'h2b == io_resp_1_4_r2 ? meta_array_43_4 : _GEN_901; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_903 = 6'h2c == io_resp_1_4_r2 ? meta_array_44_4 : _GEN_902; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_904 = 6'h2d == io_resp_1_4_r2 ? meta_array_45_4 : _GEN_903; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_905 = 6'h2e == io_resp_1_4_r2 ? meta_array_46_4 : _GEN_904; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_906 = 6'h2f == io_resp_1_4_r2 ? meta_array_47_4 : _GEN_905; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_907 = 6'h30 == io_resp_1_4_r2 ? meta_array_48_4 : _GEN_906; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_908 = 6'h31 == io_resp_1_4_r2 ? meta_array_49_4 : _GEN_907; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_909 = 6'h32 == io_resp_1_4_r2 ? meta_array_50_4 : _GEN_908; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_910 = 6'h33 == io_resp_1_4_r2 ? meta_array_51_4 : _GEN_909; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_911 = 6'h34 == io_resp_1_4_r2 ? meta_array_52_4 : _GEN_910; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_912 = 6'h35 == io_resp_1_4_r2 ? meta_array_53_4 : _GEN_911; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_913 = 6'h36 == io_resp_1_4_r2 ? meta_array_54_4 : _GEN_912; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_914 = 6'h37 == io_resp_1_4_r2 ? meta_array_55_4 : _GEN_913; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_915 = 6'h38 == io_resp_1_4_r2 ? meta_array_56_4 : _GEN_914; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_916 = 6'h39 == io_resp_1_4_r2 ? meta_array_57_4 : _GEN_915; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_917 = 6'h3a == io_resp_1_4_r2 ? meta_array_58_4 : _GEN_916; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_918 = 6'h3b == io_resp_1_4_r2 ? meta_array_59_4 : _GEN_917; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_919 = 6'h3c == io_resp_1_4_r2 ? meta_array_60_4 : _GEN_918; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_920 = 6'h3d == io_resp_1_4_r2 ? meta_array_61_4 : _GEN_919; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_921 = 6'h3e == io_resp_1_4_r2 ? meta_array_62_4 : _GEN_920; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_922 = 6'h3f == io_resp_1_4_r2 ? meta_array_63_4 : _GEN_921; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  read_way_bypass_13 = s1_way_wen_5_1_REG & s1_way_waddr_5_1_r == io_read_1_bits_idx | s1_way_wen_5_0_REG &
    s1_way_waddr_5_0_r == io_read_1_bits_idx; // @[AsynchronousMetaArray.scala 134:85 135:29]
  reg  io_resp_1_5_r; // @[Reg.scala 16:16]
  reg  io_resp_1_5_r1; // @[Reg.scala 16:16]
  reg [5:0] io_resp_1_5_r2; // @[Reg.scala 16:16]
  wire  _GEN_931 = 6'h1 == io_resp_1_5_r2 ? meta_array_1_5 : meta_array_0_5; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_932 = 6'h2 == io_resp_1_5_r2 ? meta_array_2_5 : _GEN_931; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_933 = 6'h3 == io_resp_1_5_r2 ? meta_array_3_5 : _GEN_932; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_934 = 6'h4 == io_resp_1_5_r2 ? meta_array_4_5 : _GEN_933; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_935 = 6'h5 == io_resp_1_5_r2 ? meta_array_5_5 : _GEN_934; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_936 = 6'h6 == io_resp_1_5_r2 ? meta_array_6_5 : _GEN_935; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_937 = 6'h7 == io_resp_1_5_r2 ? meta_array_7_5 : _GEN_936; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_938 = 6'h8 == io_resp_1_5_r2 ? meta_array_8_5 : _GEN_937; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_939 = 6'h9 == io_resp_1_5_r2 ? meta_array_9_5 : _GEN_938; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_940 = 6'ha == io_resp_1_5_r2 ? meta_array_10_5 : _GEN_939; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_941 = 6'hb == io_resp_1_5_r2 ? meta_array_11_5 : _GEN_940; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_942 = 6'hc == io_resp_1_5_r2 ? meta_array_12_5 : _GEN_941; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_943 = 6'hd == io_resp_1_5_r2 ? meta_array_13_5 : _GEN_942; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_944 = 6'he == io_resp_1_5_r2 ? meta_array_14_5 : _GEN_943; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_945 = 6'hf == io_resp_1_5_r2 ? meta_array_15_5 : _GEN_944; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_946 = 6'h10 == io_resp_1_5_r2 ? meta_array_16_5 : _GEN_945; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_947 = 6'h11 == io_resp_1_5_r2 ? meta_array_17_5 : _GEN_946; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_948 = 6'h12 == io_resp_1_5_r2 ? meta_array_18_5 : _GEN_947; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_949 = 6'h13 == io_resp_1_5_r2 ? meta_array_19_5 : _GEN_948; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_950 = 6'h14 == io_resp_1_5_r2 ? meta_array_20_5 : _GEN_949; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_951 = 6'h15 == io_resp_1_5_r2 ? meta_array_21_5 : _GEN_950; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_952 = 6'h16 == io_resp_1_5_r2 ? meta_array_22_5 : _GEN_951; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_953 = 6'h17 == io_resp_1_5_r2 ? meta_array_23_5 : _GEN_952; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_954 = 6'h18 == io_resp_1_5_r2 ? meta_array_24_5 : _GEN_953; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_955 = 6'h19 == io_resp_1_5_r2 ? meta_array_25_5 : _GEN_954; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_956 = 6'h1a == io_resp_1_5_r2 ? meta_array_26_5 : _GEN_955; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_957 = 6'h1b == io_resp_1_5_r2 ? meta_array_27_5 : _GEN_956; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_958 = 6'h1c == io_resp_1_5_r2 ? meta_array_28_5 : _GEN_957; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_959 = 6'h1d == io_resp_1_5_r2 ? meta_array_29_5 : _GEN_958; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_960 = 6'h1e == io_resp_1_5_r2 ? meta_array_30_5 : _GEN_959; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_961 = 6'h1f == io_resp_1_5_r2 ? meta_array_31_5 : _GEN_960; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_962 = 6'h20 == io_resp_1_5_r2 ? meta_array_32_5 : _GEN_961; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_963 = 6'h21 == io_resp_1_5_r2 ? meta_array_33_5 : _GEN_962; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_964 = 6'h22 == io_resp_1_5_r2 ? meta_array_34_5 : _GEN_963; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_965 = 6'h23 == io_resp_1_5_r2 ? meta_array_35_5 : _GEN_964; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_966 = 6'h24 == io_resp_1_5_r2 ? meta_array_36_5 : _GEN_965; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_967 = 6'h25 == io_resp_1_5_r2 ? meta_array_37_5 : _GEN_966; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_968 = 6'h26 == io_resp_1_5_r2 ? meta_array_38_5 : _GEN_967; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_969 = 6'h27 == io_resp_1_5_r2 ? meta_array_39_5 : _GEN_968; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_970 = 6'h28 == io_resp_1_5_r2 ? meta_array_40_5 : _GEN_969; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_971 = 6'h29 == io_resp_1_5_r2 ? meta_array_41_5 : _GEN_970; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_972 = 6'h2a == io_resp_1_5_r2 ? meta_array_42_5 : _GEN_971; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_973 = 6'h2b == io_resp_1_5_r2 ? meta_array_43_5 : _GEN_972; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_974 = 6'h2c == io_resp_1_5_r2 ? meta_array_44_5 : _GEN_973; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_975 = 6'h2d == io_resp_1_5_r2 ? meta_array_45_5 : _GEN_974; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_976 = 6'h2e == io_resp_1_5_r2 ? meta_array_46_5 : _GEN_975; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_977 = 6'h2f == io_resp_1_5_r2 ? meta_array_47_5 : _GEN_976; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_978 = 6'h30 == io_resp_1_5_r2 ? meta_array_48_5 : _GEN_977; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_979 = 6'h31 == io_resp_1_5_r2 ? meta_array_49_5 : _GEN_978; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_980 = 6'h32 == io_resp_1_5_r2 ? meta_array_50_5 : _GEN_979; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_981 = 6'h33 == io_resp_1_5_r2 ? meta_array_51_5 : _GEN_980; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_982 = 6'h34 == io_resp_1_5_r2 ? meta_array_52_5 : _GEN_981; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_983 = 6'h35 == io_resp_1_5_r2 ? meta_array_53_5 : _GEN_982; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_984 = 6'h36 == io_resp_1_5_r2 ? meta_array_54_5 : _GEN_983; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_985 = 6'h37 == io_resp_1_5_r2 ? meta_array_55_5 : _GEN_984; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_986 = 6'h38 == io_resp_1_5_r2 ? meta_array_56_5 : _GEN_985; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_987 = 6'h39 == io_resp_1_5_r2 ? meta_array_57_5 : _GEN_986; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_988 = 6'h3a == io_resp_1_5_r2 ? meta_array_58_5 : _GEN_987; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_989 = 6'h3b == io_resp_1_5_r2 ? meta_array_59_5 : _GEN_988; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_990 = 6'h3c == io_resp_1_5_r2 ? meta_array_60_5 : _GEN_989; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_991 = 6'h3d == io_resp_1_5_r2 ? meta_array_61_5 : _GEN_990; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_992 = 6'h3e == io_resp_1_5_r2 ? meta_array_62_5 : _GEN_991; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_993 = 6'h3f == io_resp_1_5_r2 ? meta_array_63_5 : _GEN_992; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  read_way_bypass_14 = s1_way_wen_6_1_REG & s1_way_waddr_6_1_r == io_read_1_bits_idx | s1_way_wen_6_0_REG &
    s1_way_waddr_6_0_r == io_read_1_bits_idx; // @[AsynchronousMetaArray.scala 134:85 135:29]
  reg  io_resp_1_6_r; // @[Reg.scala 16:16]
  reg  io_resp_1_6_r1; // @[Reg.scala 16:16]
  reg [5:0] io_resp_1_6_r2; // @[Reg.scala 16:16]
  wire  _GEN_1002 = 6'h1 == io_resp_1_6_r2 ? meta_array_1_6 : meta_array_0_6; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1003 = 6'h2 == io_resp_1_6_r2 ? meta_array_2_6 : _GEN_1002; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1004 = 6'h3 == io_resp_1_6_r2 ? meta_array_3_6 : _GEN_1003; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1005 = 6'h4 == io_resp_1_6_r2 ? meta_array_4_6 : _GEN_1004; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1006 = 6'h5 == io_resp_1_6_r2 ? meta_array_5_6 : _GEN_1005; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1007 = 6'h6 == io_resp_1_6_r2 ? meta_array_6_6 : _GEN_1006; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1008 = 6'h7 == io_resp_1_6_r2 ? meta_array_7_6 : _GEN_1007; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1009 = 6'h8 == io_resp_1_6_r2 ? meta_array_8_6 : _GEN_1008; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1010 = 6'h9 == io_resp_1_6_r2 ? meta_array_9_6 : _GEN_1009; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1011 = 6'ha == io_resp_1_6_r2 ? meta_array_10_6 : _GEN_1010; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1012 = 6'hb == io_resp_1_6_r2 ? meta_array_11_6 : _GEN_1011; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1013 = 6'hc == io_resp_1_6_r2 ? meta_array_12_6 : _GEN_1012; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1014 = 6'hd == io_resp_1_6_r2 ? meta_array_13_6 : _GEN_1013; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1015 = 6'he == io_resp_1_6_r2 ? meta_array_14_6 : _GEN_1014; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1016 = 6'hf == io_resp_1_6_r2 ? meta_array_15_6 : _GEN_1015; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1017 = 6'h10 == io_resp_1_6_r2 ? meta_array_16_6 : _GEN_1016; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1018 = 6'h11 == io_resp_1_6_r2 ? meta_array_17_6 : _GEN_1017; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1019 = 6'h12 == io_resp_1_6_r2 ? meta_array_18_6 : _GEN_1018; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1020 = 6'h13 == io_resp_1_6_r2 ? meta_array_19_6 : _GEN_1019; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1021 = 6'h14 == io_resp_1_6_r2 ? meta_array_20_6 : _GEN_1020; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1022 = 6'h15 == io_resp_1_6_r2 ? meta_array_21_6 : _GEN_1021; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1023 = 6'h16 == io_resp_1_6_r2 ? meta_array_22_6 : _GEN_1022; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1024 = 6'h17 == io_resp_1_6_r2 ? meta_array_23_6 : _GEN_1023; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1025 = 6'h18 == io_resp_1_6_r2 ? meta_array_24_6 : _GEN_1024; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1026 = 6'h19 == io_resp_1_6_r2 ? meta_array_25_6 : _GEN_1025; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1027 = 6'h1a == io_resp_1_6_r2 ? meta_array_26_6 : _GEN_1026; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1028 = 6'h1b == io_resp_1_6_r2 ? meta_array_27_6 : _GEN_1027; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1029 = 6'h1c == io_resp_1_6_r2 ? meta_array_28_6 : _GEN_1028; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1030 = 6'h1d == io_resp_1_6_r2 ? meta_array_29_6 : _GEN_1029; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1031 = 6'h1e == io_resp_1_6_r2 ? meta_array_30_6 : _GEN_1030; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1032 = 6'h1f == io_resp_1_6_r2 ? meta_array_31_6 : _GEN_1031; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1033 = 6'h20 == io_resp_1_6_r2 ? meta_array_32_6 : _GEN_1032; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1034 = 6'h21 == io_resp_1_6_r2 ? meta_array_33_6 : _GEN_1033; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1035 = 6'h22 == io_resp_1_6_r2 ? meta_array_34_6 : _GEN_1034; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1036 = 6'h23 == io_resp_1_6_r2 ? meta_array_35_6 : _GEN_1035; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1037 = 6'h24 == io_resp_1_6_r2 ? meta_array_36_6 : _GEN_1036; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1038 = 6'h25 == io_resp_1_6_r2 ? meta_array_37_6 : _GEN_1037; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1039 = 6'h26 == io_resp_1_6_r2 ? meta_array_38_6 : _GEN_1038; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1040 = 6'h27 == io_resp_1_6_r2 ? meta_array_39_6 : _GEN_1039; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1041 = 6'h28 == io_resp_1_6_r2 ? meta_array_40_6 : _GEN_1040; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1042 = 6'h29 == io_resp_1_6_r2 ? meta_array_41_6 : _GEN_1041; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1043 = 6'h2a == io_resp_1_6_r2 ? meta_array_42_6 : _GEN_1042; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1044 = 6'h2b == io_resp_1_6_r2 ? meta_array_43_6 : _GEN_1043; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1045 = 6'h2c == io_resp_1_6_r2 ? meta_array_44_6 : _GEN_1044; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1046 = 6'h2d == io_resp_1_6_r2 ? meta_array_45_6 : _GEN_1045; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1047 = 6'h2e == io_resp_1_6_r2 ? meta_array_46_6 : _GEN_1046; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1048 = 6'h2f == io_resp_1_6_r2 ? meta_array_47_6 : _GEN_1047; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1049 = 6'h30 == io_resp_1_6_r2 ? meta_array_48_6 : _GEN_1048; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1050 = 6'h31 == io_resp_1_6_r2 ? meta_array_49_6 : _GEN_1049; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1051 = 6'h32 == io_resp_1_6_r2 ? meta_array_50_6 : _GEN_1050; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1052 = 6'h33 == io_resp_1_6_r2 ? meta_array_51_6 : _GEN_1051; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1053 = 6'h34 == io_resp_1_6_r2 ? meta_array_52_6 : _GEN_1052; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1054 = 6'h35 == io_resp_1_6_r2 ? meta_array_53_6 : _GEN_1053; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1055 = 6'h36 == io_resp_1_6_r2 ? meta_array_54_6 : _GEN_1054; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1056 = 6'h37 == io_resp_1_6_r2 ? meta_array_55_6 : _GEN_1055; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1057 = 6'h38 == io_resp_1_6_r2 ? meta_array_56_6 : _GEN_1056; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1058 = 6'h39 == io_resp_1_6_r2 ? meta_array_57_6 : _GEN_1057; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1059 = 6'h3a == io_resp_1_6_r2 ? meta_array_58_6 : _GEN_1058; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1060 = 6'h3b == io_resp_1_6_r2 ? meta_array_59_6 : _GEN_1059; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1061 = 6'h3c == io_resp_1_6_r2 ? meta_array_60_6 : _GEN_1060; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1062 = 6'h3d == io_resp_1_6_r2 ? meta_array_61_6 : _GEN_1061; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1063 = 6'h3e == io_resp_1_6_r2 ? meta_array_62_6 : _GEN_1062; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1064 = 6'h3f == io_resp_1_6_r2 ? meta_array_63_6 : _GEN_1063; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  read_way_bypass_15 = s1_way_wen_7_1_REG & s1_way_waddr_7_1_r == io_read_1_bits_idx | s1_way_wen_7_0_REG &
    s1_way_waddr_7_0_r == io_read_1_bits_idx; // @[AsynchronousMetaArray.scala 134:85 135:29]
  reg  io_resp_1_7_r; // @[Reg.scala 16:16]
  reg  io_resp_1_7_r1; // @[Reg.scala 16:16]
  reg [5:0] io_resp_1_7_r2; // @[Reg.scala 16:16]
  wire  _GEN_1073 = 6'h1 == io_resp_1_7_r2 ? meta_array_1_7 : meta_array_0_7; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1074 = 6'h2 == io_resp_1_7_r2 ? meta_array_2_7 : _GEN_1073; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1075 = 6'h3 == io_resp_1_7_r2 ? meta_array_3_7 : _GEN_1074; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1076 = 6'h4 == io_resp_1_7_r2 ? meta_array_4_7 : _GEN_1075; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1077 = 6'h5 == io_resp_1_7_r2 ? meta_array_5_7 : _GEN_1076; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1078 = 6'h6 == io_resp_1_7_r2 ? meta_array_6_7 : _GEN_1077; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1079 = 6'h7 == io_resp_1_7_r2 ? meta_array_7_7 : _GEN_1078; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1080 = 6'h8 == io_resp_1_7_r2 ? meta_array_8_7 : _GEN_1079; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1081 = 6'h9 == io_resp_1_7_r2 ? meta_array_9_7 : _GEN_1080; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1082 = 6'ha == io_resp_1_7_r2 ? meta_array_10_7 : _GEN_1081; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1083 = 6'hb == io_resp_1_7_r2 ? meta_array_11_7 : _GEN_1082; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1084 = 6'hc == io_resp_1_7_r2 ? meta_array_12_7 : _GEN_1083; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1085 = 6'hd == io_resp_1_7_r2 ? meta_array_13_7 : _GEN_1084; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1086 = 6'he == io_resp_1_7_r2 ? meta_array_14_7 : _GEN_1085; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1087 = 6'hf == io_resp_1_7_r2 ? meta_array_15_7 : _GEN_1086; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1088 = 6'h10 == io_resp_1_7_r2 ? meta_array_16_7 : _GEN_1087; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1089 = 6'h11 == io_resp_1_7_r2 ? meta_array_17_7 : _GEN_1088; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1090 = 6'h12 == io_resp_1_7_r2 ? meta_array_18_7 : _GEN_1089; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1091 = 6'h13 == io_resp_1_7_r2 ? meta_array_19_7 : _GEN_1090; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1092 = 6'h14 == io_resp_1_7_r2 ? meta_array_20_7 : _GEN_1091; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1093 = 6'h15 == io_resp_1_7_r2 ? meta_array_21_7 : _GEN_1092; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1094 = 6'h16 == io_resp_1_7_r2 ? meta_array_22_7 : _GEN_1093; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1095 = 6'h17 == io_resp_1_7_r2 ? meta_array_23_7 : _GEN_1094; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1096 = 6'h18 == io_resp_1_7_r2 ? meta_array_24_7 : _GEN_1095; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1097 = 6'h19 == io_resp_1_7_r2 ? meta_array_25_7 : _GEN_1096; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1098 = 6'h1a == io_resp_1_7_r2 ? meta_array_26_7 : _GEN_1097; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1099 = 6'h1b == io_resp_1_7_r2 ? meta_array_27_7 : _GEN_1098; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1100 = 6'h1c == io_resp_1_7_r2 ? meta_array_28_7 : _GEN_1099; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1101 = 6'h1d == io_resp_1_7_r2 ? meta_array_29_7 : _GEN_1100; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1102 = 6'h1e == io_resp_1_7_r2 ? meta_array_30_7 : _GEN_1101; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1103 = 6'h1f == io_resp_1_7_r2 ? meta_array_31_7 : _GEN_1102; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1104 = 6'h20 == io_resp_1_7_r2 ? meta_array_32_7 : _GEN_1103; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1105 = 6'h21 == io_resp_1_7_r2 ? meta_array_33_7 : _GEN_1104; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1106 = 6'h22 == io_resp_1_7_r2 ? meta_array_34_7 : _GEN_1105; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1107 = 6'h23 == io_resp_1_7_r2 ? meta_array_35_7 : _GEN_1106; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1108 = 6'h24 == io_resp_1_7_r2 ? meta_array_36_7 : _GEN_1107; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1109 = 6'h25 == io_resp_1_7_r2 ? meta_array_37_7 : _GEN_1108; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1110 = 6'h26 == io_resp_1_7_r2 ? meta_array_38_7 : _GEN_1109; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1111 = 6'h27 == io_resp_1_7_r2 ? meta_array_39_7 : _GEN_1110; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1112 = 6'h28 == io_resp_1_7_r2 ? meta_array_40_7 : _GEN_1111; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1113 = 6'h29 == io_resp_1_7_r2 ? meta_array_41_7 : _GEN_1112; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1114 = 6'h2a == io_resp_1_7_r2 ? meta_array_42_7 : _GEN_1113; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1115 = 6'h2b == io_resp_1_7_r2 ? meta_array_43_7 : _GEN_1114; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1116 = 6'h2c == io_resp_1_7_r2 ? meta_array_44_7 : _GEN_1115; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1117 = 6'h2d == io_resp_1_7_r2 ? meta_array_45_7 : _GEN_1116; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1118 = 6'h2e == io_resp_1_7_r2 ? meta_array_46_7 : _GEN_1117; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1119 = 6'h2f == io_resp_1_7_r2 ? meta_array_47_7 : _GEN_1118; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1120 = 6'h30 == io_resp_1_7_r2 ? meta_array_48_7 : _GEN_1119; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1121 = 6'h31 == io_resp_1_7_r2 ? meta_array_49_7 : _GEN_1120; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1122 = 6'h32 == io_resp_1_7_r2 ? meta_array_50_7 : _GEN_1121; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1123 = 6'h33 == io_resp_1_7_r2 ? meta_array_51_7 : _GEN_1122; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1124 = 6'h34 == io_resp_1_7_r2 ? meta_array_52_7 : _GEN_1123; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1125 = 6'h35 == io_resp_1_7_r2 ? meta_array_53_7 : _GEN_1124; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1126 = 6'h36 == io_resp_1_7_r2 ? meta_array_54_7 : _GEN_1125; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1127 = 6'h37 == io_resp_1_7_r2 ? meta_array_55_7 : _GEN_1126; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1128 = 6'h38 == io_resp_1_7_r2 ? meta_array_56_7 : _GEN_1127; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1129 = 6'h39 == io_resp_1_7_r2 ? meta_array_57_7 : _GEN_1128; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1130 = 6'h3a == io_resp_1_7_r2 ? meta_array_58_7 : _GEN_1129; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1131 = 6'h3b == io_resp_1_7_r2 ? meta_array_59_7 : _GEN_1130; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1132 = 6'h3c == io_resp_1_7_r2 ? meta_array_60_7 : _GEN_1131; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1133 = 6'h3d == io_resp_1_7_r2 ? meta_array_61_7 : _GEN_1132; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1134 = 6'h3e == io_resp_1_7_r2 ? meta_array_62_7 : _GEN_1133; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1135 = 6'h3f == io_resp_1_7_r2 ? meta_array_63_7 : _GEN_1134; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  read_way_bypass_16 = s1_way_wen_0_1_REG & s1_way_waddr_0_1_r == io_read_2_bits_idx | s1_way_wen_0_0_REG &
    s1_way_waddr_0_0_r == io_read_2_bits_idx; // @[AsynchronousMetaArray.scala 134:85 135:29]
  reg  io_resp_2_0_r; // @[Reg.scala 16:16]
  reg  io_resp_2_0_r1; // @[Reg.scala 16:16]
  reg [5:0] io_resp_2_0_r2; // @[Reg.scala 16:16]
  wire  _GEN_1144 = 6'h1 == io_resp_2_0_r2 ? meta_array_1_0 : meta_array_0_0; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1145 = 6'h2 == io_resp_2_0_r2 ? meta_array_2_0 : _GEN_1144; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1146 = 6'h3 == io_resp_2_0_r2 ? meta_array_3_0 : _GEN_1145; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1147 = 6'h4 == io_resp_2_0_r2 ? meta_array_4_0 : _GEN_1146; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1148 = 6'h5 == io_resp_2_0_r2 ? meta_array_5_0 : _GEN_1147; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1149 = 6'h6 == io_resp_2_0_r2 ? meta_array_6_0 : _GEN_1148; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1150 = 6'h7 == io_resp_2_0_r2 ? meta_array_7_0 : _GEN_1149; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1151 = 6'h8 == io_resp_2_0_r2 ? meta_array_8_0 : _GEN_1150; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1152 = 6'h9 == io_resp_2_0_r2 ? meta_array_9_0 : _GEN_1151; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1153 = 6'ha == io_resp_2_0_r2 ? meta_array_10_0 : _GEN_1152; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1154 = 6'hb == io_resp_2_0_r2 ? meta_array_11_0 : _GEN_1153; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1155 = 6'hc == io_resp_2_0_r2 ? meta_array_12_0 : _GEN_1154; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1156 = 6'hd == io_resp_2_0_r2 ? meta_array_13_0 : _GEN_1155; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1157 = 6'he == io_resp_2_0_r2 ? meta_array_14_0 : _GEN_1156; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1158 = 6'hf == io_resp_2_0_r2 ? meta_array_15_0 : _GEN_1157; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1159 = 6'h10 == io_resp_2_0_r2 ? meta_array_16_0 : _GEN_1158; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1160 = 6'h11 == io_resp_2_0_r2 ? meta_array_17_0 : _GEN_1159; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1161 = 6'h12 == io_resp_2_0_r2 ? meta_array_18_0 : _GEN_1160; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1162 = 6'h13 == io_resp_2_0_r2 ? meta_array_19_0 : _GEN_1161; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1163 = 6'h14 == io_resp_2_0_r2 ? meta_array_20_0 : _GEN_1162; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1164 = 6'h15 == io_resp_2_0_r2 ? meta_array_21_0 : _GEN_1163; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1165 = 6'h16 == io_resp_2_0_r2 ? meta_array_22_0 : _GEN_1164; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1166 = 6'h17 == io_resp_2_0_r2 ? meta_array_23_0 : _GEN_1165; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1167 = 6'h18 == io_resp_2_0_r2 ? meta_array_24_0 : _GEN_1166; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1168 = 6'h19 == io_resp_2_0_r2 ? meta_array_25_0 : _GEN_1167; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1169 = 6'h1a == io_resp_2_0_r2 ? meta_array_26_0 : _GEN_1168; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1170 = 6'h1b == io_resp_2_0_r2 ? meta_array_27_0 : _GEN_1169; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1171 = 6'h1c == io_resp_2_0_r2 ? meta_array_28_0 : _GEN_1170; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1172 = 6'h1d == io_resp_2_0_r2 ? meta_array_29_0 : _GEN_1171; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1173 = 6'h1e == io_resp_2_0_r2 ? meta_array_30_0 : _GEN_1172; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1174 = 6'h1f == io_resp_2_0_r2 ? meta_array_31_0 : _GEN_1173; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1175 = 6'h20 == io_resp_2_0_r2 ? meta_array_32_0 : _GEN_1174; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1176 = 6'h21 == io_resp_2_0_r2 ? meta_array_33_0 : _GEN_1175; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1177 = 6'h22 == io_resp_2_0_r2 ? meta_array_34_0 : _GEN_1176; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1178 = 6'h23 == io_resp_2_0_r2 ? meta_array_35_0 : _GEN_1177; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1179 = 6'h24 == io_resp_2_0_r2 ? meta_array_36_0 : _GEN_1178; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1180 = 6'h25 == io_resp_2_0_r2 ? meta_array_37_0 : _GEN_1179; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1181 = 6'h26 == io_resp_2_0_r2 ? meta_array_38_0 : _GEN_1180; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1182 = 6'h27 == io_resp_2_0_r2 ? meta_array_39_0 : _GEN_1181; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1183 = 6'h28 == io_resp_2_0_r2 ? meta_array_40_0 : _GEN_1182; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1184 = 6'h29 == io_resp_2_0_r2 ? meta_array_41_0 : _GEN_1183; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1185 = 6'h2a == io_resp_2_0_r2 ? meta_array_42_0 : _GEN_1184; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1186 = 6'h2b == io_resp_2_0_r2 ? meta_array_43_0 : _GEN_1185; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1187 = 6'h2c == io_resp_2_0_r2 ? meta_array_44_0 : _GEN_1186; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1188 = 6'h2d == io_resp_2_0_r2 ? meta_array_45_0 : _GEN_1187; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1189 = 6'h2e == io_resp_2_0_r2 ? meta_array_46_0 : _GEN_1188; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1190 = 6'h2f == io_resp_2_0_r2 ? meta_array_47_0 : _GEN_1189; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1191 = 6'h30 == io_resp_2_0_r2 ? meta_array_48_0 : _GEN_1190; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1192 = 6'h31 == io_resp_2_0_r2 ? meta_array_49_0 : _GEN_1191; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1193 = 6'h32 == io_resp_2_0_r2 ? meta_array_50_0 : _GEN_1192; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1194 = 6'h33 == io_resp_2_0_r2 ? meta_array_51_0 : _GEN_1193; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1195 = 6'h34 == io_resp_2_0_r2 ? meta_array_52_0 : _GEN_1194; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1196 = 6'h35 == io_resp_2_0_r2 ? meta_array_53_0 : _GEN_1195; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1197 = 6'h36 == io_resp_2_0_r2 ? meta_array_54_0 : _GEN_1196; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1198 = 6'h37 == io_resp_2_0_r2 ? meta_array_55_0 : _GEN_1197; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1199 = 6'h38 == io_resp_2_0_r2 ? meta_array_56_0 : _GEN_1198; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1200 = 6'h39 == io_resp_2_0_r2 ? meta_array_57_0 : _GEN_1199; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1201 = 6'h3a == io_resp_2_0_r2 ? meta_array_58_0 : _GEN_1200; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1202 = 6'h3b == io_resp_2_0_r2 ? meta_array_59_0 : _GEN_1201; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1203 = 6'h3c == io_resp_2_0_r2 ? meta_array_60_0 : _GEN_1202; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1204 = 6'h3d == io_resp_2_0_r2 ? meta_array_61_0 : _GEN_1203; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1205 = 6'h3e == io_resp_2_0_r2 ? meta_array_62_0 : _GEN_1204; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1206 = 6'h3f == io_resp_2_0_r2 ? meta_array_63_0 : _GEN_1205; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  read_way_bypass_17 = s1_way_wen_1_1_REG & s1_way_waddr_1_1_r == io_read_2_bits_idx | s1_way_wen_1_0_REG &
    s1_way_waddr_1_0_r == io_read_2_bits_idx; // @[AsynchronousMetaArray.scala 134:85 135:29]
  reg  io_resp_2_1_r; // @[Reg.scala 16:16]
  reg  io_resp_2_1_r1; // @[Reg.scala 16:16]
  reg [5:0] io_resp_2_1_r2; // @[Reg.scala 16:16]
  wire  _GEN_1215 = 6'h1 == io_resp_2_1_r2 ? meta_array_1_1 : meta_array_0_1; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1216 = 6'h2 == io_resp_2_1_r2 ? meta_array_2_1 : _GEN_1215; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1217 = 6'h3 == io_resp_2_1_r2 ? meta_array_3_1 : _GEN_1216; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1218 = 6'h4 == io_resp_2_1_r2 ? meta_array_4_1 : _GEN_1217; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1219 = 6'h5 == io_resp_2_1_r2 ? meta_array_5_1 : _GEN_1218; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1220 = 6'h6 == io_resp_2_1_r2 ? meta_array_6_1 : _GEN_1219; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1221 = 6'h7 == io_resp_2_1_r2 ? meta_array_7_1 : _GEN_1220; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1222 = 6'h8 == io_resp_2_1_r2 ? meta_array_8_1 : _GEN_1221; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1223 = 6'h9 == io_resp_2_1_r2 ? meta_array_9_1 : _GEN_1222; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1224 = 6'ha == io_resp_2_1_r2 ? meta_array_10_1 : _GEN_1223; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1225 = 6'hb == io_resp_2_1_r2 ? meta_array_11_1 : _GEN_1224; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1226 = 6'hc == io_resp_2_1_r2 ? meta_array_12_1 : _GEN_1225; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1227 = 6'hd == io_resp_2_1_r2 ? meta_array_13_1 : _GEN_1226; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1228 = 6'he == io_resp_2_1_r2 ? meta_array_14_1 : _GEN_1227; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1229 = 6'hf == io_resp_2_1_r2 ? meta_array_15_1 : _GEN_1228; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1230 = 6'h10 == io_resp_2_1_r2 ? meta_array_16_1 : _GEN_1229; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1231 = 6'h11 == io_resp_2_1_r2 ? meta_array_17_1 : _GEN_1230; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1232 = 6'h12 == io_resp_2_1_r2 ? meta_array_18_1 : _GEN_1231; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1233 = 6'h13 == io_resp_2_1_r2 ? meta_array_19_1 : _GEN_1232; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1234 = 6'h14 == io_resp_2_1_r2 ? meta_array_20_1 : _GEN_1233; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1235 = 6'h15 == io_resp_2_1_r2 ? meta_array_21_1 : _GEN_1234; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1236 = 6'h16 == io_resp_2_1_r2 ? meta_array_22_1 : _GEN_1235; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1237 = 6'h17 == io_resp_2_1_r2 ? meta_array_23_1 : _GEN_1236; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1238 = 6'h18 == io_resp_2_1_r2 ? meta_array_24_1 : _GEN_1237; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1239 = 6'h19 == io_resp_2_1_r2 ? meta_array_25_1 : _GEN_1238; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1240 = 6'h1a == io_resp_2_1_r2 ? meta_array_26_1 : _GEN_1239; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1241 = 6'h1b == io_resp_2_1_r2 ? meta_array_27_1 : _GEN_1240; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1242 = 6'h1c == io_resp_2_1_r2 ? meta_array_28_1 : _GEN_1241; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1243 = 6'h1d == io_resp_2_1_r2 ? meta_array_29_1 : _GEN_1242; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1244 = 6'h1e == io_resp_2_1_r2 ? meta_array_30_1 : _GEN_1243; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1245 = 6'h1f == io_resp_2_1_r2 ? meta_array_31_1 : _GEN_1244; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1246 = 6'h20 == io_resp_2_1_r2 ? meta_array_32_1 : _GEN_1245; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1247 = 6'h21 == io_resp_2_1_r2 ? meta_array_33_1 : _GEN_1246; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1248 = 6'h22 == io_resp_2_1_r2 ? meta_array_34_1 : _GEN_1247; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1249 = 6'h23 == io_resp_2_1_r2 ? meta_array_35_1 : _GEN_1248; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1250 = 6'h24 == io_resp_2_1_r2 ? meta_array_36_1 : _GEN_1249; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1251 = 6'h25 == io_resp_2_1_r2 ? meta_array_37_1 : _GEN_1250; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1252 = 6'h26 == io_resp_2_1_r2 ? meta_array_38_1 : _GEN_1251; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1253 = 6'h27 == io_resp_2_1_r2 ? meta_array_39_1 : _GEN_1252; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1254 = 6'h28 == io_resp_2_1_r2 ? meta_array_40_1 : _GEN_1253; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1255 = 6'h29 == io_resp_2_1_r2 ? meta_array_41_1 : _GEN_1254; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1256 = 6'h2a == io_resp_2_1_r2 ? meta_array_42_1 : _GEN_1255; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1257 = 6'h2b == io_resp_2_1_r2 ? meta_array_43_1 : _GEN_1256; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1258 = 6'h2c == io_resp_2_1_r2 ? meta_array_44_1 : _GEN_1257; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1259 = 6'h2d == io_resp_2_1_r2 ? meta_array_45_1 : _GEN_1258; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1260 = 6'h2e == io_resp_2_1_r2 ? meta_array_46_1 : _GEN_1259; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1261 = 6'h2f == io_resp_2_1_r2 ? meta_array_47_1 : _GEN_1260; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1262 = 6'h30 == io_resp_2_1_r2 ? meta_array_48_1 : _GEN_1261; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1263 = 6'h31 == io_resp_2_1_r2 ? meta_array_49_1 : _GEN_1262; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1264 = 6'h32 == io_resp_2_1_r2 ? meta_array_50_1 : _GEN_1263; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1265 = 6'h33 == io_resp_2_1_r2 ? meta_array_51_1 : _GEN_1264; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1266 = 6'h34 == io_resp_2_1_r2 ? meta_array_52_1 : _GEN_1265; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1267 = 6'h35 == io_resp_2_1_r2 ? meta_array_53_1 : _GEN_1266; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1268 = 6'h36 == io_resp_2_1_r2 ? meta_array_54_1 : _GEN_1267; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1269 = 6'h37 == io_resp_2_1_r2 ? meta_array_55_1 : _GEN_1268; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1270 = 6'h38 == io_resp_2_1_r2 ? meta_array_56_1 : _GEN_1269; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1271 = 6'h39 == io_resp_2_1_r2 ? meta_array_57_1 : _GEN_1270; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1272 = 6'h3a == io_resp_2_1_r2 ? meta_array_58_1 : _GEN_1271; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1273 = 6'h3b == io_resp_2_1_r2 ? meta_array_59_1 : _GEN_1272; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1274 = 6'h3c == io_resp_2_1_r2 ? meta_array_60_1 : _GEN_1273; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1275 = 6'h3d == io_resp_2_1_r2 ? meta_array_61_1 : _GEN_1274; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1276 = 6'h3e == io_resp_2_1_r2 ? meta_array_62_1 : _GEN_1275; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1277 = 6'h3f == io_resp_2_1_r2 ? meta_array_63_1 : _GEN_1276; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  read_way_bypass_18 = s1_way_wen_2_1_REG & s1_way_waddr_2_1_r == io_read_2_bits_idx | s1_way_wen_2_0_REG &
    s1_way_waddr_2_0_r == io_read_2_bits_idx; // @[AsynchronousMetaArray.scala 134:85 135:29]
  reg  io_resp_2_2_r; // @[Reg.scala 16:16]
  reg  io_resp_2_2_r1; // @[Reg.scala 16:16]
  reg [5:0] io_resp_2_2_r2; // @[Reg.scala 16:16]
  wire  _GEN_1286 = 6'h1 == io_resp_2_2_r2 ? meta_array_1_2 : meta_array_0_2; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1287 = 6'h2 == io_resp_2_2_r2 ? meta_array_2_2 : _GEN_1286; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1288 = 6'h3 == io_resp_2_2_r2 ? meta_array_3_2 : _GEN_1287; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1289 = 6'h4 == io_resp_2_2_r2 ? meta_array_4_2 : _GEN_1288; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1290 = 6'h5 == io_resp_2_2_r2 ? meta_array_5_2 : _GEN_1289; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1291 = 6'h6 == io_resp_2_2_r2 ? meta_array_6_2 : _GEN_1290; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1292 = 6'h7 == io_resp_2_2_r2 ? meta_array_7_2 : _GEN_1291; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1293 = 6'h8 == io_resp_2_2_r2 ? meta_array_8_2 : _GEN_1292; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1294 = 6'h9 == io_resp_2_2_r2 ? meta_array_9_2 : _GEN_1293; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1295 = 6'ha == io_resp_2_2_r2 ? meta_array_10_2 : _GEN_1294; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1296 = 6'hb == io_resp_2_2_r2 ? meta_array_11_2 : _GEN_1295; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1297 = 6'hc == io_resp_2_2_r2 ? meta_array_12_2 : _GEN_1296; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1298 = 6'hd == io_resp_2_2_r2 ? meta_array_13_2 : _GEN_1297; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1299 = 6'he == io_resp_2_2_r2 ? meta_array_14_2 : _GEN_1298; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1300 = 6'hf == io_resp_2_2_r2 ? meta_array_15_2 : _GEN_1299; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1301 = 6'h10 == io_resp_2_2_r2 ? meta_array_16_2 : _GEN_1300; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1302 = 6'h11 == io_resp_2_2_r2 ? meta_array_17_2 : _GEN_1301; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1303 = 6'h12 == io_resp_2_2_r2 ? meta_array_18_2 : _GEN_1302; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1304 = 6'h13 == io_resp_2_2_r2 ? meta_array_19_2 : _GEN_1303; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1305 = 6'h14 == io_resp_2_2_r2 ? meta_array_20_2 : _GEN_1304; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1306 = 6'h15 == io_resp_2_2_r2 ? meta_array_21_2 : _GEN_1305; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1307 = 6'h16 == io_resp_2_2_r2 ? meta_array_22_2 : _GEN_1306; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1308 = 6'h17 == io_resp_2_2_r2 ? meta_array_23_2 : _GEN_1307; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1309 = 6'h18 == io_resp_2_2_r2 ? meta_array_24_2 : _GEN_1308; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1310 = 6'h19 == io_resp_2_2_r2 ? meta_array_25_2 : _GEN_1309; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1311 = 6'h1a == io_resp_2_2_r2 ? meta_array_26_2 : _GEN_1310; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1312 = 6'h1b == io_resp_2_2_r2 ? meta_array_27_2 : _GEN_1311; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1313 = 6'h1c == io_resp_2_2_r2 ? meta_array_28_2 : _GEN_1312; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1314 = 6'h1d == io_resp_2_2_r2 ? meta_array_29_2 : _GEN_1313; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1315 = 6'h1e == io_resp_2_2_r2 ? meta_array_30_2 : _GEN_1314; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1316 = 6'h1f == io_resp_2_2_r2 ? meta_array_31_2 : _GEN_1315; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1317 = 6'h20 == io_resp_2_2_r2 ? meta_array_32_2 : _GEN_1316; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1318 = 6'h21 == io_resp_2_2_r2 ? meta_array_33_2 : _GEN_1317; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1319 = 6'h22 == io_resp_2_2_r2 ? meta_array_34_2 : _GEN_1318; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1320 = 6'h23 == io_resp_2_2_r2 ? meta_array_35_2 : _GEN_1319; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1321 = 6'h24 == io_resp_2_2_r2 ? meta_array_36_2 : _GEN_1320; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1322 = 6'h25 == io_resp_2_2_r2 ? meta_array_37_2 : _GEN_1321; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1323 = 6'h26 == io_resp_2_2_r2 ? meta_array_38_2 : _GEN_1322; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1324 = 6'h27 == io_resp_2_2_r2 ? meta_array_39_2 : _GEN_1323; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1325 = 6'h28 == io_resp_2_2_r2 ? meta_array_40_2 : _GEN_1324; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1326 = 6'h29 == io_resp_2_2_r2 ? meta_array_41_2 : _GEN_1325; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1327 = 6'h2a == io_resp_2_2_r2 ? meta_array_42_2 : _GEN_1326; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1328 = 6'h2b == io_resp_2_2_r2 ? meta_array_43_2 : _GEN_1327; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1329 = 6'h2c == io_resp_2_2_r2 ? meta_array_44_2 : _GEN_1328; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1330 = 6'h2d == io_resp_2_2_r2 ? meta_array_45_2 : _GEN_1329; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1331 = 6'h2e == io_resp_2_2_r2 ? meta_array_46_2 : _GEN_1330; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1332 = 6'h2f == io_resp_2_2_r2 ? meta_array_47_2 : _GEN_1331; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1333 = 6'h30 == io_resp_2_2_r2 ? meta_array_48_2 : _GEN_1332; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1334 = 6'h31 == io_resp_2_2_r2 ? meta_array_49_2 : _GEN_1333; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1335 = 6'h32 == io_resp_2_2_r2 ? meta_array_50_2 : _GEN_1334; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1336 = 6'h33 == io_resp_2_2_r2 ? meta_array_51_2 : _GEN_1335; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1337 = 6'h34 == io_resp_2_2_r2 ? meta_array_52_2 : _GEN_1336; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1338 = 6'h35 == io_resp_2_2_r2 ? meta_array_53_2 : _GEN_1337; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1339 = 6'h36 == io_resp_2_2_r2 ? meta_array_54_2 : _GEN_1338; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1340 = 6'h37 == io_resp_2_2_r2 ? meta_array_55_2 : _GEN_1339; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1341 = 6'h38 == io_resp_2_2_r2 ? meta_array_56_2 : _GEN_1340; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1342 = 6'h39 == io_resp_2_2_r2 ? meta_array_57_2 : _GEN_1341; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1343 = 6'h3a == io_resp_2_2_r2 ? meta_array_58_2 : _GEN_1342; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1344 = 6'h3b == io_resp_2_2_r2 ? meta_array_59_2 : _GEN_1343; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1345 = 6'h3c == io_resp_2_2_r2 ? meta_array_60_2 : _GEN_1344; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1346 = 6'h3d == io_resp_2_2_r2 ? meta_array_61_2 : _GEN_1345; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1347 = 6'h3e == io_resp_2_2_r2 ? meta_array_62_2 : _GEN_1346; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1348 = 6'h3f == io_resp_2_2_r2 ? meta_array_63_2 : _GEN_1347; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  read_way_bypass_19 = s1_way_wen_3_1_REG & s1_way_waddr_3_1_r == io_read_2_bits_idx | s1_way_wen_3_0_REG &
    s1_way_waddr_3_0_r == io_read_2_bits_idx; // @[AsynchronousMetaArray.scala 134:85 135:29]
  reg  io_resp_2_3_r; // @[Reg.scala 16:16]
  reg  io_resp_2_3_r1; // @[Reg.scala 16:16]
  reg [5:0] io_resp_2_3_r2; // @[Reg.scala 16:16]
  wire  _GEN_1357 = 6'h1 == io_resp_2_3_r2 ? meta_array_1_3 : meta_array_0_3; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1358 = 6'h2 == io_resp_2_3_r2 ? meta_array_2_3 : _GEN_1357; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1359 = 6'h3 == io_resp_2_3_r2 ? meta_array_3_3 : _GEN_1358; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1360 = 6'h4 == io_resp_2_3_r2 ? meta_array_4_3 : _GEN_1359; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1361 = 6'h5 == io_resp_2_3_r2 ? meta_array_5_3 : _GEN_1360; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1362 = 6'h6 == io_resp_2_3_r2 ? meta_array_6_3 : _GEN_1361; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1363 = 6'h7 == io_resp_2_3_r2 ? meta_array_7_3 : _GEN_1362; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1364 = 6'h8 == io_resp_2_3_r2 ? meta_array_8_3 : _GEN_1363; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1365 = 6'h9 == io_resp_2_3_r2 ? meta_array_9_3 : _GEN_1364; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1366 = 6'ha == io_resp_2_3_r2 ? meta_array_10_3 : _GEN_1365; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1367 = 6'hb == io_resp_2_3_r2 ? meta_array_11_3 : _GEN_1366; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1368 = 6'hc == io_resp_2_3_r2 ? meta_array_12_3 : _GEN_1367; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1369 = 6'hd == io_resp_2_3_r2 ? meta_array_13_3 : _GEN_1368; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1370 = 6'he == io_resp_2_3_r2 ? meta_array_14_3 : _GEN_1369; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1371 = 6'hf == io_resp_2_3_r2 ? meta_array_15_3 : _GEN_1370; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1372 = 6'h10 == io_resp_2_3_r2 ? meta_array_16_3 : _GEN_1371; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1373 = 6'h11 == io_resp_2_3_r2 ? meta_array_17_3 : _GEN_1372; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1374 = 6'h12 == io_resp_2_3_r2 ? meta_array_18_3 : _GEN_1373; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1375 = 6'h13 == io_resp_2_3_r2 ? meta_array_19_3 : _GEN_1374; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1376 = 6'h14 == io_resp_2_3_r2 ? meta_array_20_3 : _GEN_1375; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1377 = 6'h15 == io_resp_2_3_r2 ? meta_array_21_3 : _GEN_1376; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1378 = 6'h16 == io_resp_2_3_r2 ? meta_array_22_3 : _GEN_1377; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1379 = 6'h17 == io_resp_2_3_r2 ? meta_array_23_3 : _GEN_1378; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1380 = 6'h18 == io_resp_2_3_r2 ? meta_array_24_3 : _GEN_1379; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1381 = 6'h19 == io_resp_2_3_r2 ? meta_array_25_3 : _GEN_1380; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1382 = 6'h1a == io_resp_2_3_r2 ? meta_array_26_3 : _GEN_1381; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1383 = 6'h1b == io_resp_2_3_r2 ? meta_array_27_3 : _GEN_1382; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1384 = 6'h1c == io_resp_2_3_r2 ? meta_array_28_3 : _GEN_1383; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1385 = 6'h1d == io_resp_2_3_r2 ? meta_array_29_3 : _GEN_1384; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1386 = 6'h1e == io_resp_2_3_r2 ? meta_array_30_3 : _GEN_1385; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1387 = 6'h1f == io_resp_2_3_r2 ? meta_array_31_3 : _GEN_1386; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1388 = 6'h20 == io_resp_2_3_r2 ? meta_array_32_3 : _GEN_1387; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1389 = 6'h21 == io_resp_2_3_r2 ? meta_array_33_3 : _GEN_1388; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1390 = 6'h22 == io_resp_2_3_r2 ? meta_array_34_3 : _GEN_1389; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1391 = 6'h23 == io_resp_2_3_r2 ? meta_array_35_3 : _GEN_1390; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1392 = 6'h24 == io_resp_2_3_r2 ? meta_array_36_3 : _GEN_1391; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1393 = 6'h25 == io_resp_2_3_r2 ? meta_array_37_3 : _GEN_1392; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1394 = 6'h26 == io_resp_2_3_r2 ? meta_array_38_3 : _GEN_1393; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1395 = 6'h27 == io_resp_2_3_r2 ? meta_array_39_3 : _GEN_1394; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1396 = 6'h28 == io_resp_2_3_r2 ? meta_array_40_3 : _GEN_1395; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1397 = 6'h29 == io_resp_2_3_r2 ? meta_array_41_3 : _GEN_1396; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1398 = 6'h2a == io_resp_2_3_r2 ? meta_array_42_3 : _GEN_1397; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1399 = 6'h2b == io_resp_2_3_r2 ? meta_array_43_3 : _GEN_1398; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1400 = 6'h2c == io_resp_2_3_r2 ? meta_array_44_3 : _GEN_1399; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1401 = 6'h2d == io_resp_2_3_r2 ? meta_array_45_3 : _GEN_1400; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1402 = 6'h2e == io_resp_2_3_r2 ? meta_array_46_3 : _GEN_1401; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1403 = 6'h2f == io_resp_2_3_r2 ? meta_array_47_3 : _GEN_1402; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1404 = 6'h30 == io_resp_2_3_r2 ? meta_array_48_3 : _GEN_1403; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1405 = 6'h31 == io_resp_2_3_r2 ? meta_array_49_3 : _GEN_1404; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1406 = 6'h32 == io_resp_2_3_r2 ? meta_array_50_3 : _GEN_1405; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1407 = 6'h33 == io_resp_2_3_r2 ? meta_array_51_3 : _GEN_1406; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1408 = 6'h34 == io_resp_2_3_r2 ? meta_array_52_3 : _GEN_1407; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1409 = 6'h35 == io_resp_2_3_r2 ? meta_array_53_3 : _GEN_1408; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1410 = 6'h36 == io_resp_2_3_r2 ? meta_array_54_3 : _GEN_1409; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1411 = 6'h37 == io_resp_2_3_r2 ? meta_array_55_3 : _GEN_1410; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1412 = 6'h38 == io_resp_2_3_r2 ? meta_array_56_3 : _GEN_1411; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1413 = 6'h39 == io_resp_2_3_r2 ? meta_array_57_3 : _GEN_1412; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1414 = 6'h3a == io_resp_2_3_r2 ? meta_array_58_3 : _GEN_1413; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1415 = 6'h3b == io_resp_2_3_r2 ? meta_array_59_3 : _GEN_1414; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1416 = 6'h3c == io_resp_2_3_r2 ? meta_array_60_3 : _GEN_1415; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1417 = 6'h3d == io_resp_2_3_r2 ? meta_array_61_3 : _GEN_1416; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1418 = 6'h3e == io_resp_2_3_r2 ? meta_array_62_3 : _GEN_1417; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1419 = 6'h3f == io_resp_2_3_r2 ? meta_array_63_3 : _GEN_1418; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  read_way_bypass_20 = s1_way_wen_4_1_REG & s1_way_waddr_4_1_r == io_read_2_bits_idx | s1_way_wen_4_0_REG &
    s1_way_waddr_4_0_r == io_read_2_bits_idx; // @[AsynchronousMetaArray.scala 134:85 135:29]
  reg  io_resp_2_4_r; // @[Reg.scala 16:16]
  reg  io_resp_2_4_r1; // @[Reg.scala 16:16]
  reg [5:0] io_resp_2_4_r2; // @[Reg.scala 16:16]
  wire  _GEN_1428 = 6'h1 == io_resp_2_4_r2 ? meta_array_1_4 : meta_array_0_4; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1429 = 6'h2 == io_resp_2_4_r2 ? meta_array_2_4 : _GEN_1428; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1430 = 6'h3 == io_resp_2_4_r2 ? meta_array_3_4 : _GEN_1429; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1431 = 6'h4 == io_resp_2_4_r2 ? meta_array_4_4 : _GEN_1430; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1432 = 6'h5 == io_resp_2_4_r2 ? meta_array_5_4 : _GEN_1431; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1433 = 6'h6 == io_resp_2_4_r2 ? meta_array_6_4 : _GEN_1432; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1434 = 6'h7 == io_resp_2_4_r2 ? meta_array_7_4 : _GEN_1433; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1435 = 6'h8 == io_resp_2_4_r2 ? meta_array_8_4 : _GEN_1434; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1436 = 6'h9 == io_resp_2_4_r2 ? meta_array_9_4 : _GEN_1435; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1437 = 6'ha == io_resp_2_4_r2 ? meta_array_10_4 : _GEN_1436; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1438 = 6'hb == io_resp_2_4_r2 ? meta_array_11_4 : _GEN_1437; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1439 = 6'hc == io_resp_2_4_r2 ? meta_array_12_4 : _GEN_1438; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1440 = 6'hd == io_resp_2_4_r2 ? meta_array_13_4 : _GEN_1439; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1441 = 6'he == io_resp_2_4_r2 ? meta_array_14_4 : _GEN_1440; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1442 = 6'hf == io_resp_2_4_r2 ? meta_array_15_4 : _GEN_1441; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1443 = 6'h10 == io_resp_2_4_r2 ? meta_array_16_4 : _GEN_1442; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1444 = 6'h11 == io_resp_2_4_r2 ? meta_array_17_4 : _GEN_1443; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1445 = 6'h12 == io_resp_2_4_r2 ? meta_array_18_4 : _GEN_1444; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1446 = 6'h13 == io_resp_2_4_r2 ? meta_array_19_4 : _GEN_1445; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1447 = 6'h14 == io_resp_2_4_r2 ? meta_array_20_4 : _GEN_1446; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1448 = 6'h15 == io_resp_2_4_r2 ? meta_array_21_4 : _GEN_1447; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1449 = 6'h16 == io_resp_2_4_r2 ? meta_array_22_4 : _GEN_1448; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1450 = 6'h17 == io_resp_2_4_r2 ? meta_array_23_4 : _GEN_1449; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1451 = 6'h18 == io_resp_2_4_r2 ? meta_array_24_4 : _GEN_1450; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1452 = 6'h19 == io_resp_2_4_r2 ? meta_array_25_4 : _GEN_1451; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1453 = 6'h1a == io_resp_2_4_r2 ? meta_array_26_4 : _GEN_1452; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1454 = 6'h1b == io_resp_2_4_r2 ? meta_array_27_4 : _GEN_1453; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1455 = 6'h1c == io_resp_2_4_r2 ? meta_array_28_4 : _GEN_1454; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1456 = 6'h1d == io_resp_2_4_r2 ? meta_array_29_4 : _GEN_1455; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1457 = 6'h1e == io_resp_2_4_r2 ? meta_array_30_4 : _GEN_1456; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1458 = 6'h1f == io_resp_2_4_r2 ? meta_array_31_4 : _GEN_1457; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1459 = 6'h20 == io_resp_2_4_r2 ? meta_array_32_4 : _GEN_1458; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1460 = 6'h21 == io_resp_2_4_r2 ? meta_array_33_4 : _GEN_1459; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1461 = 6'h22 == io_resp_2_4_r2 ? meta_array_34_4 : _GEN_1460; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1462 = 6'h23 == io_resp_2_4_r2 ? meta_array_35_4 : _GEN_1461; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1463 = 6'h24 == io_resp_2_4_r2 ? meta_array_36_4 : _GEN_1462; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1464 = 6'h25 == io_resp_2_4_r2 ? meta_array_37_4 : _GEN_1463; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1465 = 6'h26 == io_resp_2_4_r2 ? meta_array_38_4 : _GEN_1464; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1466 = 6'h27 == io_resp_2_4_r2 ? meta_array_39_4 : _GEN_1465; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1467 = 6'h28 == io_resp_2_4_r2 ? meta_array_40_4 : _GEN_1466; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1468 = 6'h29 == io_resp_2_4_r2 ? meta_array_41_4 : _GEN_1467; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1469 = 6'h2a == io_resp_2_4_r2 ? meta_array_42_4 : _GEN_1468; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1470 = 6'h2b == io_resp_2_4_r2 ? meta_array_43_4 : _GEN_1469; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1471 = 6'h2c == io_resp_2_4_r2 ? meta_array_44_4 : _GEN_1470; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1472 = 6'h2d == io_resp_2_4_r2 ? meta_array_45_4 : _GEN_1471; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1473 = 6'h2e == io_resp_2_4_r2 ? meta_array_46_4 : _GEN_1472; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1474 = 6'h2f == io_resp_2_4_r2 ? meta_array_47_4 : _GEN_1473; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1475 = 6'h30 == io_resp_2_4_r2 ? meta_array_48_4 : _GEN_1474; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1476 = 6'h31 == io_resp_2_4_r2 ? meta_array_49_4 : _GEN_1475; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1477 = 6'h32 == io_resp_2_4_r2 ? meta_array_50_4 : _GEN_1476; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1478 = 6'h33 == io_resp_2_4_r2 ? meta_array_51_4 : _GEN_1477; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1479 = 6'h34 == io_resp_2_4_r2 ? meta_array_52_4 : _GEN_1478; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1480 = 6'h35 == io_resp_2_4_r2 ? meta_array_53_4 : _GEN_1479; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1481 = 6'h36 == io_resp_2_4_r2 ? meta_array_54_4 : _GEN_1480; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1482 = 6'h37 == io_resp_2_4_r2 ? meta_array_55_4 : _GEN_1481; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1483 = 6'h38 == io_resp_2_4_r2 ? meta_array_56_4 : _GEN_1482; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1484 = 6'h39 == io_resp_2_4_r2 ? meta_array_57_4 : _GEN_1483; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1485 = 6'h3a == io_resp_2_4_r2 ? meta_array_58_4 : _GEN_1484; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1486 = 6'h3b == io_resp_2_4_r2 ? meta_array_59_4 : _GEN_1485; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1487 = 6'h3c == io_resp_2_4_r2 ? meta_array_60_4 : _GEN_1486; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1488 = 6'h3d == io_resp_2_4_r2 ? meta_array_61_4 : _GEN_1487; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1489 = 6'h3e == io_resp_2_4_r2 ? meta_array_62_4 : _GEN_1488; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1490 = 6'h3f == io_resp_2_4_r2 ? meta_array_63_4 : _GEN_1489; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  read_way_bypass_21 = s1_way_wen_5_1_REG & s1_way_waddr_5_1_r == io_read_2_bits_idx | s1_way_wen_5_0_REG &
    s1_way_waddr_5_0_r == io_read_2_bits_idx; // @[AsynchronousMetaArray.scala 134:85 135:29]
  reg  io_resp_2_5_r; // @[Reg.scala 16:16]
  reg  io_resp_2_5_r1; // @[Reg.scala 16:16]
  reg [5:0] io_resp_2_5_r2; // @[Reg.scala 16:16]
  wire  _GEN_1499 = 6'h1 == io_resp_2_5_r2 ? meta_array_1_5 : meta_array_0_5; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1500 = 6'h2 == io_resp_2_5_r2 ? meta_array_2_5 : _GEN_1499; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1501 = 6'h3 == io_resp_2_5_r2 ? meta_array_3_5 : _GEN_1500; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1502 = 6'h4 == io_resp_2_5_r2 ? meta_array_4_5 : _GEN_1501; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1503 = 6'h5 == io_resp_2_5_r2 ? meta_array_5_5 : _GEN_1502; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1504 = 6'h6 == io_resp_2_5_r2 ? meta_array_6_5 : _GEN_1503; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1505 = 6'h7 == io_resp_2_5_r2 ? meta_array_7_5 : _GEN_1504; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1506 = 6'h8 == io_resp_2_5_r2 ? meta_array_8_5 : _GEN_1505; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1507 = 6'h9 == io_resp_2_5_r2 ? meta_array_9_5 : _GEN_1506; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1508 = 6'ha == io_resp_2_5_r2 ? meta_array_10_5 : _GEN_1507; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1509 = 6'hb == io_resp_2_5_r2 ? meta_array_11_5 : _GEN_1508; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1510 = 6'hc == io_resp_2_5_r2 ? meta_array_12_5 : _GEN_1509; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1511 = 6'hd == io_resp_2_5_r2 ? meta_array_13_5 : _GEN_1510; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1512 = 6'he == io_resp_2_5_r2 ? meta_array_14_5 : _GEN_1511; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1513 = 6'hf == io_resp_2_5_r2 ? meta_array_15_5 : _GEN_1512; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1514 = 6'h10 == io_resp_2_5_r2 ? meta_array_16_5 : _GEN_1513; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1515 = 6'h11 == io_resp_2_5_r2 ? meta_array_17_5 : _GEN_1514; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1516 = 6'h12 == io_resp_2_5_r2 ? meta_array_18_5 : _GEN_1515; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1517 = 6'h13 == io_resp_2_5_r2 ? meta_array_19_5 : _GEN_1516; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1518 = 6'h14 == io_resp_2_5_r2 ? meta_array_20_5 : _GEN_1517; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1519 = 6'h15 == io_resp_2_5_r2 ? meta_array_21_5 : _GEN_1518; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1520 = 6'h16 == io_resp_2_5_r2 ? meta_array_22_5 : _GEN_1519; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1521 = 6'h17 == io_resp_2_5_r2 ? meta_array_23_5 : _GEN_1520; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1522 = 6'h18 == io_resp_2_5_r2 ? meta_array_24_5 : _GEN_1521; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1523 = 6'h19 == io_resp_2_5_r2 ? meta_array_25_5 : _GEN_1522; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1524 = 6'h1a == io_resp_2_5_r2 ? meta_array_26_5 : _GEN_1523; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1525 = 6'h1b == io_resp_2_5_r2 ? meta_array_27_5 : _GEN_1524; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1526 = 6'h1c == io_resp_2_5_r2 ? meta_array_28_5 : _GEN_1525; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1527 = 6'h1d == io_resp_2_5_r2 ? meta_array_29_5 : _GEN_1526; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1528 = 6'h1e == io_resp_2_5_r2 ? meta_array_30_5 : _GEN_1527; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1529 = 6'h1f == io_resp_2_5_r2 ? meta_array_31_5 : _GEN_1528; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1530 = 6'h20 == io_resp_2_5_r2 ? meta_array_32_5 : _GEN_1529; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1531 = 6'h21 == io_resp_2_5_r2 ? meta_array_33_5 : _GEN_1530; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1532 = 6'h22 == io_resp_2_5_r2 ? meta_array_34_5 : _GEN_1531; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1533 = 6'h23 == io_resp_2_5_r2 ? meta_array_35_5 : _GEN_1532; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1534 = 6'h24 == io_resp_2_5_r2 ? meta_array_36_5 : _GEN_1533; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1535 = 6'h25 == io_resp_2_5_r2 ? meta_array_37_5 : _GEN_1534; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1536 = 6'h26 == io_resp_2_5_r2 ? meta_array_38_5 : _GEN_1535; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1537 = 6'h27 == io_resp_2_5_r2 ? meta_array_39_5 : _GEN_1536; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1538 = 6'h28 == io_resp_2_5_r2 ? meta_array_40_5 : _GEN_1537; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1539 = 6'h29 == io_resp_2_5_r2 ? meta_array_41_5 : _GEN_1538; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1540 = 6'h2a == io_resp_2_5_r2 ? meta_array_42_5 : _GEN_1539; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1541 = 6'h2b == io_resp_2_5_r2 ? meta_array_43_5 : _GEN_1540; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1542 = 6'h2c == io_resp_2_5_r2 ? meta_array_44_5 : _GEN_1541; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1543 = 6'h2d == io_resp_2_5_r2 ? meta_array_45_5 : _GEN_1542; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1544 = 6'h2e == io_resp_2_5_r2 ? meta_array_46_5 : _GEN_1543; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1545 = 6'h2f == io_resp_2_5_r2 ? meta_array_47_5 : _GEN_1544; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1546 = 6'h30 == io_resp_2_5_r2 ? meta_array_48_5 : _GEN_1545; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1547 = 6'h31 == io_resp_2_5_r2 ? meta_array_49_5 : _GEN_1546; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1548 = 6'h32 == io_resp_2_5_r2 ? meta_array_50_5 : _GEN_1547; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1549 = 6'h33 == io_resp_2_5_r2 ? meta_array_51_5 : _GEN_1548; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1550 = 6'h34 == io_resp_2_5_r2 ? meta_array_52_5 : _GEN_1549; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1551 = 6'h35 == io_resp_2_5_r2 ? meta_array_53_5 : _GEN_1550; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1552 = 6'h36 == io_resp_2_5_r2 ? meta_array_54_5 : _GEN_1551; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1553 = 6'h37 == io_resp_2_5_r2 ? meta_array_55_5 : _GEN_1552; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1554 = 6'h38 == io_resp_2_5_r2 ? meta_array_56_5 : _GEN_1553; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1555 = 6'h39 == io_resp_2_5_r2 ? meta_array_57_5 : _GEN_1554; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1556 = 6'h3a == io_resp_2_5_r2 ? meta_array_58_5 : _GEN_1555; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1557 = 6'h3b == io_resp_2_5_r2 ? meta_array_59_5 : _GEN_1556; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1558 = 6'h3c == io_resp_2_5_r2 ? meta_array_60_5 : _GEN_1557; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1559 = 6'h3d == io_resp_2_5_r2 ? meta_array_61_5 : _GEN_1558; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1560 = 6'h3e == io_resp_2_5_r2 ? meta_array_62_5 : _GEN_1559; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1561 = 6'h3f == io_resp_2_5_r2 ? meta_array_63_5 : _GEN_1560; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  read_way_bypass_22 = s1_way_wen_6_1_REG & s1_way_waddr_6_1_r == io_read_2_bits_idx | s1_way_wen_6_0_REG &
    s1_way_waddr_6_0_r == io_read_2_bits_idx; // @[AsynchronousMetaArray.scala 134:85 135:29]
  reg  io_resp_2_6_r; // @[Reg.scala 16:16]
  reg  io_resp_2_6_r1; // @[Reg.scala 16:16]
  reg [5:0] io_resp_2_6_r2; // @[Reg.scala 16:16]
  wire  _GEN_1570 = 6'h1 == io_resp_2_6_r2 ? meta_array_1_6 : meta_array_0_6; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1571 = 6'h2 == io_resp_2_6_r2 ? meta_array_2_6 : _GEN_1570; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1572 = 6'h3 == io_resp_2_6_r2 ? meta_array_3_6 : _GEN_1571; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1573 = 6'h4 == io_resp_2_6_r2 ? meta_array_4_6 : _GEN_1572; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1574 = 6'h5 == io_resp_2_6_r2 ? meta_array_5_6 : _GEN_1573; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1575 = 6'h6 == io_resp_2_6_r2 ? meta_array_6_6 : _GEN_1574; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1576 = 6'h7 == io_resp_2_6_r2 ? meta_array_7_6 : _GEN_1575; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1577 = 6'h8 == io_resp_2_6_r2 ? meta_array_8_6 : _GEN_1576; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1578 = 6'h9 == io_resp_2_6_r2 ? meta_array_9_6 : _GEN_1577; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1579 = 6'ha == io_resp_2_6_r2 ? meta_array_10_6 : _GEN_1578; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1580 = 6'hb == io_resp_2_6_r2 ? meta_array_11_6 : _GEN_1579; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1581 = 6'hc == io_resp_2_6_r2 ? meta_array_12_6 : _GEN_1580; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1582 = 6'hd == io_resp_2_6_r2 ? meta_array_13_6 : _GEN_1581; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1583 = 6'he == io_resp_2_6_r2 ? meta_array_14_6 : _GEN_1582; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1584 = 6'hf == io_resp_2_6_r2 ? meta_array_15_6 : _GEN_1583; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1585 = 6'h10 == io_resp_2_6_r2 ? meta_array_16_6 : _GEN_1584; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1586 = 6'h11 == io_resp_2_6_r2 ? meta_array_17_6 : _GEN_1585; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1587 = 6'h12 == io_resp_2_6_r2 ? meta_array_18_6 : _GEN_1586; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1588 = 6'h13 == io_resp_2_6_r2 ? meta_array_19_6 : _GEN_1587; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1589 = 6'h14 == io_resp_2_6_r2 ? meta_array_20_6 : _GEN_1588; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1590 = 6'h15 == io_resp_2_6_r2 ? meta_array_21_6 : _GEN_1589; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1591 = 6'h16 == io_resp_2_6_r2 ? meta_array_22_6 : _GEN_1590; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1592 = 6'h17 == io_resp_2_6_r2 ? meta_array_23_6 : _GEN_1591; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1593 = 6'h18 == io_resp_2_6_r2 ? meta_array_24_6 : _GEN_1592; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1594 = 6'h19 == io_resp_2_6_r2 ? meta_array_25_6 : _GEN_1593; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1595 = 6'h1a == io_resp_2_6_r2 ? meta_array_26_6 : _GEN_1594; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1596 = 6'h1b == io_resp_2_6_r2 ? meta_array_27_6 : _GEN_1595; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1597 = 6'h1c == io_resp_2_6_r2 ? meta_array_28_6 : _GEN_1596; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1598 = 6'h1d == io_resp_2_6_r2 ? meta_array_29_6 : _GEN_1597; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1599 = 6'h1e == io_resp_2_6_r2 ? meta_array_30_6 : _GEN_1598; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1600 = 6'h1f == io_resp_2_6_r2 ? meta_array_31_6 : _GEN_1599; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1601 = 6'h20 == io_resp_2_6_r2 ? meta_array_32_6 : _GEN_1600; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1602 = 6'h21 == io_resp_2_6_r2 ? meta_array_33_6 : _GEN_1601; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1603 = 6'h22 == io_resp_2_6_r2 ? meta_array_34_6 : _GEN_1602; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1604 = 6'h23 == io_resp_2_6_r2 ? meta_array_35_6 : _GEN_1603; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1605 = 6'h24 == io_resp_2_6_r2 ? meta_array_36_6 : _GEN_1604; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1606 = 6'h25 == io_resp_2_6_r2 ? meta_array_37_6 : _GEN_1605; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1607 = 6'h26 == io_resp_2_6_r2 ? meta_array_38_6 : _GEN_1606; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1608 = 6'h27 == io_resp_2_6_r2 ? meta_array_39_6 : _GEN_1607; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1609 = 6'h28 == io_resp_2_6_r2 ? meta_array_40_6 : _GEN_1608; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1610 = 6'h29 == io_resp_2_6_r2 ? meta_array_41_6 : _GEN_1609; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1611 = 6'h2a == io_resp_2_6_r2 ? meta_array_42_6 : _GEN_1610; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1612 = 6'h2b == io_resp_2_6_r2 ? meta_array_43_6 : _GEN_1611; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1613 = 6'h2c == io_resp_2_6_r2 ? meta_array_44_6 : _GEN_1612; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1614 = 6'h2d == io_resp_2_6_r2 ? meta_array_45_6 : _GEN_1613; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1615 = 6'h2e == io_resp_2_6_r2 ? meta_array_46_6 : _GEN_1614; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1616 = 6'h2f == io_resp_2_6_r2 ? meta_array_47_6 : _GEN_1615; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1617 = 6'h30 == io_resp_2_6_r2 ? meta_array_48_6 : _GEN_1616; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1618 = 6'h31 == io_resp_2_6_r2 ? meta_array_49_6 : _GEN_1617; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1619 = 6'h32 == io_resp_2_6_r2 ? meta_array_50_6 : _GEN_1618; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1620 = 6'h33 == io_resp_2_6_r2 ? meta_array_51_6 : _GEN_1619; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1621 = 6'h34 == io_resp_2_6_r2 ? meta_array_52_6 : _GEN_1620; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1622 = 6'h35 == io_resp_2_6_r2 ? meta_array_53_6 : _GEN_1621; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1623 = 6'h36 == io_resp_2_6_r2 ? meta_array_54_6 : _GEN_1622; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1624 = 6'h37 == io_resp_2_6_r2 ? meta_array_55_6 : _GEN_1623; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1625 = 6'h38 == io_resp_2_6_r2 ? meta_array_56_6 : _GEN_1624; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1626 = 6'h39 == io_resp_2_6_r2 ? meta_array_57_6 : _GEN_1625; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1627 = 6'h3a == io_resp_2_6_r2 ? meta_array_58_6 : _GEN_1626; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1628 = 6'h3b == io_resp_2_6_r2 ? meta_array_59_6 : _GEN_1627; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1629 = 6'h3c == io_resp_2_6_r2 ? meta_array_60_6 : _GEN_1628; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1630 = 6'h3d == io_resp_2_6_r2 ? meta_array_61_6 : _GEN_1629; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1631 = 6'h3e == io_resp_2_6_r2 ? meta_array_62_6 : _GEN_1630; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1632 = 6'h3f == io_resp_2_6_r2 ? meta_array_63_6 : _GEN_1631; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  read_way_bypass_23 = s1_way_wen_7_1_REG & s1_way_waddr_7_1_r == io_read_2_bits_idx | s1_way_wen_7_0_REG &
    s1_way_waddr_7_0_r == io_read_2_bits_idx; // @[AsynchronousMetaArray.scala 134:85 135:29]
  reg  io_resp_2_7_r; // @[Reg.scala 16:16]
  reg  io_resp_2_7_r1; // @[Reg.scala 16:16]
  reg [5:0] io_resp_2_7_r2; // @[Reg.scala 16:16]
  wire  _GEN_1641 = 6'h1 == io_resp_2_7_r2 ? meta_array_1_7 : meta_array_0_7; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1642 = 6'h2 == io_resp_2_7_r2 ? meta_array_2_7 : _GEN_1641; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1643 = 6'h3 == io_resp_2_7_r2 ? meta_array_3_7 : _GEN_1642; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1644 = 6'h4 == io_resp_2_7_r2 ? meta_array_4_7 : _GEN_1643; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1645 = 6'h5 == io_resp_2_7_r2 ? meta_array_5_7 : _GEN_1644; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1646 = 6'h6 == io_resp_2_7_r2 ? meta_array_6_7 : _GEN_1645; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1647 = 6'h7 == io_resp_2_7_r2 ? meta_array_7_7 : _GEN_1646; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1648 = 6'h8 == io_resp_2_7_r2 ? meta_array_8_7 : _GEN_1647; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1649 = 6'h9 == io_resp_2_7_r2 ? meta_array_9_7 : _GEN_1648; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1650 = 6'ha == io_resp_2_7_r2 ? meta_array_10_7 : _GEN_1649; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1651 = 6'hb == io_resp_2_7_r2 ? meta_array_11_7 : _GEN_1650; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1652 = 6'hc == io_resp_2_7_r2 ? meta_array_12_7 : _GEN_1651; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1653 = 6'hd == io_resp_2_7_r2 ? meta_array_13_7 : _GEN_1652; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1654 = 6'he == io_resp_2_7_r2 ? meta_array_14_7 : _GEN_1653; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1655 = 6'hf == io_resp_2_7_r2 ? meta_array_15_7 : _GEN_1654; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1656 = 6'h10 == io_resp_2_7_r2 ? meta_array_16_7 : _GEN_1655; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1657 = 6'h11 == io_resp_2_7_r2 ? meta_array_17_7 : _GEN_1656; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1658 = 6'h12 == io_resp_2_7_r2 ? meta_array_18_7 : _GEN_1657; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1659 = 6'h13 == io_resp_2_7_r2 ? meta_array_19_7 : _GEN_1658; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1660 = 6'h14 == io_resp_2_7_r2 ? meta_array_20_7 : _GEN_1659; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1661 = 6'h15 == io_resp_2_7_r2 ? meta_array_21_7 : _GEN_1660; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1662 = 6'h16 == io_resp_2_7_r2 ? meta_array_22_7 : _GEN_1661; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1663 = 6'h17 == io_resp_2_7_r2 ? meta_array_23_7 : _GEN_1662; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1664 = 6'h18 == io_resp_2_7_r2 ? meta_array_24_7 : _GEN_1663; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1665 = 6'h19 == io_resp_2_7_r2 ? meta_array_25_7 : _GEN_1664; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1666 = 6'h1a == io_resp_2_7_r2 ? meta_array_26_7 : _GEN_1665; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1667 = 6'h1b == io_resp_2_7_r2 ? meta_array_27_7 : _GEN_1666; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1668 = 6'h1c == io_resp_2_7_r2 ? meta_array_28_7 : _GEN_1667; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1669 = 6'h1d == io_resp_2_7_r2 ? meta_array_29_7 : _GEN_1668; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1670 = 6'h1e == io_resp_2_7_r2 ? meta_array_30_7 : _GEN_1669; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1671 = 6'h1f == io_resp_2_7_r2 ? meta_array_31_7 : _GEN_1670; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1672 = 6'h20 == io_resp_2_7_r2 ? meta_array_32_7 : _GEN_1671; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1673 = 6'h21 == io_resp_2_7_r2 ? meta_array_33_7 : _GEN_1672; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1674 = 6'h22 == io_resp_2_7_r2 ? meta_array_34_7 : _GEN_1673; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1675 = 6'h23 == io_resp_2_7_r2 ? meta_array_35_7 : _GEN_1674; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1676 = 6'h24 == io_resp_2_7_r2 ? meta_array_36_7 : _GEN_1675; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1677 = 6'h25 == io_resp_2_7_r2 ? meta_array_37_7 : _GEN_1676; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1678 = 6'h26 == io_resp_2_7_r2 ? meta_array_38_7 : _GEN_1677; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1679 = 6'h27 == io_resp_2_7_r2 ? meta_array_39_7 : _GEN_1678; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1680 = 6'h28 == io_resp_2_7_r2 ? meta_array_40_7 : _GEN_1679; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1681 = 6'h29 == io_resp_2_7_r2 ? meta_array_41_7 : _GEN_1680; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1682 = 6'h2a == io_resp_2_7_r2 ? meta_array_42_7 : _GEN_1681; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1683 = 6'h2b == io_resp_2_7_r2 ? meta_array_43_7 : _GEN_1682; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1684 = 6'h2c == io_resp_2_7_r2 ? meta_array_44_7 : _GEN_1683; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1685 = 6'h2d == io_resp_2_7_r2 ? meta_array_45_7 : _GEN_1684; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1686 = 6'h2e == io_resp_2_7_r2 ? meta_array_46_7 : _GEN_1685; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1687 = 6'h2f == io_resp_2_7_r2 ? meta_array_47_7 : _GEN_1686; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1688 = 6'h30 == io_resp_2_7_r2 ? meta_array_48_7 : _GEN_1687; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1689 = 6'h31 == io_resp_2_7_r2 ? meta_array_49_7 : _GEN_1688; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1690 = 6'h32 == io_resp_2_7_r2 ? meta_array_50_7 : _GEN_1689; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1691 = 6'h33 == io_resp_2_7_r2 ? meta_array_51_7 : _GEN_1690; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1692 = 6'h34 == io_resp_2_7_r2 ? meta_array_52_7 : _GEN_1691; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1693 = 6'h35 == io_resp_2_7_r2 ? meta_array_53_7 : _GEN_1692; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1694 = 6'h36 == io_resp_2_7_r2 ? meta_array_54_7 : _GEN_1693; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1695 = 6'h37 == io_resp_2_7_r2 ? meta_array_55_7 : _GEN_1694; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1696 = 6'h38 == io_resp_2_7_r2 ? meta_array_56_7 : _GEN_1695; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1697 = 6'h39 == io_resp_2_7_r2 ? meta_array_57_7 : _GEN_1696; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1698 = 6'h3a == io_resp_2_7_r2 ? meta_array_58_7 : _GEN_1697; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1699 = 6'h3b == io_resp_2_7_r2 ? meta_array_59_7 : _GEN_1698; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1700 = 6'h3c == io_resp_2_7_r2 ? meta_array_60_7 : _GEN_1699; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1701 = 6'h3d == io_resp_2_7_r2 ? meta_array_61_7 : _GEN_1700; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1702 = 6'h3e == io_resp_2_7_r2 ? meta_array_62_7 : _GEN_1701; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  _GEN_1703 = 6'h3f == io_resp_2_7_r2 ? meta_array_63_7 : _GEN_1702; // @[AsynchronousMetaArray.scala 139:{25,25}]
  wire  s0_way_wen_0_0 = io_write_0_valid & io_write_0_bits_way_en[0]; // @[AsynchronousMetaArray.scala 152:49]
  wire  _GEN_1706 = 6'h0 == s1_way_waddr_0_0_r ? s1_way_wdata_0_0_r : meta_array_0_0; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1707 = 6'h1 == s1_way_waddr_0_0_r ? s1_way_wdata_0_0_r : meta_array_1_0; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1708 = 6'h2 == s1_way_waddr_0_0_r ? s1_way_wdata_0_0_r : meta_array_2_0; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1709 = 6'h3 == s1_way_waddr_0_0_r ? s1_way_wdata_0_0_r : meta_array_3_0; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1710 = 6'h4 == s1_way_waddr_0_0_r ? s1_way_wdata_0_0_r : meta_array_4_0; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1711 = 6'h5 == s1_way_waddr_0_0_r ? s1_way_wdata_0_0_r : meta_array_5_0; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1712 = 6'h6 == s1_way_waddr_0_0_r ? s1_way_wdata_0_0_r : meta_array_6_0; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1713 = 6'h7 == s1_way_waddr_0_0_r ? s1_way_wdata_0_0_r : meta_array_7_0; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1714 = 6'h8 == s1_way_waddr_0_0_r ? s1_way_wdata_0_0_r : meta_array_8_0; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1715 = 6'h9 == s1_way_waddr_0_0_r ? s1_way_wdata_0_0_r : meta_array_9_0; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1716 = 6'ha == s1_way_waddr_0_0_r ? s1_way_wdata_0_0_r : meta_array_10_0; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1717 = 6'hb == s1_way_waddr_0_0_r ? s1_way_wdata_0_0_r : meta_array_11_0; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1718 = 6'hc == s1_way_waddr_0_0_r ? s1_way_wdata_0_0_r : meta_array_12_0; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1719 = 6'hd == s1_way_waddr_0_0_r ? s1_way_wdata_0_0_r : meta_array_13_0; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1720 = 6'he == s1_way_waddr_0_0_r ? s1_way_wdata_0_0_r : meta_array_14_0; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1721 = 6'hf == s1_way_waddr_0_0_r ? s1_way_wdata_0_0_r : meta_array_15_0; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1722 = 6'h10 == s1_way_waddr_0_0_r ? s1_way_wdata_0_0_r : meta_array_16_0; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1723 = 6'h11 == s1_way_waddr_0_0_r ? s1_way_wdata_0_0_r : meta_array_17_0; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1724 = 6'h12 == s1_way_waddr_0_0_r ? s1_way_wdata_0_0_r : meta_array_18_0; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1725 = 6'h13 == s1_way_waddr_0_0_r ? s1_way_wdata_0_0_r : meta_array_19_0; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1726 = 6'h14 == s1_way_waddr_0_0_r ? s1_way_wdata_0_0_r : meta_array_20_0; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1727 = 6'h15 == s1_way_waddr_0_0_r ? s1_way_wdata_0_0_r : meta_array_21_0; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1728 = 6'h16 == s1_way_waddr_0_0_r ? s1_way_wdata_0_0_r : meta_array_22_0; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1729 = 6'h17 == s1_way_waddr_0_0_r ? s1_way_wdata_0_0_r : meta_array_23_0; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1730 = 6'h18 == s1_way_waddr_0_0_r ? s1_way_wdata_0_0_r : meta_array_24_0; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1731 = 6'h19 == s1_way_waddr_0_0_r ? s1_way_wdata_0_0_r : meta_array_25_0; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1732 = 6'h1a == s1_way_waddr_0_0_r ? s1_way_wdata_0_0_r : meta_array_26_0; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1733 = 6'h1b == s1_way_waddr_0_0_r ? s1_way_wdata_0_0_r : meta_array_27_0; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1734 = 6'h1c == s1_way_waddr_0_0_r ? s1_way_wdata_0_0_r : meta_array_28_0; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1735 = 6'h1d == s1_way_waddr_0_0_r ? s1_way_wdata_0_0_r : meta_array_29_0; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1736 = 6'h1e == s1_way_waddr_0_0_r ? s1_way_wdata_0_0_r : meta_array_30_0; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1737 = 6'h1f == s1_way_waddr_0_0_r ? s1_way_wdata_0_0_r : meta_array_31_0; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1738 = 6'h20 == s1_way_waddr_0_0_r ? s1_way_wdata_0_0_r : meta_array_32_0; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1739 = 6'h21 == s1_way_waddr_0_0_r ? s1_way_wdata_0_0_r : meta_array_33_0; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1740 = 6'h22 == s1_way_waddr_0_0_r ? s1_way_wdata_0_0_r : meta_array_34_0; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1741 = 6'h23 == s1_way_waddr_0_0_r ? s1_way_wdata_0_0_r : meta_array_35_0; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1742 = 6'h24 == s1_way_waddr_0_0_r ? s1_way_wdata_0_0_r : meta_array_36_0; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1743 = 6'h25 == s1_way_waddr_0_0_r ? s1_way_wdata_0_0_r : meta_array_37_0; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1744 = 6'h26 == s1_way_waddr_0_0_r ? s1_way_wdata_0_0_r : meta_array_38_0; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1745 = 6'h27 == s1_way_waddr_0_0_r ? s1_way_wdata_0_0_r : meta_array_39_0; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1746 = 6'h28 == s1_way_waddr_0_0_r ? s1_way_wdata_0_0_r : meta_array_40_0; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1747 = 6'h29 == s1_way_waddr_0_0_r ? s1_way_wdata_0_0_r : meta_array_41_0; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1748 = 6'h2a == s1_way_waddr_0_0_r ? s1_way_wdata_0_0_r : meta_array_42_0; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1749 = 6'h2b == s1_way_waddr_0_0_r ? s1_way_wdata_0_0_r : meta_array_43_0; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1750 = 6'h2c == s1_way_waddr_0_0_r ? s1_way_wdata_0_0_r : meta_array_44_0; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1751 = 6'h2d == s1_way_waddr_0_0_r ? s1_way_wdata_0_0_r : meta_array_45_0; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1752 = 6'h2e == s1_way_waddr_0_0_r ? s1_way_wdata_0_0_r : meta_array_46_0; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1753 = 6'h2f == s1_way_waddr_0_0_r ? s1_way_wdata_0_0_r : meta_array_47_0; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1754 = 6'h30 == s1_way_waddr_0_0_r ? s1_way_wdata_0_0_r : meta_array_48_0; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1755 = 6'h31 == s1_way_waddr_0_0_r ? s1_way_wdata_0_0_r : meta_array_49_0; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1756 = 6'h32 == s1_way_waddr_0_0_r ? s1_way_wdata_0_0_r : meta_array_50_0; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1757 = 6'h33 == s1_way_waddr_0_0_r ? s1_way_wdata_0_0_r : meta_array_51_0; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1758 = 6'h34 == s1_way_waddr_0_0_r ? s1_way_wdata_0_0_r : meta_array_52_0; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1759 = 6'h35 == s1_way_waddr_0_0_r ? s1_way_wdata_0_0_r : meta_array_53_0; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1760 = 6'h36 == s1_way_waddr_0_0_r ? s1_way_wdata_0_0_r : meta_array_54_0; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1761 = 6'h37 == s1_way_waddr_0_0_r ? s1_way_wdata_0_0_r : meta_array_55_0; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1762 = 6'h38 == s1_way_waddr_0_0_r ? s1_way_wdata_0_0_r : meta_array_56_0; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1763 = 6'h39 == s1_way_waddr_0_0_r ? s1_way_wdata_0_0_r : meta_array_57_0; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1764 = 6'h3a == s1_way_waddr_0_0_r ? s1_way_wdata_0_0_r : meta_array_58_0; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1765 = 6'h3b == s1_way_waddr_0_0_r ? s1_way_wdata_0_0_r : meta_array_59_0; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1766 = 6'h3c == s1_way_waddr_0_0_r ? s1_way_wdata_0_0_r : meta_array_60_0; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1767 = 6'h3d == s1_way_waddr_0_0_r ? s1_way_wdata_0_0_r : meta_array_61_0; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1768 = 6'h3e == s1_way_waddr_0_0_r ? s1_way_wdata_0_0_r : meta_array_62_0; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1769 = 6'h3f == s1_way_waddr_0_0_r ? s1_way_wdata_0_0_r : meta_array_63_0; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1770 = s1_way_wen_0_0_REG ? _GEN_1706 : meta_array_0_0; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1771 = s1_way_wen_0_0_REG ? _GEN_1707 : meta_array_1_0; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1772 = s1_way_wen_0_0_REG ? _GEN_1708 : meta_array_2_0; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1773 = s1_way_wen_0_0_REG ? _GEN_1709 : meta_array_3_0; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1774 = s1_way_wen_0_0_REG ? _GEN_1710 : meta_array_4_0; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1775 = s1_way_wen_0_0_REG ? _GEN_1711 : meta_array_5_0; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1776 = s1_way_wen_0_0_REG ? _GEN_1712 : meta_array_6_0; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1777 = s1_way_wen_0_0_REG ? _GEN_1713 : meta_array_7_0; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1778 = s1_way_wen_0_0_REG ? _GEN_1714 : meta_array_8_0; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1779 = s1_way_wen_0_0_REG ? _GEN_1715 : meta_array_9_0; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1780 = s1_way_wen_0_0_REG ? _GEN_1716 : meta_array_10_0; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1781 = s1_way_wen_0_0_REG ? _GEN_1717 : meta_array_11_0; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1782 = s1_way_wen_0_0_REG ? _GEN_1718 : meta_array_12_0; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1783 = s1_way_wen_0_0_REG ? _GEN_1719 : meta_array_13_0; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1784 = s1_way_wen_0_0_REG ? _GEN_1720 : meta_array_14_0; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1785 = s1_way_wen_0_0_REG ? _GEN_1721 : meta_array_15_0; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1786 = s1_way_wen_0_0_REG ? _GEN_1722 : meta_array_16_0; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1787 = s1_way_wen_0_0_REG ? _GEN_1723 : meta_array_17_0; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1788 = s1_way_wen_0_0_REG ? _GEN_1724 : meta_array_18_0; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1789 = s1_way_wen_0_0_REG ? _GEN_1725 : meta_array_19_0; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1790 = s1_way_wen_0_0_REG ? _GEN_1726 : meta_array_20_0; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1791 = s1_way_wen_0_0_REG ? _GEN_1727 : meta_array_21_0; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1792 = s1_way_wen_0_0_REG ? _GEN_1728 : meta_array_22_0; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1793 = s1_way_wen_0_0_REG ? _GEN_1729 : meta_array_23_0; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1794 = s1_way_wen_0_0_REG ? _GEN_1730 : meta_array_24_0; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1795 = s1_way_wen_0_0_REG ? _GEN_1731 : meta_array_25_0; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1796 = s1_way_wen_0_0_REG ? _GEN_1732 : meta_array_26_0; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1797 = s1_way_wen_0_0_REG ? _GEN_1733 : meta_array_27_0; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1798 = s1_way_wen_0_0_REG ? _GEN_1734 : meta_array_28_0; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1799 = s1_way_wen_0_0_REG ? _GEN_1735 : meta_array_29_0; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1800 = s1_way_wen_0_0_REG ? _GEN_1736 : meta_array_30_0; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1801 = s1_way_wen_0_0_REG ? _GEN_1737 : meta_array_31_0; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1802 = s1_way_wen_0_0_REG ? _GEN_1738 : meta_array_32_0; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1803 = s1_way_wen_0_0_REG ? _GEN_1739 : meta_array_33_0; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1804 = s1_way_wen_0_0_REG ? _GEN_1740 : meta_array_34_0; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1805 = s1_way_wen_0_0_REG ? _GEN_1741 : meta_array_35_0; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1806 = s1_way_wen_0_0_REG ? _GEN_1742 : meta_array_36_0; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1807 = s1_way_wen_0_0_REG ? _GEN_1743 : meta_array_37_0; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1808 = s1_way_wen_0_0_REG ? _GEN_1744 : meta_array_38_0; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1809 = s1_way_wen_0_0_REG ? _GEN_1745 : meta_array_39_0; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1810 = s1_way_wen_0_0_REG ? _GEN_1746 : meta_array_40_0; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1811 = s1_way_wen_0_0_REG ? _GEN_1747 : meta_array_41_0; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1812 = s1_way_wen_0_0_REG ? _GEN_1748 : meta_array_42_0; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1813 = s1_way_wen_0_0_REG ? _GEN_1749 : meta_array_43_0; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1814 = s1_way_wen_0_0_REG ? _GEN_1750 : meta_array_44_0; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1815 = s1_way_wen_0_0_REG ? _GEN_1751 : meta_array_45_0; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1816 = s1_way_wen_0_0_REG ? _GEN_1752 : meta_array_46_0; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1817 = s1_way_wen_0_0_REG ? _GEN_1753 : meta_array_47_0; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1818 = s1_way_wen_0_0_REG ? _GEN_1754 : meta_array_48_0; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1819 = s1_way_wen_0_0_REG ? _GEN_1755 : meta_array_49_0; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1820 = s1_way_wen_0_0_REG ? _GEN_1756 : meta_array_50_0; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1821 = s1_way_wen_0_0_REG ? _GEN_1757 : meta_array_51_0; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1822 = s1_way_wen_0_0_REG ? _GEN_1758 : meta_array_52_0; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1823 = s1_way_wen_0_0_REG ? _GEN_1759 : meta_array_53_0; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1824 = s1_way_wen_0_0_REG ? _GEN_1760 : meta_array_54_0; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1825 = s1_way_wen_0_0_REG ? _GEN_1761 : meta_array_55_0; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1826 = s1_way_wen_0_0_REG ? _GEN_1762 : meta_array_56_0; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1827 = s1_way_wen_0_0_REG ? _GEN_1763 : meta_array_57_0; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1828 = s1_way_wen_0_0_REG ? _GEN_1764 : meta_array_58_0; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1829 = s1_way_wen_0_0_REG ? _GEN_1765 : meta_array_59_0; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1830 = s1_way_wen_0_0_REG ? _GEN_1766 : meta_array_60_0; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1831 = s1_way_wen_0_0_REG ? _GEN_1767 : meta_array_61_0; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1832 = s1_way_wen_0_0_REG ? _GEN_1768 : meta_array_62_0; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1833 = s1_way_wen_0_0_REG ? _GEN_1769 : meta_array_63_0; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  s0_way_wen_1_0 = io_write_0_valid & io_write_0_bits_way_en[1]; // @[AsynchronousMetaArray.scala 152:49]
  wire  _GEN_1836 = 6'h0 == s1_way_waddr_1_0_r ? s1_way_wdata_1_0_r : meta_array_0_1; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1837 = 6'h1 == s1_way_waddr_1_0_r ? s1_way_wdata_1_0_r : meta_array_1_1; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1838 = 6'h2 == s1_way_waddr_1_0_r ? s1_way_wdata_1_0_r : meta_array_2_1; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1839 = 6'h3 == s1_way_waddr_1_0_r ? s1_way_wdata_1_0_r : meta_array_3_1; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1840 = 6'h4 == s1_way_waddr_1_0_r ? s1_way_wdata_1_0_r : meta_array_4_1; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1841 = 6'h5 == s1_way_waddr_1_0_r ? s1_way_wdata_1_0_r : meta_array_5_1; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1842 = 6'h6 == s1_way_waddr_1_0_r ? s1_way_wdata_1_0_r : meta_array_6_1; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1843 = 6'h7 == s1_way_waddr_1_0_r ? s1_way_wdata_1_0_r : meta_array_7_1; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1844 = 6'h8 == s1_way_waddr_1_0_r ? s1_way_wdata_1_0_r : meta_array_8_1; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1845 = 6'h9 == s1_way_waddr_1_0_r ? s1_way_wdata_1_0_r : meta_array_9_1; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1846 = 6'ha == s1_way_waddr_1_0_r ? s1_way_wdata_1_0_r : meta_array_10_1; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1847 = 6'hb == s1_way_waddr_1_0_r ? s1_way_wdata_1_0_r : meta_array_11_1; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1848 = 6'hc == s1_way_waddr_1_0_r ? s1_way_wdata_1_0_r : meta_array_12_1; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1849 = 6'hd == s1_way_waddr_1_0_r ? s1_way_wdata_1_0_r : meta_array_13_1; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1850 = 6'he == s1_way_waddr_1_0_r ? s1_way_wdata_1_0_r : meta_array_14_1; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1851 = 6'hf == s1_way_waddr_1_0_r ? s1_way_wdata_1_0_r : meta_array_15_1; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1852 = 6'h10 == s1_way_waddr_1_0_r ? s1_way_wdata_1_0_r : meta_array_16_1; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1853 = 6'h11 == s1_way_waddr_1_0_r ? s1_way_wdata_1_0_r : meta_array_17_1; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1854 = 6'h12 == s1_way_waddr_1_0_r ? s1_way_wdata_1_0_r : meta_array_18_1; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1855 = 6'h13 == s1_way_waddr_1_0_r ? s1_way_wdata_1_0_r : meta_array_19_1; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1856 = 6'h14 == s1_way_waddr_1_0_r ? s1_way_wdata_1_0_r : meta_array_20_1; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1857 = 6'h15 == s1_way_waddr_1_0_r ? s1_way_wdata_1_0_r : meta_array_21_1; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1858 = 6'h16 == s1_way_waddr_1_0_r ? s1_way_wdata_1_0_r : meta_array_22_1; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1859 = 6'h17 == s1_way_waddr_1_0_r ? s1_way_wdata_1_0_r : meta_array_23_1; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1860 = 6'h18 == s1_way_waddr_1_0_r ? s1_way_wdata_1_0_r : meta_array_24_1; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1861 = 6'h19 == s1_way_waddr_1_0_r ? s1_way_wdata_1_0_r : meta_array_25_1; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1862 = 6'h1a == s1_way_waddr_1_0_r ? s1_way_wdata_1_0_r : meta_array_26_1; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1863 = 6'h1b == s1_way_waddr_1_0_r ? s1_way_wdata_1_0_r : meta_array_27_1; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1864 = 6'h1c == s1_way_waddr_1_0_r ? s1_way_wdata_1_0_r : meta_array_28_1; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1865 = 6'h1d == s1_way_waddr_1_0_r ? s1_way_wdata_1_0_r : meta_array_29_1; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1866 = 6'h1e == s1_way_waddr_1_0_r ? s1_way_wdata_1_0_r : meta_array_30_1; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1867 = 6'h1f == s1_way_waddr_1_0_r ? s1_way_wdata_1_0_r : meta_array_31_1; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1868 = 6'h20 == s1_way_waddr_1_0_r ? s1_way_wdata_1_0_r : meta_array_32_1; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1869 = 6'h21 == s1_way_waddr_1_0_r ? s1_way_wdata_1_0_r : meta_array_33_1; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1870 = 6'h22 == s1_way_waddr_1_0_r ? s1_way_wdata_1_0_r : meta_array_34_1; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1871 = 6'h23 == s1_way_waddr_1_0_r ? s1_way_wdata_1_0_r : meta_array_35_1; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1872 = 6'h24 == s1_way_waddr_1_0_r ? s1_way_wdata_1_0_r : meta_array_36_1; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1873 = 6'h25 == s1_way_waddr_1_0_r ? s1_way_wdata_1_0_r : meta_array_37_1; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1874 = 6'h26 == s1_way_waddr_1_0_r ? s1_way_wdata_1_0_r : meta_array_38_1; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1875 = 6'h27 == s1_way_waddr_1_0_r ? s1_way_wdata_1_0_r : meta_array_39_1; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1876 = 6'h28 == s1_way_waddr_1_0_r ? s1_way_wdata_1_0_r : meta_array_40_1; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1877 = 6'h29 == s1_way_waddr_1_0_r ? s1_way_wdata_1_0_r : meta_array_41_1; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1878 = 6'h2a == s1_way_waddr_1_0_r ? s1_way_wdata_1_0_r : meta_array_42_1; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1879 = 6'h2b == s1_way_waddr_1_0_r ? s1_way_wdata_1_0_r : meta_array_43_1; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1880 = 6'h2c == s1_way_waddr_1_0_r ? s1_way_wdata_1_0_r : meta_array_44_1; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1881 = 6'h2d == s1_way_waddr_1_0_r ? s1_way_wdata_1_0_r : meta_array_45_1; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1882 = 6'h2e == s1_way_waddr_1_0_r ? s1_way_wdata_1_0_r : meta_array_46_1; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1883 = 6'h2f == s1_way_waddr_1_0_r ? s1_way_wdata_1_0_r : meta_array_47_1; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1884 = 6'h30 == s1_way_waddr_1_0_r ? s1_way_wdata_1_0_r : meta_array_48_1; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1885 = 6'h31 == s1_way_waddr_1_0_r ? s1_way_wdata_1_0_r : meta_array_49_1; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1886 = 6'h32 == s1_way_waddr_1_0_r ? s1_way_wdata_1_0_r : meta_array_50_1; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1887 = 6'h33 == s1_way_waddr_1_0_r ? s1_way_wdata_1_0_r : meta_array_51_1; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1888 = 6'h34 == s1_way_waddr_1_0_r ? s1_way_wdata_1_0_r : meta_array_52_1; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1889 = 6'h35 == s1_way_waddr_1_0_r ? s1_way_wdata_1_0_r : meta_array_53_1; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1890 = 6'h36 == s1_way_waddr_1_0_r ? s1_way_wdata_1_0_r : meta_array_54_1; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1891 = 6'h37 == s1_way_waddr_1_0_r ? s1_way_wdata_1_0_r : meta_array_55_1; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1892 = 6'h38 == s1_way_waddr_1_0_r ? s1_way_wdata_1_0_r : meta_array_56_1; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1893 = 6'h39 == s1_way_waddr_1_0_r ? s1_way_wdata_1_0_r : meta_array_57_1; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1894 = 6'h3a == s1_way_waddr_1_0_r ? s1_way_wdata_1_0_r : meta_array_58_1; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1895 = 6'h3b == s1_way_waddr_1_0_r ? s1_way_wdata_1_0_r : meta_array_59_1; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1896 = 6'h3c == s1_way_waddr_1_0_r ? s1_way_wdata_1_0_r : meta_array_60_1; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1897 = 6'h3d == s1_way_waddr_1_0_r ? s1_way_wdata_1_0_r : meta_array_61_1; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1898 = 6'h3e == s1_way_waddr_1_0_r ? s1_way_wdata_1_0_r : meta_array_62_1; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1899 = 6'h3f == s1_way_waddr_1_0_r ? s1_way_wdata_1_0_r : meta_array_63_1; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1900 = s1_way_wen_1_0_REG ? _GEN_1836 : meta_array_0_1; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1901 = s1_way_wen_1_0_REG ? _GEN_1837 : meta_array_1_1; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1902 = s1_way_wen_1_0_REG ? _GEN_1838 : meta_array_2_1; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1903 = s1_way_wen_1_0_REG ? _GEN_1839 : meta_array_3_1; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1904 = s1_way_wen_1_0_REG ? _GEN_1840 : meta_array_4_1; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1905 = s1_way_wen_1_0_REG ? _GEN_1841 : meta_array_5_1; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1906 = s1_way_wen_1_0_REG ? _GEN_1842 : meta_array_6_1; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1907 = s1_way_wen_1_0_REG ? _GEN_1843 : meta_array_7_1; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1908 = s1_way_wen_1_0_REG ? _GEN_1844 : meta_array_8_1; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1909 = s1_way_wen_1_0_REG ? _GEN_1845 : meta_array_9_1; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1910 = s1_way_wen_1_0_REG ? _GEN_1846 : meta_array_10_1; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1911 = s1_way_wen_1_0_REG ? _GEN_1847 : meta_array_11_1; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1912 = s1_way_wen_1_0_REG ? _GEN_1848 : meta_array_12_1; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1913 = s1_way_wen_1_0_REG ? _GEN_1849 : meta_array_13_1; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1914 = s1_way_wen_1_0_REG ? _GEN_1850 : meta_array_14_1; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1915 = s1_way_wen_1_0_REG ? _GEN_1851 : meta_array_15_1; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1916 = s1_way_wen_1_0_REG ? _GEN_1852 : meta_array_16_1; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1917 = s1_way_wen_1_0_REG ? _GEN_1853 : meta_array_17_1; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1918 = s1_way_wen_1_0_REG ? _GEN_1854 : meta_array_18_1; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1919 = s1_way_wen_1_0_REG ? _GEN_1855 : meta_array_19_1; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1920 = s1_way_wen_1_0_REG ? _GEN_1856 : meta_array_20_1; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1921 = s1_way_wen_1_0_REG ? _GEN_1857 : meta_array_21_1; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1922 = s1_way_wen_1_0_REG ? _GEN_1858 : meta_array_22_1; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1923 = s1_way_wen_1_0_REG ? _GEN_1859 : meta_array_23_1; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1924 = s1_way_wen_1_0_REG ? _GEN_1860 : meta_array_24_1; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1925 = s1_way_wen_1_0_REG ? _GEN_1861 : meta_array_25_1; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1926 = s1_way_wen_1_0_REG ? _GEN_1862 : meta_array_26_1; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1927 = s1_way_wen_1_0_REG ? _GEN_1863 : meta_array_27_1; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1928 = s1_way_wen_1_0_REG ? _GEN_1864 : meta_array_28_1; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1929 = s1_way_wen_1_0_REG ? _GEN_1865 : meta_array_29_1; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1930 = s1_way_wen_1_0_REG ? _GEN_1866 : meta_array_30_1; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1931 = s1_way_wen_1_0_REG ? _GEN_1867 : meta_array_31_1; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1932 = s1_way_wen_1_0_REG ? _GEN_1868 : meta_array_32_1; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1933 = s1_way_wen_1_0_REG ? _GEN_1869 : meta_array_33_1; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1934 = s1_way_wen_1_0_REG ? _GEN_1870 : meta_array_34_1; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1935 = s1_way_wen_1_0_REG ? _GEN_1871 : meta_array_35_1; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1936 = s1_way_wen_1_0_REG ? _GEN_1872 : meta_array_36_1; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1937 = s1_way_wen_1_0_REG ? _GEN_1873 : meta_array_37_1; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1938 = s1_way_wen_1_0_REG ? _GEN_1874 : meta_array_38_1; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1939 = s1_way_wen_1_0_REG ? _GEN_1875 : meta_array_39_1; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1940 = s1_way_wen_1_0_REG ? _GEN_1876 : meta_array_40_1; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1941 = s1_way_wen_1_0_REG ? _GEN_1877 : meta_array_41_1; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1942 = s1_way_wen_1_0_REG ? _GEN_1878 : meta_array_42_1; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1943 = s1_way_wen_1_0_REG ? _GEN_1879 : meta_array_43_1; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1944 = s1_way_wen_1_0_REG ? _GEN_1880 : meta_array_44_1; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1945 = s1_way_wen_1_0_REG ? _GEN_1881 : meta_array_45_1; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1946 = s1_way_wen_1_0_REG ? _GEN_1882 : meta_array_46_1; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1947 = s1_way_wen_1_0_REG ? _GEN_1883 : meta_array_47_1; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1948 = s1_way_wen_1_0_REG ? _GEN_1884 : meta_array_48_1; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1949 = s1_way_wen_1_0_REG ? _GEN_1885 : meta_array_49_1; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1950 = s1_way_wen_1_0_REG ? _GEN_1886 : meta_array_50_1; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1951 = s1_way_wen_1_0_REG ? _GEN_1887 : meta_array_51_1; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1952 = s1_way_wen_1_0_REG ? _GEN_1888 : meta_array_52_1; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1953 = s1_way_wen_1_0_REG ? _GEN_1889 : meta_array_53_1; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1954 = s1_way_wen_1_0_REG ? _GEN_1890 : meta_array_54_1; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1955 = s1_way_wen_1_0_REG ? _GEN_1891 : meta_array_55_1; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1956 = s1_way_wen_1_0_REG ? _GEN_1892 : meta_array_56_1; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1957 = s1_way_wen_1_0_REG ? _GEN_1893 : meta_array_57_1; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1958 = s1_way_wen_1_0_REG ? _GEN_1894 : meta_array_58_1; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1959 = s1_way_wen_1_0_REG ? _GEN_1895 : meta_array_59_1; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1960 = s1_way_wen_1_0_REG ? _GEN_1896 : meta_array_60_1; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1961 = s1_way_wen_1_0_REG ? _GEN_1897 : meta_array_61_1; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1962 = s1_way_wen_1_0_REG ? _GEN_1898 : meta_array_62_1; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_1963 = s1_way_wen_1_0_REG ? _GEN_1899 : meta_array_63_1; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  s0_way_wen_2_0 = io_write_0_valid & io_write_0_bits_way_en[2]; // @[AsynchronousMetaArray.scala 152:49]
  wire  _GEN_1966 = 6'h0 == s1_way_waddr_2_0_r ? s1_way_wdata_2_0_r : meta_array_0_2; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1967 = 6'h1 == s1_way_waddr_2_0_r ? s1_way_wdata_2_0_r : meta_array_1_2; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1968 = 6'h2 == s1_way_waddr_2_0_r ? s1_way_wdata_2_0_r : meta_array_2_2; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1969 = 6'h3 == s1_way_waddr_2_0_r ? s1_way_wdata_2_0_r : meta_array_3_2; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1970 = 6'h4 == s1_way_waddr_2_0_r ? s1_way_wdata_2_0_r : meta_array_4_2; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1971 = 6'h5 == s1_way_waddr_2_0_r ? s1_way_wdata_2_0_r : meta_array_5_2; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1972 = 6'h6 == s1_way_waddr_2_0_r ? s1_way_wdata_2_0_r : meta_array_6_2; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1973 = 6'h7 == s1_way_waddr_2_0_r ? s1_way_wdata_2_0_r : meta_array_7_2; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1974 = 6'h8 == s1_way_waddr_2_0_r ? s1_way_wdata_2_0_r : meta_array_8_2; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1975 = 6'h9 == s1_way_waddr_2_0_r ? s1_way_wdata_2_0_r : meta_array_9_2; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1976 = 6'ha == s1_way_waddr_2_0_r ? s1_way_wdata_2_0_r : meta_array_10_2; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1977 = 6'hb == s1_way_waddr_2_0_r ? s1_way_wdata_2_0_r : meta_array_11_2; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1978 = 6'hc == s1_way_waddr_2_0_r ? s1_way_wdata_2_0_r : meta_array_12_2; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1979 = 6'hd == s1_way_waddr_2_0_r ? s1_way_wdata_2_0_r : meta_array_13_2; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1980 = 6'he == s1_way_waddr_2_0_r ? s1_way_wdata_2_0_r : meta_array_14_2; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1981 = 6'hf == s1_way_waddr_2_0_r ? s1_way_wdata_2_0_r : meta_array_15_2; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1982 = 6'h10 == s1_way_waddr_2_0_r ? s1_way_wdata_2_0_r : meta_array_16_2; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1983 = 6'h11 == s1_way_waddr_2_0_r ? s1_way_wdata_2_0_r : meta_array_17_2; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1984 = 6'h12 == s1_way_waddr_2_0_r ? s1_way_wdata_2_0_r : meta_array_18_2; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1985 = 6'h13 == s1_way_waddr_2_0_r ? s1_way_wdata_2_0_r : meta_array_19_2; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1986 = 6'h14 == s1_way_waddr_2_0_r ? s1_way_wdata_2_0_r : meta_array_20_2; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1987 = 6'h15 == s1_way_waddr_2_0_r ? s1_way_wdata_2_0_r : meta_array_21_2; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1988 = 6'h16 == s1_way_waddr_2_0_r ? s1_way_wdata_2_0_r : meta_array_22_2; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1989 = 6'h17 == s1_way_waddr_2_0_r ? s1_way_wdata_2_0_r : meta_array_23_2; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1990 = 6'h18 == s1_way_waddr_2_0_r ? s1_way_wdata_2_0_r : meta_array_24_2; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1991 = 6'h19 == s1_way_waddr_2_0_r ? s1_way_wdata_2_0_r : meta_array_25_2; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1992 = 6'h1a == s1_way_waddr_2_0_r ? s1_way_wdata_2_0_r : meta_array_26_2; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1993 = 6'h1b == s1_way_waddr_2_0_r ? s1_way_wdata_2_0_r : meta_array_27_2; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1994 = 6'h1c == s1_way_waddr_2_0_r ? s1_way_wdata_2_0_r : meta_array_28_2; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1995 = 6'h1d == s1_way_waddr_2_0_r ? s1_way_wdata_2_0_r : meta_array_29_2; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1996 = 6'h1e == s1_way_waddr_2_0_r ? s1_way_wdata_2_0_r : meta_array_30_2; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1997 = 6'h1f == s1_way_waddr_2_0_r ? s1_way_wdata_2_0_r : meta_array_31_2; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1998 = 6'h20 == s1_way_waddr_2_0_r ? s1_way_wdata_2_0_r : meta_array_32_2; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_1999 = 6'h21 == s1_way_waddr_2_0_r ? s1_way_wdata_2_0_r : meta_array_33_2; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2000 = 6'h22 == s1_way_waddr_2_0_r ? s1_way_wdata_2_0_r : meta_array_34_2; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2001 = 6'h23 == s1_way_waddr_2_0_r ? s1_way_wdata_2_0_r : meta_array_35_2; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2002 = 6'h24 == s1_way_waddr_2_0_r ? s1_way_wdata_2_0_r : meta_array_36_2; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2003 = 6'h25 == s1_way_waddr_2_0_r ? s1_way_wdata_2_0_r : meta_array_37_2; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2004 = 6'h26 == s1_way_waddr_2_0_r ? s1_way_wdata_2_0_r : meta_array_38_2; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2005 = 6'h27 == s1_way_waddr_2_0_r ? s1_way_wdata_2_0_r : meta_array_39_2; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2006 = 6'h28 == s1_way_waddr_2_0_r ? s1_way_wdata_2_0_r : meta_array_40_2; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2007 = 6'h29 == s1_way_waddr_2_0_r ? s1_way_wdata_2_0_r : meta_array_41_2; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2008 = 6'h2a == s1_way_waddr_2_0_r ? s1_way_wdata_2_0_r : meta_array_42_2; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2009 = 6'h2b == s1_way_waddr_2_0_r ? s1_way_wdata_2_0_r : meta_array_43_2; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2010 = 6'h2c == s1_way_waddr_2_0_r ? s1_way_wdata_2_0_r : meta_array_44_2; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2011 = 6'h2d == s1_way_waddr_2_0_r ? s1_way_wdata_2_0_r : meta_array_45_2; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2012 = 6'h2e == s1_way_waddr_2_0_r ? s1_way_wdata_2_0_r : meta_array_46_2; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2013 = 6'h2f == s1_way_waddr_2_0_r ? s1_way_wdata_2_0_r : meta_array_47_2; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2014 = 6'h30 == s1_way_waddr_2_0_r ? s1_way_wdata_2_0_r : meta_array_48_2; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2015 = 6'h31 == s1_way_waddr_2_0_r ? s1_way_wdata_2_0_r : meta_array_49_2; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2016 = 6'h32 == s1_way_waddr_2_0_r ? s1_way_wdata_2_0_r : meta_array_50_2; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2017 = 6'h33 == s1_way_waddr_2_0_r ? s1_way_wdata_2_0_r : meta_array_51_2; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2018 = 6'h34 == s1_way_waddr_2_0_r ? s1_way_wdata_2_0_r : meta_array_52_2; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2019 = 6'h35 == s1_way_waddr_2_0_r ? s1_way_wdata_2_0_r : meta_array_53_2; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2020 = 6'h36 == s1_way_waddr_2_0_r ? s1_way_wdata_2_0_r : meta_array_54_2; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2021 = 6'h37 == s1_way_waddr_2_0_r ? s1_way_wdata_2_0_r : meta_array_55_2; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2022 = 6'h38 == s1_way_waddr_2_0_r ? s1_way_wdata_2_0_r : meta_array_56_2; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2023 = 6'h39 == s1_way_waddr_2_0_r ? s1_way_wdata_2_0_r : meta_array_57_2; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2024 = 6'h3a == s1_way_waddr_2_0_r ? s1_way_wdata_2_0_r : meta_array_58_2; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2025 = 6'h3b == s1_way_waddr_2_0_r ? s1_way_wdata_2_0_r : meta_array_59_2; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2026 = 6'h3c == s1_way_waddr_2_0_r ? s1_way_wdata_2_0_r : meta_array_60_2; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2027 = 6'h3d == s1_way_waddr_2_0_r ? s1_way_wdata_2_0_r : meta_array_61_2; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2028 = 6'h3e == s1_way_waddr_2_0_r ? s1_way_wdata_2_0_r : meta_array_62_2; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2029 = 6'h3f == s1_way_waddr_2_0_r ? s1_way_wdata_2_0_r : meta_array_63_2; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2030 = s1_way_wen_2_0_REG ? _GEN_1966 : meta_array_0_2; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2031 = s1_way_wen_2_0_REG ? _GEN_1967 : meta_array_1_2; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2032 = s1_way_wen_2_0_REG ? _GEN_1968 : meta_array_2_2; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2033 = s1_way_wen_2_0_REG ? _GEN_1969 : meta_array_3_2; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2034 = s1_way_wen_2_0_REG ? _GEN_1970 : meta_array_4_2; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2035 = s1_way_wen_2_0_REG ? _GEN_1971 : meta_array_5_2; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2036 = s1_way_wen_2_0_REG ? _GEN_1972 : meta_array_6_2; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2037 = s1_way_wen_2_0_REG ? _GEN_1973 : meta_array_7_2; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2038 = s1_way_wen_2_0_REG ? _GEN_1974 : meta_array_8_2; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2039 = s1_way_wen_2_0_REG ? _GEN_1975 : meta_array_9_2; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2040 = s1_way_wen_2_0_REG ? _GEN_1976 : meta_array_10_2; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2041 = s1_way_wen_2_0_REG ? _GEN_1977 : meta_array_11_2; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2042 = s1_way_wen_2_0_REG ? _GEN_1978 : meta_array_12_2; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2043 = s1_way_wen_2_0_REG ? _GEN_1979 : meta_array_13_2; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2044 = s1_way_wen_2_0_REG ? _GEN_1980 : meta_array_14_2; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2045 = s1_way_wen_2_0_REG ? _GEN_1981 : meta_array_15_2; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2046 = s1_way_wen_2_0_REG ? _GEN_1982 : meta_array_16_2; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2047 = s1_way_wen_2_0_REG ? _GEN_1983 : meta_array_17_2; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2048 = s1_way_wen_2_0_REG ? _GEN_1984 : meta_array_18_2; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2049 = s1_way_wen_2_0_REG ? _GEN_1985 : meta_array_19_2; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2050 = s1_way_wen_2_0_REG ? _GEN_1986 : meta_array_20_2; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2051 = s1_way_wen_2_0_REG ? _GEN_1987 : meta_array_21_2; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2052 = s1_way_wen_2_0_REG ? _GEN_1988 : meta_array_22_2; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2053 = s1_way_wen_2_0_REG ? _GEN_1989 : meta_array_23_2; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2054 = s1_way_wen_2_0_REG ? _GEN_1990 : meta_array_24_2; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2055 = s1_way_wen_2_0_REG ? _GEN_1991 : meta_array_25_2; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2056 = s1_way_wen_2_0_REG ? _GEN_1992 : meta_array_26_2; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2057 = s1_way_wen_2_0_REG ? _GEN_1993 : meta_array_27_2; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2058 = s1_way_wen_2_0_REG ? _GEN_1994 : meta_array_28_2; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2059 = s1_way_wen_2_0_REG ? _GEN_1995 : meta_array_29_2; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2060 = s1_way_wen_2_0_REG ? _GEN_1996 : meta_array_30_2; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2061 = s1_way_wen_2_0_REG ? _GEN_1997 : meta_array_31_2; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2062 = s1_way_wen_2_0_REG ? _GEN_1998 : meta_array_32_2; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2063 = s1_way_wen_2_0_REG ? _GEN_1999 : meta_array_33_2; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2064 = s1_way_wen_2_0_REG ? _GEN_2000 : meta_array_34_2; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2065 = s1_way_wen_2_0_REG ? _GEN_2001 : meta_array_35_2; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2066 = s1_way_wen_2_0_REG ? _GEN_2002 : meta_array_36_2; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2067 = s1_way_wen_2_0_REG ? _GEN_2003 : meta_array_37_2; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2068 = s1_way_wen_2_0_REG ? _GEN_2004 : meta_array_38_2; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2069 = s1_way_wen_2_0_REG ? _GEN_2005 : meta_array_39_2; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2070 = s1_way_wen_2_0_REG ? _GEN_2006 : meta_array_40_2; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2071 = s1_way_wen_2_0_REG ? _GEN_2007 : meta_array_41_2; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2072 = s1_way_wen_2_0_REG ? _GEN_2008 : meta_array_42_2; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2073 = s1_way_wen_2_0_REG ? _GEN_2009 : meta_array_43_2; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2074 = s1_way_wen_2_0_REG ? _GEN_2010 : meta_array_44_2; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2075 = s1_way_wen_2_0_REG ? _GEN_2011 : meta_array_45_2; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2076 = s1_way_wen_2_0_REG ? _GEN_2012 : meta_array_46_2; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2077 = s1_way_wen_2_0_REG ? _GEN_2013 : meta_array_47_2; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2078 = s1_way_wen_2_0_REG ? _GEN_2014 : meta_array_48_2; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2079 = s1_way_wen_2_0_REG ? _GEN_2015 : meta_array_49_2; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2080 = s1_way_wen_2_0_REG ? _GEN_2016 : meta_array_50_2; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2081 = s1_way_wen_2_0_REG ? _GEN_2017 : meta_array_51_2; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2082 = s1_way_wen_2_0_REG ? _GEN_2018 : meta_array_52_2; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2083 = s1_way_wen_2_0_REG ? _GEN_2019 : meta_array_53_2; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2084 = s1_way_wen_2_0_REG ? _GEN_2020 : meta_array_54_2; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2085 = s1_way_wen_2_0_REG ? _GEN_2021 : meta_array_55_2; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2086 = s1_way_wen_2_0_REG ? _GEN_2022 : meta_array_56_2; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2087 = s1_way_wen_2_0_REG ? _GEN_2023 : meta_array_57_2; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2088 = s1_way_wen_2_0_REG ? _GEN_2024 : meta_array_58_2; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2089 = s1_way_wen_2_0_REG ? _GEN_2025 : meta_array_59_2; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2090 = s1_way_wen_2_0_REG ? _GEN_2026 : meta_array_60_2; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2091 = s1_way_wen_2_0_REG ? _GEN_2027 : meta_array_61_2; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2092 = s1_way_wen_2_0_REG ? _GEN_2028 : meta_array_62_2; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2093 = s1_way_wen_2_0_REG ? _GEN_2029 : meta_array_63_2; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  s0_way_wen_3_0 = io_write_0_valid & io_write_0_bits_way_en[3]; // @[AsynchronousMetaArray.scala 152:49]
  wire  _GEN_2096 = 6'h0 == s1_way_waddr_3_0_r ? s1_way_wdata_3_0_r : meta_array_0_3; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2097 = 6'h1 == s1_way_waddr_3_0_r ? s1_way_wdata_3_0_r : meta_array_1_3; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2098 = 6'h2 == s1_way_waddr_3_0_r ? s1_way_wdata_3_0_r : meta_array_2_3; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2099 = 6'h3 == s1_way_waddr_3_0_r ? s1_way_wdata_3_0_r : meta_array_3_3; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2100 = 6'h4 == s1_way_waddr_3_0_r ? s1_way_wdata_3_0_r : meta_array_4_3; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2101 = 6'h5 == s1_way_waddr_3_0_r ? s1_way_wdata_3_0_r : meta_array_5_3; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2102 = 6'h6 == s1_way_waddr_3_0_r ? s1_way_wdata_3_0_r : meta_array_6_3; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2103 = 6'h7 == s1_way_waddr_3_0_r ? s1_way_wdata_3_0_r : meta_array_7_3; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2104 = 6'h8 == s1_way_waddr_3_0_r ? s1_way_wdata_3_0_r : meta_array_8_3; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2105 = 6'h9 == s1_way_waddr_3_0_r ? s1_way_wdata_3_0_r : meta_array_9_3; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2106 = 6'ha == s1_way_waddr_3_0_r ? s1_way_wdata_3_0_r : meta_array_10_3; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2107 = 6'hb == s1_way_waddr_3_0_r ? s1_way_wdata_3_0_r : meta_array_11_3; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2108 = 6'hc == s1_way_waddr_3_0_r ? s1_way_wdata_3_0_r : meta_array_12_3; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2109 = 6'hd == s1_way_waddr_3_0_r ? s1_way_wdata_3_0_r : meta_array_13_3; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2110 = 6'he == s1_way_waddr_3_0_r ? s1_way_wdata_3_0_r : meta_array_14_3; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2111 = 6'hf == s1_way_waddr_3_0_r ? s1_way_wdata_3_0_r : meta_array_15_3; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2112 = 6'h10 == s1_way_waddr_3_0_r ? s1_way_wdata_3_0_r : meta_array_16_3; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2113 = 6'h11 == s1_way_waddr_3_0_r ? s1_way_wdata_3_0_r : meta_array_17_3; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2114 = 6'h12 == s1_way_waddr_3_0_r ? s1_way_wdata_3_0_r : meta_array_18_3; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2115 = 6'h13 == s1_way_waddr_3_0_r ? s1_way_wdata_3_0_r : meta_array_19_3; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2116 = 6'h14 == s1_way_waddr_3_0_r ? s1_way_wdata_3_0_r : meta_array_20_3; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2117 = 6'h15 == s1_way_waddr_3_0_r ? s1_way_wdata_3_0_r : meta_array_21_3; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2118 = 6'h16 == s1_way_waddr_3_0_r ? s1_way_wdata_3_0_r : meta_array_22_3; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2119 = 6'h17 == s1_way_waddr_3_0_r ? s1_way_wdata_3_0_r : meta_array_23_3; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2120 = 6'h18 == s1_way_waddr_3_0_r ? s1_way_wdata_3_0_r : meta_array_24_3; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2121 = 6'h19 == s1_way_waddr_3_0_r ? s1_way_wdata_3_0_r : meta_array_25_3; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2122 = 6'h1a == s1_way_waddr_3_0_r ? s1_way_wdata_3_0_r : meta_array_26_3; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2123 = 6'h1b == s1_way_waddr_3_0_r ? s1_way_wdata_3_0_r : meta_array_27_3; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2124 = 6'h1c == s1_way_waddr_3_0_r ? s1_way_wdata_3_0_r : meta_array_28_3; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2125 = 6'h1d == s1_way_waddr_3_0_r ? s1_way_wdata_3_0_r : meta_array_29_3; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2126 = 6'h1e == s1_way_waddr_3_0_r ? s1_way_wdata_3_0_r : meta_array_30_3; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2127 = 6'h1f == s1_way_waddr_3_0_r ? s1_way_wdata_3_0_r : meta_array_31_3; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2128 = 6'h20 == s1_way_waddr_3_0_r ? s1_way_wdata_3_0_r : meta_array_32_3; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2129 = 6'h21 == s1_way_waddr_3_0_r ? s1_way_wdata_3_0_r : meta_array_33_3; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2130 = 6'h22 == s1_way_waddr_3_0_r ? s1_way_wdata_3_0_r : meta_array_34_3; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2131 = 6'h23 == s1_way_waddr_3_0_r ? s1_way_wdata_3_0_r : meta_array_35_3; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2132 = 6'h24 == s1_way_waddr_3_0_r ? s1_way_wdata_3_0_r : meta_array_36_3; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2133 = 6'h25 == s1_way_waddr_3_0_r ? s1_way_wdata_3_0_r : meta_array_37_3; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2134 = 6'h26 == s1_way_waddr_3_0_r ? s1_way_wdata_3_0_r : meta_array_38_3; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2135 = 6'h27 == s1_way_waddr_3_0_r ? s1_way_wdata_3_0_r : meta_array_39_3; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2136 = 6'h28 == s1_way_waddr_3_0_r ? s1_way_wdata_3_0_r : meta_array_40_3; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2137 = 6'h29 == s1_way_waddr_3_0_r ? s1_way_wdata_3_0_r : meta_array_41_3; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2138 = 6'h2a == s1_way_waddr_3_0_r ? s1_way_wdata_3_0_r : meta_array_42_3; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2139 = 6'h2b == s1_way_waddr_3_0_r ? s1_way_wdata_3_0_r : meta_array_43_3; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2140 = 6'h2c == s1_way_waddr_3_0_r ? s1_way_wdata_3_0_r : meta_array_44_3; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2141 = 6'h2d == s1_way_waddr_3_0_r ? s1_way_wdata_3_0_r : meta_array_45_3; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2142 = 6'h2e == s1_way_waddr_3_0_r ? s1_way_wdata_3_0_r : meta_array_46_3; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2143 = 6'h2f == s1_way_waddr_3_0_r ? s1_way_wdata_3_0_r : meta_array_47_3; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2144 = 6'h30 == s1_way_waddr_3_0_r ? s1_way_wdata_3_0_r : meta_array_48_3; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2145 = 6'h31 == s1_way_waddr_3_0_r ? s1_way_wdata_3_0_r : meta_array_49_3; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2146 = 6'h32 == s1_way_waddr_3_0_r ? s1_way_wdata_3_0_r : meta_array_50_3; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2147 = 6'h33 == s1_way_waddr_3_0_r ? s1_way_wdata_3_0_r : meta_array_51_3; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2148 = 6'h34 == s1_way_waddr_3_0_r ? s1_way_wdata_3_0_r : meta_array_52_3; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2149 = 6'h35 == s1_way_waddr_3_0_r ? s1_way_wdata_3_0_r : meta_array_53_3; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2150 = 6'h36 == s1_way_waddr_3_0_r ? s1_way_wdata_3_0_r : meta_array_54_3; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2151 = 6'h37 == s1_way_waddr_3_0_r ? s1_way_wdata_3_0_r : meta_array_55_3; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2152 = 6'h38 == s1_way_waddr_3_0_r ? s1_way_wdata_3_0_r : meta_array_56_3; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2153 = 6'h39 == s1_way_waddr_3_0_r ? s1_way_wdata_3_0_r : meta_array_57_3; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2154 = 6'h3a == s1_way_waddr_3_0_r ? s1_way_wdata_3_0_r : meta_array_58_3; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2155 = 6'h3b == s1_way_waddr_3_0_r ? s1_way_wdata_3_0_r : meta_array_59_3; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2156 = 6'h3c == s1_way_waddr_3_0_r ? s1_way_wdata_3_0_r : meta_array_60_3; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2157 = 6'h3d == s1_way_waddr_3_0_r ? s1_way_wdata_3_0_r : meta_array_61_3; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2158 = 6'h3e == s1_way_waddr_3_0_r ? s1_way_wdata_3_0_r : meta_array_62_3; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2159 = 6'h3f == s1_way_waddr_3_0_r ? s1_way_wdata_3_0_r : meta_array_63_3; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2160 = s1_way_wen_3_0_REG ? _GEN_2096 : meta_array_0_3; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2161 = s1_way_wen_3_0_REG ? _GEN_2097 : meta_array_1_3; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2162 = s1_way_wen_3_0_REG ? _GEN_2098 : meta_array_2_3; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2163 = s1_way_wen_3_0_REG ? _GEN_2099 : meta_array_3_3; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2164 = s1_way_wen_3_0_REG ? _GEN_2100 : meta_array_4_3; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2165 = s1_way_wen_3_0_REG ? _GEN_2101 : meta_array_5_3; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2166 = s1_way_wen_3_0_REG ? _GEN_2102 : meta_array_6_3; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2167 = s1_way_wen_3_0_REG ? _GEN_2103 : meta_array_7_3; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2168 = s1_way_wen_3_0_REG ? _GEN_2104 : meta_array_8_3; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2169 = s1_way_wen_3_0_REG ? _GEN_2105 : meta_array_9_3; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2170 = s1_way_wen_3_0_REG ? _GEN_2106 : meta_array_10_3; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2171 = s1_way_wen_3_0_REG ? _GEN_2107 : meta_array_11_3; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2172 = s1_way_wen_3_0_REG ? _GEN_2108 : meta_array_12_3; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2173 = s1_way_wen_3_0_REG ? _GEN_2109 : meta_array_13_3; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2174 = s1_way_wen_3_0_REG ? _GEN_2110 : meta_array_14_3; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2175 = s1_way_wen_3_0_REG ? _GEN_2111 : meta_array_15_3; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2176 = s1_way_wen_3_0_REG ? _GEN_2112 : meta_array_16_3; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2177 = s1_way_wen_3_0_REG ? _GEN_2113 : meta_array_17_3; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2178 = s1_way_wen_3_0_REG ? _GEN_2114 : meta_array_18_3; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2179 = s1_way_wen_3_0_REG ? _GEN_2115 : meta_array_19_3; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2180 = s1_way_wen_3_0_REG ? _GEN_2116 : meta_array_20_3; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2181 = s1_way_wen_3_0_REG ? _GEN_2117 : meta_array_21_3; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2182 = s1_way_wen_3_0_REG ? _GEN_2118 : meta_array_22_3; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2183 = s1_way_wen_3_0_REG ? _GEN_2119 : meta_array_23_3; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2184 = s1_way_wen_3_0_REG ? _GEN_2120 : meta_array_24_3; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2185 = s1_way_wen_3_0_REG ? _GEN_2121 : meta_array_25_3; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2186 = s1_way_wen_3_0_REG ? _GEN_2122 : meta_array_26_3; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2187 = s1_way_wen_3_0_REG ? _GEN_2123 : meta_array_27_3; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2188 = s1_way_wen_3_0_REG ? _GEN_2124 : meta_array_28_3; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2189 = s1_way_wen_3_0_REG ? _GEN_2125 : meta_array_29_3; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2190 = s1_way_wen_3_0_REG ? _GEN_2126 : meta_array_30_3; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2191 = s1_way_wen_3_0_REG ? _GEN_2127 : meta_array_31_3; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2192 = s1_way_wen_3_0_REG ? _GEN_2128 : meta_array_32_3; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2193 = s1_way_wen_3_0_REG ? _GEN_2129 : meta_array_33_3; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2194 = s1_way_wen_3_0_REG ? _GEN_2130 : meta_array_34_3; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2195 = s1_way_wen_3_0_REG ? _GEN_2131 : meta_array_35_3; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2196 = s1_way_wen_3_0_REG ? _GEN_2132 : meta_array_36_3; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2197 = s1_way_wen_3_0_REG ? _GEN_2133 : meta_array_37_3; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2198 = s1_way_wen_3_0_REG ? _GEN_2134 : meta_array_38_3; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2199 = s1_way_wen_3_0_REG ? _GEN_2135 : meta_array_39_3; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2200 = s1_way_wen_3_0_REG ? _GEN_2136 : meta_array_40_3; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2201 = s1_way_wen_3_0_REG ? _GEN_2137 : meta_array_41_3; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2202 = s1_way_wen_3_0_REG ? _GEN_2138 : meta_array_42_3; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2203 = s1_way_wen_3_0_REG ? _GEN_2139 : meta_array_43_3; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2204 = s1_way_wen_3_0_REG ? _GEN_2140 : meta_array_44_3; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2205 = s1_way_wen_3_0_REG ? _GEN_2141 : meta_array_45_3; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2206 = s1_way_wen_3_0_REG ? _GEN_2142 : meta_array_46_3; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2207 = s1_way_wen_3_0_REG ? _GEN_2143 : meta_array_47_3; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2208 = s1_way_wen_3_0_REG ? _GEN_2144 : meta_array_48_3; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2209 = s1_way_wen_3_0_REG ? _GEN_2145 : meta_array_49_3; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2210 = s1_way_wen_3_0_REG ? _GEN_2146 : meta_array_50_3; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2211 = s1_way_wen_3_0_REG ? _GEN_2147 : meta_array_51_3; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2212 = s1_way_wen_3_0_REG ? _GEN_2148 : meta_array_52_3; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2213 = s1_way_wen_3_0_REG ? _GEN_2149 : meta_array_53_3; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2214 = s1_way_wen_3_0_REG ? _GEN_2150 : meta_array_54_3; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2215 = s1_way_wen_3_0_REG ? _GEN_2151 : meta_array_55_3; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2216 = s1_way_wen_3_0_REG ? _GEN_2152 : meta_array_56_3; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2217 = s1_way_wen_3_0_REG ? _GEN_2153 : meta_array_57_3; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2218 = s1_way_wen_3_0_REG ? _GEN_2154 : meta_array_58_3; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2219 = s1_way_wen_3_0_REG ? _GEN_2155 : meta_array_59_3; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2220 = s1_way_wen_3_0_REG ? _GEN_2156 : meta_array_60_3; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2221 = s1_way_wen_3_0_REG ? _GEN_2157 : meta_array_61_3; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2222 = s1_way_wen_3_0_REG ? _GEN_2158 : meta_array_62_3; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2223 = s1_way_wen_3_0_REG ? _GEN_2159 : meta_array_63_3; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  s0_way_wen_4_0 = io_write_0_valid & io_write_0_bits_way_en[4]; // @[AsynchronousMetaArray.scala 152:49]
  wire  _GEN_2226 = 6'h0 == s1_way_waddr_4_0_r ? s1_way_wdata_4_0_r : meta_array_0_4; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2227 = 6'h1 == s1_way_waddr_4_0_r ? s1_way_wdata_4_0_r : meta_array_1_4; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2228 = 6'h2 == s1_way_waddr_4_0_r ? s1_way_wdata_4_0_r : meta_array_2_4; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2229 = 6'h3 == s1_way_waddr_4_0_r ? s1_way_wdata_4_0_r : meta_array_3_4; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2230 = 6'h4 == s1_way_waddr_4_0_r ? s1_way_wdata_4_0_r : meta_array_4_4; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2231 = 6'h5 == s1_way_waddr_4_0_r ? s1_way_wdata_4_0_r : meta_array_5_4; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2232 = 6'h6 == s1_way_waddr_4_0_r ? s1_way_wdata_4_0_r : meta_array_6_4; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2233 = 6'h7 == s1_way_waddr_4_0_r ? s1_way_wdata_4_0_r : meta_array_7_4; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2234 = 6'h8 == s1_way_waddr_4_0_r ? s1_way_wdata_4_0_r : meta_array_8_4; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2235 = 6'h9 == s1_way_waddr_4_0_r ? s1_way_wdata_4_0_r : meta_array_9_4; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2236 = 6'ha == s1_way_waddr_4_0_r ? s1_way_wdata_4_0_r : meta_array_10_4; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2237 = 6'hb == s1_way_waddr_4_0_r ? s1_way_wdata_4_0_r : meta_array_11_4; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2238 = 6'hc == s1_way_waddr_4_0_r ? s1_way_wdata_4_0_r : meta_array_12_4; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2239 = 6'hd == s1_way_waddr_4_0_r ? s1_way_wdata_4_0_r : meta_array_13_4; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2240 = 6'he == s1_way_waddr_4_0_r ? s1_way_wdata_4_0_r : meta_array_14_4; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2241 = 6'hf == s1_way_waddr_4_0_r ? s1_way_wdata_4_0_r : meta_array_15_4; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2242 = 6'h10 == s1_way_waddr_4_0_r ? s1_way_wdata_4_0_r : meta_array_16_4; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2243 = 6'h11 == s1_way_waddr_4_0_r ? s1_way_wdata_4_0_r : meta_array_17_4; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2244 = 6'h12 == s1_way_waddr_4_0_r ? s1_way_wdata_4_0_r : meta_array_18_4; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2245 = 6'h13 == s1_way_waddr_4_0_r ? s1_way_wdata_4_0_r : meta_array_19_4; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2246 = 6'h14 == s1_way_waddr_4_0_r ? s1_way_wdata_4_0_r : meta_array_20_4; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2247 = 6'h15 == s1_way_waddr_4_0_r ? s1_way_wdata_4_0_r : meta_array_21_4; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2248 = 6'h16 == s1_way_waddr_4_0_r ? s1_way_wdata_4_0_r : meta_array_22_4; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2249 = 6'h17 == s1_way_waddr_4_0_r ? s1_way_wdata_4_0_r : meta_array_23_4; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2250 = 6'h18 == s1_way_waddr_4_0_r ? s1_way_wdata_4_0_r : meta_array_24_4; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2251 = 6'h19 == s1_way_waddr_4_0_r ? s1_way_wdata_4_0_r : meta_array_25_4; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2252 = 6'h1a == s1_way_waddr_4_0_r ? s1_way_wdata_4_0_r : meta_array_26_4; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2253 = 6'h1b == s1_way_waddr_4_0_r ? s1_way_wdata_4_0_r : meta_array_27_4; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2254 = 6'h1c == s1_way_waddr_4_0_r ? s1_way_wdata_4_0_r : meta_array_28_4; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2255 = 6'h1d == s1_way_waddr_4_0_r ? s1_way_wdata_4_0_r : meta_array_29_4; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2256 = 6'h1e == s1_way_waddr_4_0_r ? s1_way_wdata_4_0_r : meta_array_30_4; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2257 = 6'h1f == s1_way_waddr_4_0_r ? s1_way_wdata_4_0_r : meta_array_31_4; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2258 = 6'h20 == s1_way_waddr_4_0_r ? s1_way_wdata_4_0_r : meta_array_32_4; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2259 = 6'h21 == s1_way_waddr_4_0_r ? s1_way_wdata_4_0_r : meta_array_33_4; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2260 = 6'h22 == s1_way_waddr_4_0_r ? s1_way_wdata_4_0_r : meta_array_34_4; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2261 = 6'h23 == s1_way_waddr_4_0_r ? s1_way_wdata_4_0_r : meta_array_35_4; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2262 = 6'h24 == s1_way_waddr_4_0_r ? s1_way_wdata_4_0_r : meta_array_36_4; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2263 = 6'h25 == s1_way_waddr_4_0_r ? s1_way_wdata_4_0_r : meta_array_37_4; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2264 = 6'h26 == s1_way_waddr_4_0_r ? s1_way_wdata_4_0_r : meta_array_38_4; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2265 = 6'h27 == s1_way_waddr_4_0_r ? s1_way_wdata_4_0_r : meta_array_39_4; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2266 = 6'h28 == s1_way_waddr_4_0_r ? s1_way_wdata_4_0_r : meta_array_40_4; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2267 = 6'h29 == s1_way_waddr_4_0_r ? s1_way_wdata_4_0_r : meta_array_41_4; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2268 = 6'h2a == s1_way_waddr_4_0_r ? s1_way_wdata_4_0_r : meta_array_42_4; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2269 = 6'h2b == s1_way_waddr_4_0_r ? s1_way_wdata_4_0_r : meta_array_43_4; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2270 = 6'h2c == s1_way_waddr_4_0_r ? s1_way_wdata_4_0_r : meta_array_44_4; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2271 = 6'h2d == s1_way_waddr_4_0_r ? s1_way_wdata_4_0_r : meta_array_45_4; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2272 = 6'h2e == s1_way_waddr_4_0_r ? s1_way_wdata_4_0_r : meta_array_46_4; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2273 = 6'h2f == s1_way_waddr_4_0_r ? s1_way_wdata_4_0_r : meta_array_47_4; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2274 = 6'h30 == s1_way_waddr_4_0_r ? s1_way_wdata_4_0_r : meta_array_48_4; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2275 = 6'h31 == s1_way_waddr_4_0_r ? s1_way_wdata_4_0_r : meta_array_49_4; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2276 = 6'h32 == s1_way_waddr_4_0_r ? s1_way_wdata_4_0_r : meta_array_50_4; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2277 = 6'h33 == s1_way_waddr_4_0_r ? s1_way_wdata_4_0_r : meta_array_51_4; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2278 = 6'h34 == s1_way_waddr_4_0_r ? s1_way_wdata_4_0_r : meta_array_52_4; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2279 = 6'h35 == s1_way_waddr_4_0_r ? s1_way_wdata_4_0_r : meta_array_53_4; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2280 = 6'h36 == s1_way_waddr_4_0_r ? s1_way_wdata_4_0_r : meta_array_54_4; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2281 = 6'h37 == s1_way_waddr_4_0_r ? s1_way_wdata_4_0_r : meta_array_55_4; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2282 = 6'h38 == s1_way_waddr_4_0_r ? s1_way_wdata_4_0_r : meta_array_56_4; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2283 = 6'h39 == s1_way_waddr_4_0_r ? s1_way_wdata_4_0_r : meta_array_57_4; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2284 = 6'h3a == s1_way_waddr_4_0_r ? s1_way_wdata_4_0_r : meta_array_58_4; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2285 = 6'h3b == s1_way_waddr_4_0_r ? s1_way_wdata_4_0_r : meta_array_59_4; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2286 = 6'h3c == s1_way_waddr_4_0_r ? s1_way_wdata_4_0_r : meta_array_60_4; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2287 = 6'h3d == s1_way_waddr_4_0_r ? s1_way_wdata_4_0_r : meta_array_61_4; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2288 = 6'h3e == s1_way_waddr_4_0_r ? s1_way_wdata_4_0_r : meta_array_62_4; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2289 = 6'h3f == s1_way_waddr_4_0_r ? s1_way_wdata_4_0_r : meta_array_63_4; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2290 = s1_way_wen_4_0_REG ? _GEN_2226 : meta_array_0_4; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2291 = s1_way_wen_4_0_REG ? _GEN_2227 : meta_array_1_4; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2292 = s1_way_wen_4_0_REG ? _GEN_2228 : meta_array_2_4; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2293 = s1_way_wen_4_0_REG ? _GEN_2229 : meta_array_3_4; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2294 = s1_way_wen_4_0_REG ? _GEN_2230 : meta_array_4_4; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2295 = s1_way_wen_4_0_REG ? _GEN_2231 : meta_array_5_4; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2296 = s1_way_wen_4_0_REG ? _GEN_2232 : meta_array_6_4; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2297 = s1_way_wen_4_0_REG ? _GEN_2233 : meta_array_7_4; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2298 = s1_way_wen_4_0_REG ? _GEN_2234 : meta_array_8_4; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2299 = s1_way_wen_4_0_REG ? _GEN_2235 : meta_array_9_4; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2300 = s1_way_wen_4_0_REG ? _GEN_2236 : meta_array_10_4; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2301 = s1_way_wen_4_0_REG ? _GEN_2237 : meta_array_11_4; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2302 = s1_way_wen_4_0_REG ? _GEN_2238 : meta_array_12_4; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2303 = s1_way_wen_4_0_REG ? _GEN_2239 : meta_array_13_4; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2304 = s1_way_wen_4_0_REG ? _GEN_2240 : meta_array_14_4; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2305 = s1_way_wen_4_0_REG ? _GEN_2241 : meta_array_15_4; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2306 = s1_way_wen_4_0_REG ? _GEN_2242 : meta_array_16_4; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2307 = s1_way_wen_4_0_REG ? _GEN_2243 : meta_array_17_4; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2308 = s1_way_wen_4_0_REG ? _GEN_2244 : meta_array_18_4; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2309 = s1_way_wen_4_0_REG ? _GEN_2245 : meta_array_19_4; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2310 = s1_way_wen_4_0_REG ? _GEN_2246 : meta_array_20_4; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2311 = s1_way_wen_4_0_REG ? _GEN_2247 : meta_array_21_4; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2312 = s1_way_wen_4_0_REG ? _GEN_2248 : meta_array_22_4; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2313 = s1_way_wen_4_0_REG ? _GEN_2249 : meta_array_23_4; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2314 = s1_way_wen_4_0_REG ? _GEN_2250 : meta_array_24_4; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2315 = s1_way_wen_4_0_REG ? _GEN_2251 : meta_array_25_4; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2316 = s1_way_wen_4_0_REG ? _GEN_2252 : meta_array_26_4; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2317 = s1_way_wen_4_0_REG ? _GEN_2253 : meta_array_27_4; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2318 = s1_way_wen_4_0_REG ? _GEN_2254 : meta_array_28_4; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2319 = s1_way_wen_4_0_REG ? _GEN_2255 : meta_array_29_4; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2320 = s1_way_wen_4_0_REG ? _GEN_2256 : meta_array_30_4; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2321 = s1_way_wen_4_0_REG ? _GEN_2257 : meta_array_31_4; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2322 = s1_way_wen_4_0_REG ? _GEN_2258 : meta_array_32_4; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2323 = s1_way_wen_4_0_REG ? _GEN_2259 : meta_array_33_4; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2324 = s1_way_wen_4_0_REG ? _GEN_2260 : meta_array_34_4; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2325 = s1_way_wen_4_0_REG ? _GEN_2261 : meta_array_35_4; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2326 = s1_way_wen_4_0_REG ? _GEN_2262 : meta_array_36_4; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2327 = s1_way_wen_4_0_REG ? _GEN_2263 : meta_array_37_4; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2328 = s1_way_wen_4_0_REG ? _GEN_2264 : meta_array_38_4; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2329 = s1_way_wen_4_0_REG ? _GEN_2265 : meta_array_39_4; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2330 = s1_way_wen_4_0_REG ? _GEN_2266 : meta_array_40_4; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2331 = s1_way_wen_4_0_REG ? _GEN_2267 : meta_array_41_4; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2332 = s1_way_wen_4_0_REG ? _GEN_2268 : meta_array_42_4; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2333 = s1_way_wen_4_0_REG ? _GEN_2269 : meta_array_43_4; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2334 = s1_way_wen_4_0_REG ? _GEN_2270 : meta_array_44_4; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2335 = s1_way_wen_4_0_REG ? _GEN_2271 : meta_array_45_4; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2336 = s1_way_wen_4_0_REG ? _GEN_2272 : meta_array_46_4; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2337 = s1_way_wen_4_0_REG ? _GEN_2273 : meta_array_47_4; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2338 = s1_way_wen_4_0_REG ? _GEN_2274 : meta_array_48_4; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2339 = s1_way_wen_4_0_REG ? _GEN_2275 : meta_array_49_4; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2340 = s1_way_wen_4_0_REG ? _GEN_2276 : meta_array_50_4; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2341 = s1_way_wen_4_0_REG ? _GEN_2277 : meta_array_51_4; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2342 = s1_way_wen_4_0_REG ? _GEN_2278 : meta_array_52_4; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2343 = s1_way_wen_4_0_REG ? _GEN_2279 : meta_array_53_4; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2344 = s1_way_wen_4_0_REG ? _GEN_2280 : meta_array_54_4; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2345 = s1_way_wen_4_0_REG ? _GEN_2281 : meta_array_55_4; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2346 = s1_way_wen_4_0_REG ? _GEN_2282 : meta_array_56_4; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2347 = s1_way_wen_4_0_REG ? _GEN_2283 : meta_array_57_4; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2348 = s1_way_wen_4_0_REG ? _GEN_2284 : meta_array_58_4; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2349 = s1_way_wen_4_0_REG ? _GEN_2285 : meta_array_59_4; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2350 = s1_way_wen_4_0_REG ? _GEN_2286 : meta_array_60_4; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2351 = s1_way_wen_4_0_REG ? _GEN_2287 : meta_array_61_4; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2352 = s1_way_wen_4_0_REG ? _GEN_2288 : meta_array_62_4; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2353 = s1_way_wen_4_0_REG ? _GEN_2289 : meta_array_63_4; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  s0_way_wen_5_0 = io_write_0_valid & io_write_0_bits_way_en[5]; // @[AsynchronousMetaArray.scala 152:49]
  wire  _GEN_2356 = 6'h0 == s1_way_waddr_5_0_r ? s1_way_wdata_5_0_r : meta_array_0_5; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2357 = 6'h1 == s1_way_waddr_5_0_r ? s1_way_wdata_5_0_r : meta_array_1_5; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2358 = 6'h2 == s1_way_waddr_5_0_r ? s1_way_wdata_5_0_r : meta_array_2_5; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2359 = 6'h3 == s1_way_waddr_5_0_r ? s1_way_wdata_5_0_r : meta_array_3_5; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2360 = 6'h4 == s1_way_waddr_5_0_r ? s1_way_wdata_5_0_r : meta_array_4_5; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2361 = 6'h5 == s1_way_waddr_5_0_r ? s1_way_wdata_5_0_r : meta_array_5_5; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2362 = 6'h6 == s1_way_waddr_5_0_r ? s1_way_wdata_5_0_r : meta_array_6_5; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2363 = 6'h7 == s1_way_waddr_5_0_r ? s1_way_wdata_5_0_r : meta_array_7_5; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2364 = 6'h8 == s1_way_waddr_5_0_r ? s1_way_wdata_5_0_r : meta_array_8_5; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2365 = 6'h9 == s1_way_waddr_5_0_r ? s1_way_wdata_5_0_r : meta_array_9_5; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2366 = 6'ha == s1_way_waddr_5_0_r ? s1_way_wdata_5_0_r : meta_array_10_5; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2367 = 6'hb == s1_way_waddr_5_0_r ? s1_way_wdata_5_0_r : meta_array_11_5; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2368 = 6'hc == s1_way_waddr_5_0_r ? s1_way_wdata_5_0_r : meta_array_12_5; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2369 = 6'hd == s1_way_waddr_5_0_r ? s1_way_wdata_5_0_r : meta_array_13_5; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2370 = 6'he == s1_way_waddr_5_0_r ? s1_way_wdata_5_0_r : meta_array_14_5; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2371 = 6'hf == s1_way_waddr_5_0_r ? s1_way_wdata_5_0_r : meta_array_15_5; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2372 = 6'h10 == s1_way_waddr_5_0_r ? s1_way_wdata_5_0_r : meta_array_16_5; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2373 = 6'h11 == s1_way_waddr_5_0_r ? s1_way_wdata_5_0_r : meta_array_17_5; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2374 = 6'h12 == s1_way_waddr_5_0_r ? s1_way_wdata_5_0_r : meta_array_18_5; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2375 = 6'h13 == s1_way_waddr_5_0_r ? s1_way_wdata_5_0_r : meta_array_19_5; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2376 = 6'h14 == s1_way_waddr_5_0_r ? s1_way_wdata_5_0_r : meta_array_20_5; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2377 = 6'h15 == s1_way_waddr_5_0_r ? s1_way_wdata_5_0_r : meta_array_21_5; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2378 = 6'h16 == s1_way_waddr_5_0_r ? s1_way_wdata_5_0_r : meta_array_22_5; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2379 = 6'h17 == s1_way_waddr_5_0_r ? s1_way_wdata_5_0_r : meta_array_23_5; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2380 = 6'h18 == s1_way_waddr_5_0_r ? s1_way_wdata_5_0_r : meta_array_24_5; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2381 = 6'h19 == s1_way_waddr_5_0_r ? s1_way_wdata_5_0_r : meta_array_25_5; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2382 = 6'h1a == s1_way_waddr_5_0_r ? s1_way_wdata_5_0_r : meta_array_26_5; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2383 = 6'h1b == s1_way_waddr_5_0_r ? s1_way_wdata_5_0_r : meta_array_27_5; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2384 = 6'h1c == s1_way_waddr_5_0_r ? s1_way_wdata_5_0_r : meta_array_28_5; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2385 = 6'h1d == s1_way_waddr_5_0_r ? s1_way_wdata_5_0_r : meta_array_29_5; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2386 = 6'h1e == s1_way_waddr_5_0_r ? s1_way_wdata_5_0_r : meta_array_30_5; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2387 = 6'h1f == s1_way_waddr_5_0_r ? s1_way_wdata_5_0_r : meta_array_31_5; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2388 = 6'h20 == s1_way_waddr_5_0_r ? s1_way_wdata_5_0_r : meta_array_32_5; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2389 = 6'h21 == s1_way_waddr_5_0_r ? s1_way_wdata_5_0_r : meta_array_33_5; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2390 = 6'h22 == s1_way_waddr_5_0_r ? s1_way_wdata_5_0_r : meta_array_34_5; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2391 = 6'h23 == s1_way_waddr_5_0_r ? s1_way_wdata_5_0_r : meta_array_35_5; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2392 = 6'h24 == s1_way_waddr_5_0_r ? s1_way_wdata_5_0_r : meta_array_36_5; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2393 = 6'h25 == s1_way_waddr_5_0_r ? s1_way_wdata_5_0_r : meta_array_37_5; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2394 = 6'h26 == s1_way_waddr_5_0_r ? s1_way_wdata_5_0_r : meta_array_38_5; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2395 = 6'h27 == s1_way_waddr_5_0_r ? s1_way_wdata_5_0_r : meta_array_39_5; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2396 = 6'h28 == s1_way_waddr_5_0_r ? s1_way_wdata_5_0_r : meta_array_40_5; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2397 = 6'h29 == s1_way_waddr_5_0_r ? s1_way_wdata_5_0_r : meta_array_41_5; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2398 = 6'h2a == s1_way_waddr_5_0_r ? s1_way_wdata_5_0_r : meta_array_42_5; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2399 = 6'h2b == s1_way_waddr_5_0_r ? s1_way_wdata_5_0_r : meta_array_43_5; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2400 = 6'h2c == s1_way_waddr_5_0_r ? s1_way_wdata_5_0_r : meta_array_44_5; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2401 = 6'h2d == s1_way_waddr_5_0_r ? s1_way_wdata_5_0_r : meta_array_45_5; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2402 = 6'h2e == s1_way_waddr_5_0_r ? s1_way_wdata_5_0_r : meta_array_46_5; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2403 = 6'h2f == s1_way_waddr_5_0_r ? s1_way_wdata_5_0_r : meta_array_47_5; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2404 = 6'h30 == s1_way_waddr_5_0_r ? s1_way_wdata_5_0_r : meta_array_48_5; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2405 = 6'h31 == s1_way_waddr_5_0_r ? s1_way_wdata_5_0_r : meta_array_49_5; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2406 = 6'h32 == s1_way_waddr_5_0_r ? s1_way_wdata_5_0_r : meta_array_50_5; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2407 = 6'h33 == s1_way_waddr_5_0_r ? s1_way_wdata_5_0_r : meta_array_51_5; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2408 = 6'h34 == s1_way_waddr_5_0_r ? s1_way_wdata_5_0_r : meta_array_52_5; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2409 = 6'h35 == s1_way_waddr_5_0_r ? s1_way_wdata_5_0_r : meta_array_53_5; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2410 = 6'h36 == s1_way_waddr_5_0_r ? s1_way_wdata_5_0_r : meta_array_54_5; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2411 = 6'h37 == s1_way_waddr_5_0_r ? s1_way_wdata_5_0_r : meta_array_55_5; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2412 = 6'h38 == s1_way_waddr_5_0_r ? s1_way_wdata_5_0_r : meta_array_56_5; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2413 = 6'h39 == s1_way_waddr_5_0_r ? s1_way_wdata_5_0_r : meta_array_57_5; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2414 = 6'h3a == s1_way_waddr_5_0_r ? s1_way_wdata_5_0_r : meta_array_58_5; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2415 = 6'h3b == s1_way_waddr_5_0_r ? s1_way_wdata_5_0_r : meta_array_59_5; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2416 = 6'h3c == s1_way_waddr_5_0_r ? s1_way_wdata_5_0_r : meta_array_60_5; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2417 = 6'h3d == s1_way_waddr_5_0_r ? s1_way_wdata_5_0_r : meta_array_61_5; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2418 = 6'h3e == s1_way_waddr_5_0_r ? s1_way_wdata_5_0_r : meta_array_62_5; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2419 = 6'h3f == s1_way_waddr_5_0_r ? s1_way_wdata_5_0_r : meta_array_63_5; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2420 = s1_way_wen_5_0_REG ? _GEN_2356 : meta_array_0_5; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2421 = s1_way_wen_5_0_REG ? _GEN_2357 : meta_array_1_5; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2422 = s1_way_wen_5_0_REG ? _GEN_2358 : meta_array_2_5; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2423 = s1_way_wen_5_0_REG ? _GEN_2359 : meta_array_3_5; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2424 = s1_way_wen_5_0_REG ? _GEN_2360 : meta_array_4_5; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2425 = s1_way_wen_5_0_REG ? _GEN_2361 : meta_array_5_5; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2426 = s1_way_wen_5_0_REG ? _GEN_2362 : meta_array_6_5; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2427 = s1_way_wen_5_0_REG ? _GEN_2363 : meta_array_7_5; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2428 = s1_way_wen_5_0_REG ? _GEN_2364 : meta_array_8_5; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2429 = s1_way_wen_5_0_REG ? _GEN_2365 : meta_array_9_5; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2430 = s1_way_wen_5_0_REG ? _GEN_2366 : meta_array_10_5; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2431 = s1_way_wen_5_0_REG ? _GEN_2367 : meta_array_11_5; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2432 = s1_way_wen_5_0_REG ? _GEN_2368 : meta_array_12_5; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2433 = s1_way_wen_5_0_REG ? _GEN_2369 : meta_array_13_5; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2434 = s1_way_wen_5_0_REG ? _GEN_2370 : meta_array_14_5; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2435 = s1_way_wen_5_0_REG ? _GEN_2371 : meta_array_15_5; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2436 = s1_way_wen_5_0_REG ? _GEN_2372 : meta_array_16_5; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2437 = s1_way_wen_5_0_REG ? _GEN_2373 : meta_array_17_5; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2438 = s1_way_wen_5_0_REG ? _GEN_2374 : meta_array_18_5; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2439 = s1_way_wen_5_0_REG ? _GEN_2375 : meta_array_19_5; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2440 = s1_way_wen_5_0_REG ? _GEN_2376 : meta_array_20_5; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2441 = s1_way_wen_5_0_REG ? _GEN_2377 : meta_array_21_5; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2442 = s1_way_wen_5_0_REG ? _GEN_2378 : meta_array_22_5; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2443 = s1_way_wen_5_0_REG ? _GEN_2379 : meta_array_23_5; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2444 = s1_way_wen_5_0_REG ? _GEN_2380 : meta_array_24_5; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2445 = s1_way_wen_5_0_REG ? _GEN_2381 : meta_array_25_5; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2446 = s1_way_wen_5_0_REG ? _GEN_2382 : meta_array_26_5; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2447 = s1_way_wen_5_0_REG ? _GEN_2383 : meta_array_27_5; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2448 = s1_way_wen_5_0_REG ? _GEN_2384 : meta_array_28_5; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2449 = s1_way_wen_5_0_REG ? _GEN_2385 : meta_array_29_5; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2450 = s1_way_wen_5_0_REG ? _GEN_2386 : meta_array_30_5; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2451 = s1_way_wen_5_0_REG ? _GEN_2387 : meta_array_31_5; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2452 = s1_way_wen_5_0_REG ? _GEN_2388 : meta_array_32_5; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2453 = s1_way_wen_5_0_REG ? _GEN_2389 : meta_array_33_5; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2454 = s1_way_wen_5_0_REG ? _GEN_2390 : meta_array_34_5; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2455 = s1_way_wen_5_0_REG ? _GEN_2391 : meta_array_35_5; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2456 = s1_way_wen_5_0_REG ? _GEN_2392 : meta_array_36_5; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2457 = s1_way_wen_5_0_REG ? _GEN_2393 : meta_array_37_5; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2458 = s1_way_wen_5_0_REG ? _GEN_2394 : meta_array_38_5; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2459 = s1_way_wen_5_0_REG ? _GEN_2395 : meta_array_39_5; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2460 = s1_way_wen_5_0_REG ? _GEN_2396 : meta_array_40_5; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2461 = s1_way_wen_5_0_REG ? _GEN_2397 : meta_array_41_5; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2462 = s1_way_wen_5_0_REG ? _GEN_2398 : meta_array_42_5; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2463 = s1_way_wen_5_0_REG ? _GEN_2399 : meta_array_43_5; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2464 = s1_way_wen_5_0_REG ? _GEN_2400 : meta_array_44_5; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2465 = s1_way_wen_5_0_REG ? _GEN_2401 : meta_array_45_5; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2466 = s1_way_wen_5_0_REG ? _GEN_2402 : meta_array_46_5; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2467 = s1_way_wen_5_0_REG ? _GEN_2403 : meta_array_47_5; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2468 = s1_way_wen_5_0_REG ? _GEN_2404 : meta_array_48_5; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2469 = s1_way_wen_5_0_REG ? _GEN_2405 : meta_array_49_5; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2470 = s1_way_wen_5_0_REG ? _GEN_2406 : meta_array_50_5; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2471 = s1_way_wen_5_0_REG ? _GEN_2407 : meta_array_51_5; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2472 = s1_way_wen_5_0_REG ? _GEN_2408 : meta_array_52_5; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2473 = s1_way_wen_5_0_REG ? _GEN_2409 : meta_array_53_5; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2474 = s1_way_wen_5_0_REG ? _GEN_2410 : meta_array_54_5; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2475 = s1_way_wen_5_0_REG ? _GEN_2411 : meta_array_55_5; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2476 = s1_way_wen_5_0_REG ? _GEN_2412 : meta_array_56_5; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2477 = s1_way_wen_5_0_REG ? _GEN_2413 : meta_array_57_5; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2478 = s1_way_wen_5_0_REG ? _GEN_2414 : meta_array_58_5; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2479 = s1_way_wen_5_0_REG ? _GEN_2415 : meta_array_59_5; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2480 = s1_way_wen_5_0_REG ? _GEN_2416 : meta_array_60_5; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2481 = s1_way_wen_5_0_REG ? _GEN_2417 : meta_array_61_5; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2482 = s1_way_wen_5_0_REG ? _GEN_2418 : meta_array_62_5; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2483 = s1_way_wen_5_0_REG ? _GEN_2419 : meta_array_63_5; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  s0_way_wen_6_0 = io_write_0_valid & io_write_0_bits_way_en[6]; // @[AsynchronousMetaArray.scala 152:49]
  wire  _GEN_2486 = 6'h0 == s1_way_waddr_6_0_r ? s1_way_wdata_6_0_r : meta_array_0_6; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2487 = 6'h1 == s1_way_waddr_6_0_r ? s1_way_wdata_6_0_r : meta_array_1_6; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2488 = 6'h2 == s1_way_waddr_6_0_r ? s1_way_wdata_6_0_r : meta_array_2_6; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2489 = 6'h3 == s1_way_waddr_6_0_r ? s1_way_wdata_6_0_r : meta_array_3_6; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2490 = 6'h4 == s1_way_waddr_6_0_r ? s1_way_wdata_6_0_r : meta_array_4_6; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2491 = 6'h5 == s1_way_waddr_6_0_r ? s1_way_wdata_6_0_r : meta_array_5_6; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2492 = 6'h6 == s1_way_waddr_6_0_r ? s1_way_wdata_6_0_r : meta_array_6_6; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2493 = 6'h7 == s1_way_waddr_6_0_r ? s1_way_wdata_6_0_r : meta_array_7_6; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2494 = 6'h8 == s1_way_waddr_6_0_r ? s1_way_wdata_6_0_r : meta_array_8_6; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2495 = 6'h9 == s1_way_waddr_6_0_r ? s1_way_wdata_6_0_r : meta_array_9_6; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2496 = 6'ha == s1_way_waddr_6_0_r ? s1_way_wdata_6_0_r : meta_array_10_6; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2497 = 6'hb == s1_way_waddr_6_0_r ? s1_way_wdata_6_0_r : meta_array_11_6; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2498 = 6'hc == s1_way_waddr_6_0_r ? s1_way_wdata_6_0_r : meta_array_12_6; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2499 = 6'hd == s1_way_waddr_6_0_r ? s1_way_wdata_6_0_r : meta_array_13_6; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2500 = 6'he == s1_way_waddr_6_0_r ? s1_way_wdata_6_0_r : meta_array_14_6; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2501 = 6'hf == s1_way_waddr_6_0_r ? s1_way_wdata_6_0_r : meta_array_15_6; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2502 = 6'h10 == s1_way_waddr_6_0_r ? s1_way_wdata_6_0_r : meta_array_16_6; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2503 = 6'h11 == s1_way_waddr_6_0_r ? s1_way_wdata_6_0_r : meta_array_17_6; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2504 = 6'h12 == s1_way_waddr_6_0_r ? s1_way_wdata_6_0_r : meta_array_18_6; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2505 = 6'h13 == s1_way_waddr_6_0_r ? s1_way_wdata_6_0_r : meta_array_19_6; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2506 = 6'h14 == s1_way_waddr_6_0_r ? s1_way_wdata_6_0_r : meta_array_20_6; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2507 = 6'h15 == s1_way_waddr_6_0_r ? s1_way_wdata_6_0_r : meta_array_21_6; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2508 = 6'h16 == s1_way_waddr_6_0_r ? s1_way_wdata_6_0_r : meta_array_22_6; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2509 = 6'h17 == s1_way_waddr_6_0_r ? s1_way_wdata_6_0_r : meta_array_23_6; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2510 = 6'h18 == s1_way_waddr_6_0_r ? s1_way_wdata_6_0_r : meta_array_24_6; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2511 = 6'h19 == s1_way_waddr_6_0_r ? s1_way_wdata_6_0_r : meta_array_25_6; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2512 = 6'h1a == s1_way_waddr_6_0_r ? s1_way_wdata_6_0_r : meta_array_26_6; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2513 = 6'h1b == s1_way_waddr_6_0_r ? s1_way_wdata_6_0_r : meta_array_27_6; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2514 = 6'h1c == s1_way_waddr_6_0_r ? s1_way_wdata_6_0_r : meta_array_28_6; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2515 = 6'h1d == s1_way_waddr_6_0_r ? s1_way_wdata_6_0_r : meta_array_29_6; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2516 = 6'h1e == s1_way_waddr_6_0_r ? s1_way_wdata_6_0_r : meta_array_30_6; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2517 = 6'h1f == s1_way_waddr_6_0_r ? s1_way_wdata_6_0_r : meta_array_31_6; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2518 = 6'h20 == s1_way_waddr_6_0_r ? s1_way_wdata_6_0_r : meta_array_32_6; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2519 = 6'h21 == s1_way_waddr_6_0_r ? s1_way_wdata_6_0_r : meta_array_33_6; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2520 = 6'h22 == s1_way_waddr_6_0_r ? s1_way_wdata_6_0_r : meta_array_34_6; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2521 = 6'h23 == s1_way_waddr_6_0_r ? s1_way_wdata_6_0_r : meta_array_35_6; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2522 = 6'h24 == s1_way_waddr_6_0_r ? s1_way_wdata_6_0_r : meta_array_36_6; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2523 = 6'h25 == s1_way_waddr_6_0_r ? s1_way_wdata_6_0_r : meta_array_37_6; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2524 = 6'h26 == s1_way_waddr_6_0_r ? s1_way_wdata_6_0_r : meta_array_38_6; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2525 = 6'h27 == s1_way_waddr_6_0_r ? s1_way_wdata_6_0_r : meta_array_39_6; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2526 = 6'h28 == s1_way_waddr_6_0_r ? s1_way_wdata_6_0_r : meta_array_40_6; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2527 = 6'h29 == s1_way_waddr_6_0_r ? s1_way_wdata_6_0_r : meta_array_41_6; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2528 = 6'h2a == s1_way_waddr_6_0_r ? s1_way_wdata_6_0_r : meta_array_42_6; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2529 = 6'h2b == s1_way_waddr_6_0_r ? s1_way_wdata_6_0_r : meta_array_43_6; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2530 = 6'h2c == s1_way_waddr_6_0_r ? s1_way_wdata_6_0_r : meta_array_44_6; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2531 = 6'h2d == s1_way_waddr_6_0_r ? s1_way_wdata_6_0_r : meta_array_45_6; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2532 = 6'h2e == s1_way_waddr_6_0_r ? s1_way_wdata_6_0_r : meta_array_46_6; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2533 = 6'h2f == s1_way_waddr_6_0_r ? s1_way_wdata_6_0_r : meta_array_47_6; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2534 = 6'h30 == s1_way_waddr_6_0_r ? s1_way_wdata_6_0_r : meta_array_48_6; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2535 = 6'h31 == s1_way_waddr_6_0_r ? s1_way_wdata_6_0_r : meta_array_49_6; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2536 = 6'h32 == s1_way_waddr_6_0_r ? s1_way_wdata_6_0_r : meta_array_50_6; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2537 = 6'h33 == s1_way_waddr_6_0_r ? s1_way_wdata_6_0_r : meta_array_51_6; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2538 = 6'h34 == s1_way_waddr_6_0_r ? s1_way_wdata_6_0_r : meta_array_52_6; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2539 = 6'h35 == s1_way_waddr_6_0_r ? s1_way_wdata_6_0_r : meta_array_53_6; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2540 = 6'h36 == s1_way_waddr_6_0_r ? s1_way_wdata_6_0_r : meta_array_54_6; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2541 = 6'h37 == s1_way_waddr_6_0_r ? s1_way_wdata_6_0_r : meta_array_55_6; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2542 = 6'h38 == s1_way_waddr_6_0_r ? s1_way_wdata_6_0_r : meta_array_56_6; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2543 = 6'h39 == s1_way_waddr_6_0_r ? s1_way_wdata_6_0_r : meta_array_57_6; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2544 = 6'h3a == s1_way_waddr_6_0_r ? s1_way_wdata_6_0_r : meta_array_58_6; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2545 = 6'h3b == s1_way_waddr_6_0_r ? s1_way_wdata_6_0_r : meta_array_59_6; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2546 = 6'h3c == s1_way_waddr_6_0_r ? s1_way_wdata_6_0_r : meta_array_60_6; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2547 = 6'h3d == s1_way_waddr_6_0_r ? s1_way_wdata_6_0_r : meta_array_61_6; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2548 = 6'h3e == s1_way_waddr_6_0_r ? s1_way_wdata_6_0_r : meta_array_62_6; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2549 = 6'h3f == s1_way_waddr_6_0_r ? s1_way_wdata_6_0_r : meta_array_63_6; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2550 = s1_way_wen_6_0_REG ? _GEN_2486 : meta_array_0_6; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2551 = s1_way_wen_6_0_REG ? _GEN_2487 : meta_array_1_6; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2552 = s1_way_wen_6_0_REG ? _GEN_2488 : meta_array_2_6; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2553 = s1_way_wen_6_0_REG ? _GEN_2489 : meta_array_3_6; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2554 = s1_way_wen_6_0_REG ? _GEN_2490 : meta_array_4_6; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2555 = s1_way_wen_6_0_REG ? _GEN_2491 : meta_array_5_6; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2556 = s1_way_wen_6_0_REG ? _GEN_2492 : meta_array_6_6; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2557 = s1_way_wen_6_0_REG ? _GEN_2493 : meta_array_7_6; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2558 = s1_way_wen_6_0_REG ? _GEN_2494 : meta_array_8_6; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2559 = s1_way_wen_6_0_REG ? _GEN_2495 : meta_array_9_6; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2560 = s1_way_wen_6_0_REG ? _GEN_2496 : meta_array_10_6; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2561 = s1_way_wen_6_0_REG ? _GEN_2497 : meta_array_11_6; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2562 = s1_way_wen_6_0_REG ? _GEN_2498 : meta_array_12_6; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2563 = s1_way_wen_6_0_REG ? _GEN_2499 : meta_array_13_6; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2564 = s1_way_wen_6_0_REG ? _GEN_2500 : meta_array_14_6; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2565 = s1_way_wen_6_0_REG ? _GEN_2501 : meta_array_15_6; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2566 = s1_way_wen_6_0_REG ? _GEN_2502 : meta_array_16_6; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2567 = s1_way_wen_6_0_REG ? _GEN_2503 : meta_array_17_6; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2568 = s1_way_wen_6_0_REG ? _GEN_2504 : meta_array_18_6; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2569 = s1_way_wen_6_0_REG ? _GEN_2505 : meta_array_19_6; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2570 = s1_way_wen_6_0_REG ? _GEN_2506 : meta_array_20_6; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2571 = s1_way_wen_6_0_REG ? _GEN_2507 : meta_array_21_6; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2572 = s1_way_wen_6_0_REG ? _GEN_2508 : meta_array_22_6; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2573 = s1_way_wen_6_0_REG ? _GEN_2509 : meta_array_23_6; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2574 = s1_way_wen_6_0_REG ? _GEN_2510 : meta_array_24_6; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2575 = s1_way_wen_6_0_REG ? _GEN_2511 : meta_array_25_6; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2576 = s1_way_wen_6_0_REG ? _GEN_2512 : meta_array_26_6; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2577 = s1_way_wen_6_0_REG ? _GEN_2513 : meta_array_27_6; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2578 = s1_way_wen_6_0_REG ? _GEN_2514 : meta_array_28_6; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2579 = s1_way_wen_6_0_REG ? _GEN_2515 : meta_array_29_6; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2580 = s1_way_wen_6_0_REG ? _GEN_2516 : meta_array_30_6; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2581 = s1_way_wen_6_0_REG ? _GEN_2517 : meta_array_31_6; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2582 = s1_way_wen_6_0_REG ? _GEN_2518 : meta_array_32_6; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2583 = s1_way_wen_6_0_REG ? _GEN_2519 : meta_array_33_6; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2584 = s1_way_wen_6_0_REG ? _GEN_2520 : meta_array_34_6; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2585 = s1_way_wen_6_0_REG ? _GEN_2521 : meta_array_35_6; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2586 = s1_way_wen_6_0_REG ? _GEN_2522 : meta_array_36_6; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2587 = s1_way_wen_6_0_REG ? _GEN_2523 : meta_array_37_6; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2588 = s1_way_wen_6_0_REG ? _GEN_2524 : meta_array_38_6; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2589 = s1_way_wen_6_0_REG ? _GEN_2525 : meta_array_39_6; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2590 = s1_way_wen_6_0_REG ? _GEN_2526 : meta_array_40_6; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2591 = s1_way_wen_6_0_REG ? _GEN_2527 : meta_array_41_6; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2592 = s1_way_wen_6_0_REG ? _GEN_2528 : meta_array_42_6; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2593 = s1_way_wen_6_0_REG ? _GEN_2529 : meta_array_43_6; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2594 = s1_way_wen_6_0_REG ? _GEN_2530 : meta_array_44_6; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2595 = s1_way_wen_6_0_REG ? _GEN_2531 : meta_array_45_6; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2596 = s1_way_wen_6_0_REG ? _GEN_2532 : meta_array_46_6; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2597 = s1_way_wen_6_0_REG ? _GEN_2533 : meta_array_47_6; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2598 = s1_way_wen_6_0_REG ? _GEN_2534 : meta_array_48_6; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2599 = s1_way_wen_6_0_REG ? _GEN_2535 : meta_array_49_6; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2600 = s1_way_wen_6_0_REG ? _GEN_2536 : meta_array_50_6; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2601 = s1_way_wen_6_0_REG ? _GEN_2537 : meta_array_51_6; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2602 = s1_way_wen_6_0_REG ? _GEN_2538 : meta_array_52_6; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2603 = s1_way_wen_6_0_REG ? _GEN_2539 : meta_array_53_6; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2604 = s1_way_wen_6_0_REG ? _GEN_2540 : meta_array_54_6; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2605 = s1_way_wen_6_0_REG ? _GEN_2541 : meta_array_55_6; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2606 = s1_way_wen_6_0_REG ? _GEN_2542 : meta_array_56_6; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2607 = s1_way_wen_6_0_REG ? _GEN_2543 : meta_array_57_6; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2608 = s1_way_wen_6_0_REG ? _GEN_2544 : meta_array_58_6; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2609 = s1_way_wen_6_0_REG ? _GEN_2545 : meta_array_59_6; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2610 = s1_way_wen_6_0_REG ? _GEN_2546 : meta_array_60_6; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2611 = s1_way_wen_6_0_REG ? _GEN_2547 : meta_array_61_6; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2612 = s1_way_wen_6_0_REG ? _GEN_2548 : meta_array_62_6; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2613 = s1_way_wen_6_0_REG ? _GEN_2549 : meta_array_63_6; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  s0_way_wen_7_0 = io_write_0_valid & io_write_0_bits_way_en[7]; // @[AsynchronousMetaArray.scala 152:49]
  wire  _GEN_2616 = 6'h0 == s1_way_waddr_7_0_r ? s1_way_wdata_7_0_r : meta_array_0_7; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2617 = 6'h1 == s1_way_waddr_7_0_r ? s1_way_wdata_7_0_r : meta_array_1_7; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2618 = 6'h2 == s1_way_waddr_7_0_r ? s1_way_wdata_7_0_r : meta_array_2_7; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2619 = 6'h3 == s1_way_waddr_7_0_r ? s1_way_wdata_7_0_r : meta_array_3_7; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2620 = 6'h4 == s1_way_waddr_7_0_r ? s1_way_wdata_7_0_r : meta_array_4_7; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2621 = 6'h5 == s1_way_waddr_7_0_r ? s1_way_wdata_7_0_r : meta_array_5_7; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2622 = 6'h6 == s1_way_waddr_7_0_r ? s1_way_wdata_7_0_r : meta_array_6_7; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2623 = 6'h7 == s1_way_waddr_7_0_r ? s1_way_wdata_7_0_r : meta_array_7_7; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2624 = 6'h8 == s1_way_waddr_7_0_r ? s1_way_wdata_7_0_r : meta_array_8_7; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2625 = 6'h9 == s1_way_waddr_7_0_r ? s1_way_wdata_7_0_r : meta_array_9_7; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2626 = 6'ha == s1_way_waddr_7_0_r ? s1_way_wdata_7_0_r : meta_array_10_7; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2627 = 6'hb == s1_way_waddr_7_0_r ? s1_way_wdata_7_0_r : meta_array_11_7; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2628 = 6'hc == s1_way_waddr_7_0_r ? s1_way_wdata_7_0_r : meta_array_12_7; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2629 = 6'hd == s1_way_waddr_7_0_r ? s1_way_wdata_7_0_r : meta_array_13_7; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2630 = 6'he == s1_way_waddr_7_0_r ? s1_way_wdata_7_0_r : meta_array_14_7; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2631 = 6'hf == s1_way_waddr_7_0_r ? s1_way_wdata_7_0_r : meta_array_15_7; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2632 = 6'h10 == s1_way_waddr_7_0_r ? s1_way_wdata_7_0_r : meta_array_16_7; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2633 = 6'h11 == s1_way_waddr_7_0_r ? s1_way_wdata_7_0_r : meta_array_17_7; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2634 = 6'h12 == s1_way_waddr_7_0_r ? s1_way_wdata_7_0_r : meta_array_18_7; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2635 = 6'h13 == s1_way_waddr_7_0_r ? s1_way_wdata_7_0_r : meta_array_19_7; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2636 = 6'h14 == s1_way_waddr_7_0_r ? s1_way_wdata_7_0_r : meta_array_20_7; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2637 = 6'h15 == s1_way_waddr_7_0_r ? s1_way_wdata_7_0_r : meta_array_21_7; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2638 = 6'h16 == s1_way_waddr_7_0_r ? s1_way_wdata_7_0_r : meta_array_22_7; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2639 = 6'h17 == s1_way_waddr_7_0_r ? s1_way_wdata_7_0_r : meta_array_23_7; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2640 = 6'h18 == s1_way_waddr_7_0_r ? s1_way_wdata_7_0_r : meta_array_24_7; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2641 = 6'h19 == s1_way_waddr_7_0_r ? s1_way_wdata_7_0_r : meta_array_25_7; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2642 = 6'h1a == s1_way_waddr_7_0_r ? s1_way_wdata_7_0_r : meta_array_26_7; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2643 = 6'h1b == s1_way_waddr_7_0_r ? s1_way_wdata_7_0_r : meta_array_27_7; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2644 = 6'h1c == s1_way_waddr_7_0_r ? s1_way_wdata_7_0_r : meta_array_28_7; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2645 = 6'h1d == s1_way_waddr_7_0_r ? s1_way_wdata_7_0_r : meta_array_29_7; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2646 = 6'h1e == s1_way_waddr_7_0_r ? s1_way_wdata_7_0_r : meta_array_30_7; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2647 = 6'h1f == s1_way_waddr_7_0_r ? s1_way_wdata_7_0_r : meta_array_31_7; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2648 = 6'h20 == s1_way_waddr_7_0_r ? s1_way_wdata_7_0_r : meta_array_32_7; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2649 = 6'h21 == s1_way_waddr_7_0_r ? s1_way_wdata_7_0_r : meta_array_33_7; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2650 = 6'h22 == s1_way_waddr_7_0_r ? s1_way_wdata_7_0_r : meta_array_34_7; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2651 = 6'h23 == s1_way_waddr_7_0_r ? s1_way_wdata_7_0_r : meta_array_35_7; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2652 = 6'h24 == s1_way_waddr_7_0_r ? s1_way_wdata_7_0_r : meta_array_36_7; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2653 = 6'h25 == s1_way_waddr_7_0_r ? s1_way_wdata_7_0_r : meta_array_37_7; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2654 = 6'h26 == s1_way_waddr_7_0_r ? s1_way_wdata_7_0_r : meta_array_38_7; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2655 = 6'h27 == s1_way_waddr_7_0_r ? s1_way_wdata_7_0_r : meta_array_39_7; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2656 = 6'h28 == s1_way_waddr_7_0_r ? s1_way_wdata_7_0_r : meta_array_40_7; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2657 = 6'h29 == s1_way_waddr_7_0_r ? s1_way_wdata_7_0_r : meta_array_41_7; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2658 = 6'h2a == s1_way_waddr_7_0_r ? s1_way_wdata_7_0_r : meta_array_42_7; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2659 = 6'h2b == s1_way_waddr_7_0_r ? s1_way_wdata_7_0_r : meta_array_43_7; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2660 = 6'h2c == s1_way_waddr_7_0_r ? s1_way_wdata_7_0_r : meta_array_44_7; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2661 = 6'h2d == s1_way_waddr_7_0_r ? s1_way_wdata_7_0_r : meta_array_45_7; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2662 = 6'h2e == s1_way_waddr_7_0_r ? s1_way_wdata_7_0_r : meta_array_46_7; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2663 = 6'h2f == s1_way_waddr_7_0_r ? s1_way_wdata_7_0_r : meta_array_47_7; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2664 = 6'h30 == s1_way_waddr_7_0_r ? s1_way_wdata_7_0_r : meta_array_48_7; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2665 = 6'h31 == s1_way_waddr_7_0_r ? s1_way_wdata_7_0_r : meta_array_49_7; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2666 = 6'h32 == s1_way_waddr_7_0_r ? s1_way_wdata_7_0_r : meta_array_50_7; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2667 = 6'h33 == s1_way_waddr_7_0_r ? s1_way_wdata_7_0_r : meta_array_51_7; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2668 = 6'h34 == s1_way_waddr_7_0_r ? s1_way_wdata_7_0_r : meta_array_52_7; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2669 = 6'h35 == s1_way_waddr_7_0_r ? s1_way_wdata_7_0_r : meta_array_53_7; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2670 = 6'h36 == s1_way_waddr_7_0_r ? s1_way_wdata_7_0_r : meta_array_54_7; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2671 = 6'h37 == s1_way_waddr_7_0_r ? s1_way_wdata_7_0_r : meta_array_55_7; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2672 = 6'h38 == s1_way_waddr_7_0_r ? s1_way_wdata_7_0_r : meta_array_56_7; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2673 = 6'h39 == s1_way_waddr_7_0_r ? s1_way_wdata_7_0_r : meta_array_57_7; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2674 = 6'h3a == s1_way_waddr_7_0_r ? s1_way_wdata_7_0_r : meta_array_58_7; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2675 = 6'h3b == s1_way_waddr_7_0_r ? s1_way_wdata_7_0_r : meta_array_59_7; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2676 = 6'h3c == s1_way_waddr_7_0_r ? s1_way_wdata_7_0_r : meta_array_60_7; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2677 = 6'h3d == s1_way_waddr_7_0_r ? s1_way_wdata_7_0_r : meta_array_61_7; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2678 = 6'h3e == s1_way_waddr_7_0_r ? s1_way_wdata_7_0_r : meta_array_62_7; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2679 = 6'h3f == s1_way_waddr_7_0_r ? s1_way_wdata_7_0_r : meta_array_63_7; // @[AsynchronousMetaArray.scala 115:27 157:{55,55}]
  wire  _GEN_2680 = s1_way_wen_7_0_REG ? _GEN_2616 : meta_array_0_7; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2681 = s1_way_wen_7_0_REG ? _GEN_2617 : meta_array_1_7; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2682 = s1_way_wen_7_0_REG ? _GEN_2618 : meta_array_2_7; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2683 = s1_way_wen_7_0_REG ? _GEN_2619 : meta_array_3_7; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2684 = s1_way_wen_7_0_REG ? _GEN_2620 : meta_array_4_7; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2685 = s1_way_wen_7_0_REG ? _GEN_2621 : meta_array_5_7; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2686 = s1_way_wen_7_0_REG ? _GEN_2622 : meta_array_6_7; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2687 = s1_way_wen_7_0_REG ? _GEN_2623 : meta_array_7_7; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2688 = s1_way_wen_7_0_REG ? _GEN_2624 : meta_array_8_7; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2689 = s1_way_wen_7_0_REG ? _GEN_2625 : meta_array_9_7; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2690 = s1_way_wen_7_0_REG ? _GEN_2626 : meta_array_10_7; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2691 = s1_way_wen_7_0_REG ? _GEN_2627 : meta_array_11_7; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2692 = s1_way_wen_7_0_REG ? _GEN_2628 : meta_array_12_7; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2693 = s1_way_wen_7_0_REG ? _GEN_2629 : meta_array_13_7; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2694 = s1_way_wen_7_0_REG ? _GEN_2630 : meta_array_14_7; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2695 = s1_way_wen_7_0_REG ? _GEN_2631 : meta_array_15_7; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2696 = s1_way_wen_7_0_REG ? _GEN_2632 : meta_array_16_7; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2697 = s1_way_wen_7_0_REG ? _GEN_2633 : meta_array_17_7; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2698 = s1_way_wen_7_0_REG ? _GEN_2634 : meta_array_18_7; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2699 = s1_way_wen_7_0_REG ? _GEN_2635 : meta_array_19_7; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2700 = s1_way_wen_7_0_REG ? _GEN_2636 : meta_array_20_7; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2701 = s1_way_wen_7_0_REG ? _GEN_2637 : meta_array_21_7; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2702 = s1_way_wen_7_0_REG ? _GEN_2638 : meta_array_22_7; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2703 = s1_way_wen_7_0_REG ? _GEN_2639 : meta_array_23_7; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2704 = s1_way_wen_7_0_REG ? _GEN_2640 : meta_array_24_7; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2705 = s1_way_wen_7_0_REG ? _GEN_2641 : meta_array_25_7; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2706 = s1_way_wen_7_0_REG ? _GEN_2642 : meta_array_26_7; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2707 = s1_way_wen_7_0_REG ? _GEN_2643 : meta_array_27_7; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2708 = s1_way_wen_7_0_REG ? _GEN_2644 : meta_array_28_7; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2709 = s1_way_wen_7_0_REG ? _GEN_2645 : meta_array_29_7; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2710 = s1_way_wen_7_0_REG ? _GEN_2646 : meta_array_30_7; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2711 = s1_way_wen_7_0_REG ? _GEN_2647 : meta_array_31_7; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2712 = s1_way_wen_7_0_REG ? _GEN_2648 : meta_array_32_7; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2713 = s1_way_wen_7_0_REG ? _GEN_2649 : meta_array_33_7; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2714 = s1_way_wen_7_0_REG ? _GEN_2650 : meta_array_34_7; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2715 = s1_way_wen_7_0_REG ? _GEN_2651 : meta_array_35_7; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2716 = s1_way_wen_7_0_REG ? _GEN_2652 : meta_array_36_7; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2717 = s1_way_wen_7_0_REG ? _GEN_2653 : meta_array_37_7; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2718 = s1_way_wen_7_0_REG ? _GEN_2654 : meta_array_38_7; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2719 = s1_way_wen_7_0_REG ? _GEN_2655 : meta_array_39_7; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2720 = s1_way_wen_7_0_REG ? _GEN_2656 : meta_array_40_7; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2721 = s1_way_wen_7_0_REG ? _GEN_2657 : meta_array_41_7; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2722 = s1_way_wen_7_0_REG ? _GEN_2658 : meta_array_42_7; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2723 = s1_way_wen_7_0_REG ? _GEN_2659 : meta_array_43_7; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2724 = s1_way_wen_7_0_REG ? _GEN_2660 : meta_array_44_7; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2725 = s1_way_wen_7_0_REG ? _GEN_2661 : meta_array_45_7; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2726 = s1_way_wen_7_0_REG ? _GEN_2662 : meta_array_46_7; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2727 = s1_way_wen_7_0_REG ? _GEN_2663 : meta_array_47_7; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2728 = s1_way_wen_7_0_REG ? _GEN_2664 : meta_array_48_7; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2729 = s1_way_wen_7_0_REG ? _GEN_2665 : meta_array_49_7; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2730 = s1_way_wen_7_0_REG ? _GEN_2666 : meta_array_50_7; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2731 = s1_way_wen_7_0_REG ? _GEN_2667 : meta_array_51_7; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2732 = s1_way_wen_7_0_REG ? _GEN_2668 : meta_array_52_7; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2733 = s1_way_wen_7_0_REG ? _GEN_2669 : meta_array_53_7; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2734 = s1_way_wen_7_0_REG ? _GEN_2670 : meta_array_54_7; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2735 = s1_way_wen_7_0_REG ? _GEN_2671 : meta_array_55_7; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2736 = s1_way_wen_7_0_REG ? _GEN_2672 : meta_array_56_7; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2737 = s1_way_wen_7_0_REG ? _GEN_2673 : meta_array_57_7; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2738 = s1_way_wen_7_0_REG ? _GEN_2674 : meta_array_58_7; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2739 = s1_way_wen_7_0_REG ? _GEN_2675 : meta_array_59_7; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2740 = s1_way_wen_7_0_REG ? _GEN_2676 : meta_array_60_7; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2741 = s1_way_wen_7_0_REG ? _GEN_2677 : meta_array_61_7; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2742 = s1_way_wen_7_0_REG ? _GEN_2678 : meta_array_62_7; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  _GEN_2743 = s1_way_wen_7_0_REG ? _GEN_2679 : meta_array_63_7; // @[AsynchronousMetaArray.scala 115:27 156:41]
  wire  s0_way_wen_0_1 = io_write_1_valid & io_write_1_bits_way_en[0]; // @[AsynchronousMetaArray.scala 152:49]
  wire  s0_way_wen_1_1 = io_write_1_valid & io_write_1_bits_way_en[1]; // @[AsynchronousMetaArray.scala 152:49]
  wire  s0_way_wen_2_1 = io_write_1_valid & io_write_1_bits_way_en[2]; // @[AsynchronousMetaArray.scala 152:49]
  wire  s0_way_wen_3_1 = io_write_1_valid & io_write_1_bits_way_en[3]; // @[AsynchronousMetaArray.scala 152:49]
  wire  s0_way_wen_4_1 = io_write_1_valid & io_write_1_bits_way_en[4]; // @[AsynchronousMetaArray.scala 152:49]
  wire  s0_way_wen_5_1 = io_write_1_valid & io_write_1_bits_way_en[5]; // @[AsynchronousMetaArray.scala 152:49]
  wire  s0_way_wen_6_1 = io_write_1_valid & io_write_1_bits_way_en[6]; // @[AsynchronousMetaArray.scala 152:49]
  wire  s0_way_wen_7_1 = io_write_1_valid & io_write_1_bits_way_en[7]; // @[AsynchronousMetaArray.scala 152:49]
  assign io_resp_0_0 = io_resp_0_0_r ? io_resp_0_0_r1 : _GEN_70; // @[AsynchronousMetaArray.scala 139:25]
  assign io_resp_0_1 = io_resp_0_1_r ? io_resp_0_1_r1 : _GEN_141; // @[AsynchronousMetaArray.scala 139:25]
  assign io_resp_0_2 = io_resp_0_2_r ? io_resp_0_2_r1 : _GEN_212; // @[AsynchronousMetaArray.scala 139:25]
  assign io_resp_0_3 = io_resp_0_3_r ? io_resp_0_3_r1 : _GEN_283; // @[AsynchronousMetaArray.scala 139:25]
  assign io_resp_0_4 = io_resp_0_4_r ? io_resp_0_4_r1 : _GEN_354; // @[AsynchronousMetaArray.scala 139:25]
  assign io_resp_0_5 = io_resp_0_5_r ? io_resp_0_5_r1 : _GEN_425; // @[AsynchronousMetaArray.scala 139:25]
  assign io_resp_0_6 = io_resp_0_6_r ? io_resp_0_6_r1 : _GEN_496; // @[AsynchronousMetaArray.scala 139:25]
  assign io_resp_0_7 = io_resp_0_7_r ? io_resp_0_7_r1 : _GEN_567; // @[AsynchronousMetaArray.scala 139:25]
  assign io_resp_1_0 = io_resp_1_0_r ? io_resp_1_0_r1 : _GEN_638; // @[AsynchronousMetaArray.scala 139:25]
  assign io_resp_1_1 = io_resp_1_1_r ? io_resp_1_1_r1 : _GEN_709; // @[AsynchronousMetaArray.scala 139:25]
  assign io_resp_1_2 = io_resp_1_2_r ? io_resp_1_2_r1 : _GEN_780; // @[AsynchronousMetaArray.scala 139:25]
  assign io_resp_1_3 = io_resp_1_3_r ? io_resp_1_3_r1 : _GEN_851; // @[AsynchronousMetaArray.scala 139:25]
  assign io_resp_1_4 = io_resp_1_4_r ? io_resp_1_4_r1 : _GEN_922; // @[AsynchronousMetaArray.scala 139:25]
  assign io_resp_1_5 = io_resp_1_5_r ? io_resp_1_5_r1 : _GEN_993; // @[AsynchronousMetaArray.scala 139:25]
  assign io_resp_1_6 = io_resp_1_6_r ? io_resp_1_6_r1 : _GEN_1064; // @[AsynchronousMetaArray.scala 139:25]
  assign io_resp_1_7 = io_resp_1_7_r ? io_resp_1_7_r1 : _GEN_1135; // @[AsynchronousMetaArray.scala 139:25]
  assign io_resp_2_0 = io_resp_2_0_r ? io_resp_2_0_r1 : _GEN_1206; // @[AsynchronousMetaArray.scala 139:25]
  assign io_resp_2_1 = io_resp_2_1_r ? io_resp_2_1_r1 : _GEN_1277; // @[AsynchronousMetaArray.scala 139:25]
  assign io_resp_2_2 = io_resp_2_2_r ? io_resp_2_2_r1 : _GEN_1348; // @[AsynchronousMetaArray.scala 139:25]
  assign io_resp_2_3 = io_resp_2_3_r ? io_resp_2_3_r1 : _GEN_1419; // @[AsynchronousMetaArray.scala 139:25]
  assign io_resp_2_4 = io_resp_2_4_r ? io_resp_2_4_r1 : _GEN_1490; // @[AsynchronousMetaArray.scala 139:25]
  assign io_resp_2_5 = io_resp_2_5_r ? io_resp_2_5_r1 : _GEN_1561; // @[AsynchronousMetaArray.scala 139:25]
  assign io_resp_2_6 = io_resp_2_6_r ? io_resp_2_6_r1 : _GEN_1632; // @[AsynchronousMetaArray.scala 139:25]
  assign io_resp_2_7 = io_resp_2_7_r ? io_resp_2_7_r1 : _GEN_1703; // @[AsynchronousMetaArray.scala 139:25]
  always @(posedge clock) begin
    if (s0_way_wen_0_0) begin // @[Reg.scala 17:18]
      s1_way_waddr_0_0_r <= io_write_0_bits_idx; // @[Reg.scala 17:22]
    end
    s1_way_wen_0_0_REG <= io_write_0_valid & io_write_0_bits_way_en[0]; // @[AsynchronousMetaArray.scala 152:49]
    if (s0_way_wen_0_0) begin // @[Reg.scala 17:18]
      s1_way_wdata_0_0_r <= io_write_0_bits_flag; // @[Reg.scala 17:22]
    end
    if (s0_way_wen_0_1) begin // @[Reg.scala 17:18]
      s1_way_waddr_0_1_r <= io_write_1_bits_idx; // @[Reg.scala 17:22]
    end
    s1_way_wen_0_1_REG <= io_write_1_valid & io_write_1_bits_way_en[0]; // @[AsynchronousMetaArray.scala 152:49]
    if (s0_way_wen_0_1) begin // @[Reg.scala 17:18]
      s1_way_wdata_0_1_r <= io_write_1_bits_flag; // @[Reg.scala 17:22]
    end
    if (io_read_0_valid) begin // @[Reg.scala 17:18]
      io_resp_0_0_r <= read_way_bypass; // @[Reg.scala 17:22]
    end
    if (read_way_bypass) begin // @[Reg.scala 17:18]
      if (s1_way_wen_0_1_REG & s1_way_waddr_0_1_r == io_read_0_bits_idx) begin // @[AsynchronousMetaArray.scala 134:85]
        io_resp_0_0_r1 <= s1_way_wdata_0_1_r; // @[AsynchronousMetaArray.scala 136:25]
      end else begin
        io_resp_0_0_r1 <= s1_way_wdata_0_0_r;
      end
    end
    if (io_read_0_valid) begin // @[Reg.scala 17:18]
      io_resp_0_0_r2 <= io_read_0_bits_idx; // @[Reg.scala 17:22]
    end
    if (s0_way_wen_1_0) begin // @[Reg.scala 17:18]
      s1_way_waddr_1_0_r <= io_write_0_bits_idx; // @[Reg.scala 17:22]
    end
    s1_way_wen_1_0_REG <= io_write_0_valid & io_write_0_bits_way_en[1]; // @[AsynchronousMetaArray.scala 152:49]
    if (s0_way_wen_1_0) begin // @[Reg.scala 17:18]
      s1_way_wdata_1_0_r <= io_write_0_bits_flag; // @[Reg.scala 17:22]
    end
    if (s0_way_wen_1_1) begin // @[Reg.scala 17:18]
      s1_way_waddr_1_1_r <= io_write_1_bits_idx; // @[Reg.scala 17:22]
    end
    s1_way_wen_1_1_REG <= io_write_1_valid & io_write_1_bits_way_en[1]; // @[AsynchronousMetaArray.scala 152:49]
    if (s0_way_wen_1_1) begin // @[Reg.scala 17:18]
      s1_way_wdata_1_1_r <= io_write_1_bits_flag; // @[Reg.scala 17:22]
    end
    if (io_read_0_valid) begin // @[Reg.scala 17:18]
      io_resp_0_1_r <= read_way_bypass_1; // @[Reg.scala 17:22]
    end
    if (read_way_bypass_1) begin // @[Reg.scala 17:18]
      if (s1_way_wen_1_1_REG & s1_way_waddr_1_1_r == io_read_0_bits_idx) begin // @[AsynchronousMetaArray.scala 134:85]
        io_resp_0_1_r1 <= s1_way_wdata_1_1_r; // @[AsynchronousMetaArray.scala 136:25]
      end else begin
        io_resp_0_1_r1 <= s1_way_wdata_1_0_r;
      end
    end
    if (io_read_0_valid) begin // @[Reg.scala 17:18]
      io_resp_0_1_r2 <= io_read_0_bits_idx; // @[Reg.scala 17:22]
    end
    if (s0_way_wen_2_0) begin // @[Reg.scala 17:18]
      s1_way_waddr_2_0_r <= io_write_0_bits_idx; // @[Reg.scala 17:22]
    end
    s1_way_wen_2_0_REG <= io_write_0_valid & io_write_0_bits_way_en[2]; // @[AsynchronousMetaArray.scala 152:49]
    if (s0_way_wen_2_0) begin // @[Reg.scala 17:18]
      s1_way_wdata_2_0_r <= io_write_0_bits_flag; // @[Reg.scala 17:22]
    end
    if (s0_way_wen_2_1) begin // @[Reg.scala 17:18]
      s1_way_waddr_2_1_r <= io_write_1_bits_idx; // @[Reg.scala 17:22]
    end
    s1_way_wen_2_1_REG <= io_write_1_valid & io_write_1_bits_way_en[2]; // @[AsynchronousMetaArray.scala 152:49]
    if (s0_way_wen_2_1) begin // @[Reg.scala 17:18]
      s1_way_wdata_2_1_r <= io_write_1_bits_flag; // @[Reg.scala 17:22]
    end
    if (io_read_0_valid) begin // @[Reg.scala 17:18]
      io_resp_0_2_r <= read_way_bypass_2; // @[Reg.scala 17:22]
    end
    if (read_way_bypass_2) begin // @[Reg.scala 17:18]
      if (s1_way_wen_2_1_REG & s1_way_waddr_2_1_r == io_read_0_bits_idx) begin // @[AsynchronousMetaArray.scala 134:85]
        io_resp_0_2_r1 <= s1_way_wdata_2_1_r; // @[AsynchronousMetaArray.scala 136:25]
      end else begin
        io_resp_0_2_r1 <= s1_way_wdata_2_0_r;
      end
    end
    if (io_read_0_valid) begin // @[Reg.scala 17:18]
      io_resp_0_2_r2 <= io_read_0_bits_idx; // @[Reg.scala 17:22]
    end
    if (s0_way_wen_3_0) begin // @[Reg.scala 17:18]
      s1_way_waddr_3_0_r <= io_write_0_bits_idx; // @[Reg.scala 17:22]
    end
    s1_way_wen_3_0_REG <= io_write_0_valid & io_write_0_bits_way_en[3]; // @[AsynchronousMetaArray.scala 152:49]
    if (s0_way_wen_3_0) begin // @[Reg.scala 17:18]
      s1_way_wdata_3_0_r <= io_write_0_bits_flag; // @[Reg.scala 17:22]
    end
    if (s0_way_wen_3_1) begin // @[Reg.scala 17:18]
      s1_way_waddr_3_1_r <= io_write_1_bits_idx; // @[Reg.scala 17:22]
    end
    s1_way_wen_3_1_REG <= io_write_1_valid & io_write_1_bits_way_en[3]; // @[AsynchronousMetaArray.scala 152:49]
    if (s0_way_wen_3_1) begin // @[Reg.scala 17:18]
      s1_way_wdata_3_1_r <= io_write_1_bits_flag; // @[Reg.scala 17:22]
    end
    if (io_read_0_valid) begin // @[Reg.scala 17:18]
      io_resp_0_3_r <= read_way_bypass_3; // @[Reg.scala 17:22]
    end
    if (read_way_bypass_3) begin // @[Reg.scala 17:18]
      if (s1_way_wen_3_1_REG & s1_way_waddr_3_1_r == io_read_0_bits_idx) begin // @[AsynchronousMetaArray.scala 134:85]
        io_resp_0_3_r1 <= s1_way_wdata_3_1_r; // @[AsynchronousMetaArray.scala 136:25]
      end else begin
        io_resp_0_3_r1 <= s1_way_wdata_3_0_r;
      end
    end
    if (io_read_0_valid) begin // @[Reg.scala 17:18]
      io_resp_0_3_r2 <= io_read_0_bits_idx; // @[Reg.scala 17:22]
    end
    if (s0_way_wen_4_0) begin // @[Reg.scala 17:18]
      s1_way_waddr_4_0_r <= io_write_0_bits_idx; // @[Reg.scala 17:22]
    end
    s1_way_wen_4_0_REG <= io_write_0_valid & io_write_0_bits_way_en[4]; // @[AsynchronousMetaArray.scala 152:49]
    if (s0_way_wen_4_0) begin // @[Reg.scala 17:18]
      s1_way_wdata_4_0_r <= io_write_0_bits_flag; // @[Reg.scala 17:22]
    end
    if (s0_way_wen_4_1) begin // @[Reg.scala 17:18]
      s1_way_waddr_4_1_r <= io_write_1_bits_idx; // @[Reg.scala 17:22]
    end
    s1_way_wen_4_1_REG <= io_write_1_valid & io_write_1_bits_way_en[4]; // @[AsynchronousMetaArray.scala 152:49]
    if (s0_way_wen_4_1) begin // @[Reg.scala 17:18]
      s1_way_wdata_4_1_r <= io_write_1_bits_flag; // @[Reg.scala 17:22]
    end
    if (io_read_0_valid) begin // @[Reg.scala 17:18]
      io_resp_0_4_r <= read_way_bypass_4; // @[Reg.scala 17:22]
    end
    if (read_way_bypass_4) begin // @[Reg.scala 17:18]
      if (s1_way_wen_4_1_REG & s1_way_waddr_4_1_r == io_read_0_bits_idx) begin // @[AsynchronousMetaArray.scala 134:85]
        io_resp_0_4_r1 <= s1_way_wdata_4_1_r; // @[AsynchronousMetaArray.scala 136:25]
      end else begin
        io_resp_0_4_r1 <= s1_way_wdata_4_0_r;
      end
    end
    if (io_read_0_valid) begin // @[Reg.scala 17:18]
      io_resp_0_4_r2 <= io_read_0_bits_idx; // @[Reg.scala 17:22]
    end
    if (s0_way_wen_5_0) begin // @[Reg.scala 17:18]
      s1_way_waddr_5_0_r <= io_write_0_bits_idx; // @[Reg.scala 17:22]
    end
    s1_way_wen_5_0_REG <= io_write_0_valid & io_write_0_bits_way_en[5]; // @[AsynchronousMetaArray.scala 152:49]
    if (s0_way_wen_5_0) begin // @[Reg.scala 17:18]
      s1_way_wdata_5_0_r <= io_write_0_bits_flag; // @[Reg.scala 17:22]
    end
    if (s0_way_wen_5_1) begin // @[Reg.scala 17:18]
      s1_way_waddr_5_1_r <= io_write_1_bits_idx; // @[Reg.scala 17:22]
    end
    s1_way_wen_5_1_REG <= io_write_1_valid & io_write_1_bits_way_en[5]; // @[AsynchronousMetaArray.scala 152:49]
    if (s0_way_wen_5_1) begin // @[Reg.scala 17:18]
      s1_way_wdata_5_1_r <= io_write_1_bits_flag; // @[Reg.scala 17:22]
    end
    if (io_read_0_valid) begin // @[Reg.scala 17:18]
      io_resp_0_5_r <= read_way_bypass_5; // @[Reg.scala 17:22]
    end
    if (read_way_bypass_5) begin // @[Reg.scala 17:18]
      if (s1_way_wen_5_1_REG & s1_way_waddr_5_1_r == io_read_0_bits_idx) begin // @[AsynchronousMetaArray.scala 134:85]
        io_resp_0_5_r1 <= s1_way_wdata_5_1_r; // @[AsynchronousMetaArray.scala 136:25]
      end else begin
        io_resp_0_5_r1 <= s1_way_wdata_5_0_r;
      end
    end
    if (io_read_0_valid) begin // @[Reg.scala 17:18]
      io_resp_0_5_r2 <= io_read_0_bits_idx; // @[Reg.scala 17:22]
    end
    if (s0_way_wen_6_0) begin // @[Reg.scala 17:18]
      s1_way_waddr_6_0_r <= io_write_0_bits_idx; // @[Reg.scala 17:22]
    end
    s1_way_wen_6_0_REG <= io_write_0_valid & io_write_0_bits_way_en[6]; // @[AsynchronousMetaArray.scala 152:49]
    if (s0_way_wen_6_0) begin // @[Reg.scala 17:18]
      s1_way_wdata_6_0_r <= io_write_0_bits_flag; // @[Reg.scala 17:22]
    end
    if (s0_way_wen_6_1) begin // @[Reg.scala 17:18]
      s1_way_waddr_6_1_r <= io_write_1_bits_idx; // @[Reg.scala 17:22]
    end
    s1_way_wen_6_1_REG <= io_write_1_valid & io_write_1_bits_way_en[6]; // @[AsynchronousMetaArray.scala 152:49]
    if (s0_way_wen_6_1) begin // @[Reg.scala 17:18]
      s1_way_wdata_6_1_r <= io_write_1_bits_flag; // @[Reg.scala 17:22]
    end
    if (io_read_0_valid) begin // @[Reg.scala 17:18]
      io_resp_0_6_r <= read_way_bypass_6; // @[Reg.scala 17:22]
    end
    if (read_way_bypass_6) begin // @[Reg.scala 17:18]
      if (s1_way_wen_6_1_REG & s1_way_waddr_6_1_r == io_read_0_bits_idx) begin // @[AsynchronousMetaArray.scala 134:85]
        io_resp_0_6_r1 <= s1_way_wdata_6_1_r; // @[AsynchronousMetaArray.scala 136:25]
      end else begin
        io_resp_0_6_r1 <= s1_way_wdata_6_0_r;
      end
    end
    if (io_read_0_valid) begin // @[Reg.scala 17:18]
      io_resp_0_6_r2 <= io_read_0_bits_idx; // @[Reg.scala 17:22]
    end
    if (s0_way_wen_7_0) begin // @[Reg.scala 17:18]
      s1_way_waddr_7_0_r <= io_write_0_bits_idx; // @[Reg.scala 17:22]
    end
    s1_way_wen_7_0_REG <= io_write_0_valid & io_write_0_bits_way_en[7]; // @[AsynchronousMetaArray.scala 152:49]
    if (s0_way_wen_7_0) begin // @[Reg.scala 17:18]
      s1_way_wdata_7_0_r <= io_write_0_bits_flag; // @[Reg.scala 17:22]
    end
    if (s0_way_wen_7_1) begin // @[Reg.scala 17:18]
      s1_way_waddr_7_1_r <= io_write_1_bits_idx; // @[Reg.scala 17:22]
    end
    s1_way_wen_7_1_REG <= io_write_1_valid & io_write_1_bits_way_en[7]; // @[AsynchronousMetaArray.scala 152:49]
    if (s0_way_wen_7_1) begin // @[Reg.scala 17:18]
      s1_way_wdata_7_1_r <= io_write_1_bits_flag; // @[Reg.scala 17:22]
    end
    if (io_read_0_valid) begin // @[Reg.scala 17:18]
      io_resp_0_7_r <= read_way_bypass_7; // @[Reg.scala 17:22]
    end
    if (read_way_bypass_7) begin // @[Reg.scala 17:18]
      if (s1_way_wen_7_1_REG & s1_way_waddr_7_1_r == io_read_0_bits_idx) begin // @[AsynchronousMetaArray.scala 134:85]
        io_resp_0_7_r1 <= s1_way_wdata_7_1_r; // @[AsynchronousMetaArray.scala 136:25]
      end else begin
        io_resp_0_7_r1 <= s1_way_wdata_7_0_r;
      end
    end
    if (io_read_0_valid) begin // @[Reg.scala 17:18]
      io_resp_0_7_r2 <= io_read_0_bits_idx; // @[Reg.scala 17:22]
    end
    if (io_read_1_valid) begin // @[Reg.scala 17:18]
      io_resp_1_0_r <= read_way_bypass_8; // @[Reg.scala 17:22]
    end
    if (read_way_bypass_8) begin // @[Reg.scala 17:18]
      if (s1_way_wen_0_1_REG & s1_way_waddr_0_1_r == io_read_1_bits_idx) begin // @[AsynchronousMetaArray.scala 134:85]
        io_resp_1_0_r1 <= s1_way_wdata_0_1_r; // @[AsynchronousMetaArray.scala 136:25]
      end else begin
        io_resp_1_0_r1 <= s1_way_wdata_0_0_r;
      end
    end
    if (io_read_1_valid) begin // @[Reg.scala 17:18]
      io_resp_1_0_r2 <= io_read_1_bits_idx; // @[Reg.scala 17:22]
    end
    if (io_read_1_valid) begin // @[Reg.scala 17:18]
      io_resp_1_1_r <= read_way_bypass_9; // @[Reg.scala 17:22]
    end
    if (read_way_bypass_9) begin // @[Reg.scala 17:18]
      if (s1_way_wen_1_1_REG & s1_way_waddr_1_1_r == io_read_1_bits_idx) begin // @[AsynchronousMetaArray.scala 134:85]
        io_resp_1_1_r1 <= s1_way_wdata_1_1_r; // @[AsynchronousMetaArray.scala 136:25]
      end else begin
        io_resp_1_1_r1 <= s1_way_wdata_1_0_r;
      end
    end
    if (io_read_1_valid) begin // @[Reg.scala 17:18]
      io_resp_1_1_r2 <= io_read_1_bits_idx; // @[Reg.scala 17:22]
    end
    if (io_read_1_valid) begin // @[Reg.scala 17:18]
      io_resp_1_2_r <= read_way_bypass_10; // @[Reg.scala 17:22]
    end
    if (read_way_bypass_10) begin // @[Reg.scala 17:18]
      if (s1_way_wen_2_1_REG & s1_way_waddr_2_1_r == io_read_1_bits_idx) begin // @[AsynchronousMetaArray.scala 134:85]
        io_resp_1_2_r1 <= s1_way_wdata_2_1_r; // @[AsynchronousMetaArray.scala 136:25]
      end else begin
        io_resp_1_2_r1 <= s1_way_wdata_2_0_r;
      end
    end
    if (io_read_1_valid) begin // @[Reg.scala 17:18]
      io_resp_1_2_r2 <= io_read_1_bits_idx; // @[Reg.scala 17:22]
    end
    if (io_read_1_valid) begin // @[Reg.scala 17:18]
      io_resp_1_3_r <= read_way_bypass_11; // @[Reg.scala 17:22]
    end
    if (read_way_bypass_11) begin // @[Reg.scala 17:18]
      if (s1_way_wen_3_1_REG & s1_way_waddr_3_1_r == io_read_1_bits_idx) begin // @[AsynchronousMetaArray.scala 134:85]
        io_resp_1_3_r1 <= s1_way_wdata_3_1_r; // @[AsynchronousMetaArray.scala 136:25]
      end else begin
        io_resp_1_3_r1 <= s1_way_wdata_3_0_r;
      end
    end
    if (io_read_1_valid) begin // @[Reg.scala 17:18]
      io_resp_1_3_r2 <= io_read_1_bits_idx; // @[Reg.scala 17:22]
    end
    if (io_read_1_valid) begin // @[Reg.scala 17:18]
      io_resp_1_4_r <= read_way_bypass_12; // @[Reg.scala 17:22]
    end
    if (read_way_bypass_12) begin // @[Reg.scala 17:18]
      if (s1_way_wen_4_1_REG & s1_way_waddr_4_1_r == io_read_1_bits_idx) begin // @[AsynchronousMetaArray.scala 134:85]
        io_resp_1_4_r1 <= s1_way_wdata_4_1_r; // @[AsynchronousMetaArray.scala 136:25]
      end else begin
        io_resp_1_4_r1 <= s1_way_wdata_4_0_r;
      end
    end
    if (io_read_1_valid) begin // @[Reg.scala 17:18]
      io_resp_1_4_r2 <= io_read_1_bits_idx; // @[Reg.scala 17:22]
    end
    if (io_read_1_valid) begin // @[Reg.scala 17:18]
      io_resp_1_5_r <= read_way_bypass_13; // @[Reg.scala 17:22]
    end
    if (read_way_bypass_13) begin // @[Reg.scala 17:18]
      if (s1_way_wen_5_1_REG & s1_way_waddr_5_1_r == io_read_1_bits_idx) begin // @[AsynchronousMetaArray.scala 134:85]
        io_resp_1_5_r1 <= s1_way_wdata_5_1_r; // @[AsynchronousMetaArray.scala 136:25]
      end else begin
        io_resp_1_5_r1 <= s1_way_wdata_5_0_r;
      end
    end
    if (io_read_1_valid) begin // @[Reg.scala 17:18]
      io_resp_1_5_r2 <= io_read_1_bits_idx; // @[Reg.scala 17:22]
    end
    if (io_read_1_valid) begin // @[Reg.scala 17:18]
      io_resp_1_6_r <= read_way_bypass_14; // @[Reg.scala 17:22]
    end
    if (read_way_bypass_14) begin // @[Reg.scala 17:18]
      if (s1_way_wen_6_1_REG & s1_way_waddr_6_1_r == io_read_1_bits_idx) begin // @[AsynchronousMetaArray.scala 134:85]
        io_resp_1_6_r1 <= s1_way_wdata_6_1_r; // @[AsynchronousMetaArray.scala 136:25]
      end else begin
        io_resp_1_6_r1 <= s1_way_wdata_6_0_r;
      end
    end
    if (io_read_1_valid) begin // @[Reg.scala 17:18]
      io_resp_1_6_r2 <= io_read_1_bits_idx; // @[Reg.scala 17:22]
    end
    if (io_read_1_valid) begin // @[Reg.scala 17:18]
      io_resp_1_7_r <= read_way_bypass_15; // @[Reg.scala 17:22]
    end
    if (read_way_bypass_15) begin // @[Reg.scala 17:18]
      if (s1_way_wen_7_1_REG & s1_way_waddr_7_1_r == io_read_1_bits_idx) begin // @[AsynchronousMetaArray.scala 134:85]
        io_resp_1_7_r1 <= s1_way_wdata_7_1_r; // @[AsynchronousMetaArray.scala 136:25]
      end else begin
        io_resp_1_7_r1 <= s1_way_wdata_7_0_r;
      end
    end
    if (io_read_1_valid) begin // @[Reg.scala 17:18]
      io_resp_1_7_r2 <= io_read_1_bits_idx; // @[Reg.scala 17:22]
    end
    if (io_read_2_valid) begin // @[Reg.scala 17:18]
      io_resp_2_0_r <= read_way_bypass_16; // @[Reg.scala 17:22]
    end
    if (read_way_bypass_16) begin // @[Reg.scala 17:18]
      if (s1_way_wen_0_1_REG & s1_way_waddr_0_1_r == io_read_2_bits_idx) begin // @[AsynchronousMetaArray.scala 134:85]
        io_resp_2_0_r1 <= s1_way_wdata_0_1_r; // @[AsynchronousMetaArray.scala 136:25]
      end else begin
        io_resp_2_0_r1 <= s1_way_wdata_0_0_r;
      end
    end
    if (io_read_2_valid) begin // @[Reg.scala 17:18]
      io_resp_2_0_r2 <= io_read_2_bits_idx; // @[Reg.scala 17:22]
    end
    if (io_read_2_valid) begin // @[Reg.scala 17:18]
      io_resp_2_1_r <= read_way_bypass_17; // @[Reg.scala 17:22]
    end
    if (read_way_bypass_17) begin // @[Reg.scala 17:18]
      if (s1_way_wen_1_1_REG & s1_way_waddr_1_1_r == io_read_2_bits_idx) begin // @[AsynchronousMetaArray.scala 134:85]
        io_resp_2_1_r1 <= s1_way_wdata_1_1_r; // @[AsynchronousMetaArray.scala 136:25]
      end else begin
        io_resp_2_1_r1 <= s1_way_wdata_1_0_r;
      end
    end
    if (io_read_2_valid) begin // @[Reg.scala 17:18]
      io_resp_2_1_r2 <= io_read_2_bits_idx; // @[Reg.scala 17:22]
    end
    if (io_read_2_valid) begin // @[Reg.scala 17:18]
      io_resp_2_2_r <= read_way_bypass_18; // @[Reg.scala 17:22]
    end
    if (read_way_bypass_18) begin // @[Reg.scala 17:18]
      if (s1_way_wen_2_1_REG & s1_way_waddr_2_1_r == io_read_2_bits_idx) begin // @[AsynchronousMetaArray.scala 134:85]
        io_resp_2_2_r1 <= s1_way_wdata_2_1_r; // @[AsynchronousMetaArray.scala 136:25]
      end else begin
        io_resp_2_2_r1 <= s1_way_wdata_2_0_r;
      end
    end
    if (io_read_2_valid) begin // @[Reg.scala 17:18]
      io_resp_2_2_r2 <= io_read_2_bits_idx; // @[Reg.scala 17:22]
    end
    if (io_read_2_valid) begin // @[Reg.scala 17:18]
      io_resp_2_3_r <= read_way_bypass_19; // @[Reg.scala 17:22]
    end
    if (read_way_bypass_19) begin // @[Reg.scala 17:18]
      if (s1_way_wen_3_1_REG & s1_way_waddr_3_1_r == io_read_2_bits_idx) begin // @[AsynchronousMetaArray.scala 134:85]
        io_resp_2_3_r1 <= s1_way_wdata_3_1_r; // @[AsynchronousMetaArray.scala 136:25]
      end else begin
        io_resp_2_3_r1 <= s1_way_wdata_3_0_r;
      end
    end
    if (io_read_2_valid) begin // @[Reg.scala 17:18]
      io_resp_2_3_r2 <= io_read_2_bits_idx; // @[Reg.scala 17:22]
    end
    if (io_read_2_valid) begin // @[Reg.scala 17:18]
      io_resp_2_4_r <= read_way_bypass_20; // @[Reg.scala 17:22]
    end
    if (read_way_bypass_20) begin // @[Reg.scala 17:18]
      if (s1_way_wen_4_1_REG & s1_way_waddr_4_1_r == io_read_2_bits_idx) begin // @[AsynchronousMetaArray.scala 134:85]
        io_resp_2_4_r1 <= s1_way_wdata_4_1_r; // @[AsynchronousMetaArray.scala 136:25]
      end else begin
        io_resp_2_4_r1 <= s1_way_wdata_4_0_r;
      end
    end
    if (io_read_2_valid) begin // @[Reg.scala 17:18]
      io_resp_2_4_r2 <= io_read_2_bits_idx; // @[Reg.scala 17:22]
    end
    if (io_read_2_valid) begin // @[Reg.scala 17:18]
      io_resp_2_5_r <= read_way_bypass_21; // @[Reg.scala 17:22]
    end
    if (read_way_bypass_21) begin // @[Reg.scala 17:18]
      if (s1_way_wen_5_1_REG & s1_way_waddr_5_1_r == io_read_2_bits_idx) begin // @[AsynchronousMetaArray.scala 134:85]
        io_resp_2_5_r1 <= s1_way_wdata_5_1_r; // @[AsynchronousMetaArray.scala 136:25]
      end else begin
        io_resp_2_5_r1 <= s1_way_wdata_5_0_r;
      end
    end
    if (io_read_2_valid) begin // @[Reg.scala 17:18]
      io_resp_2_5_r2 <= io_read_2_bits_idx; // @[Reg.scala 17:22]
    end
    if (io_read_2_valid) begin // @[Reg.scala 17:18]
      io_resp_2_6_r <= read_way_bypass_22; // @[Reg.scala 17:22]
    end
    if (read_way_bypass_22) begin // @[Reg.scala 17:18]
      if (s1_way_wen_6_1_REG & s1_way_waddr_6_1_r == io_read_2_bits_idx) begin // @[AsynchronousMetaArray.scala 134:85]
        io_resp_2_6_r1 <= s1_way_wdata_6_1_r; // @[AsynchronousMetaArray.scala 136:25]
      end else begin
        io_resp_2_6_r1 <= s1_way_wdata_6_0_r;
      end
    end
    if (io_read_2_valid) begin // @[Reg.scala 17:18]
      io_resp_2_6_r2 <= io_read_2_bits_idx; // @[Reg.scala 17:22]
    end
    if (io_read_2_valid) begin // @[Reg.scala 17:18]
      io_resp_2_7_r <= read_way_bypass_23; // @[Reg.scala 17:22]
    end
    if (read_way_bypass_23) begin // @[Reg.scala 17:18]
      if (s1_way_wen_7_1_REG & s1_way_waddr_7_1_r == io_read_2_bits_idx) begin // @[AsynchronousMetaArray.scala 134:85]
        io_resp_2_7_r1 <= s1_way_wdata_7_1_r; // @[AsynchronousMetaArray.scala 136:25]
      end else begin
        io_resp_2_7_r1 <= s1_way_wdata_7_0_r;
      end
    end
    if (io_read_2_valid) begin // @[Reg.scala 17:18]
      io_resp_2_7_r2 <= io_read_2_bits_idx; // @[Reg.scala 17:22]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_0_0 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_0_1_REG) begin
      if (6'h0 == s1_way_waddr_0_1_r) begin
        meta_array_0_0 <= s1_way_wdata_0_1_r;
      end else begin
        meta_array_0_0 <= _GEN_1770;
      end
    end else begin
      meta_array_0_0 <= _GEN_1770;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_0_1 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_1_1_REG) begin
      if (6'h0 == s1_way_waddr_1_1_r) begin
        meta_array_0_1 <= s1_way_wdata_1_1_r;
      end else begin
        meta_array_0_1 <= _GEN_1900;
      end
    end else begin
      meta_array_0_1 <= _GEN_1900;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_0_2 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_2_1_REG) begin
      if (6'h0 == s1_way_waddr_2_1_r) begin
        meta_array_0_2 <= s1_way_wdata_2_1_r;
      end else begin
        meta_array_0_2 <= _GEN_2030;
      end
    end else begin
      meta_array_0_2 <= _GEN_2030;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_0_3 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_3_1_REG) begin
      if (6'h0 == s1_way_waddr_3_1_r) begin
        meta_array_0_3 <= s1_way_wdata_3_1_r;
      end else begin
        meta_array_0_3 <= _GEN_2160;
      end
    end else begin
      meta_array_0_3 <= _GEN_2160;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_0_4 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_4_1_REG) begin
      if (6'h0 == s1_way_waddr_4_1_r) begin
        meta_array_0_4 <= s1_way_wdata_4_1_r;
      end else begin
        meta_array_0_4 <= _GEN_2290;
      end
    end else begin
      meta_array_0_4 <= _GEN_2290;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_0_5 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_5_1_REG) begin
      if (6'h0 == s1_way_waddr_5_1_r) begin
        meta_array_0_5 <= s1_way_wdata_5_1_r;
      end else begin
        meta_array_0_5 <= _GEN_2420;
      end
    end else begin
      meta_array_0_5 <= _GEN_2420;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_0_6 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_6_1_REG) begin
      if (6'h0 == s1_way_waddr_6_1_r) begin
        meta_array_0_6 <= s1_way_wdata_6_1_r;
      end else begin
        meta_array_0_6 <= _GEN_2550;
      end
    end else begin
      meta_array_0_6 <= _GEN_2550;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_0_7 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_7_1_REG) begin
      if (6'h0 == s1_way_waddr_7_1_r) begin
        meta_array_0_7 <= s1_way_wdata_7_1_r;
      end else begin
        meta_array_0_7 <= _GEN_2680;
      end
    end else begin
      meta_array_0_7 <= _GEN_2680;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_1_0 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_0_1_REG) begin
      if (6'h1 == s1_way_waddr_0_1_r) begin
        meta_array_1_0 <= s1_way_wdata_0_1_r;
      end else begin
        meta_array_1_0 <= _GEN_1771;
      end
    end else begin
      meta_array_1_0 <= _GEN_1771;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_1_1 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_1_1_REG) begin
      if (6'h1 == s1_way_waddr_1_1_r) begin
        meta_array_1_1 <= s1_way_wdata_1_1_r;
      end else begin
        meta_array_1_1 <= _GEN_1901;
      end
    end else begin
      meta_array_1_1 <= _GEN_1901;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_1_2 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_2_1_REG) begin
      if (6'h1 == s1_way_waddr_2_1_r) begin
        meta_array_1_2 <= s1_way_wdata_2_1_r;
      end else begin
        meta_array_1_2 <= _GEN_2031;
      end
    end else begin
      meta_array_1_2 <= _GEN_2031;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_1_3 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_3_1_REG) begin
      if (6'h1 == s1_way_waddr_3_1_r) begin
        meta_array_1_3 <= s1_way_wdata_3_1_r;
      end else begin
        meta_array_1_3 <= _GEN_2161;
      end
    end else begin
      meta_array_1_3 <= _GEN_2161;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_1_4 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_4_1_REG) begin
      if (6'h1 == s1_way_waddr_4_1_r) begin
        meta_array_1_4 <= s1_way_wdata_4_1_r;
      end else begin
        meta_array_1_4 <= _GEN_2291;
      end
    end else begin
      meta_array_1_4 <= _GEN_2291;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_1_5 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_5_1_REG) begin
      if (6'h1 == s1_way_waddr_5_1_r) begin
        meta_array_1_5 <= s1_way_wdata_5_1_r;
      end else begin
        meta_array_1_5 <= _GEN_2421;
      end
    end else begin
      meta_array_1_5 <= _GEN_2421;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_1_6 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_6_1_REG) begin
      if (6'h1 == s1_way_waddr_6_1_r) begin
        meta_array_1_6 <= s1_way_wdata_6_1_r;
      end else begin
        meta_array_1_6 <= _GEN_2551;
      end
    end else begin
      meta_array_1_6 <= _GEN_2551;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_1_7 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_7_1_REG) begin
      if (6'h1 == s1_way_waddr_7_1_r) begin
        meta_array_1_7 <= s1_way_wdata_7_1_r;
      end else begin
        meta_array_1_7 <= _GEN_2681;
      end
    end else begin
      meta_array_1_7 <= _GEN_2681;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_2_0 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_0_1_REG) begin
      if (6'h2 == s1_way_waddr_0_1_r) begin
        meta_array_2_0 <= s1_way_wdata_0_1_r;
      end else begin
        meta_array_2_0 <= _GEN_1772;
      end
    end else begin
      meta_array_2_0 <= _GEN_1772;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_2_1 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_1_1_REG) begin
      if (6'h2 == s1_way_waddr_1_1_r) begin
        meta_array_2_1 <= s1_way_wdata_1_1_r;
      end else begin
        meta_array_2_1 <= _GEN_1902;
      end
    end else begin
      meta_array_2_1 <= _GEN_1902;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_2_2 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_2_1_REG) begin
      if (6'h2 == s1_way_waddr_2_1_r) begin
        meta_array_2_2 <= s1_way_wdata_2_1_r;
      end else begin
        meta_array_2_2 <= _GEN_2032;
      end
    end else begin
      meta_array_2_2 <= _GEN_2032;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_2_3 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_3_1_REG) begin
      if (6'h2 == s1_way_waddr_3_1_r) begin
        meta_array_2_3 <= s1_way_wdata_3_1_r;
      end else begin
        meta_array_2_3 <= _GEN_2162;
      end
    end else begin
      meta_array_2_3 <= _GEN_2162;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_2_4 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_4_1_REG) begin
      if (6'h2 == s1_way_waddr_4_1_r) begin
        meta_array_2_4 <= s1_way_wdata_4_1_r;
      end else begin
        meta_array_2_4 <= _GEN_2292;
      end
    end else begin
      meta_array_2_4 <= _GEN_2292;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_2_5 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_5_1_REG) begin
      if (6'h2 == s1_way_waddr_5_1_r) begin
        meta_array_2_5 <= s1_way_wdata_5_1_r;
      end else begin
        meta_array_2_5 <= _GEN_2422;
      end
    end else begin
      meta_array_2_5 <= _GEN_2422;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_2_6 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_6_1_REG) begin
      if (6'h2 == s1_way_waddr_6_1_r) begin
        meta_array_2_6 <= s1_way_wdata_6_1_r;
      end else begin
        meta_array_2_6 <= _GEN_2552;
      end
    end else begin
      meta_array_2_6 <= _GEN_2552;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_2_7 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_7_1_REG) begin
      if (6'h2 == s1_way_waddr_7_1_r) begin
        meta_array_2_7 <= s1_way_wdata_7_1_r;
      end else begin
        meta_array_2_7 <= _GEN_2682;
      end
    end else begin
      meta_array_2_7 <= _GEN_2682;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_3_0 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_0_1_REG) begin
      if (6'h3 == s1_way_waddr_0_1_r) begin
        meta_array_3_0 <= s1_way_wdata_0_1_r;
      end else begin
        meta_array_3_0 <= _GEN_1773;
      end
    end else begin
      meta_array_3_0 <= _GEN_1773;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_3_1 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_1_1_REG) begin
      if (6'h3 == s1_way_waddr_1_1_r) begin
        meta_array_3_1 <= s1_way_wdata_1_1_r;
      end else begin
        meta_array_3_1 <= _GEN_1903;
      end
    end else begin
      meta_array_3_1 <= _GEN_1903;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_3_2 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_2_1_REG) begin
      if (6'h3 == s1_way_waddr_2_1_r) begin
        meta_array_3_2 <= s1_way_wdata_2_1_r;
      end else begin
        meta_array_3_2 <= _GEN_2033;
      end
    end else begin
      meta_array_3_2 <= _GEN_2033;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_3_3 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_3_1_REG) begin
      if (6'h3 == s1_way_waddr_3_1_r) begin
        meta_array_3_3 <= s1_way_wdata_3_1_r;
      end else begin
        meta_array_3_3 <= _GEN_2163;
      end
    end else begin
      meta_array_3_3 <= _GEN_2163;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_3_4 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_4_1_REG) begin
      if (6'h3 == s1_way_waddr_4_1_r) begin
        meta_array_3_4 <= s1_way_wdata_4_1_r;
      end else begin
        meta_array_3_4 <= _GEN_2293;
      end
    end else begin
      meta_array_3_4 <= _GEN_2293;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_3_5 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_5_1_REG) begin
      if (6'h3 == s1_way_waddr_5_1_r) begin
        meta_array_3_5 <= s1_way_wdata_5_1_r;
      end else begin
        meta_array_3_5 <= _GEN_2423;
      end
    end else begin
      meta_array_3_5 <= _GEN_2423;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_3_6 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_6_1_REG) begin
      if (6'h3 == s1_way_waddr_6_1_r) begin
        meta_array_3_6 <= s1_way_wdata_6_1_r;
      end else begin
        meta_array_3_6 <= _GEN_2553;
      end
    end else begin
      meta_array_3_6 <= _GEN_2553;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_3_7 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_7_1_REG) begin
      if (6'h3 == s1_way_waddr_7_1_r) begin
        meta_array_3_7 <= s1_way_wdata_7_1_r;
      end else begin
        meta_array_3_7 <= _GEN_2683;
      end
    end else begin
      meta_array_3_7 <= _GEN_2683;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_4_0 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_0_1_REG) begin
      if (6'h4 == s1_way_waddr_0_1_r) begin
        meta_array_4_0 <= s1_way_wdata_0_1_r;
      end else begin
        meta_array_4_0 <= _GEN_1774;
      end
    end else begin
      meta_array_4_0 <= _GEN_1774;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_4_1 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_1_1_REG) begin
      if (6'h4 == s1_way_waddr_1_1_r) begin
        meta_array_4_1 <= s1_way_wdata_1_1_r;
      end else begin
        meta_array_4_1 <= _GEN_1904;
      end
    end else begin
      meta_array_4_1 <= _GEN_1904;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_4_2 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_2_1_REG) begin
      if (6'h4 == s1_way_waddr_2_1_r) begin
        meta_array_4_2 <= s1_way_wdata_2_1_r;
      end else begin
        meta_array_4_2 <= _GEN_2034;
      end
    end else begin
      meta_array_4_2 <= _GEN_2034;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_4_3 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_3_1_REG) begin
      if (6'h4 == s1_way_waddr_3_1_r) begin
        meta_array_4_3 <= s1_way_wdata_3_1_r;
      end else begin
        meta_array_4_3 <= _GEN_2164;
      end
    end else begin
      meta_array_4_3 <= _GEN_2164;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_4_4 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_4_1_REG) begin
      if (6'h4 == s1_way_waddr_4_1_r) begin
        meta_array_4_4 <= s1_way_wdata_4_1_r;
      end else begin
        meta_array_4_4 <= _GEN_2294;
      end
    end else begin
      meta_array_4_4 <= _GEN_2294;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_4_5 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_5_1_REG) begin
      if (6'h4 == s1_way_waddr_5_1_r) begin
        meta_array_4_5 <= s1_way_wdata_5_1_r;
      end else begin
        meta_array_4_5 <= _GEN_2424;
      end
    end else begin
      meta_array_4_5 <= _GEN_2424;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_4_6 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_6_1_REG) begin
      if (6'h4 == s1_way_waddr_6_1_r) begin
        meta_array_4_6 <= s1_way_wdata_6_1_r;
      end else begin
        meta_array_4_6 <= _GEN_2554;
      end
    end else begin
      meta_array_4_6 <= _GEN_2554;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_4_7 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_7_1_REG) begin
      if (6'h4 == s1_way_waddr_7_1_r) begin
        meta_array_4_7 <= s1_way_wdata_7_1_r;
      end else begin
        meta_array_4_7 <= _GEN_2684;
      end
    end else begin
      meta_array_4_7 <= _GEN_2684;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_5_0 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_0_1_REG) begin
      if (6'h5 == s1_way_waddr_0_1_r) begin
        meta_array_5_0 <= s1_way_wdata_0_1_r;
      end else begin
        meta_array_5_0 <= _GEN_1775;
      end
    end else begin
      meta_array_5_0 <= _GEN_1775;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_5_1 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_1_1_REG) begin
      if (6'h5 == s1_way_waddr_1_1_r) begin
        meta_array_5_1 <= s1_way_wdata_1_1_r;
      end else begin
        meta_array_5_1 <= _GEN_1905;
      end
    end else begin
      meta_array_5_1 <= _GEN_1905;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_5_2 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_2_1_REG) begin
      if (6'h5 == s1_way_waddr_2_1_r) begin
        meta_array_5_2 <= s1_way_wdata_2_1_r;
      end else begin
        meta_array_5_2 <= _GEN_2035;
      end
    end else begin
      meta_array_5_2 <= _GEN_2035;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_5_3 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_3_1_REG) begin
      if (6'h5 == s1_way_waddr_3_1_r) begin
        meta_array_5_3 <= s1_way_wdata_3_1_r;
      end else begin
        meta_array_5_3 <= _GEN_2165;
      end
    end else begin
      meta_array_5_3 <= _GEN_2165;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_5_4 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_4_1_REG) begin
      if (6'h5 == s1_way_waddr_4_1_r) begin
        meta_array_5_4 <= s1_way_wdata_4_1_r;
      end else begin
        meta_array_5_4 <= _GEN_2295;
      end
    end else begin
      meta_array_5_4 <= _GEN_2295;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_5_5 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_5_1_REG) begin
      if (6'h5 == s1_way_waddr_5_1_r) begin
        meta_array_5_5 <= s1_way_wdata_5_1_r;
      end else begin
        meta_array_5_5 <= _GEN_2425;
      end
    end else begin
      meta_array_5_5 <= _GEN_2425;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_5_6 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_6_1_REG) begin
      if (6'h5 == s1_way_waddr_6_1_r) begin
        meta_array_5_6 <= s1_way_wdata_6_1_r;
      end else begin
        meta_array_5_6 <= _GEN_2555;
      end
    end else begin
      meta_array_5_6 <= _GEN_2555;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_5_7 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_7_1_REG) begin
      if (6'h5 == s1_way_waddr_7_1_r) begin
        meta_array_5_7 <= s1_way_wdata_7_1_r;
      end else begin
        meta_array_5_7 <= _GEN_2685;
      end
    end else begin
      meta_array_5_7 <= _GEN_2685;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_6_0 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_0_1_REG) begin
      if (6'h6 == s1_way_waddr_0_1_r) begin
        meta_array_6_0 <= s1_way_wdata_0_1_r;
      end else begin
        meta_array_6_0 <= _GEN_1776;
      end
    end else begin
      meta_array_6_0 <= _GEN_1776;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_6_1 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_1_1_REG) begin
      if (6'h6 == s1_way_waddr_1_1_r) begin
        meta_array_6_1 <= s1_way_wdata_1_1_r;
      end else begin
        meta_array_6_1 <= _GEN_1906;
      end
    end else begin
      meta_array_6_1 <= _GEN_1906;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_6_2 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_2_1_REG) begin
      if (6'h6 == s1_way_waddr_2_1_r) begin
        meta_array_6_2 <= s1_way_wdata_2_1_r;
      end else begin
        meta_array_6_2 <= _GEN_2036;
      end
    end else begin
      meta_array_6_2 <= _GEN_2036;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_6_3 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_3_1_REG) begin
      if (6'h6 == s1_way_waddr_3_1_r) begin
        meta_array_6_3 <= s1_way_wdata_3_1_r;
      end else begin
        meta_array_6_3 <= _GEN_2166;
      end
    end else begin
      meta_array_6_3 <= _GEN_2166;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_6_4 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_4_1_REG) begin
      if (6'h6 == s1_way_waddr_4_1_r) begin
        meta_array_6_4 <= s1_way_wdata_4_1_r;
      end else begin
        meta_array_6_4 <= _GEN_2296;
      end
    end else begin
      meta_array_6_4 <= _GEN_2296;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_6_5 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_5_1_REG) begin
      if (6'h6 == s1_way_waddr_5_1_r) begin
        meta_array_6_5 <= s1_way_wdata_5_1_r;
      end else begin
        meta_array_6_5 <= _GEN_2426;
      end
    end else begin
      meta_array_6_5 <= _GEN_2426;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_6_6 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_6_1_REG) begin
      if (6'h6 == s1_way_waddr_6_1_r) begin
        meta_array_6_6 <= s1_way_wdata_6_1_r;
      end else begin
        meta_array_6_6 <= _GEN_2556;
      end
    end else begin
      meta_array_6_6 <= _GEN_2556;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_6_7 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_7_1_REG) begin
      if (6'h6 == s1_way_waddr_7_1_r) begin
        meta_array_6_7 <= s1_way_wdata_7_1_r;
      end else begin
        meta_array_6_7 <= _GEN_2686;
      end
    end else begin
      meta_array_6_7 <= _GEN_2686;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_7_0 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_0_1_REG) begin
      if (6'h7 == s1_way_waddr_0_1_r) begin
        meta_array_7_0 <= s1_way_wdata_0_1_r;
      end else begin
        meta_array_7_0 <= _GEN_1777;
      end
    end else begin
      meta_array_7_0 <= _GEN_1777;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_7_1 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_1_1_REG) begin
      if (6'h7 == s1_way_waddr_1_1_r) begin
        meta_array_7_1 <= s1_way_wdata_1_1_r;
      end else begin
        meta_array_7_1 <= _GEN_1907;
      end
    end else begin
      meta_array_7_1 <= _GEN_1907;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_7_2 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_2_1_REG) begin
      if (6'h7 == s1_way_waddr_2_1_r) begin
        meta_array_7_2 <= s1_way_wdata_2_1_r;
      end else begin
        meta_array_7_2 <= _GEN_2037;
      end
    end else begin
      meta_array_7_2 <= _GEN_2037;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_7_3 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_3_1_REG) begin
      if (6'h7 == s1_way_waddr_3_1_r) begin
        meta_array_7_3 <= s1_way_wdata_3_1_r;
      end else begin
        meta_array_7_3 <= _GEN_2167;
      end
    end else begin
      meta_array_7_3 <= _GEN_2167;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_7_4 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_4_1_REG) begin
      if (6'h7 == s1_way_waddr_4_1_r) begin
        meta_array_7_4 <= s1_way_wdata_4_1_r;
      end else begin
        meta_array_7_4 <= _GEN_2297;
      end
    end else begin
      meta_array_7_4 <= _GEN_2297;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_7_5 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_5_1_REG) begin
      if (6'h7 == s1_way_waddr_5_1_r) begin
        meta_array_7_5 <= s1_way_wdata_5_1_r;
      end else begin
        meta_array_7_5 <= _GEN_2427;
      end
    end else begin
      meta_array_7_5 <= _GEN_2427;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_7_6 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_6_1_REG) begin
      if (6'h7 == s1_way_waddr_6_1_r) begin
        meta_array_7_6 <= s1_way_wdata_6_1_r;
      end else begin
        meta_array_7_6 <= _GEN_2557;
      end
    end else begin
      meta_array_7_6 <= _GEN_2557;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_7_7 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_7_1_REG) begin
      if (6'h7 == s1_way_waddr_7_1_r) begin
        meta_array_7_7 <= s1_way_wdata_7_1_r;
      end else begin
        meta_array_7_7 <= _GEN_2687;
      end
    end else begin
      meta_array_7_7 <= _GEN_2687;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_8_0 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_0_1_REG) begin
      if (6'h8 == s1_way_waddr_0_1_r) begin
        meta_array_8_0 <= s1_way_wdata_0_1_r;
      end else begin
        meta_array_8_0 <= _GEN_1778;
      end
    end else begin
      meta_array_8_0 <= _GEN_1778;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_8_1 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_1_1_REG) begin
      if (6'h8 == s1_way_waddr_1_1_r) begin
        meta_array_8_1 <= s1_way_wdata_1_1_r;
      end else begin
        meta_array_8_1 <= _GEN_1908;
      end
    end else begin
      meta_array_8_1 <= _GEN_1908;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_8_2 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_2_1_REG) begin
      if (6'h8 == s1_way_waddr_2_1_r) begin
        meta_array_8_2 <= s1_way_wdata_2_1_r;
      end else begin
        meta_array_8_2 <= _GEN_2038;
      end
    end else begin
      meta_array_8_2 <= _GEN_2038;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_8_3 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_3_1_REG) begin
      if (6'h8 == s1_way_waddr_3_1_r) begin
        meta_array_8_3 <= s1_way_wdata_3_1_r;
      end else begin
        meta_array_8_3 <= _GEN_2168;
      end
    end else begin
      meta_array_8_3 <= _GEN_2168;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_8_4 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_4_1_REG) begin
      if (6'h8 == s1_way_waddr_4_1_r) begin
        meta_array_8_4 <= s1_way_wdata_4_1_r;
      end else begin
        meta_array_8_4 <= _GEN_2298;
      end
    end else begin
      meta_array_8_4 <= _GEN_2298;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_8_5 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_5_1_REG) begin
      if (6'h8 == s1_way_waddr_5_1_r) begin
        meta_array_8_5 <= s1_way_wdata_5_1_r;
      end else begin
        meta_array_8_5 <= _GEN_2428;
      end
    end else begin
      meta_array_8_5 <= _GEN_2428;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_8_6 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_6_1_REG) begin
      if (6'h8 == s1_way_waddr_6_1_r) begin
        meta_array_8_6 <= s1_way_wdata_6_1_r;
      end else begin
        meta_array_8_6 <= _GEN_2558;
      end
    end else begin
      meta_array_8_6 <= _GEN_2558;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_8_7 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_7_1_REG) begin
      if (6'h8 == s1_way_waddr_7_1_r) begin
        meta_array_8_7 <= s1_way_wdata_7_1_r;
      end else begin
        meta_array_8_7 <= _GEN_2688;
      end
    end else begin
      meta_array_8_7 <= _GEN_2688;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_9_0 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_0_1_REG) begin
      if (6'h9 == s1_way_waddr_0_1_r) begin
        meta_array_9_0 <= s1_way_wdata_0_1_r;
      end else begin
        meta_array_9_0 <= _GEN_1779;
      end
    end else begin
      meta_array_9_0 <= _GEN_1779;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_9_1 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_1_1_REG) begin
      if (6'h9 == s1_way_waddr_1_1_r) begin
        meta_array_9_1 <= s1_way_wdata_1_1_r;
      end else begin
        meta_array_9_1 <= _GEN_1909;
      end
    end else begin
      meta_array_9_1 <= _GEN_1909;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_9_2 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_2_1_REG) begin
      if (6'h9 == s1_way_waddr_2_1_r) begin
        meta_array_9_2 <= s1_way_wdata_2_1_r;
      end else begin
        meta_array_9_2 <= _GEN_2039;
      end
    end else begin
      meta_array_9_2 <= _GEN_2039;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_9_3 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_3_1_REG) begin
      if (6'h9 == s1_way_waddr_3_1_r) begin
        meta_array_9_3 <= s1_way_wdata_3_1_r;
      end else begin
        meta_array_9_3 <= _GEN_2169;
      end
    end else begin
      meta_array_9_3 <= _GEN_2169;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_9_4 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_4_1_REG) begin
      if (6'h9 == s1_way_waddr_4_1_r) begin
        meta_array_9_4 <= s1_way_wdata_4_1_r;
      end else begin
        meta_array_9_4 <= _GEN_2299;
      end
    end else begin
      meta_array_9_4 <= _GEN_2299;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_9_5 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_5_1_REG) begin
      if (6'h9 == s1_way_waddr_5_1_r) begin
        meta_array_9_5 <= s1_way_wdata_5_1_r;
      end else begin
        meta_array_9_5 <= _GEN_2429;
      end
    end else begin
      meta_array_9_5 <= _GEN_2429;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_9_6 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_6_1_REG) begin
      if (6'h9 == s1_way_waddr_6_1_r) begin
        meta_array_9_6 <= s1_way_wdata_6_1_r;
      end else begin
        meta_array_9_6 <= _GEN_2559;
      end
    end else begin
      meta_array_9_6 <= _GEN_2559;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_9_7 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_7_1_REG) begin
      if (6'h9 == s1_way_waddr_7_1_r) begin
        meta_array_9_7 <= s1_way_wdata_7_1_r;
      end else begin
        meta_array_9_7 <= _GEN_2689;
      end
    end else begin
      meta_array_9_7 <= _GEN_2689;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_10_0 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_0_1_REG) begin
      if (6'ha == s1_way_waddr_0_1_r) begin
        meta_array_10_0 <= s1_way_wdata_0_1_r;
      end else begin
        meta_array_10_0 <= _GEN_1780;
      end
    end else begin
      meta_array_10_0 <= _GEN_1780;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_10_1 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_1_1_REG) begin
      if (6'ha == s1_way_waddr_1_1_r) begin
        meta_array_10_1 <= s1_way_wdata_1_1_r;
      end else begin
        meta_array_10_1 <= _GEN_1910;
      end
    end else begin
      meta_array_10_1 <= _GEN_1910;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_10_2 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_2_1_REG) begin
      if (6'ha == s1_way_waddr_2_1_r) begin
        meta_array_10_2 <= s1_way_wdata_2_1_r;
      end else begin
        meta_array_10_2 <= _GEN_2040;
      end
    end else begin
      meta_array_10_2 <= _GEN_2040;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_10_3 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_3_1_REG) begin
      if (6'ha == s1_way_waddr_3_1_r) begin
        meta_array_10_3 <= s1_way_wdata_3_1_r;
      end else begin
        meta_array_10_3 <= _GEN_2170;
      end
    end else begin
      meta_array_10_3 <= _GEN_2170;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_10_4 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_4_1_REG) begin
      if (6'ha == s1_way_waddr_4_1_r) begin
        meta_array_10_4 <= s1_way_wdata_4_1_r;
      end else begin
        meta_array_10_4 <= _GEN_2300;
      end
    end else begin
      meta_array_10_4 <= _GEN_2300;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_10_5 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_5_1_REG) begin
      if (6'ha == s1_way_waddr_5_1_r) begin
        meta_array_10_5 <= s1_way_wdata_5_1_r;
      end else begin
        meta_array_10_5 <= _GEN_2430;
      end
    end else begin
      meta_array_10_5 <= _GEN_2430;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_10_6 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_6_1_REG) begin
      if (6'ha == s1_way_waddr_6_1_r) begin
        meta_array_10_6 <= s1_way_wdata_6_1_r;
      end else begin
        meta_array_10_6 <= _GEN_2560;
      end
    end else begin
      meta_array_10_6 <= _GEN_2560;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_10_7 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_7_1_REG) begin
      if (6'ha == s1_way_waddr_7_1_r) begin
        meta_array_10_7 <= s1_way_wdata_7_1_r;
      end else begin
        meta_array_10_7 <= _GEN_2690;
      end
    end else begin
      meta_array_10_7 <= _GEN_2690;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_11_0 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_0_1_REG) begin
      if (6'hb == s1_way_waddr_0_1_r) begin
        meta_array_11_0 <= s1_way_wdata_0_1_r;
      end else begin
        meta_array_11_0 <= _GEN_1781;
      end
    end else begin
      meta_array_11_0 <= _GEN_1781;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_11_1 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_1_1_REG) begin
      if (6'hb == s1_way_waddr_1_1_r) begin
        meta_array_11_1 <= s1_way_wdata_1_1_r;
      end else begin
        meta_array_11_1 <= _GEN_1911;
      end
    end else begin
      meta_array_11_1 <= _GEN_1911;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_11_2 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_2_1_REG) begin
      if (6'hb == s1_way_waddr_2_1_r) begin
        meta_array_11_2 <= s1_way_wdata_2_1_r;
      end else begin
        meta_array_11_2 <= _GEN_2041;
      end
    end else begin
      meta_array_11_2 <= _GEN_2041;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_11_3 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_3_1_REG) begin
      if (6'hb == s1_way_waddr_3_1_r) begin
        meta_array_11_3 <= s1_way_wdata_3_1_r;
      end else begin
        meta_array_11_3 <= _GEN_2171;
      end
    end else begin
      meta_array_11_3 <= _GEN_2171;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_11_4 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_4_1_REG) begin
      if (6'hb == s1_way_waddr_4_1_r) begin
        meta_array_11_4 <= s1_way_wdata_4_1_r;
      end else begin
        meta_array_11_4 <= _GEN_2301;
      end
    end else begin
      meta_array_11_4 <= _GEN_2301;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_11_5 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_5_1_REG) begin
      if (6'hb == s1_way_waddr_5_1_r) begin
        meta_array_11_5 <= s1_way_wdata_5_1_r;
      end else begin
        meta_array_11_5 <= _GEN_2431;
      end
    end else begin
      meta_array_11_5 <= _GEN_2431;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_11_6 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_6_1_REG) begin
      if (6'hb == s1_way_waddr_6_1_r) begin
        meta_array_11_6 <= s1_way_wdata_6_1_r;
      end else begin
        meta_array_11_6 <= _GEN_2561;
      end
    end else begin
      meta_array_11_6 <= _GEN_2561;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_11_7 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_7_1_REG) begin
      if (6'hb == s1_way_waddr_7_1_r) begin
        meta_array_11_7 <= s1_way_wdata_7_1_r;
      end else begin
        meta_array_11_7 <= _GEN_2691;
      end
    end else begin
      meta_array_11_7 <= _GEN_2691;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_12_0 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_0_1_REG) begin
      if (6'hc == s1_way_waddr_0_1_r) begin
        meta_array_12_0 <= s1_way_wdata_0_1_r;
      end else begin
        meta_array_12_0 <= _GEN_1782;
      end
    end else begin
      meta_array_12_0 <= _GEN_1782;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_12_1 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_1_1_REG) begin
      if (6'hc == s1_way_waddr_1_1_r) begin
        meta_array_12_1 <= s1_way_wdata_1_1_r;
      end else begin
        meta_array_12_1 <= _GEN_1912;
      end
    end else begin
      meta_array_12_1 <= _GEN_1912;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_12_2 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_2_1_REG) begin
      if (6'hc == s1_way_waddr_2_1_r) begin
        meta_array_12_2 <= s1_way_wdata_2_1_r;
      end else begin
        meta_array_12_2 <= _GEN_2042;
      end
    end else begin
      meta_array_12_2 <= _GEN_2042;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_12_3 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_3_1_REG) begin
      if (6'hc == s1_way_waddr_3_1_r) begin
        meta_array_12_3 <= s1_way_wdata_3_1_r;
      end else begin
        meta_array_12_3 <= _GEN_2172;
      end
    end else begin
      meta_array_12_3 <= _GEN_2172;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_12_4 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_4_1_REG) begin
      if (6'hc == s1_way_waddr_4_1_r) begin
        meta_array_12_4 <= s1_way_wdata_4_1_r;
      end else begin
        meta_array_12_4 <= _GEN_2302;
      end
    end else begin
      meta_array_12_4 <= _GEN_2302;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_12_5 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_5_1_REG) begin
      if (6'hc == s1_way_waddr_5_1_r) begin
        meta_array_12_5 <= s1_way_wdata_5_1_r;
      end else begin
        meta_array_12_5 <= _GEN_2432;
      end
    end else begin
      meta_array_12_5 <= _GEN_2432;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_12_6 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_6_1_REG) begin
      if (6'hc == s1_way_waddr_6_1_r) begin
        meta_array_12_6 <= s1_way_wdata_6_1_r;
      end else begin
        meta_array_12_6 <= _GEN_2562;
      end
    end else begin
      meta_array_12_6 <= _GEN_2562;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_12_7 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_7_1_REG) begin
      if (6'hc == s1_way_waddr_7_1_r) begin
        meta_array_12_7 <= s1_way_wdata_7_1_r;
      end else begin
        meta_array_12_7 <= _GEN_2692;
      end
    end else begin
      meta_array_12_7 <= _GEN_2692;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_13_0 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_0_1_REG) begin
      if (6'hd == s1_way_waddr_0_1_r) begin
        meta_array_13_0 <= s1_way_wdata_0_1_r;
      end else begin
        meta_array_13_0 <= _GEN_1783;
      end
    end else begin
      meta_array_13_0 <= _GEN_1783;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_13_1 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_1_1_REG) begin
      if (6'hd == s1_way_waddr_1_1_r) begin
        meta_array_13_1 <= s1_way_wdata_1_1_r;
      end else begin
        meta_array_13_1 <= _GEN_1913;
      end
    end else begin
      meta_array_13_1 <= _GEN_1913;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_13_2 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_2_1_REG) begin
      if (6'hd == s1_way_waddr_2_1_r) begin
        meta_array_13_2 <= s1_way_wdata_2_1_r;
      end else begin
        meta_array_13_2 <= _GEN_2043;
      end
    end else begin
      meta_array_13_2 <= _GEN_2043;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_13_3 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_3_1_REG) begin
      if (6'hd == s1_way_waddr_3_1_r) begin
        meta_array_13_3 <= s1_way_wdata_3_1_r;
      end else begin
        meta_array_13_3 <= _GEN_2173;
      end
    end else begin
      meta_array_13_3 <= _GEN_2173;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_13_4 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_4_1_REG) begin
      if (6'hd == s1_way_waddr_4_1_r) begin
        meta_array_13_4 <= s1_way_wdata_4_1_r;
      end else begin
        meta_array_13_4 <= _GEN_2303;
      end
    end else begin
      meta_array_13_4 <= _GEN_2303;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_13_5 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_5_1_REG) begin
      if (6'hd == s1_way_waddr_5_1_r) begin
        meta_array_13_5 <= s1_way_wdata_5_1_r;
      end else begin
        meta_array_13_5 <= _GEN_2433;
      end
    end else begin
      meta_array_13_5 <= _GEN_2433;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_13_6 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_6_1_REG) begin
      if (6'hd == s1_way_waddr_6_1_r) begin
        meta_array_13_6 <= s1_way_wdata_6_1_r;
      end else begin
        meta_array_13_6 <= _GEN_2563;
      end
    end else begin
      meta_array_13_6 <= _GEN_2563;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_13_7 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_7_1_REG) begin
      if (6'hd == s1_way_waddr_7_1_r) begin
        meta_array_13_7 <= s1_way_wdata_7_1_r;
      end else begin
        meta_array_13_7 <= _GEN_2693;
      end
    end else begin
      meta_array_13_7 <= _GEN_2693;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_14_0 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_0_1_REG) begin
      if (6'he == s1_way_waddr_0_1_r) begin
        meta_array_14_0 <= s1_way_wdata_0_1_r;
      end else begin
        meta_array_14_0 <= _GEN_1784;
      end
    end else begin
      meta_array_14_0 <= _GEN_1784;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_14_1 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_1_1_REG) begin
      if (6'he == s1_way_waddr_1_1_r) begin
        meta_array_14_1 <= s1_way_wdata_1_1_r;
      end else begin
        meta_array_14_1 <= _GEN_1914;
      end
    end else begin
      meta_array_14_1 <= _GEN_1914;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_14_2 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_2_1_REG) begin
      if (6'he == s1_way_waddr_2_1_r) begin
        meta_array_14_2 <= s1_way_wdata_2_1_r;
      end else begin
        meta_array_14_2 <= _GEN_2044;
      end
    end else begin
      meta_array_14_2 <= _GEN_2044;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_14_3 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_3_1_REG) begin
      if (6'he == s1_way_waddr_3_1_r) begin
        meta_array_14_3 <= s1_way_wdata_3_1_r;
      end else begin
        meta_array_14_3 <= _GEN_2174;
      end
    end else begin
      meta_array_14_3 <= _GEN_2174;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_14_4 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_4_1_REG) begin
      if (6'he == s1_way_waddr_4_1_r) begin
        meta_array_14_4 <= s1_way_wdata_4_1_r;
      end else begin
        meta_array_14_4 <= _GEN_2304;
      end
    end else begin
      meta_array_14_4 <= _GEN_2304;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_14_5 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_5_1_REG) begin
      if (6'he == s1_way_waddr_5_1_r) begin
        meta_array_14_5 <= s1_way_wdata_5_1_r;
      end else begin
        meta_array_14_5 <= _GEN_2434;
      end
    end else begin
      meta_array_14_5 <= _GEN_2434;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_14_6 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_6_1_REG) begin
      if (6'he == s1_way_waddr_6_1_r) begin
        meta_array_14_6 <= s1_way_wdata_6_1_r;
      end else begin
        meta_array_14_6 <= _GEN_2564;
      end
    end else begin
      meta_array_14_6 <= _GEN_2564;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_14_7 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_7_1_REG) begin
      if (6'he == s1_way_waddr_7_1_r) begin
        meta_array_14_7 <= s1_way_wdata_7_1_r;
      end else begin
        meta_array_14_7 <= _GEN_2694;
      end
    end else begin
      meta_array_14_7 <= _GEN_2694;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_15_0 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_0_1_REG) begin
      if (6'hf == s1_way_waddr_0_1_r) begin
        meta_array_15_0 <= s1_way_wdata_0_1_r;
      end else begin
        meta_array_15_0 <= _GEN_1785;
      end
    end else begin
      meta_array_15_0 <= _GEN_1785;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_15_1 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_1_1_REG) begin
      if (6'hf == s1_way_waddr_1_1_r) begin
        meta_array_15_1 <= s1_way_wdata_1_1_r;
      end else begin
        meta_array_15_1 <= _GEN_1915;
      end
    end else begin
      meta_array_15_1 <= _GEN_1915;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_15_2 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_2_1_REG) begin
      if (6'hf == s1_way_waddr_2_1_r) begin
        meta_array_15_2 <= s1_way_wdata_2_1_r;
      end else begin
        meta_array_15_2 <= _GEN_2045;
      end
    end else begin
      meta_array_15_2 <= _GEN_2045;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_15_3 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_3_1_REG) begin
      if (6'hf == s1_way_waddr_3_1_r) begin
        meta_array_15_3 <= s1_way_wdata_3_1_r;
      end else begin
        meta_array_15_3 <= _GEN_2175;
      end
    end else begin
      meta_array_15_3 <= _GEN_2175;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_15_4 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_4_1_REG) begin
      if (6'hf == s1_way_waddr_4_1_r) begin
        meta_array_15_4 <= s1_way_wdata_4_1_r;
      end else begin
        meta_array_15_4 <= _GEN_2305;
      end
    end else begin
      meta_array_15_4 <= _GEN_2305;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_15_5 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_5_1_REG) begin
      if (6'hf == s1_way_waddr_5_1_r) begin
        meta_array_15_5 <= s1_way_wdata_5_1_r;
      end else begin
        meta_array_15_5 <= _GEN_2435;
      end
    end else begin
      meta_array_15_5 <= _GEN_2435;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_15_6 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_6_1_REG) begin
      if (6'hf == s1_way_waddr_6_1_r) begin
        meta_array_15_6 <= s1_way_wdata_6_1_r;
      end else begin
        meta_array_15_6 <= _GEN_2565;
      end
    end else begin
      meta_array_15_6 <= _GEN_2565;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_15_7 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_7_1_REG) begin
      if (6'hf == s1_way_waddr_7_1_r) begin
        meta_array_15_7 <= s1_way_wdata_7_1_r;
      end else begin
        meta_array_15_7 <= _GEN_2695;
      end
    end else begin
      meta_array_15_7 <= _GEN_2695;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_16_0 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_0_1_REG) begin
      if (6'h10 == s1_way_waddr_0_1_r) begin
        meta_array_16_0 <= s1_way_wdata_0_1_r;
      end else begin
        meta_array_16_0 <= _GEN_1786;
      end
    end else begin
      meta_array_16_0 <= _GEN_1786;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_16_1 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_1_1_REG) begin
      if (6'h10 == s1_way_waddr_1_1_r) begin
        meta_array_16_1 <= s1_way_wdata_1_1_r;
      end else begin
        meta_array_16_1 <= _GEN_1916;
      end
    end else begin
      meta_array_16_1 <= _GEN_1916;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_16_2 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_2_1_REG) begin
      if (6'h10 == s1_way_waddr_2_1_r) begin
        meta_array_16_2 <= s1_way_wdata_2_1_r;
      end else begin
        meta_array_16_2 <= _GEN_2046;
      end
    end else begin
      meta_array_16_2 <= _GEN_2046;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_16_3 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_3_1_REG) begin
      if (6'h10 == s1_way_waddr_3_1_r) begin
        meta_array_16_3 <= s1_way_wdata_3_1_r;
      end else begin
        meta_array_16_3 <= _GEN_2176;
      end
    end else begin
      meta_array_16_3 <= _GEN_2176;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_16_4 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_4_1_REG) begin
      if (6'h10 == s1_way_waddr_4_1_r) begin
        meta_array_16_4 <= s1_way_wdata_4_1_r;
      end else begin
        meta_array_16_4 <= _GEN_2306;
      end
    end else begin
      meta_array_16_4 <= _GEN_2306;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_16_5 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_5_1_REG) begin
      if (6'h10 == s1_way_waddr_5_1_r) begin
        meta_array_16_5 <= s1_way_wdata_5_1_r;
      end else begin
        meta_array_16_5 <= _GEN_2436;
      end
    end else begin
      meta_array_16_5 <= _GEN_2436;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_16_6 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_6_1_REG) begin
      if (6'h10 == s1_way_waddr_6_1_r) begin
        meta_array_16_6 <= s1_way_wdata_6_1_r;
      end else begin
        meta_array_16_6 <= _GEN_2566;
      end
    end else begin
      meta_array_16_6 <= _GEN_2566;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_16_7 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_7_1_REG) begin
      if (6'h10 == s1_way_waddr_7_1_r) begin
        meta_array_16_7 <= s1_way_wdata_7_1_r;
      end else begin
        meta_array_16_7 <= _GEN_2696;
      end
    end else begin
      meta_array_16_7 <= _GEN_2696;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_17_0 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_0_1_REG) begin
      if (6'h11 == s1_way_waddr_0_1_r) begin
        meta_array_17_0 <= s1_way_wdata_0_1_r;
      end else begin
        meta_array_17_0 <= _GEN_1787;
      end
    end else begin
      meta_array_17_0 <= _GEN_1787;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_17_1 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_1_1_REG) begin
      if (6'h11 == s1_way_waddr_1_1_r) begin
        meta_array_17_1 <= s1_way_wdata_1_1_r;
      end else begin
        meta_array_17_1 <= _GEN_1917;
      end
    end else begin
      meta_array_17_1 <= _GEN_1917;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_17_2 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_2_1_REG) begin
      if (6'h11 == s1_way_waddr_2_1_r) begin
        meta_array_17_2 <= s1_way_wdata_2_1_r;
      end else begin
        meta_array_17_2 <= _GEN_2047;
      end
    end else begin
      meta_array_17_2 <= _GEN_2047;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_17_3 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_3_1_REG) begin
      if (6'h11 == s1_way_waddr_3_1_r) begin
        meta_array_17_3 <= s1_way_wdata_3_1_r;
      end else begin
        meta_array_17_3 <= _GEN_2177;
      end
    end else begin
      meta_array_17_3 <= _GEN_2177;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_17_4 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_4_1_REG) begin
      if (6'h11 == s1_way_waddr_4_1_r) begin
        meta_array_17_4 <= s1_way_wdata_4_1_r;
      end else begin
        meta_array_17_4 <= _GEN_2307;
      end
    end else begin
      meta_array_17_4 <= _GEN_2307;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_17_5 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_5_1_REG) begin
      if (6'h11 == s1_way_waddr_5_1_r) begin
        meta_array_17_5 <= s1_way_wdata_5_1_r;
      end else begin
        meta_array_17_5 <= _GEN_2437;
      end
    end else begin
      meta_array_17_5 <= _GEN_2437;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_17_6 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_6_1_REG) begin
      if (6'h11 == s1_way_waddr_6_1_r) begin
        meta_array_17_6 <= s1_way_wdata_6_1_r;
      end else begin
        meta_array_17_6 <= _GEN_2567;
      end
    end else begin
      meta_array_17_6 <= _GEN_2567;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_17_7 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_7_1_REG) begin
      if (6'h11 == s1_way_waddr_7_1_r) begin
        meta_array_17_7 <= s1_way_wdata_7_1_r;
      end else begin
        meta_array_17_7 <= _GEN_2697;
      end
    end else begin
      meta_array_17_7 <= _GEN_2697;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_18_0 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_0_1_REG) begin
      if (6'h12 == s1_way_waddr_0_1_r) begin
        meta_array_18_0 <= s1_way_wdata_0_1_r;
      end else begin
        meta_array_18_0 <= _GEN_1788;
      end
    end else begin
      meta_array_18_0 <= _GEN_1788;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_18_1 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_1_1_REG) begin
      if (6'h12 == s1_way_waddr_1_1_r) begin
        meta_array_18_1 <= s1_way_wdata_1_1_r;
      end else begin
        meta_array_18_1 <= _GEN_1918;
      end
    end else begin
      meta_array_18_1 <= _GEN_1918;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_18_2 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_2_1_REG) begin
      if (6'h12 == s1_way_waddr_2_1_r) begin
        meta_array_18_2 <= s1_way_wdata_2_1_r;
      end else begin
        meta_array_18_2 <= _GEN_2048;
      end
    end else begin
      meta_array_18_2 <= _GEN_2048;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_18_3 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_3_1_REG) begin
      if (6'h12 == s1_way_waddr_3_1_r) begin
        meta_array_18_3 <= s1_way_wdata_3_1_r;
      end else begin
        meta_array_18_3 <= _GEN_2178;
      end
    end else begin
      meta_array_18_3 <= _GEN_2178;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_18_4 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_4_1_REG) begin
      if (6'h12 == s1_way_waddr_4_1_r) begin
        meta_array_18_4 <= s1_way_wdata_4_1_r;
      end else begin
        meta_array_18_4 <= _GEN_2308;
      end
    end else begin
      meta_array_18_4 <= _GEN_2308;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_18_5 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_5_1_REG) begin
      if (6'h12 == s1_way_waddr_5_1_r) begin
        meta_array_18_5 <= s1_way_wdata_5_1_r;
      end else begin
        meta_array_18_5 <= _GEN_2438;
      end
    end else begin
      meta_array_18_5 <= _GEN_2438;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_18_6 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_6_1_REG) begin
      if (6'h12 == s1_way_waddr_6_1_r) begin
        meta_array_18_6 <= s1_way_wdata_6_1_r;
      end else begin
        meta_array_18_6 <= _GEN_2568;
      end
    end else begin
      meta_array_18_6 <= _GEN_2568;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_18_7 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_7_1_REG) begin
      if (6'h12 == s1_way_waddr_7_1_r) begin
        meta_array_18_7 <= s1_way_wdata_7_1_r;
      end else begin
        meta_array_18_7 <= _GEN_2698;
      end
    end else begin
      meta_array_18_7 <= _GEN_2698;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_19_0 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_0_1_REG) begin
      if (6'h13 == s1_way_waddr_0_1_r) begin
        meta_array_19_0 <= s1_way_wdata_0_1_r;
      end else begin
        meta_array_19_0 <= _GEN_1789;
      end
    end else begin
      meta_array_19_0 <= _GEN_1789;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_19_1 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_1_1_REG) begin
      if (6'h13 == s1_way_waddr_1_1_r) begin
        meta_array_19_1 <= s1_way_wdata_1_1_r;
      end else begin
        meta_array_19_1 <= _GEN_1919;
      end
    end else begin
      meta_array_19_1 <= _GEN_1919;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_19_2 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_2_1_REG) begin
      if (6'h13 == s1_way_waddr_2_1_r) begin
        meta_array_19_2 <= s1_way_wdata_2_1_r;
      end else begin
        meta_array_19_2 <= _GEN_2049;
      end
    end else begin
      meta_array_19_2 <= _GEN_2049;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_19_3 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_3_1_REG) begin
      if (6'h13 == s1_way_waddr_3_1_r) begin
        meta_array_19_3 <= s1_way_wdata_3_1_r;
      end else begin
        meta_array_19_3 <= _GEN_2179;
      end
    end else begin
      meta_array_19_3 <= _GEN_2179;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_19_4 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_4_1_REG) begin
      if (6'h13 == s1_way_waddr_4_1_r) begin
        meta_array_19_4 <= s1_way_wdata_4_1_r;
      end else begin
        meta_array_19_4 <= _GEN_2309;
      end
    end else begin
      meta_array_19_4 <= _GEN_2309;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_19_5 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_5_1_REG) begin
      if (6'h13 == s1_way_waddr_5_1_r) begin
        meta_array_19_5 <= s1_way_wdata_5_1_r;
      end else begin
        meta_array_19_5 <= _GEN_2439;
      end
    end else begin
      meta_array_19_5 <= _GEN_2439;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_19_6 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_6_1_REG) begin
      if (6'h13 == s1_way_waddr_6_1_r) begin
        meta_array_19_6 <= s1_way_wdata_6_1_r;
      end else begin
        meta_array_19_6 <= _GEN_2569;
      end
    end else begin
      meta_array_19_6 <= _GEN_2569;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_19_7 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_7_1_REG) begin
      if (6'h13 == s1_way_waddr_7_1_r) begin
        meta_array_19_7 <= s1_way_wdata_7_1_r;
      end else begin
        meta_array_19_7 <= _GEN_2699;
      end
    end else begin
      meta_array_19_7 <= _GEN_2699;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_20_0 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_0_1_REG) begin
      if (6'h14 == s1_way_waddr_0_1_r) begin
        meta_array_20_0 <= s1_way_wdata_0_1_r;
      end else begin
        meta_array_20_0 <= _GEN_1790;
      end
    end else begin
      meta_array_20_0 <= _GEN_1790;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_20_1 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_1_1_REG) begin
      if (6'h14 == s1_way_waddr_1_1_r) begin
        meta_array_20_1 <= s1_way_wdata_1_1_r;
      end else begin
        meta_array_20_1 <= _GEN_1920;
      end
    end else begin
      meta_array_20_1 <= _GEN_1920;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_20_2 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_2_1_REG) begin
      if (6'h14 == s1_way_waddr_2_1_r) begin
        meta_array_20_2 <= s1_way_wdata_2_1_r;
      end else begin
        meta_array_20_2 <= _GEN_2050;
      end
    end else begin
      meta_array_20_2 <= _GEN_2050;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_20_3 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_3_1_REG) begin
      if (6'h14 == s1_way_waddr_3_1_r) begin
        meta_array_20_3 <= s1_way_wdata_3_1_r;
      end else begin
        meta_array_20_3 <= _GEN_2180;
      end
    end else begin
      meta_array_20_3 <= _GEN_2180;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_20_4 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_4_1_REG) begin
      if (6'h14 == s1_way_waddr_4_1_r) begin
        meta_array_20_4 <= s1_way_wdata_4_1_r;
      end else begin
        meta_array_20_4 <= _GEN_2310;
      end
    end else begin
      meta_array_20_4 <= _GEN_2310;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_20_5 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_5_1_REG) begin
      if (6'h14 == s1_way_waddr_5_1_r) begin
        meta_array_20_5 <= s1_way_wdata_5_1_r;
      end else begin
        meta_array_20_5 <= _GEN_2440;
      end
    end else begin
      meta_array_20_5 <= _GEN_2440;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_20_6 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_6_1_REG) begin
      if (6'h14 == s1_way_waddr_6_1_r) begin
        meta_array_20_6 <= s1_way_wdata_6_1_r;
      end else begin
        meta_array_20_6 <= _GEN_2570;
      end
    end else begin
      meta_array_20_6 <= _GEN_2570;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_20_7 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_7_1_REG) begin
      if (6'h14 == s1_way_waddr_7_1_r) begin
        meta_array_20_7 <= s1_way_wdata_7_1_r;
      end else begin
        meta_array_20_7 <= _GEN_2700;
      end
    end else begin
      meta_array_20_7 <= _GEN_2700;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_21_0 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_0_1_REG) begin
      if (6'h15 == s1_way_waddr_0_1_r) begin
        meta_array_21_0 <= s1_way_wdata_0_1_r;
      end else begin
        meta_array_21_0 <= _GEN_1791;
      end
    end else begin
      meta_array_21_0 <= _GEN_1791;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_21_1 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_1_1_REG) begin
      if (6'h15 == s1_way_waddr_1_1_r) begin
        meta_array_21_1 <= s1_way_wdata_1_1_r;
      end else begin
        meta_array_21_1 <= _GEN_1921;
      end
    end else begin
      meta_array_21_1 <= _GEN_1921;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_21_2 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_2_1_REG) begin
      if (6'h15 == s1_way_waddr_2_1_r) begin
        meta_array_21_2 <= s1_way_wdata_2_1_r;
      end else begin
        meta_array_21_2 <= _GEN_2051;
      end
    end else begin
      meta_array_21_2 <= _GEN_2051;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_21_3 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_3_1_REG) begin
      if (6'h15 == s1_way_waddr_3_1_r) begin
        meta_array_21_3 <= s1_way_wdata_3_1_r;
      end else begin
        meta_array_21_3 <= _GEN_2181;
      end
    end else begin
      meta_array_21_3 <= _GEN_2181;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_21_4 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_4_1_REG) begin
      if (6'h15 == s1_way_waddr_4_1_r) begin
        meta_array_21_4 <= s1_way_wdata_4_1_r;
      end else begin
        meta_array_21_4 <= _GEN_2311;
      end
    end else begin
      meta_array_21_4 <= _GEN_2311;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_21_5 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_5_1_REG) begin
      if (6'h15 == s1_way_waddr_5_1_r) begin
        meta_array_21_5 <= s1_way_wdata_5_1_r;
      end else begin
        meta_array_21_5 <= _GEN_2441;
      end
    end else begin
      meta_array_21_5 <= _GEN_2441;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_21_6 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_6_1_REG) begin
      if (6'h15 == s1_way_waddr_6_1_r) begin
        meta_array_21_6 <= s1_way_wdata_6_1_r;
      end else begin
        meta_array_21_6 <= _GEN_2571;
      end
    end else begin
      meta_array_21_6 <= _GEN_2571;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_21_7 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_7_1_REG) begin
      if (6'h15 == s1_way_waddr_7_1_r) begin
        meta_array_21_7 <= s1_way_wdata_7_1_r;
      end else begin
        meta_array_21_7 <= _GEN_2701;
      end
    end else begin
      meta_array_21_7 <= _GEN_2701;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_22_0 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_0_1_REG) begin
      if (6'h16 == s1_way_waddr_0_1_r) begin
        meta_array_22_0 <= s1_way_wdata_0_1_r;
      end else begin
        meta_array_22_0 <= _GEN_1792;
      end
    end else begin
      meta_array_22_0 <= _GEN_1792;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_22_1 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_1_1_REG) begin
      if (6'h16 == s1_way_waddr_1_1_r) begin
        meta_array_22_1 <= s1_way_wdata_1_1_r;
      end else begin
        meta_array_22_1 <= _GEN_1922;
      end
    end else begin
      meta_array_22_1 <= _GEN_1922;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_22_2 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_2_1_REG) begin
      if (6'h16 == s1_way_waddr_2_1_r) begin
        meta_array_22_2 <= s1_way_wdata_2_1_r;
      end else begin
        meta_array_22_2 <= _GEN_2052;
      end
    end else begin
      meta_array_22_2 <= _GEN_2052;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_22_3 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_3_1_REG) begin
      if (6'h16 == s1_way_waddr_3_1_r) begin
        meta_array_22_3 <= s1_way_wdata_3_1_r;
      end else begin
        meta_array_22_3 <= _GEN_2182;
      end
    end else begin
      meta_array_22_3 <= _GEN_2182;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_22_4 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_4_1_REG) begin
      if (6'h16 == s1_way_waddr_4_1_r) begin
        meta_array_22_4 <= s1_way_wdata_4_1_r;
      end else begin
        meta_array_22_4 <= _GEN_2312;
      end
    end else begin
      meta_array_22_4 <= _GEN_2312;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_22_5 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_5_1_REG) begin
      if (6'h16 == s1_way_waddr_5_1_r) begin
        meta_array_22_5 <= s1_way_wdata_5_1_r;
      end else begin
        meta_array_22_5 <= _GEN_2442;
      end
    end else begin
      meta_array_22_5 <= _GEN_2442;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_22_6 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_6_1_REG) begin
      if (6'h16 == s1_way_waddr_6_1_r) begin
        meta_array_22_6 <= s1_way_wdata_6_1_r;
      end else begin
        meta_array_22_6 <= _GEN_2572;
      end
    end else begin
      meta_array_22_6 <= _GEN_2572;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_22_7 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_7_1_REG) begin
      if (6'h16 == s1_way_waddr_7_1_r) begin
        meta_array_22_7 <= s1_way_wdata_7_1_r;
      end else begin
        meta_array_22_7 <= _GEN_2702;
      end
    end else begin
      meta_array_22_7 <= _GEN_2702;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_23_0 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_0_1_REG) begin
      if (6'h17 == s1_way_waddr_0_1_r) begin
        meta_array_23_0 <= s1_way_wdata_0_1_r;
      end else begin
        meta_array_23_0 <= _GEN_1793;
      end
    end else begin
      meta_array_23_0 <= _GEN_1793;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_23_1 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_1_1_REG) begin
      if (6'h17 == s1_way_waddr_1_1_r) begin
        meta_array_23_1 <= s1_way_wdata_1_1_r;
      end else begin
        meta_array_23_1 <= _GEN_1923;
      end
    end else begin
      meta_array_23_1 <= _GEN_1923;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_23_2 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_2_1_REG) begin
      if (6'h17 == s1_way_waddr_2_1_r) begin
        meta_array_23_2 <= s1_way_wdata_2_1_r;
      end else begin
        meta_array_23_2 <= _GEN_2053;
      end
    end else begin
      meta_array_23_2 <= _GEN_2053;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_23_3 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_3_1_REG) begin
      if (6'h17 == s1_way_waddr_3_1_r) begin
        meta_array_23_3 <= s1_way_wdata_3_1_r;
      end else begin
        meta_array_23_3 <= _GEN_2183;
      end
    end else begin
      meta_array_23_3 <= _GEN_2183;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_23_4 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_4_1_REG) begin
      if (6'h17 == s1_way_waddr_4_1_r) begin
        meta_array_23_4 <= s1_way_wdata_4_1_r;
      end else begin
        meta_array_23_4 <= _GEN_2313;
      end
    end else begin
      meta_array_23_4 <= _GEN_2313;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_23_5 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_5_1_REG) begin
      if (6'h17 == s1_way_waddr_5_1_r) begin
        meta_array_23_5 <= s1_way_wdata_5_1_r;
      end else begin
        meta_array_23_5 <= _GEN_2443;
      end
    end else begin
      meta_array_23_5 <= _GEN_2443;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_23_6 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_6_1_REG) begin
      if (6'h17 == s1_way_waddr_6_1_r) begin
        meta_array_23_6 <= s1_way_wdata_6_1_r;
      end else begin
        meta_array_23_6 <= _GEN_2573;
      end
    end else begin
      meta_array_23_6 <= _GEN_2573;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_23_7 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_7_1_REG) begin
      if (6'h17 == s1_way_waddr_7_1_r) begin
        meta_array_23_7 <= s1_way_wdata_7_1_r;
      end else begin
        meta_array_23_7 <= _GEN_2703;
      end
    end else begin
      meta_array_23_7 <= _GEN_2703;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_24_0 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_0_1_REG) begin
      if (6'h18 == s1_way_waddr_0_1_r) begin
        meta_array_24_0 <= s1_way_wdata_0_1_r;
      end else begin
        meta_array_24_0 <= _GEN_1794;
      end
    end else begin
      meta_array_24_0 <= _GEN_1794;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_24_1 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_1_1_REG) begin
      if (6'h18 == s1_way_waddr_1_1_r) begin
        meta_array_24_1 <= s1_way_wdata_1_1_r;
      end else begin
        meta_array_24_1 <= _GEN_1924;
      end
    end else begin
      meta_array_24_1 <= _GEN_1924;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_24_2 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_2_1_REG) begin
      if (6'h18 == s1_way_waddr_2_1_r) begin
        meta_array_24_2 <= s1_way_wdata_2_1_r;
      end else begin
        meta_array_24_2 <= _GEN_2054;
      end
    end else begin
      meta_array_24_2 <= _GEN_2054;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_24_3 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_3_1_REG) begin
      if (6'h18 == s1_way_waddr_3_1_r) begin
        meta_array_24_3 <= s1_way_wdata_3_1_r;
      end else begin
        meta_array_24_3 <= _GEN_2184;
      end
    end else begin
      meta_array_24_3 <= _GEN_2184;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_24_4 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_4_1_REG) begin
      if (6'h18 == s1_way_waddr_4_1_r) begin
        meta_array_24_4 <= s1_way_wdata_4_1_r;
      end else begin
        meta_array_24_4 <= _GEN_2314;
      end
    end else begin
      meta_array_24_4 <= _GEN_2314;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_24_5 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_5_1_REG) begin
      if (6'h18 == s1_way_waddr_5_1_r) begin
        meta_array_24_5 <= s1_way_wdata_5_1_r;
      end else begin
        meta_array_24_5 <= _GEN_2444;
      end
    end else begin
      meta_array_24_5 <= _GEN_2444;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_24_6 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_6_1_REG) begin
      if (6'h18 == s1_way_waddr_6_1_r) begin
        meta_array_24_6 <= s1_way_wdata_6_1_r;
      end else begin
        meta_array_24_6 <= _GEN_2574;
      end
    end else begin
      meta_array_24_6 <= _GEN_2574;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_24_7 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_7_1_REG) begin
      if (6'h18 == s1_way_waddr_7_1_r) begin
        meta_array_24_7 <= s1_way_wdata_7_1_r;
      end else begin
        meta_array_24_7 <= _GEN_2704;
      end
    end else begin
      meta_array_24_7 <= _GEN_2704;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_25_0 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_0_1_REG) begin
      if (6'h19 == s1_way_waddr_0_1_r) begin
        meta_array_25_0 <= s1_way_wdata_0_1_r;
      end else begin
        meta_array_25_0 <= _GEN_1795;
      end
    end else begin
      meta_array_25_0 <= _GEN_1795;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_25_1 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_1_1_REG) begin
      if (6'h19 == s1_way_waddr_1_1_r) begin
        meta_array_25_1 <= s1_way_wdata_1_1_r;
      end else begin
        meta_array_25_1 <= _GEN_1925;
      end
    end else begin
      meta_array_25_1 <= _GEN_1925;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_25_2 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_2_1_REG) begin
      if (6'h19 == s1_way_waddr_2_1_r) begin
        meta_array_25_2 <= s1_way_wdata_2_1_r;
      end else begin
        meta_array_25_2 <= _GEN_2055;
      end
    end else begin
      meta_array_25_2 <= _GEN_2055;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_25_3 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_3_1_REG) begin
      if (6'h19 == s1_way_waddr_3_1_r) begin
        meta_array_25_3 <= s1_way_wdata_3_1_r;
      end else begin
        meta_array_25_3 <= _GEN_2185;
      end
    end else begin
      meta_array_25_3 <= _GEN_2185;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_25_4 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_4_1_REG) begin
      if (6'h19 == s1_way_waddr_4_1_r) begin
        meta_array_25_4 <= s1_way_wdata_4_1_r;
      end else begin
        meta_array_25_4 <= _GEN_2315;
      end
    end else begin
      meta_array_25_4 <= _GEN_2315;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_25_5 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_5_1_REG) begin
      if (6'h19 == s1_way_waddr_5_1_r) begin
        meta_array_25_5 <= s1_way_wdata_5_1_r;
      end else begin
        meta_array_25_5 <= _GEN_2445;
      end
    end else begin
      meta_array_25_5 <= _GEN_2445;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_25_6 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_6_1_REG) begin
      if (6'h19 == s1_way_waddr_6_1_r) begin
        meta_array_25_6 <= s1_way_wdata_6_1_r;
      end else begin
        meta_array_25_6 <= _GEN_2575;
      end
    end else begin
      meta_array_25_6 <= _GEN_2575;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_25_7 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_7_1_REG) begin
      if (6'h19 == s1_way_waddr_7_1_r) begin
        meta_array_25_7 <= s1_way_wdata_7_1_r;
      end else begin
        meta_array_25_7 <= _GEN_2705;
      end
    end else begin
      meta_array_25_7 <= _GEN_2705;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_26_0 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_0_1_REG) begin
      if (6'h1a == s1_way_waddr_0_1_r) begin
        meta_array_26_0 <= s1_way_wdata_0_1_r;
      end else begin
        meta_array_26_0 <= _GEN_1796;
      end
    end else begin
      meta_array_26_0 <= _GEN_1796;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_26_1 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_1_1_REG) begin
      if (6'h1a == s1_way_waddr_1_1_r) begin
        meta_array_26_1 <= s1_way_wdata_1_1_r;
      end else begin
        meta_array_26_1 <= _GEN_1926;
      end
    end else begin
      meta_array_26_1 <= _GEN_1926;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_26_2 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_2_1_REG) begin
      if (6'h1a == s1_way_waddr_2_1_r) begin
        meta_array_26_2 <= s1_way_wdata_2_1_r;
      end else begin
        meta_array_26_2 <= _GEN_2056;
      end
    end else begin
      meta_array_26_2 <= _GEN_2056;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_26_3 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_3_1_REG) begin
      if (6'h1a == s1_way_waddr_3_1_r) begin
        meta_array_26_3 <= s1_way_wdata_3_1_r;
      end else begin
        meta_array_26_3 <= _GEN_2186;
      end
    end else begin
      meta_array_26_3 <= _GEN_2186;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_26_4 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_4_1_REG) begin
      if (6'h1a == s1_way_waddr_4_1_r) begin
        meta_array_26_4 <= s1_way_wdata_4_1_r;
      end else begin
        meta_array_26_4 <= _GEN_2316;
      end
    end else begin
      meta_array_26_4 <= _GEN_2316;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_26_5 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_5_1_REG) begin
      if (6'h1a == s1_way_waddr_5_1_r) begin
        meta_array_26_5 <= s1_way_wdata_5_1_r;
      end else begin
        meta_array_26_5 <= _GEN_2446;
      end
    end else begin
      meta_array_26_5 <= _GEN_2446;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_26_6 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_6_1_REG) begin
      if (6'h1a == s1_way_waddr_6_1_r) begin
        meta_array_26_6 <= s1_way_wdata_6_1_r;
      end else begin
        meta_array_26_6 <= _GEN_2576;
      end
    end else begin
      meta_array_26_6 <= _GEN_2576;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_26_7 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_7_1_REG) begin
      if (6'h1a == s1_way_waddr_7_1_r) begin
        meta_array_26_7 <= s1_way_wdata_7_1_r;
      end else begin
        meta_array_26_7 <= _GEN_2706;
      end
    end else begin
      meta_array_26_7 <= _GEN_2706;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_27_0 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_0_1_REG) begin
      if (6'h1b == s1_way_waddr_0_1_r) begin
        meta_array_27_0 <= s1_way_wdata_0_1_r;
      end else begin
        meta_array_27_0 <= _GEN_1797;
      end
    end else begin
      meta_array_27_0 <= _GEN_1797;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_27_1 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_1_1_REG) begin
      if (6'h1b == s1_way_waddr_1_1_r) begin
        meta_array_27_1 <= s1_way_wdata_1_1_r;
      end else begin
        meta_array_27_1 <= _GEN_1927;
      end
    end else begin
      meta_array_27_1 <= _GEN_1927;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_27_2 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_2_1_REG) begin
      if (6'h1b == s1_way_waddr_2_1_r) begin
        meta_array_27_2 <= s1_way_wdata_2_1_r;
      end else begin
        meta_array_27_2 <= _GEN_2057;
      end
    end else begin
      meta_array_27_2 <= _GEN_2057;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_27_3 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_3_1_REG) begin
      if (6'h1b == s1_way_waddr_3_1_r) begin
        meta_array_27_3 <= s1_way_wdata_3_1_r;
      end else begin
        meta_array_27_3 <= _GEN_2187;
      end
    end else begin
      meta_array_27_3 <= _GEN_2187;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_27_4 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_4_1_REG) begin
      if (6'h1b == s1_way_waddr_4_1_r) begin
        meta_array_27_4 <= s1_way_wdata_4_1_r;
      end else begin
        meta_array_27_4 <= _GEN_2317;
      end
    end else begin
      meta_array_27_4 <= _GEN_2317;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_27_5 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_5_1_REG) begin
      if (6'h1b == s1_way_waddr_5_1_r) begin
        meta_array_27_5 <= s1_way_wdata_5_1_r;
      end else begin
        meta_array_27_5 <= _GEN_2447;
      end
    end else begin
      meta_array_27_5 <= _GEN_2447;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_27_6 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_6_1_REG) begin
      if (6'h1b == s1_way_waddr_6_1_r) begin
        meta_array_27_6 <= s1_way_wdata_6_1_r;
      end else begin
        meta_array_27_6 <= _GEN_2577;
      end
    end else begin
      meta_array_27_6 <= _GEN_2577;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_27_7 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_7_1_REG) begin
      if (6'h1b == s1_way_waddr_7_1_r) begin
        meta_array_27_7 <= s1_way_wdata_7_1_r;
      end else begin
        meta_array_27_7 <= _GEN_2707;
      end
    end else begin
      meta_array_27_7 <= _GEN_2707;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_28_0 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_0_1_REG) begin
      if (6'h1c == s1_way_waddr_0_1_r) begin
        meta_array_28_0 <= s1_way_wdata_0_1_r;
      end else begin
        meta_array_28_0 <= _GEN_1798;
      end
    end else begin
      meta_array_28_0 <= _GEN_1798;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_28_1 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_1_1_REG) begin
      if (6'h1c == s1_way_waddr_1_1_r) begin
        meta_array_28_1 <= s1_way_wdata_1_1_r;
      end else begin
        meta_array_28_1 <= _GEN_1928;
      end
    end else begin
      meta_array_28_1 <= _GEN_1928;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_28_2 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_2_1_REG) begin
      if (6'h1c == s1_way_waddr_2_1_r) begin
        meta_array_28_2 <= s1_way_wdata_2_1_r;
      end else begin
        meta_array_28_2 <= _GEN_2058;
      end
    end else begin
      meta_array_28_2 <= _GEN_2058;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_28_3 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_3_1_REG) begin
      if (6'h1c == s1_way_waddr_3_1_r) begin
        meta_array_28_3 <= s1_way_wdata_3_1_r;
      end else begin
        meta_array_28_3 <= _GEN_2188;
      end
    end else begin
      meta_array_28_3 <= _GEN_2188;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_28_4 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_4_1_REG) begin
      if (6'h1c == s1_way_waddr_4_1_r) begin
        meta_array_28_4 <= s1_way_wdata_4_1_r;
      end else begin
        meta_array_28_4 <= _GEN_2318;
      end
    end else begin
      meta_array_28_4 <= _GEN_2318;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_28_5 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_5_1_REG) begin
      if (6'h1c == s1_way_waddr_5_1_r) begin
        meta_array_28_5 <= s1_way_wdata_5_1_r;
      end else begin
        meta_array_28_5 <= _GEN_2448;
      end
    end else begin
      meta_array_28_5 <= _GEN_2448;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_28_6 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_6_1_REG) begin
      if (6'h1c == s1_way_waddr_6_1_r) begin
        meta_array_28_6 <= s1_way_wdata_6_1_r;
      end else begin
        meta_array_28_6 <= _GEN_2578;
      end
    end else begin
      meta_array_28_6 <= _GEN_2578;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_28_7 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_7_1_REG) begin
      if (6'h1c == s1_way_waddr_7_1_r) begin
        meta_array_28_7 <= s1_way_wdata_7_1_r;
      end else begin
        meta_array_28_7 <= _GEN_2708;
      end
    end else begin
      meta_array_28_7 <= _GEN_2708;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_29_0 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_0_1_REG) begin
      if (6'h1d == s1_way_waddr_0_1_r) begin
        meta_array_29_0 <= s1_way_wdata_0_1_r;
      end else begin
        meta_array_29_0 <= _GEN_1799;
      end
    end else begin
      meta_array_29_0 <= _GEN_1799;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_29_1 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_1_1_REG) begin
      if (6'h1d == s1_way_waddr_1_1_r) begin
        meta_array_29_1 <= s1_way_wdata_1_1_r;
      end else begin
        meta_array_29_1 <= _GEN_1929;
      end
    end else begin
      meta_array_29_1 <= _GEN_1929;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_29_2 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_2_1_REG) begin
      if (6'h1d == s1_way_waddr_2_1_r) begin
        meta_array_29_2 <= s1_way_wdata_2_1_r;
      end else begin
        meta_array_29_2 <= _GEN_2059;
      end
    end else begin
      meta_array_29_2 <= _GEN_2059;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_29_3 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_3_1_REG) begin
      if (6'h1d == s1_way_waddr_3_1_r) begin
        meta_array_29_3 <= s1_way_wdata_3_1_r;
      end else begin
        meta_array_29_3 <= _GEN_2189;
      end
    end else begin
      meta_array_29_3 <= _GEN_2189;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_29_4 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_4_1_REG) begin
      if (6'h1d == s1_way_waddr_4_1_r) begin
        meta_array_29_4 <= s1_way_wdata_4_1_r;
      end else begin
        meta_array_29_4 <= _GEN_2319;
      end
    end else begin
      meta_array_29_4 <= _GEN_2319;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_29_5 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_5_1_REG) begin
      if (6'h1d == s1_way_waddr_5_1_r) begin
        meta_array_29_5 <= s1_way_wdata_5_1_r;
      end else begin
        meta_array_29_5 <= _GEN_2449;
      end
    end else begin
      meta_array_29_5 <= _GEN_2449;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_29_6 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_6_1_REG) begin
      if (6'h1d == s1_way_waddr_6_1_r) begin
        meta_array_29_6 <= s1_way_wdata_6_1_r;
      end else begin
        meta_array_29_6 <= _GEN_2579;
      end
    end else begin
      meta_array_29_6 <= _GEN_2579;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_29_7 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_7_1_REG) begin
      if (6'h1d == s1_way_waddr_7_1_r) begin
        meta_array_29_7 <= s1_way_wdata_7_1_r;
      end else begin
        meta_array_29_7 <= _GEN_2709;
      end
    end else begin
      meta_array_29_7 <= _GEN_2709;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_30_0 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_0_1_REG) begin
      if (6'h1e == s1_way_waddr_0_1_r) begin
        meta_array_30_0 <= s1_way_wdata_0_1_r;
      end else begin
        meta_array_30_0 <= _GEN_1800;
      end
    end else begin
      meta_array_30_0 <= _GEN_1800;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_30_1 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_1_1_REG) begin
      if (6'h1e == s1_way_waddr_1_1_r) begin
        meta_array_30_1 <= s1_way_wdata_1_1_r;
      end else begin
        meta_array_30_1 <= _GEN_1930;
      end
    end else begin
      meta_array_30_1 <= _GEN_1930;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_30_2 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_2_1_REG) begin
      if (6'h1e == s1_way_waddr_2_1_r) begin
        meta_array_30_2 <= s1_way_wdata_2_1_r;
      end else begin
        meta_array_30_2 <= _GEN_2060;
      end
    end else begin
      meta_array_30_2 <= _GEN_2060;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_30_3 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_3_1_REG) begin
      if (6'h1e == s1_way_waddr_3_1_r) begin
        meta_array_30_3 <= s1_way_wdata_3_1_r;
      end else begin
        meta_array_30_3 <= _GEN_2190;
      end
    end else begin
      meta_array_30_3 <= _GEN_2190;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_30_4 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_4_1_REG) begin
      if (6'h1e == s1_way_waddr_4_1_r) begin
        meta_array_30_4 <= s1_way_wdata_4_1_r;
      end else begin
        meta_array_30_4 <= _GEN_2320;
      end
    end else begin
      meta_array_30_4 <= _GEN_2320;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_30_5 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_5_1_REG) begin
      if (6'h1e == s1_way_waddr_5_1_r) begin
        meta_array_30_5 <= s1_way_wdata_5_1_r;
      end else begin
        meta_array_30_5 <= _GEN_2450;
      end
    end else begin
      meta_array_30_5 <= _GEN_2450;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_30_6 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_6_1_REG) begin
      if (6'h1e == s1_way_waddr_6_1_r) begin
        meta_array_30_6 <= s1_way_wdata_6_1_r;
      end else begin
        meta_array_30_6 <= _GEN_2580;
      end
    end else begin
      meta_array_30_6 <= _GEN_2580;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_30_7 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_7_1_REG) begin
      if (6'h1e == s1_way_waddr_7_1_r) begin
        meta_array_30_7 <= s1_way_wdata_7_1_r;
      end else begin
        meta_array_30_7 <= _GEN_2710;
      end
    end else begin
      meta_array_30_7 <= _GEN_2710;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_31_0 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_0_1_REG) begin
      if (6'h1f == s1_way_waddr_0_1_r) begin
        meta_array_31_0 <= s1_way_wdata_0_1_r;
      end else begin
        meta_array_31_0 <= _GEN_1801;
      end
    end else begin
      meta_array_31_0 <= _GEN_1801;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_31_1 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_1_1_REG) begin
      if (6'h1f == s1_way_waddr_1_1_r) begin
        meta_array_31_1 <= s1_way_wdata_1_1_r;
      end else begin
        meta_array_31_1 <= _GEN_1931;
      end
    end else begin
      meta_array_31_1 <= _GEN_1931;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_31_2 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_2_1_REG) begin
      if (6'h1f == s1_way_waddr_2_1_r) begin
        meta_array_31_2 <= s1_way_wdata_2_1_r;
      end else begin
        meta_array_31_2 <= _GEN_2061;
      end
    end else begin
      meta_array_31_2 <= _GEN_2061;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_31_3 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_3_1_REG) begin
      if (6'h1f == s1_way_waddr_3_1_r) begin
        meta_array_31_3 <= s1_way_wdata_3_1_r;
      end else begin
        meta_array_31_3 <= _GEN_2191;
      end
    end else begin
      meta_array_31_3 <= _GEN_2191;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_31_4 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_4_1_REG) begin
      if (6'h1f == s1_way_waddr_4_1_r) begin
        meta_array_31_4 <= s1_way_wdata_4_1_r;
      end else begin
        meta_array_31_4 <= _GEN_2321;
      end
    end else begin
      meta_array_31_4 <= _GEN_2321;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_31_5 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_5_1_REG) begin
      if (6'h1f == s1_way_waddr_5_1_r) begin
        meta_array_31_5 <= s1_way_wdata_5_1_r;
      end else begin
        meta_array_31_5 <= _GEN_2451;
      end
    end else begin
      meta_array_31_5 <= _GEN_2451;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_31_6 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_6_1_REG) begin
      if (6'h1f == s1_way_waddr_6_1_r) begin
        meta_array_31_6 <= s1_way_wdata_6_1_r;
      end else begin
        meta_array_31_6 <= _GEN_2581;
      end
    end else begin
      meta_array_31_6 <= _GEN_2581;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_31_7 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_7_1_REG) begin
      if (6'h1f == s1_way_waddr_7_1_r) begin
        meta_array_31_7 <= s1_way_wdata_7_1_r;
      end else begin
        meta_array_31_7 <= _GEN_2711;
      end
    end else begin
      meta_array_31_7 <= _GEN_2711;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_32_0 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_0_1_REG) begin
      if (6'h20 == s1_way_waddr_0_1_r) begin
        meta_array_32_0 <= s1_way_wdata_0_1_r;
      end else begin
        meta_array_32_0 <= _GEN_1802;
      end
    end else begin
      meta_array_32_0 <= _GEN_1802;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_32_1 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_1_1_REG) begin
      if (6'h20 == s1_way_waddr_1_1_r) begin
        meta_array_32_1 <= s1_way_wdata_1_1_r;
      end else begin
        meta_array_32_1 <= _GEN_1932;
      end
    end else begin
      meta_array_32_1 <= _GEN_1932;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_32_2 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_2_1_REG) begin
      if (6'h20 == s1_way_waddr_2_1_r) begin
        meta_array_32_2 <= s1_way_wdata_2_1_r;
      end else begin
        meta_array_32_2 <= _GEN_2062;
      end
    end else begin
      meta_array_32_2 <= _GEN_2062;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_32_3 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_3_1_REG) begin
      if (6'h20 == s1_way_waddr_3_1_r) begin
        meta_array_32_3 <= s1_way_wdata_3_1_r;
      end else begin
        meta_array_32_3 <= _GEN_2192;
      end
    end else begin
      meta_array_32_3 <= _GEN_2192;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_32_4 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_4_1_REG) begin
      if (6'h20 == s1_way_waddr_4_1_r) begin
        meta_array_32_4 <= s1_way_wdata_4_1_r;
      end else begin
        meta_array_32_4 <= _GEN_2322;
      end
    end else begin
      meta_array_32_4 <= _GEN_2322;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_32_5 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_5_1_REG) begin
      if (6'h20 == s1_way_waddr_5_1_r) begin
        meta_array_32_5 <= s1_way_wdata_5_1_r;
      end else begin
        meta_array_32_5 <= _GEN_2452;
      end
    end else begin
      meta_array_32_5 <= _GEN_2452;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_32_6 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_6_1_REG) begin
      if (6'h20 == s1_way_waddr_6_1_r) begin
        meta_array_32_6 <= s1_way_wdata_6_1_r;
      end else begin
        meta_array_32_6 <= _GEN_2582;
      end
    end else begin
      meta_array_32_6 <= _GEN_2582;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_32_7 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_7_1_REG) begin
      if (6'h20 == s1_way_waddr_7_1_r) begin
        meta_array_32_7 <= s1_way_wdata_7_1_r;
      end else begin
        meta_array_32_7 <= _GEN_2712;
      end
    end else begin
      meta_array_32_7 <= _GEN_2712;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_33_0 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_0_1_REG) begin
      if (6'h21 == s1_way_waddr_0_1_r) begin
        meta_array_33_0 <= s1_way_wdata_0_1_r;
      end else begin
        meta_array_33_0 <= _GEN_1803;
      end
    end else begin
      meta_array_33_0 <= _GEN_1803;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_33_1 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_1_1_REG) begin
      if (6'h21 == s1_way_waddr_1_1_r) begin
        meta_array_33_1 <= s1_way_wdata_1_1_r;
      end else begin
        meta_array_33_1 <= _GEN_1933;
      end
    end else begin
      meta_array_33_1 <= _GEN_1933;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_33_2 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_2_1_REG) begin
      if (6'h21 == s1_way_waddr_2_1_r) begin
        meta_array_33_2 <= s1_way_wdata_2_1_r;
      end else begin
        meta_array_33_2 <= _GEN_2063;
      end
    end else begin
      meta_array_33_2 <= _GEN_2063;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_33_3 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_3_1_REG) begin
      if (6'h21 == s1_way_waddr_3_1_r) begin
        meta_array_33_3 <= s1_way_wdata_3_1_r;
      end else begin
        meta_array_33_3 <= _GEN_2193;
      end
    end else begin
      meta_array_33_3 <= _GEN_2193;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_33_4 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_4_1_REG) begin
      if (6'h21 == s1_way_waddr_4_1_r) begin
        meta_array_33_4 <= s1_way_wdata_4_1_r;
      end else begin
        meta_array_33_4 <= _GEN_2323;
      end
    end else begin
      meta_array_33_4 <= _GEN_2323;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_33_5 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_5_1_REG) begin
      if (6'h21 == s1_way_waddr_5_1_r) begin
        meta_array_33_5 <= s1_way_wdata_5_1_r;
      end else begin
        meta_array_33_5 <= _GEN_2453;
      end
    end else begin
      meta_array_33_5 <= _GEN_2453;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_33_6 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_6_1_REG) begin
      if (6'h21 == s1_way_waddr_6_1_r) begin
        meta_array_33_6 <= s1_way_wdata_6_1_r;
      end else begin
        meta_array_33_6 <= _GEN_2583;
      end
    end else begin
      meta_array_33_6 <= _GEN_2583;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_33_7 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_7_1_REG) begin
      if (6'h21 == s1_way_waddr_7_1_r) begin
        meta_array_33_7 <= s1_way_wdata_7_1_r;
      end else begin
        meta_array_33_7 <= _GEN_2713;
      end
    end else begin
      meta_array_33_7 <= _GEN_2713;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_34_0 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_0_1_REG) begin
      if (6'h22 == s1_way_waddr_0_1_r) begin
        meta_array_34_0 <= s1_way_wdata_0_1_r;
      end else begin
        meta_array_34_0 <= _GEN_1804;
      end
    end else begin
      meta_array_34_0 <= _GEN_1804;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_34_1 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_1_1_REG) begin
      if (6'h22 == s1_way_waddr_1_1_r) begin
        meta_array_34_1 <= s1_way_wdata_1_1_r;
      end else begin
        meta_array_34_1 <= _GEN_1934;
      end
    end else begin
      meta_array_34_1 <= _GEN_1934;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_34_2 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_2_1_REG) begin
      if (6'h22 == s1_way_waddr_2_1_r) begin
        meta_array_34_2 <= s1_way_wdata_2_1_r;
      end else begin
        meta_array_34_2 <= _GEN_2064;
      end
    end else begin
      meta_array_34_2 <= _GEN_2064;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_34_3 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_3_1_REG) begin
      if (6'h22 == s1_way_waddr_3_1_r) begin
        meta_array_34_3 <= s1_way_wdata_3_1_r;
      end else begin
        meta_array_34_3 <= _GEN_2194;
      end
    end else begin
      meta_array_34_3 <= _GEN_2194;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_34_4 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_4_1_REG) begin
      if (6'h22 == s1_way_waddr_4_1_r) begin
        meta_array_34_4 <= s1_way_wdata_4_1_r;
      end else begin
        meta_array_34_4 <= _GEN_2324;
      end
    end else begin
      meta_array_34_4 <= _GEN_2324;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_34_5 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_5_1_REG) begin
      if (6'h22 == s1_way_waddr_5_1_r) begin
        meta_array_34_5 <= s1_way_wdata_5_1_r;
      end else begin
        meta_array_34_5 <= _GEN_2454;
      end
    end else begin
      meta_array_34_5 <= _GEN_2454;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_34_6 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_6_1_REG) begin
      if (6'h22 == s1_way_waddr_6_1_r) begin
        meta_array_34_6 <= s1_way_wdata_6_1_r;
      end else begin
        meta_array_34_6 <= _GEN_2584;
      end
    end else begin
      meta_array_34_6 <= _GEN_2584;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_34_7 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_7_1_REG) begin
      if (6'h22 == s1_way_waddr_7_1_r) begin
        meta_array_34_7 <= s1_way_wdata_7_1_r;
      end else begin
        meta_array_34_7 <= _GEN_2714;
      end
    end else begin
      meta_array_34_7 <= _GEN_2714;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_35_0 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_0_1_REG) begin
      if (6'h23 == s1_way_waddr_0_1_r) begin
        meta_array_35_0 <= s1_way_wdata_0_1_r;
      end else begin
        meta_array_35_0 <= _GEN_1805;
      end
    end else begin
      meta_array_35_0 <= _GEN_1805;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_35_1 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_1_1_REG) begin
      if (6'h23 == s1_way_waddr_1_1_r) begin
        meta_array_35_1 <= s1_way_wdata_1_1_r;
      end else begin
        meta_array_35_1 <= _GEN_1935;
      end
    end else begin
      meta_array_35_1 <= _GEN_1935;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_35_2 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_2_1_REG) begin
      if (6'h23 == s1_way_waddr_2_1_r) begin
        meta_array_35_2 <= s1_way_wdata_2_1_r;
      end else begin
        meta_array_35_2 <= _GEN_2065;
      end
    end else begin
      meta_array_35_2 <= _GEN_2065;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_35_3 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_3_1_REG) begin
      if (6'h23 == s1_way_waddr_3_1_r) begin
        meta_array_35_3 <= s1_way_wdata_3_1_r;
      end else begin
        meta_array_35_3 <= _GEN_2195;
      end
    end else begin
      meta_array_35_3 <= _GEN_2195;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_35_4 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_4_1_REG) begin
      if (6'h23 == s1_way_waddr_4_1_r) begin
        meta_array_35_4 <= s1_way_wdata_4_1_r;
      end else begin
        meta_array_35_4 <= _GEN_2325;
      end
    end else begin
      meta_array_35_4 <= _GEN_2325;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_35_5 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_5_1_REG) begin
      if (6'h23 == s1_way_waddr_5_1_r) begin
        meta_array_35_5 <= s1_way_wdata_5_1_r;
      end else begin
        meta_array_35_5 <= _GEN_2455;
      end
    end else begin
      meta_array_35_5 <= _GEN_2455;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_35_6 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_6_1_REG) begin
      if (6'h23 == s1_way_waddr_6_1_r) begin
        meta_array_35_6 <= s1_way_wdata_6_1_r;
      end else begin
        meta_array_35_6 <= _GEN_2585;
      end
    end else begin
      meta_array_35_6 <= _GEN_2585;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_35_7 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_7_1_REG) begin
      if (6'h23 == s1_way_waddr_7_1_r) begin
        meta_array_35_7 <= s1_way_wdata_7_1_r;
      end else begin
        meta_array_35_7 <= _GEN_2715;
      end
    end else begin
      meta_array_35_7 <= _GEN_2715;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_36_0 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_0_1_REG) begin
      if (6'h24 == s1_way_waddr_0_1_r) begin
        meta_array_36_0 <= s1_way_wdata_0_1_r;
      end else begin
        meta_array_36_0 <= _GEN_1806;
      end
    end else begin
      meta_array_36_0 <= _GEN_1806;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_36_1 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_1_1_REG) begin
      if (6'h24 == s1_way_waddr_1_1_r) begin
        meta_array_36_1 <= s1_way_wdata_1_1_r;
      end else begin
        meta_array_36_1 <= _GEN_1936;
      end
    end else begin
      meta_array_36_1 <= _GEN_1936;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_36_2 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_2_1_REG) begin
      if (6'h24 == s1_way_waddr_2_1_r) begin
        meta_array_36_2 <= s1_way_wdata_2_1_r;
      end else begin
        meta_array_36_2 <= _GEN_2066;
      end
    end else begin
      meta_array_36_2 <= _GEN_2066;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_36_3 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_3_1_REG) begin
      if (6'h24 == s1_way_waddr_3_1_r) begin
        meta_array_36_3 <= s1_way_wdata_3_1_r;
      end else begin
        meta_array_36_3 <= _GEN_2196;
      end
    end else begin
      meta_array_36_3 <= _GEN_2196;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_36_4 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_4_1_REG) begin
      if (6'h24 == s1_way_waddr_4_1_r) begin
        meta_array_36_4 <= s1_way_wdata_4_1_r;
      end else begin
        meta_array_36_4 <= _GEN_2326;
      end
    end else begin
      meta_array_36_4 <= _GEN_2326;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_36_5 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_5_1_REG) begin
      if (6'h24 == s1_way_waddr_5_1_r) begin
        meta_array_36_5 <= s1_way_wdata_5_1_r;
      end else begin
        meta_array_36_5 <= _GEN_2456;
      end
    end else begin
      meta_array_36_5 <= _GEN_2456;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_36_6 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_6_1_REG) begin
      if (6'h24 == s1_way_waddr_6_1_r) begin
        meta_array_36_6 <= s1_way_wdata_6_1_r;
      end else begin
        meta_array_36_6 <= _GEN_2586;
      end
    end else begin
      meta_array_36_6 <= _GEN_2586;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_36_7 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_7_1_REG) begin
      if (6'h24 == s1_way_waddr_7_1_r) begin
        meta_array_36_7 <= s1_way_wdata_7_1_r;
      end else begin
        meta_array_36_7 <= _GEN_2716;
      end
    end else begin
      meta_array_36_7 <= _GEN_2716;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_37_0 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_0_1_REG) begin
      if (6'h25 == s1_way_waddr_0_1_r) begin
        meta_array_37_0 <= s1_way_wdata_0_1_r;
      end else begin
        meta_array_37_0 <= _GEN_1807;
      end
    end else begin
      meta_array_37_0 <= _GEN_1807;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_37_1 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_1_1_REG) begin
      if (6'h25 == s1_way_waddr_1_1_r) begin
        meta_array_37_1 <= s1_way_wdata_1_1_r;
      end else begin
        meta_array_37_1 <= _GEN_1937;
      end
    end else begin
      meta_array_37_1 <= _GEN_1937;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_37_2 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_2_1_REG) begin
      if (6'h25 == s1_way_waddr_2_1_r) begin
        meta_array_37_2 <= s1_way_wdata_2_1_r;
      end else begin
        meta_array_37_2 <= _GEN_2067;
      end
    end else begin
      meta_array_37_2 <= _GEN_2067;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_37_3 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_3_1_REG) begin
      if (6'h25 == s1_way_waddr_3_1_r) begin
        meta_array_37_3 <= s1_way_wdata_3_1_r;
      end else begin
        meta_array_37_3 <= _GEN_2197;
      end
    end else begin
      meta_array_37_3 <= _GEN_2197;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_37_4 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_4_1_REG) begin
      if (6'h25 == s1_way_waddr_4_1_r) begin
        meta_array_37_4 <= s1_way_wdata_4_1_r;
      end else begin
        meta_array_37_4 <= _GEN_2327;
      end
    end else begin
      meta_array_37_4 <= _GEN_2327;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_37_5 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_5_1_REG) begin
      if (6'h25 == s1_way_waddr_5_1_r) begin
        meta_array_37_5 <= s1_way_wdata_5_1_r;
      end else begin
        meta_array_37_5 <= _GEN_2457;
      end
    end else begin
      meta_array_37_5 <= _GEN_2457;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_37_6 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_6_1_REG) begin
      if (6'h25 == s1_way_waddr_6_1_r) begin
        meta_array_37_6 <= s1_way_wdata_6_1_r;
      end else begin
        meta_array_37_6 <= _GEN_2587;
      end
    end else begin
      meta_array_37_6 <= _GEN_2587;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_37_7 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_7_1_REG) begin
      if (6'h25 == s1_way_waddr_7_1_r) begin
        meta_array_37_7 <= s1_way_wdata_7_1_r;
      end else begin
        meta_array_37_7 <= _GEN_2717;
      end
    end else begin
      meta_array_37_7 <= _GEN_2717;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_38_0 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_0_1_REG) begin
      if (6'h26 == s1_way_waddr_0_1_r) begin
        meta_array_38_0 <= s1_way_wdata_0_1_r;
      end else begin
        meta_array_38_0 <= _GEN_1808;
      end
    end else begin
      meta_array_38_0 <= _GEN_1808;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_38_1 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_1_1_REG) begin
      if (6'h26 == s1_way_waddr_1_1_r) begin
        meta_array_38_1 <= s1_way_wdata_1_1_r;
      end else begin
        meta_array_38_1 <= _GEN_1938;
      end
    end else begin
      meta_array_38_1 <= _GEN_1938;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_38_2 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_2_1_REG) begin
      if (6'h26 == s1_way_waddr_2_1_r) begin
        meta_array_38_2 <= s1_way_wdata_2_1_r;
      end else begin
        meta_array_38_2 <= _GEN_2068;
      end
    end else begin
      meta_array_38_2 <= _GEN_2068;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_38_3 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_3_1_REG) begin
      if (6'h26 == s1_way_waddr_3_1_r) begin
        meta_array_38_3 <= s1_way_wdata_3_1_r;
      end else begin
        meta_array_38_3 <= _GEN_2198;
      end
    end else begin
      meta_array_38_3 <= _GEN_2198;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_38_4 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_4_1_REG) begin
      if (6'h26 == s1_way_waddr_4_1_r) begin
        meta_array_38_4 <= s1_way_wdata_4_1_r;
      end else begin
        meta_array_38_4 <= _GEN_2328;
      end
    end else begin
      meta_array_38_4 <= _GEN_2328;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_38_5 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_5_1_REG) begin
      if (6'h26 == s1_way_waddr_5_1_r) begin
        meta_array_38_5 <= s1_way_wdata_5_1_r;
      end else begin
        meta_array_38_5 <= _GEN_2458;
      end
    end else begin
      meta_array_38_5 <= _GEN_2458;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_38_6 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_6_1_REG) begin
      if (6'h26 == s1_way_waddr_6_1_r) begin
        meta_array_38_6 <= s1_way_wdata_6_1_r;
      end else begin
        meta_array_38_6 <= _GEN_2588;
      end
    end else begin
      meta_array_38_6 <= _GEN_2588;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_38_7 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_7_1_REG) begin
      if (6'h26 == s1_way_waddr_7_1_r) begin
        meta_array_38_7 <= s1_way_wdata_7_1_r;
      end else begin
        meta_array_38_7 <= _GEN_2718;
      end
    end else begin
      meta_array_38_7 <= _GEN_2718;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_39_0 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_0_1_REG) begin
      if (6'h27 == s1_way_waddr_0_1_r) begin
        meta_array_39_0 <= s1_way_wdata_0_1_r;
      end else begin
        meta_array_39_0 <= _GEN_1809;
      end
    end else begin
      meta_array_39_0 <= _GEN_1809;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_39_1 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_1_1_REG) begin
      if (6'h27 == s1_way_waddr_1_1_r) begin
        meta_array_39_1 <= s1_way_wdata_1_1_r;
      end else begin
        meta_array_39_1 <= _GEN_1939;
      end
    end else begin
      meta_array_39_1 <= _GEN_1939;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_39_2 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_2_1_REG) begin
      if (6'h27 == s1_way_waddr_2_1_r) begin
        meta_array_39_2 <= s1_way_wdata_2_1_r;
      end else begin
        meta_array_39_2 <= _GEN_2069;
      end
    end else begin
      meta_array_39_2 <= _GEN_2069;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_39_3 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_3_1_REG) begin
      if (6'h27 == s1_way_waddr_3_1_r) begin
        meta_array_39_3 <= s1_way_wdata_3_1_r;
      end else begin
        meta_array_39_3 <= _GEN_2199;
      end
    end else begin
      meta_array_39_3 <= _GEN_2199;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_39_4 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_4_1_REG) begin
      if (6'h27 == s1_way_waddr_4_1_r) begin
        meta_array_39_4 <= s1_way_wdata_4_1_r;
      end else begin
        meta_array_39_4 <= _GEN_2329;
      end
    end else begin
      meta_array_39_4 <= _GEN_2329;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_39_5 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_5_1_REG) begin
      if (6'h27 == s1_way_waddr_5_1_r) begin
        meta_array_39_5 <= s1_way_wdata_5_1_r;
      end else begin
        meta_array_39_5 <= _GEN_2459;
      end
    end else begin
      meta_array_39_5 <= _GEN_2459;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_39_6 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_6_1_REG) begin
      if (6'h27 == s1_way_waddr_6_1_r) begin
        meta_array_39_6 <= s1_way_wdata_6_1_r;
      end else begin
        meta_array_39_6 <= _GEN_2589;
      end
    end else begin
      meta_array_39_6 <= _GEN_2589;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_39_7 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_7_1_REG) begin
      if (6'h27 == s1_way_waddr_7_1_r) begin
        meta_array_39_7 <= s1_way_wdata_7_1_r;
      end else begin
        meta_array_39_7 <= _GEN_2719;
      end
    end else begin
      meta_array_39_7 <= _GEN_2719;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_40_0 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_0_1_REG) begin
      if (6'h28 == s1_way_waddr_0_1_r) begin
        meta_array_40_0 <= s1_way_wdata_0_1_r;
      end else begin
        meta_array_40_0 <= _GEN_1810;
      end
    end else begin
      meta_array_40_0 <= _GEN_1810;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_40_1 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_1_1_REG) begin
      if (6'h28 == s1_way_waddr_1_1_r) begin
        meta_array_40_1 <= s1_way_wdata_1_1_r;
      end else begin
        meta_array_40_1 <= _GEN_1940;
      end
    end else begin
      meta_array_40_1 <= _GEN_1940;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_40_2 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_2_1_REG) begin
      if (6'h28 == s1_way_waddr_2_1_r) begin
        meta_array_40_2 <= s1_way_wdata_2_1_r;
      end else begin
        meta_array_40_2 <= _GEN_2070;
      end
    end else begin
      meta_array_40_2 <= _GEN_2070;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_40_3 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_3_1_REG) begin
      if (6'h28 == s1_way_waddr_3_1_r) begin
        meta_array_40_3 <= s1_way_wdata_3_1_r;
      end else begin
        meta_array_40_3 <= _GEN_2200;
      end
    end else begin
      meta_array_40_3 <= _GEN_2200;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_40_4 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_4_1_REG) begin
      if (6'h28 == s1_way_waddr_4_1_r) begin
        meta_array_40_4 <= s1_way_wdata_4_1_r;
      end else begin
        meta_array_40_4 <= _GEN_2330;
      end
    end else begin
      meta_array_40_4 <= _GEN_2330;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_40_5 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_5_1_REG) begin
      if (6'h28 == s1_way_waddr_5_1_r) begin
        meta_array_40_5 <= s1_way_wdata_5_1_r;
      end else begin
        meta_array_40_5 <= _GEN_2460;
      end
    end else begin
      meta_array_40_5 <= _GEN_2460;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_40_6 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_6_1_REG) begin
      if (6'h28 == s1_way_waddr_6_1_r) begin
        meta_array_40_6 <= s1_way_wdata_6_1_r;
      end else begin
        meta_array_40_6 <= _GEN_2590;
      end
    end else begin
      meta_array_40_6 <= _GEN_2590;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_40_7 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_7_1_REG) begin
      if (6'h28 == s1_way_waddr_7_1_r) begin
        meta_array_40_7 <= s1_way_wdata_7_1_r;
      end else begin
        meta_array_40_7 <= _GEN_2720;
      end
    end else begin
      meta_array_40_7 <= _GEN_2720;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_41_0 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_0_1_REG) begin
      if (6'h29 == s1_way_waddr_0_1_r) begin
        meta_array_41_0 <= s1_way_wdata_0_1_r;
      end else begin
        meta_array_41_0 <= _GEN_1811;
      end
    end else begin
      meta_array_41_0 <= _GEN_1811;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_41_1 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_1_1_REG) begin
      if (6'h29 == s1_way_waddr_1_1_r) begin
        meta_array_41_1 <= s1_way_wdata_1_1_r;
      end else begin
        meta_array_41_1 <= _GEN_1941;
      end
    end else begin
      meta_array_41_1 <= _GEN_1941;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_41_2 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_2_1_REG) begin
      if (6'h29 == s1_way_waddr_2_1_r) begin
        meta_array_41_2 <= s1_way_wdata_2_1_r;
      end else begin
        meta_array_41_2 <= _GEN_2071;
      end
    end else begin
      meta_array_41_2 <= _GEN_2071;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_41_3 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_3_1_REG) begin
      if (6'h29 == s1_way_waddr_3_1_r) begin
        meta_array_41_3 <= s1_way_wdata_3_1_r;
      end else begin
        meta_array_41_3 <= _GEN_2201;
      end
    end else begin
      meta_array_41_3 <= _GEN_2201;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_41_4 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_4_1_REG) begin
      if (6'h29 == s1_way_waddr_4_1_r) begin
        meta_array_41_4 <= s1_way_wdata_4_1_r;
      end else begin
        meta_array_41_4 <= _GEN_2331;
      end
    end else begin
      meta_array_41_4 <= _GEN_2331;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_41_5 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_5_1_REG) begin
      if (6'h29 == s1_way_waddr_5_1_r) begin
        meta_array_41_5 <= s1_way_wdata_5_1_r;
      end else begin
        meta_array_41_5 <= _GEN_2461;
      end
    end else begin
      meta_array_41_5 <= _GEN_2461;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_41_6 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_6_1_REG) begin
      if (6'h29 == s1_way_waddr_6_1_r) begin
        meta_array_41_6 <= s1_way_wdata_6_1_r;
      end else begin
        meta_array_41_6 <= _GEN_2591;
      end
    end else begin
      meta_array_41_6 <= _GEN_2591;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_41_7 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_7_1_REG) begin
      if (6'h29 == s1_way_waddr_7_1_r) begin
        meta_array_41_7 <= s1_way_wdata_7_1_r;
      end else begin
        meta_array_41_7 <= _GEN_2721;
      end
    end else begin
      meta_array_41_7 <= _GEN_2721;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_42_0 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_0_1_REG) begin
      if (6'h2a == s1_way_waddr_0_1_r) begin
        meta_array_42_0 <= s1_way_wdata_0_1_r;
      end else begin
        meta_array_42_0 <= _GEN_1812;
      end
    end else begin
      meta_array_42_0 <= _GEN_1812;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_42_1 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_1_1_REG) begin
      if (6'h2a == s1_way_waddr_1_1_r) begin
        meta_array_42_1 <= s1_way_wdata_1_1_r;
      end else begin
        meta_array_42_1 <= _GEN_1942;
      end
    end else begin
      meta_array_42_1 <= _GEN_1942;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_42_2 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_2_1_REG) begin
      if (6'h2a == s1_way_waddr_2_1_r) begin
        meta_array_42_2 <= s1_way_wdata_2_1_r;
      end else begin
        meta_array_42_2 <= _GEN_2072;
      end
    end else begin
      meta_array_42_2 <= _GEN_2072;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_42_3 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_3_1_REG) begin
      if (6'h2a == s1_way_waddr_3_1_r) begin
        meta_array_42_3 <= s1_way_wdata_3_1_r;
      end else begin
        meta_array_42_3 <= _GEN_2202;
      end
    end else begin
      meta_array_42_3 <= _GEN_2202;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_42_4 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_4_1_REG) begin
      if (6'h2a == s1_way_waddr_4_1_r) begin
        meta_array_42_4 <= s1_way_wdata_4_1_r;
      end else begin
        meta_array_42_4 <= _GEN_2332;
      end
    end else begin
      meta_array_42_4 <= _GEN_2332;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_42_5 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_5_1_REG) begin
      if (6'h2a == s1_way_waddr_5_1_r) begin
        meta_array_42_5 <= s1_way_wdata_5_1_r;
      end else begin
        meta_array_42_5 <= _GEN_2462;
      end
    end else begin
      meta_array_42_5 <= _GEN_2462;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_42_6 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_6_1_REG) begin
      if (6'h2a == s1_way_waddr_6_1_r) begin
        meta_array_42_6 <= s1_way_wdata_6_1_r;
      end else begin
        meta_array_42_6 <= _GEN_2592;
      end
    end else begin
      meta_array_42_6 <= _GEN_2592;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_42_7 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_7_1_REG) begin
      if (6'h2a == s1_way_waddr_7_1_r) begin
        meta_array_42_7 <= s1_way_wdata_7_1_r;
      end else begin
        meta_array_42_7 <= _GEN_2722;
      end
    end else begin
      meta_array_42_7 <= _GEN_2722;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_43_0 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_0_1_REG) begin
      if (6'h2b == s1_way_waddr_0_1_r) begin
        meta_array_43_0 <= s1_way_wdata_0_1_r;
      end else begin
        meta_array_43_0 <= _GEN_1813;
      end
    end else begin
      meta_array_43_0 <= _GEN_1813;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_43_1 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_1_1_REG) begin
      if (6'h2b == s1_way_waddr_1_1_r) begin
        meta_array_43_1 <= s1_way_wdata_1_1_r;
      end else begin
        meta_array_43_1 <= _GEN_1943;
      end
    end else begin
      meta_array_43_1 <= _GEN_1943;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_43_2 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_2_1_REG) begin
      if (6'h2b == s1_way_waddr_2_1_r) begin
        meta_array_43_2 <= s1_way_wdata_2_1_r;
      end else begin
        meta_array_43_2 <= _GEN_2073;
      end
    end else begin
      meta_array_43_2 <= _GEN_2073;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_43_3 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_3_1_REG) begin
      if (6'h2b == s1_way_waddr_3_1_r) begin
        meta_array_43_3 <= s1_way_wdata_3_1_r;
      end else begin
        meta_array_43_3 <= _GEN_2203;
      end
    end else begin
      meta_array_43_3 <= _GEN_2203;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_43_4 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_4_1_REG) begin
      if (6'h2b == s1_way_waddr_4_1_r) begin
        meta_array_43_4 <= s1_way_wdata_4_1_r;
      end else begin
        meta_array_43_4 <= _GEN_2333;
      end
    end else begin
      meta_array_43_4 <= _GEN_2333;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_43_5 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_5_1_REG) begin
      if (6'h2b == s1_way_waddr_5_1_r) begin
        meta_array_43_5 <= s1_way_wdata_5_1_r;
      end else begin
        meta_array_43_5 <= _GEN_2463;
      end
    end else begin
      meta_array_43_5 <= _GEN_2463;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_43_6 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_6_1_REG) begin
      if (6'h2b == s1_way_waddr_6_1_r) begin
        meta_array_43_6 <= s1_way_wdata_6_1_r;
      end else begin
        meta_array_43_6 <= _GEN_2593;
      end
    end else begin
      meta_array_43_6 <= _GEN_2593;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_43_7 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_7_1_REG) begin
      if (6'h2b == s1_way_waddr_7_1_r) begin
        meta_array_43_7 <= s1_way_wdata_7_1_r;
      end else begin
        meta_array_43_7 <= _GEN_2723;
      end
    end else begin
      meta_array_43_7 <= _GEN_2723;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_44_0 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_0_1_REG) begin
      if (6'h2c == s1_way_waddr_0_1_r) begin
        meta_array_44_0 <= s1_way_wdata_0_1_r;
      end else begin
        meta_array_44_0 <= _GEN_1814;
      end
    end else begin
      meta_array_44_0 <= _GEN_1814;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_44_1 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_1_1_REG) begin
      if (6'h2c == s1_way_waddr_1_1_r) begin
        meta_array_44_1 <= s1_way_wdata_1_1_r;
      end else begin
        meta_array_44_1 <= _GEN_1944;
      end
    end else begin
      meta_array_44_1 <= _GEN_1944;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_44_2 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_2_1_REG) begin
      if (6'h2c == s1_way_waddr_2_1_r) begin
        meta_array_44_2 <= s1_way_wdata_2_1_r;
      end else begin
        meta_array_44_2 <= _GEN_2074;
      end
    end else begin
      meta_array_44_2 <= _GEN_2074;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_44_3 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_3_1_REG) begin
      if (6'h2c == s1_way_waddr_3_1_r) begin
        meta_array_44_3 <= s1_way_wdata_3_1_r;
      end else begin
        meta_array_44_3 <= _GEN_2204;
      end
    end else begin
      meta_array_44_3 <= _GEN_2204;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_44_4 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_4_1_REG) begin
      if (6'h2c == s1_way_waddr_4_1_r) begin
        meta_array_44_4 <= s1_way_wdata_4_1_r;
      end else begin
        meta_array_44_4 <= _GEN_2334;
      end
    end else begin
      meta_array_44_4 <= _GEN_2334;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_44_5 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_5_1_REG) begin
      if (6'h2c == s1_way_waddr_5_1_r) begin
        meta_array_44_5 <= s1_way_wdata_5_1_r;
      end else begin
        meta_array_44_5 <= _GEN_2464;
      end
    end else begin
      meta_array_44_5 <= _GEN_2464;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_44_6 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_6_1_REG) begin
      if (6'h2c == s1_way_waddr_6_1_r) begin
        meta_array_44_6 <= s1_way_wdata_6_1_r;
      end else begin
        meta_array_44_6 <= _GEN_2594;
      end
    end else begin
      meta_array_44_6 <= _GEN_2594;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_44_7 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_7_1_REG) begin
      if (6'h2c == s1_way_waddr_7_1_r) begin
        meta_array_44_7 <= s1_way_wdata_7_1_r;
      end else begin
        meta_array_44_7 <= _GEN_2724;
      end
    end else begin
      meta_array_44_7 <= _GEN_2724;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_45_0 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_0_1_REG) begin
      if (6'h2d == s1_way_waddr_0_1_r) begin
        meta_array_45_0 <= s1_way_wdata_0_1_r;
      end else begin
        meta_array_45_0 <= _GEN_1815;
      end
    end else begin
      meta_array_45_0 <= _GEN_1815;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_45_1 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_1_1_REG) begin
      if (6'h2d == s1_way_waddr_1_1_r) begin
        meta_array_45_1 <= s1_way_wdata_1_1_r;
      end else begin
        meta_array_45_1 <= _GEN_1945;
      end
    end else begin
      meta_array_45_1 <= _GEN_1945;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_45_2 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_2_1_REG) begin
      if (6'h2d == s1_way_waddr_2_1_r) begin
        meta_array_45_2 <= s1_way_wdata_2_1_r;
      end else begin
        meta_array_45_2 <= _GEN_2075;
      end
    end else begin
      meta_array_45_2 <= _GEN_2075;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_45_3 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_3_1_REG) begin
      if (6'h2d == s1_way_waddr_3_1_r) begin
        meta_array_45_3 <= s1_way_wdata_3_1_r;
      end else begin
        meta_array_45_3 <= _GEN_2205;
      end
    end else begin
      meta_array_45_3 <= _GEN_2205;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_45_4 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_4_1_REG) begin
      if (6'h2d == s1_way_waddr_4_1_r) begin
        meta_array_45_4 <= s1_way_wdata_4_1_r;
      end else begin
        meta_array_45_4 <= _GEN_2335;
      end
    end else begin
      meta_array_45_4 <= _GEN_2335;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_45_5 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_5_1_REG) begin
      if (6'h2d == s1_way_waddr_5_1_r) begin
        meta_array_45_5 <= s1_way_wdata_5_1_r;
      end else begin
        meta_array_45_5 <= _GEN_2465;
      end
    end else begin
      meta_array_45_5 <= _GEN_2465;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_45_6 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_6_1_REG) begin
      if (6'h2d == s1_way_waddr_6_1_r) begin
        meta_array_45_6 <= s1_way_wdata_6_1_r;
      end else begin
        meta_array_45_6 <= _GEN_2595;
      end
    end else begin
      meta_array_45_6 <= _GEN_2595;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_45_7 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_7_1_REG) begin
      if (6'h2d == s1_way_waddr_7_1_r) begin
        meta_array_45_7 <= s1_way_wdata_7_1_r;
      end else begin
        meta_array_45_7 <= _GEN_2725;
      end
    end else begin
      meta_array_45_7 <= _GEN_2725;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_46_0 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_0_1_REG) begin
      if (6'h2e == s1_way_waddr_0_1_r) begin
        meta_array_46_0 <= s1_way_wdata_0_1_r;
      end else begin
        meta_array_46_0 <= _GEN_1816;
      end
    end else begin
      meta_array_46_0 <= _GEN_1816;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_46_1 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_1_1_REG) begin
      if (6'h2e == s1_way_waddr_1_1_r) begin
        meta_array_46_1 <= s1_way_wdata_1_1_r;
      end else begin
        meta_array_46_1 <= _GEN_1946;
      end
    end else begin
      meta_array_46_1 <= _GEN_1946;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_46_2 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_2_1_REG) begin
      if (6'h2e == s1_way_waddr_2_1_r) begin
        meta_array_46_2 <= s1_way_wdata_2_1_r;
      end else begin
        meta_array_46_2 <= _GEN_2076;
      end
    end else begin
      meta_array_46_2 <= _GEN_2076;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_46_3 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_3_1_REG) begin
      if (6'h2e == s1_way_waddr_3_1_r) begin
        meta_array_46_3 <= s1_way_wdata_3_1_r;
      end else begin
        meta_array_46_3 <= _GEN_2206;
      end
    end else begin
      meta_array_46_3 <= _GEN_2206;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_46_4 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_4_1_REG) begin
      if (6'h2e == s1_way_waddr_4_1_r) begin
        meta_array_46_4 <= s1_way_wdata_4_1_r;
      end else begin
        meta_array_46_4 <= _GEN_2336;
      end
    end else begin
      meta_array_46_4 <= _GEN_2336;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_46_5 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_5_1_REG) begin
      if (6'h2e == s1_way_waddr_5_1_r) begin
        meta_array_46_5 <= s1_way_wdata_5_1_r;
      end else begin
        meta_array_46_5 <= _GEN_2466;
      end
    end else begin
      meta_array_46_5 <= _GEN_2466;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_46_6 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_6_1_REG) begin
      if (6'h2e == s1_way_waddr_6_1_r) begin
        meta_array_46_6 <= s1_way_wdata_6_1_r;
      end else begin
        meta_array_46_6 <= _GEN_2596;
      end
    end else begin
      meta_array_46_6 <= _GEN_2596;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_46_7 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_7_1_REG) begin
      if (6'h2e == s1_way_waddr_7_1_r) begin
        meta_array_46_7 <= s1_way_wdata_7_1_r;
      end else begin
        meta_array_46_7 <= _GEN_2726;
      end
    end else begin
      meta_array_46_7 <= _GEN_2726;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_47_0 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_0_1_REG) begin
      if (6'h2f == s1_way_waddr_0_1_r) begin
        meta_array_47_0 <= s1_way_wdata_0_1_r;
      end else begin
        meta_array_47_0 <= _GEN_1817;
      end
    end else begin
      meta_array_47_0 <= _GEN_1817;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_47_1 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_1_1_REG) begin
      if (6'h2f == s1_way_waddr_1_1_r) begin
        meta_array_47_1 <= s1_way_wdata_1_1_r;
      end else begin
        meta_array_47_1 <= _GEN_1947;
      end
    end else begin
      meta_array_47_1 <= _GEN_1947;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_47_2 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_2_1_REG) begin
      if (6'h2f == s1_way_waddr_2_1_r) begin
        meta_array_47_2 <= s1_way_wdata_2_1_r;
      end else begin
        meta_array_47_2 <= _GEN_2077;
      end
    end else begin
      meta_array_47_2 <= _GEN_2077;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_47_3 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_3_1_REG) begin
      if (6'h2f == s1_way_waddr_3_1_r) begin
        meta_array_47_3 <= s1_way_wdata_3_1_r;
      end else begin
        meta_array_47_3 <= _GEN_2207;
      end
    end else begin
      meta_array_47_3 <= _GEN_2207;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_47_4 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_4_1_REG) begin
      if (6'h2f == s1_way_waddr_4_1_r) begin
        meta_array_47_4 <= s1_way_wdata_4_1_r;
      end else begin
        meta_array_47_4 <= _GEN_2337;
      end
    end else begin
      meta_array_47_4 <= _GEN_2337;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_47_5 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_5_1_REG) begin
      if (6'h2f == s1_way_waddr_5_1_r) begin
        meta_array_47_5 <= s1_way_wdata_5_1_r;
      end else begin
        meta_array_47_5 <= _GEN_2467;
      end
    end else begin
      meta_array_47_5 <= _GEN_2467;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_47_6 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_6_1_REG) begin
      if (6'h2f == s1_way_waddr_6_1_r) begin
        meta_array_47_6 <= s1_way_wdata_6_1_r;
      end else begin
        meta_array_47_6 <= _GEN_2597;
      end
    end else begin
      meta_array_47_6 <= _GEN_2597;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_47_7 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_7_1_REG) begin
      if (6'h2f == s1_way_waddr_7_1_r) begin
        meta_array_47_7 <= s1_way_wdata_7_1_r;
      end else begin
        meta_array_47_7 <= _GEN_2727;
      end
    end else begin
      meta_array_47_7 <= _GEN_2727;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_48_0 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_0_1_REG) begin
      if (6'h30 == s1_way_waddr_0_1_r) begin
        meta_array_48_0 <= s1_way_wdata_0_1_r;
      end else begin
        meta_array_48_0 <= _GEN_1818;
      end
    end else begin
      meta_array_48_0 <= _GEN_1818;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_48_1 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_1_1_REG) begin
      if (6'h30 == s1_way_waddr_1_1_r) begin
        meta_array_48_1 <= s1_way_wdata_1_1_r;
      end else begin
        meta_array_48_1 <= _GEN_1948;
      end
    end else begin
      meta_array_48_1 <= _GEN_1948;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_48_2 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_2_1_REG) begin
      if (6'h30 == s1_way_waddr_2_1_r) begin
        meta_array_48_2 <= s1_way_wdata_2_1_r;
      end else begin
        meta_array_48_2 <= _GEN_2078;
      end
    end else begin
      meta_array_48_2 <= _GEN_2078;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_48_3 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_3_1_REG) begin
      if (6'h30 == s1_way_waddr_3_1_r) begin
        meta_array_48_3 <= s1_way_wdata_3_1_r;
      end else begin
        meta_array_48_3 <= _GEN_2208;
      end
    end else begin
      meta_array_48_3 <= _GEN_2208;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_48_4 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_4_1_REG) begin
      if (6'h30 == s1_way_waddr_4_1_r) begin
        meta_array_48_4 <= s1_way_wdata_4_1_r;
      end else begin
        meta_array_48_4 <= _GEN_2338;
      end
    end else begin
      meta_array_48_4 <= _GEN_2338;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_48_5 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_5_1_REG) begin
      if (6'h30 == s1_way_waddr_5_1_r) begin
        meta_array_48_5 <= s1_way_wdata_5_1_r;
      end else begin
        meta_array_48_5 <= _GEN_2468;
      end
    end else begin
      meta_array_48_5 <= _GEN_2468;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_48_6 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_6_1_REG) begin
      if (6'h30 == s1_way_waddr_6_1_r) begin
        meta_array_48_6 <= s1_way_wdata_6_1_r;
      end else begin
        meta_array_48_6 <= _GEN_2598;
      end
    end else begin
      meta_array_48_6 <= _GEN_2598;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_48_7 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_7_1_REG) begin
      if (6'h30 == s1_way_waddr_7_1_r) begin
        meta_array_48_7 <= s1_way_wdata_7_1_r;
      end else begin
        meta_array_48_7 <= _GEN_2728;
      end
    end else begin
      meta_array_48_7 <= _GEN_2728;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_49_0 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_0_1_REG) begin
      if (6'h31 == s1_way_waddr_0_1_r) begin
        meta_array_49_0 <= s1_way_wdata_0_1_r;
      end else begin
        meta_array_49_0 <= _GEN_1819;
      end
    end else begin
      meta_array_49_0 <= _GEN_1819;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_49_1 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_1_1_REG) begin
      if (6'h31 == s1_way_waddr_1_1_r) begin
        meta_array_49_1 <= s1_way_wdata_1_1_r;
      end else begin
        meta_array_49_1 <= _GEN_1949;
      end
    end else begin
      meta_array_49_1 <= _GEN_1949;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_49_2 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_2_1_REG) begin
      if (6'h31 == s1_way_waddr_2_1_r) begin
        meta_array_49_2 <= s1_way_wdata_2_1_r;
      end else begin
        meta_array_49_2 <= _GEN_2079;
      end
    end else begin
      meta_array_49_2 <= _GEN_2079;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_49_3 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_3_1_REG) begin
      if (6'h31 == s1_way_waddr_3_1_r) begin
        meta_array_49_3 <= s1_way_wdata_3_1_r;
      end else begin
        meta_array_49_3 <= _GEN_2209;
      end
    end else begin
      meta_array_49_3 <= _GEN_2209;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_49_4 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_4_1_REG) begin
      if (6'h31 == s1_way_waddr_4_1_r) begin
        meta_array_49_4 <= s1_way_wdata_4_1_r;
      end else begin
        meta_array_49_4 <= _GEN_2339;
      end
    end else begin
      meta_array_49_4 <= _GEN_2339;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_49_5 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_5_1_REG) begin
      if (6'h31 == s1_way_waddr_5_1_r) begin
        meta_array_49_5 <= s1_way_wdata_5_1_r;
      end else begin
        meta_array_49_5 <= _GEN_2469;
      end
    end else begin
      meta_array_49_5 <= _GEN_2469;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_49_6 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_6_1_REG) begin
      if (6'h31 == s1_way_waddr_6_1_r) begin
        meta_array_49_6 <= s1_way_wdata_6_1_r;
      end else begin
        meta_array_49_6 <= _GEN_2599;
      end
    end else begin
      meta_array_49_6 <= _GEN_2599;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_49_7 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_7_1_REG) begin
      if (6'h31 == s1_way_waddr_7_1_r) begin
        meta_array_49_7 <= s1_way_wdata_7_1_r;
      end else begin
        meta_array_49_7 <= _GEN_2729;
      end
    end else begin
      meta_array_49_7 <= _GEN_2729;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_50_0 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_0_1_REG) begin
      if (6'h32 == s1_way_waddr_0_1_r) begin
        meta_array_50_0 <= s1_way_wdata_0_1_r;
      end else begin
        meta_array_50_0 <= _GEN_1820;
      end
    end else begin
      meta_array_50_0 <= _GEN_1820;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_50_1 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_1_1_REG) begin
      if (6'h32 == s1_way_waddr_1_1_r) begin
        meta_array_50_1 <= s1_way_wdata_1_1_r;
      end else begin
        meta_array_50_1 <= _GEN_1950;
      end
    end else begin
      meta_array_50_1 <= _GEN_1950;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_50_2 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_2_1_REG) begin
      if (6'h32 == s1_way_waddr_2_1_r) begin
        meta_array_50_2 <= s1_way_wdata_2_1_r;
      end else begin
        meta_array_50_2 <= _GEN_2080;
      end
    end else begin
      meta_array_50_2 <= _GEN_2080;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_50_3 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_3_1_REG) begin
      if (6'h32 == s1_way_waddr_3_1_r) begin
        meta_array_50_3 <= s1_way_wdata_3_1_r;
      end else begin
        meta_array_50_3 <= _GEN_2210;
      end
    end else begin
      meta_array_50_3 <= _GEN_2210;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_50_4 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_4_1_REG) begin
      if (6'h32 == s1_way_waddr_4_1_r) begin
        meta_array_50_4 <= s1_way_wdata_4_1_r;
      end else begin
        meta_array_50_4 <= _GEN_2340;
      end
    end else begin
      meta_array_50_4 <= _GEN_2340;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_50_5 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_5_1_REG) begin
      if (6'h32 == s1_way_waddr_5_1_r) begin
        meta_array_50_5 <= s1_way_wdata_5_1_r;
      end else begin
        meta_array_50_5 <= _GEN_2470;
      end
    end else begin
      meta_array_50_5 <= _GEN_2470;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_50_6 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_6_1_REG) begin
      if (6'h32 == s1_way_waddr_6_1_r) begin
        meta_array_50_6 <= s1_way_wdata_6_1_r;
      end else begin
        meta_array_50_6 <= _GEN_2600;
      end
    end else begin
      meta_array_50_6 <= _GEN_2600;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_50_7 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_7_1_REG) begin
      if (6'h32 == s1_way_waddr_7_1_r) begin
        meta_array_50_7 <= s1_way_wdata_7_1_r;
      end else begin
        meta_array_50_7 <= _GEN_2730;
      end
    end else begin
      meta_array_50_7 <= _GEN_2730;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_51_0 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_0_1_REG) begin
      if (6'h33 == s1_way_waddr_0_1_r) begin
        meta_array_51_0 <= s1_way_wdata_0_1_r;
      end else begin
        meta_array_51_0 <= _GEN_1821;
      end
    end else begin
      meta_array_51_0 <= _GEN_1821;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_51_1 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_1_1_REG) begin
      if (6'h33 == s1_way_waddr_1_1_r) begin
        meta_array_51_1 <= s1_way_wdata_1_1_r;
      end else begin
        meta_array_51_1 <= _GEN_1951;
      end
    end else begin
      meta_array_51_1 <= _GEN_1951;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_51_2 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_2_1_REG) begin
      if (6'h33 == s1_way_waddr_2_1_r) begin
        meta_array_51_2 <= s1_way_wdata_2_1_r;
      end else begin
        meta_array_51_2 <= _GEN_2081;
      end
    end else begin
      meta_array_51_2 <= _GEN_2081;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_51_3 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_3_1_REG) begin
      if (6'h33 == s1_way_waddr_3_1_r) begin
        meta_array_51_3 <= s1_way_wdata_3_1_r;
      end else begin
        meta_array_51_3 <= _GEN_2211;
      end
    end else begin
      meta_array_51_3 <= _GEN_2211;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_51_4 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_4_1_REG) begin
      if (6'h33 == s1_way_waddr_4_1_r) begin
        meta_array_51_4 <= s1_way_wdata_4_1_r;
      end else begin
        meta_array_51_4 <= _GEN_2341;
      end
    end else begin
      meta_array_51_4 <= _GEN_2341;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_51_5 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_5_1_REG) begin
      if (6'h33 == s1_way_waddr_5_1_r) begin
        meta_array_51_5 <= s1_way_wdata_5_1_r;
      end else begin
        meta_array_51_5 <= _GEN_2471;
      end
    end else begin
      meta_array_51_5 <= _GEN_2471;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_51_6 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_6_1_REG) begin
      if (6'h33 == s1_way_waddr_6_1_r) begin
        meta_array_51_6 <= s1_way_wdata_6_1_r;
      end else begin
        meta_array_51_6 <= _GEN_2601;
      end
    end else begin
      meta_array_51_6 <= _GEN_2601;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_51_7 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_7_1_REG) begin
      if (6'h33 == s1_way_waddr_7_1_r) begin
        meta_array_51_7 <= s1_way_wdata_7_1_r;
      end else begin
        meta_array_51_7 <= _GEN_2731;
      end
    end else begin
      meta_array_51_7 <= _GEN_2731;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_52_0 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_0_1_REG) begin
      if (6'h34 == s1_way_waddr_0_1_r) begin
        meta_array_52_0 <= s1_way_wdata_0_1_r;
      end else begin
        meta_array_52_0 <= _GEN_1822;
      end
    end else begin
      meta_array_52_0 <= _GEN_1822;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_52_1 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_1_1_REG) begin
      if (6'h34 == s1_way_waddr_1_1_r) begin
        meta_array_52_1 <= s1_way_wdata_1_1_r;
      end else begin
        meta_array_52_1 <= _GEN_1952;
      end
    end else begin
      meta_array_52_1 <= _GEN_1952;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_52_2 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_2_1_REG) begin
      if (6'h34 == s1_way_waddr_2_1_r) begin
        meta_array_52_2 <= s1_way_wdata_2_1_r;
      end else begin
        meta_array_52_2 <= _GEN_2082;
      end
    end else begin
      meta_array_52_2 <= _GEN_2082;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_52_3 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_3_1_REG) begin
      if (6'h34 == s1_way_waddr_3_1_r) begin
        meta_array_52_3 <= s1_way_wdata_3_1_r;
      end else begin
        meta_array_52_3 <= _GEN_2212;
      end
    end else begin
      meta_array_52_3 <= _GEN_2212;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_52_4 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_4_1_REG) begin
      if (6'h34 == s1_way_waddr_4_1_r) begin
        meta_array_52_4 <= s1_way_wdata_4_1_r;
      end else begin
        meta_array_52_4 <= _GEN_2342;
      end
    end else begin
      meta_array_52_4 <= _GEN_2342;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_52_5 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_5_1_REG) begin
      if (6'h34 == s1_way_waddr_5_1_r) begin
        meta_array_52_5 <= s1_way_wdata_5_1_r;
      end else begin
        meta_array_52_5 <= _GEN_2472;
      end
    end else begin
      meta_array_52_5 <= _GEN_2472;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_52_6 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_6_1_REG) begin
      if (6'h34 == s1_way_waddr_6_1_r) begin
        meta_array_52_6 <= s1_way_wdata_6_1_r;
      end else begin
        meta_array_52_6 <= _GEN_2602;
      end
    end else begin
      meta_array_52_6 <= _GEN_2602;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_52_7 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_7_1_REG) begin
      if (6'h34 == s1_way_waddr_7_1_r) begin
        meta_array_52_7 <= s1_way_wdata_7_1_r;
      end else begin
        meta_array_52_7 <= _GEN_2732;
      end
    end else begin
      meta_array_52_7 <= _GEN_2732;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_53_0 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_0_1_REG) begin
      if (6'h35 == s1_way_waddr_0_1_r) begin
        meta_array_53_0 <= s1_way_wdata_0_1_r;
      end else begin
        meta_array_53_0 <= _GEN_1823;
      end
    end else begin
      meta_array_53_0 <= _GEN_1823;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_53_1 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_1_1_REG) begin
      if (6'h35 == s1_way_waddr_1_1_r) begin
        meta_array_53_1 <= s1_way_wdata_1_1_r;
      end else begin
        meta_array_53_1 <= _GEN_1953;
      end
    end else begin
      meta_array_53_1 <= _GEN_1953;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_53_2 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_2_1_REG) begin
      if (6'h35 == s1_way_waddr_2_1_r) begin
        meta_array_53_2 <= s1_way_wdata_2_1_r;
      end else begin
        meta_array_53_2 <= _GEN_2083;
      end
    end else begin
      meta_array_53_2 <= _GEN_2083;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_53_3 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_3_1_REG) begin
      if (6'h35 == s1_way_waddr_3_1_r) begin
        meta_array_53_3 <= s1_way_wdata_3_1_r;
      end else begin
        meta_array_53_3 <= _GEN_2213;
      end
    end else begin
      meta_array_53_3 <= _GEN_2213;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_53_4 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_4_1_REG) begin
      if (6'h35 == s1_way_waddr_4_1_r) begin
        meta_array_53_4 <= s1_way_wdata_4_1_r;
      end else begin
        meta_array_53_4 <= _GEN_2343;
      end
    end else begin
      meta_array_53_4 <= _GEN_2343;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_53_5 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_5_1_REG) begin
      if (6'h35 == s1_way_waddr_5_1_r) begin
        meta_array_53_5 <= s1_way_wdata_5_1_r;
      end else begin
        meta_array_53_5 <= _GEN_2473;
      end
    end else begin
      meta_array_53_5 <= _GEN_2473;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_53_6 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_6_1_REG) begin
      if (6'h35 == s1_way_waddr_6_1_r) begin
        meta_array_53_6 <= s1_way_wdata_6_1_r;
      end else begin
        meta_array_53_6 <= _GEN_2603;
      end
    end else begin
      meta_array_53_6 <= _GEN_2603;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_53_7 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_7_1_REG) begin
      if (6'h35 == s1_way_waddr_7_1_r) begin
        meta_array_53_7 <= s1_way_wdata_7_1_r;
      end else begin
        meta_array_53_7 <= _GEN_2733;
      end
    end else begin
      meta_array_53_7 <= _GEN_2733;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_54_0 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_0_1_REG) begin
      if (6'h36 == s1_way_waddr_0_1_r) begin
        meta_array_54_0 <= s1_way_wdata_0_1_r;
      end else begin
        meta_array_54_0 <= _GEN_1824;
      end
    end else begin
      meta_array_54_0 <= _GEN_1824;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_54_1 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_1_1_REG) begin
      if (6'h36 == s1_way_waddr_1_1_r) begin
        meta_array_54_1 <= s1_way_wdata_1_1_r;
      end else begin
        meta_array_54_1 <= _GEN_1954;
      end
    end else begin
      meta_array_54_1 <= _GEN_1954;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_54_2 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_2_1_REG) begin
      if (6'h36 == s1_way_waddr_2_1_r) begin
        meta_array_54_2 <= s1_way_wdata_2_1_r;
      end else begin
        meta_array_54_2 <= _GEN_2084;
      end
    end else begin
      meta_array_54_2 <= _GEN_2084;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_54_3 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_3_1_REG) begin
      if (6'h36 == s1_way_waddr_3_1_r) begin
        meta_array_54_3 <= s1_way_wdata_3_1_r;
      end else begin
        meta_array_54_3 <= _GEN_2214;
      end
    end else begin
      meta_array_54_3 <= _GEN_2214;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_54_4 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_4_1_REG) begin
      if (6'h36 == s1_way_waddr_4_1_r) begin
        meta_array_54_4 <= s1_way_wdata_4_1_r;
      end else begin
        meta_array_54_4 <= _GEN_2344;
      end
    end else begin
      meta_array_54_4 <= _GEN_2344;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_54_5 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_5_1_REG) begin
      if (6'h36 == s1_way_waddr_5_1_r) begin
        meta_array_54_5 <= s1_way_wdata_5_1_r;
      end else begin
        meta_array_54_5 <= _GEN_2474;
      end
    end else begin
      meta_array_54_5 <= _GEN_2474;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_54_6 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_6_1_REG) begin
      if (6'h36 == s1_way_waddr_6_1_r) begin
        meta_array_54_6 <= s1_way_wdata_6_1_r;
      end else begin
        meta_array_54_6 <= _GEN_2604;
      end
    end else begin
      meta_array_54_6 <= _GEN_2604;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_54_7 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_7_1_REG) begin
      if (6'h36 == s1_way_waddr_7_1_r) begin
        meta_array_54_7 <= s1_way_wdata_7_1_r;
      end else begin
        meta_array_54_7 <= _GEN_2734;
      end
    end else begin
      meta_array_54_7 <= _GEN_2734;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_55_0 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_0_1_REG) begin
      if (6'h37 == s1_way_waddr_0_1_r) begin
        meta_array_55_0 <= s1_way_wdata_0_1_r;
      end else begin
        meta_array_55_0 <= _GEN_1825;
      end
    end else begin
      meta_array_55_0 <= _GEN_1825;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_55_1 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_1_1_REG) begin
      if (6'h37 == s1_way_waddr_1_1_r) begin
        meta_array_55_1 <= s1_way_wdata_1_1_r;
      end else begin
        meta_array_55_1 <= _GEN_1955;
      end
    end else begin
      meta_array_55_1 <= _GEN_1955;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_55_2 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_2_1_REG) begin
      if (6'h37 == s1_way_waddr_2_1_r) begin
        meta_array_55_2 <= s1_way_wdata_2_1_r;
      end else begin
        meta_array_55_2 <= _GEN_2085;
      end
    end else begin
      meta_array_55_2 <= _GEN_2085;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_55_3 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_3_1_REG) begin
      if (6'h37 == s1_way_waddr_3_1_r) begin
        meta_array_55_3 <= s1_way_wdata_3_1_r;
      end else begin
        meta_array_55_3 <= _GEN_2215;
      end
    end else begin
      meta_array_55_3 <= _GEN_2215;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_55_4 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_4_1_REG) begin
      if (6'h37 == s1_way_waddr_4_1_r) begin
        meta_array_55_4 <= s1_way_wdata_4_1_r;
      end else begin
        meta_array_55_4 <= _GEN_2345;
      end
    end else begin
      meta_array_55_4 <= _GEN_2345;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_55_5 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_5_1_REG) begin
      if (6'h37 == s1_way_waddr_5_1_r) begin
        meta_array_55_5 <= s1_way_wdata_5_1_r;
      end else begin
        meta_array_55_5 <= _GEN_2475;
      end
    end else begin
      meta_array_55_5 <= _GEN_2475;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_55_6 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_6_1_REG) begin
      if (6'h37 == s1_way_waddr_6_1_r) begin
        meta_array_55_6 <= s1_way_wdata_6_1_r;
      end else begin
        meta_array_55_6 <= _GEN_2605;
      end
    end else begin
      meta_array_55_6 <= _GEN_2605;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_55_7 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_7_1_REG) begin
      if (6'h37 == s1_way_waddr_7_1_r) begin
        meta_array_55_7 <= s1_way_wdata_7_1_r;
      end else begin
        meta_array_55_7 <= _GEN_2735;
      end
    end else begin
      meta_array_55_7 <= _GEN_2735;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_56_0 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_0_1_REG) begin
      if (6'h38 == s1_way_waddr_0_1_r) begin
        meta_array_56_0 <= s1_way_wdata_0_1_r;
      end else begin
        meta_array_56_0 <= _GEN_1826;
      end
    end else begin
      meta_array_56_0 <= _GEN_1826;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_56_1 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_1_1_REG) begin
      if (6'h38 == s1_way_waddr_1_1_r) begin
        meta_array_56_1 <= s1_way_wdata_1_1_r;
      end else begin
        meta_array_56_1 <= _GEN_1956;
      end
    end else begin
      meta_array_56_1 <= _GEN_1956;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_56_2 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_2_1_REG) begin
      if (6'h38 == s1_way_waddr_2_1_r) begin
        meta_array_56_2 <= s1_way_wdata_2_1_r;
      end else begin
        meta_array_56_2 <= _GEN_2086;
      end
    end else begin
      meta_array_56_2 <= _GEN_2086;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_56_3 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_3_1_REG) begin
      if (6'h38 == s1_way_waddr_3_1_r) begin
        meta_array_56_3 <= s1_way_wdata_3_1_r;
      end else begin
        meta_array_56_3 <= _GEN_2216;
      end
    end else begin
      meta_array_56_3 <= _GEN_2216;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_56_4 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_4_1_REG) begin
      if (6'h38 == s1_way_waddr_4_1_r) begin
        meta_array_56_4 <= s1_way_wdata_4_1_r;
      end else begin
        meta_array_56_4 <= _GEN_2346;
      end
    end else begin
      meta_array_56_4 <= _GEN_2346;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_56_5 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_5_1_REG) begin
      if (6'h38 == s1_way_waddr_5_1_r) begin
        meta_array_56_5 <= s1_way_wdata_5_1_r;
      end else begin
        meta_array_56_5 <= _GEN_2476;
      end
    end else begin
      meta_array_56_5 <= _GEN_2476;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_56_6 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_6_1_REG) begin
      if (6'h38 == s1_way_waddr_6_1_r) begin
        meta_array_56_6 <= s1_way_wdata_6_1_r;
      end else begin
        meta_array_56_6 <= _GEN_2606;
      end
    end else begin
      meta_array_56_6 <= _GEN_2606;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_56_7 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_7_1_REG) begin
      if (6'h38 == s1_way_waddr_7_1_r) begin
        meta_array_56_7 <= s1_way_wdata_7_1_r;
      end else begin
        meta_array_56_7 <= _GEN_2736;
      end
    end else begin
      meta_array_56_7 <= _GEN_2736;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_57_0 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_0_1_REG) begin
      if (6'h39 == s1_way_waddr_0_1_r) begin
        meta_array_57_0 <= s1_way_wdata_0_1_r;
      end else begin
        meta_array_57_0 <= _GEN_1827;
      end
    end else begin
      meta_array_57_0 <= _GEN_1827;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_57_1 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_1_1_REG) begin
      if (6'h39 == s1_way_waddr_1_1_r) begin
        meta_array_57_1 <= s1_way_wdata_1_1_r;
      end else begin
        meta_array_57_1 <= _GEN_1957;
      end
    end else begin
      meta_array_57_1 <= _GEN_1957;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_57_2 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_2_1_REG) begin
      if (6'h39 == s1_way_waddr_2_1_r) begin
        meta_array_57_2 <= s1_way_wdata_2_1_r;
      end else begin
        meta_array_57_2 <= _GEN_2087;
      end
    end else begin
      meta_array_57_2 <= _GEN_2087;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_57_3 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_3_1_REG) begin
      if (6'h39 == s1_way_waddr_3_1_r) begin
        meta_array_57_3 <= s1_way_wdata_3_1_r;
      end else begin
        meta_array_57_3 <= _GEN_2217;
      end
    end else begin
      meta_array_57_3 <= _GEN_2217;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_57_4 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_4_1_REG) begin
      if (6'h39 == s1_way_waddr_4_1_r) begin
        meta_array_57_4 <= s1_way_wdata_4_1_r;
      end else begin
        meta_array_57_4 <= _GEN_2347;
      end
    end else begin
      meta_array_57_4 <= _GEN_2347;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_57_5 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_5_1_REG) begin
      if (6'h39 == s1_way_waddr_5_1_r) begin
        meta_array_57_5 <= s1_way_wdata_5_1_r;
      end else begin
        meta_array_57_5 <= _GEN_2477;
      end
    end else begin
      meta_array_57_5 <= _GEN_2477;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_57_6 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_6_1_REG) begin
      if (6'h39 == s1_way_waddr_6_1_r) begin
        meta_array_57_6 <= s1_way_wdata_6_1_r;
      end else begin
        meta_array_57_6 <= _GEN_2607;
      end
    end else begin
      meta_array_57_6 <= _GEN_2607;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_57_7 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_7_1_REG) begin
      if (6'h39 == s1_way_waddr_7_1_r) begin
        meta_array_57_7 <= s1_way_wdata_7_1_r;
      end else begin
        meta_array_57_7 <= _GEN_2737;
      end
    end else begin
      meta_array_57_7 <= _GEN_2737;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_58_0 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_0_1_REG) begin
      if (6'h3a == s1_way_waddr_0_1_r) begin
        meta_array_58_0 <= s1_way_wdata_0_1_r;
      end else begin
        meta_array_58_0 <= _GEN_1828;
      end
    end else begin
      meta_array_58_0 <= _GEN_1828;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_58_1 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_1_1_REG) begin
      if (6'h3a == s1_way_waddr_1_1_r) begin
        meta_array_58_1 <= s1_way_wdata_1_1_r;
      end else begin
        meta_array_58_1 <= _GEN_1958;
      end
    end else begin
      meta_array_58_1 <= _GEN_1958;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_58_2 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_2_1_REG) begin
      if (6'h3a == s1_way_waddr_2_1_r) begin
        meta_array_58_2 <= s1_way_wdata_2_1_r;
      end else begin
        meta_array_58_2 <= _GEN_2088;
      end
    end else begin
      meta_array_58_2 <= _GEN_2088;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_58_3 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_3_1_REG) begin
      if (6'h3a == s1_way_waddr_3_1_r) begin
        meta_array_58_3 <= s1_way_wdata_3_1_r;
      end else begin
        meta_array_58_3 <= _GEN_2218;
      end
    end else begin
      meta_array_58_3 <= _GEN_2218;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_58_4 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_4_1_REG) begin
      if (6'h3a == s1_way_waddr_4_1_r) begin
        meta_array_58_4 <= s1_way_wdata_4_1_r;
      end else begin
        meta_array_58_4 <= _GEN_2348;
      end
    end else begin
      meta_array_58_4 <= _GEN_2348;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_58_5 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_5_1_REG) begin
      if (6'h3a == s1_way_waddr_5_1_r) begin
        meta_array_58_5 <= s1_way_wdata_5_1_r;
      end else begin
        meta_array_58_5 <= _GEN_2478;
      end
    end else begin
      meta_array_58_5 <= _GEN_2478;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_58_6 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_6_1_REG) begin
      if (6'h3a == s1_way_waddr_6_1_r) begin
        meta_array_58_6 <= s1_way_wdata_6_1_r;
      end else begin
        meta_array_58_6 <= _GEN_2608;
      end
    end else begin
      meta_array_58_6 <= _GEN_2608;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_58_7 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_7_1_REG) begin
      if (6'h3a == s1_way_waddr_7_1_r) begin
        meta_array_58_7 <= s1_way_wdata_7_1_r;
      end else begin
        meta_array_58_7 <= _GEN_2738;
      end
    end else begin
      meta_array_58_7 <= _GEN_2738;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_59_0 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_0_1_REG) begin
      if (6'h3b == s1_way_waddr_0_1_r) begin
        meta_array_59_0 <= s1_way_wdata_0_1_r;
      end else begin
        meta_array_59_0 <= _GEN_1829;
      end
    end else begin
      meta_array_59_0 <= _GEN_1829;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_59_1 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_1_1_REG) begin
      if (6'h3b == s1_way_waddr_1_1_r) begin
        meta_array_59_1 <= s1_way_wdata_1_1_r;
      end else begin
        meta_array_59_1 <= _GEN_1959;
      end
    end else begin
      meta_array_59_1 <= _GEN_1959;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_59_2 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_2_1_REG) begin
      if (6'h3b == s1_way_waddr_2_1_r) begin
        meta_array_59_2 <= s1_way_wdata_2_1_r;
      end else begin
        meta_array_59_2 <= _GEN_2089;
      end
    end else begin
      meta_array_59_2 <= _GEN_2089;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_59_3 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_3_1_REG) begin
      if (6'h3b == s1_way_waddr_3_1_r) begin
        meta_array_59_3 <= s1_way_wdata_3_1_r;
      end else begin
        meta_array_59_3 <= _GEN_2219;
      end
    end else begin
      meta_array_59_3 <= _GEN_2219;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_59_4 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_4_1_REG) begin
      if (6'h3b == s1_way_waddr_4_1_r) begin
        meta_array_59_4 <= s1_way_wdata_4_1_r;
      end else begin
        meta_array_59_4 <= _GEN_2349;
      end
    end else begin
      meta_array_59_4 <= _GEN_2349;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_59_5 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_5_1_REG) begin
      if (6'h3b == s1_way_waddr_5_1_r) begin
        meta_array_59_5 <= s1_way_wdata_5_1_r;
      end else begin
        meta_array_59_5 <= _GEN_2479;
      end
    end else begin
      meta_array_59_5 <= _GEN_2479;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_59_6 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_6_1_REG) begin
      if (6'h3b == s1_way_waddr_6_1_r) begin
        meta_array_59_6 <= s1_way_wdata_6_1_r;
      end else begin
        meta_array_59_6 <= _GEN_2609;
      end
    end else begin
      meta_array_59_6 <= _GEN_2609;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_59_7 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_7_1_REG) begin
      if (6'h3b == s1_way_waddr_7_1_r) begin
        meta_array_59_7 <= s1_way_wdata_7_1_r;
      end else begin
        meta_array_59_7 <= _GEN_2739;
      end
    end else begin
      meta_array_59_7 <= _GEN_2739;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_60_0 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_0_1_REG) begin
      if (6'h3c == s1_way_waddr_0_1_r) begin
        meta_array_60_0 <= s1_way_wdata_0_1_r;
      end else begin
        meta_array_60_0 <= _GEN_1830;
      end
    end else begin
      meta_array_60_0 <= _GEN_1830;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_60_1 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_1_1_REG) begin
      if (6'h3c == s1_way_waddr_1_1_r) begin
        meta_array_60_1 <= s1_way_wdata_1_1_r;
      end else begin
        meta_array_60_1 <= _GEN_1960;
      end
    end else begin
      meta_array_60_1 <= _GEN_1960;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_60_2 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_2_1_REG) begin
      if (6'h3c == s1_way_waddr_2_1_r) begin
        meta_array_60_2 <= s1_way_wdata_2_1_r;
      end else begin
        meta_array_60_2 <= _GEN_2090;
      end
    end else begin
      meta_array_60_2 <= _GEN_2090;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_60_3 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_3_1_REG) begin
      if (6'h3c == s1_way_waddr_3_1_r) begin
        meta_array_60_3 <= s1_way_wdata_3_1_r;
      end else begin
        meta_array_60_3 <= _GEN_2220;
      end
    end else begin
      meta_array_60_3 <= _GEN_2220;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_60_4 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_4_1_REG) begin
      if (6'h3c == s1_way_waddr_4_1_r) begin
        meta_array_60_4 <= s1_way_wdata_4_1_r;
      end else begin
        meta_array_60_4 <= _GEN_2350;
      end
    end else begin
      meta_array_60_4 <= _GEN_2350;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_60_5 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_5_1_REG) begin
      if (6'h3c == s1_way_waddr_5_1_r) begin
        meta_array_60_5 <= s1_way_wdata_5_1_r;
      end else begin
        meta_array_60_5 <= _GEN_2480;
      end
    end else begin
      meta_array_60_5 <= _GEN_2480;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_60_6 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_6_1_REG) begin
      if (6'h3c == s1_way_waddr_6_1_r) begin
        meta_array_60_6 <= s1_way_wdata_6_1_r;
      end else begin
        meta_array_60_6 <= _GEN_2610;
      end
    end else begin
      meta_array_60_6 <= _GEN_2610;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_60_7 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_7_1_REG) begin
      if (6'h3c == s1_way_waddr_7_1_r) begin
        meta_array_60_7 <= s1_way_wdata_7_1_r;
      end else begin
        meta_array_60_7 <= _GEN_2740;
      end
    end else begin
      meta_array_60_7 <= _GEN_2740;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_61_0 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_0_1_REG) begin
      if (6'h3d == s1_way_waddr_0_1_r) begin
        meta_array_61_0 <= s1_way_wdata_0_1_r;
      end else begin
        meta_array_61_0 <= _GEN_1831;
      end
    end else begin
      meta_array_61_0 <= _GEN_1831;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_61_1 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_1_1_REG) begin
      if (6'h3d == s1_way_waddr_1_1_r) begin
        meta_array_61_1 <= s1_way_wdata_1_1_r;
      end else begin
        meta_array_61_1 <= _GEN_1961;
      end
    end else begin
      meta_array_61_1 <= _GEN_1961;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_61_2 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_2_1_REG) begin
      if (6'h3d == s1_way_waddr_2_1_r) begin
        meta_array_61_2 <= s1_way_wdata_2_1_r;
      end else begin
        meta_array_61_2 <= _GEN_2091;
      end
    end else begin
      meta_array_61_2 <= _GEN_2091;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_61_3 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_3_1_REG) begin
      if (6'h3d == s1_way_waddr_3_1_r) begin
        meta_array_61_3 <= s1_way_wdata_3_1_r;
      end else begin
        meta_array_61_3 <= _GEN_2221;
      end
    end else begin
      meta_array_61_3 <= _GEN_2221;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_61_4 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_4_1_REG) begin
      if (6'h3d == s1_way_waddr_4_1_r) begin
        meta_array_61_4 <= s1_way_wdata_4_1_r;
      end else begin
        meta_array_61_4 <= _GEN_2351;
      end
    end else begin
      meta_array_61_4 <= _GEN_2351;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_61_5 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_5_1_REG) begin
      if (6'h3d == s1_way_waddr_5_1_r) begin
        meta_array_61_5 <= s1_way_wdata_5_1_r;
      end else begin
        meta_array_61_5 <= _GEN_2481;
      end
    end else begin
      meta_array_61_5 <= _GEN_2481;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_61_6 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_6_1_REG) begin
      if (6'h3d == s1_way_waddr_6_1_r) begin
        meta_array_61_6 <= s1_way_wdata_6_1_r;
      end else begin
        meta_array_61_6 <= _GEN_2611;
      end
    end else begin
      meta_array_61_6 <= _GEN_2611;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_61_7 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_7_1_REG) begin
      if (6'h3d == s1_way_waddr_7_1_r) begin
        meta_array_61_7 <= s1_way_wdata_7_1_r;
      end else begin
        meta_array_61_7 <= _GEN_2741;
      end
    end else begin
      meta_array_61_7 <= _GEN_2741;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_62_0 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_0_1_REG) begin
      if (6'h3e == s1_way_waddr_0_1_r) begin
        meta_array_62_0 <= s1_way_wdata_0_1_r;
      end else begin
        meta_array_62_0 <= _GEN_1832;
      end
    end else begin
      meta_array_62_0 <= _GEN_1832;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_62_1 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_1_1_REG) begin
      if (6'h3e == s1_way_waddr_1_1_r) begin
        meta_array_62_1 <= s1_way_wdata_1_1_r;
      end else begin
        meta_array_62_1 <= _GEN_1962;
      end
    end else begin
      meta_array_62_1 <= _GEN_1962;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_62_2 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_2_1_REG) begin
      if (6'h3e == s1_way_waddr_2_1_r) begin
        meta_array_62_2 <= s1_way_wdata_2_1_r;
      end else begin
        meta_array_62_2 <= _GEN_2092;
      end
    end else begin
      meta_array_62_2 <= _GEN_2092;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_62_3 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_3_1_REG) begin
      if (6'h3e == s1_way_waddr_3_1_r) begin
        meta_array_62_3 <= s1_way_wdata_3_1_r;
      end else begin
        meta_array_62_3 <= _GEN_2222;
      end
    end else begin
      meta_array_62_3 <= _GEN_2222;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_62_4 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_4_1_REG) begin
      if (6'h3e == s1_way_waddr_4_1_r) begin
        meta_array_62_4 <= s1_way_wdata_4_1_r;
      end else begin
        meta_array_62_4 <= _GEN_2352;
      end
    end else begin
      meta_array_62_4 <= _GEN_2352;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_62_5 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_5_1_REG) begin
      if (6'h3e == s1_way_waddr_5_1_r) begin
        meta_array_62_5 <= s1_way_wdata_5_1_r;
      end else begin
        meta_array_62_5 <= _GEN_2482;
      end
    end else begin
      meta_array_62_5 <= _GEN_2482;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_62_6 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_6_1_REG) begin
      if (6'h3e == s1_way_waddr_6_1_r) begin
        meta_array_62_6 <= s1_way_wdata_6_1_r;
      end else begin
        meta_array_62_6 <= _GEN_2612;
      end
    end else begin
      meta_array_62_6 <= _GEN_2612;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_62_7 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_7_1_REG) begin
      if (6'h3e == s1_way_waddr_7_1_r) begin
        meta_array_62_7 <= s1_way_wdata_7_1_r;
      end else begin
        meta_array_62_7 <= _GEN_2742;
      end
    end else begin
      meta_array_62_7 <= _GEN_2742;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_63_0 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_0_1_REG) begin
      if (6'h3f == s1_way_waddr_0_1_r) begin
        meta_array_63_0 <= s1_way_wdata_0_1_r;
      end else begin
        meta_array_63_0 <= _GEN_1833;
      end
    end else begin
      meta_array_63_0 <= _GEN_1833;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_63_1 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_1_1_REG) begin
      if (6'h3f == s1_way_waddr_1_1_r) begin
        meta_array_63_1 <= s1_way_wdata_1_1_r;
      end else begin
        meta_array_63_1 <= _GEN_1963;
      end
    end else begin
      meta_array_63_1 <= _GEN_1963;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_63_2 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_2_1_REG) begin
      if (6'h3f == s1_way_waddr_2_1_r) begin
        meta_array_63_2 <= s1_way_wdata_2_1_r;
      end else begin
        meta_array_63_2 <= _GEN_2093;
      end
    end else begin
      meta_array_63_2 <= _GEN_2093;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_63_3 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_3_1_REG) begin
      if (6'h3f == s1_way_waddr_3_1_r) begin
        meta_array_63_3 <= s1_way_wdata_3_1_r;
      end else begin
        meta_array_63_3 <= _GEN_2223;
      end
    end else begin
      meta_array_63_3 <= _GEN_2223;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_63_4 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_4_1_REG) begin
      if (6'h3f == s1_way_waddr_4_1_r) begin
        meta_array_63_4 <= s1_way_wdata_4_1_r;
      end else begin
        meta_array_63_4 <= _GEN_2353;
      end
    end else begin
      meta_array_63_4 <= _GEN_2353;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_63_5 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_5_1_REG) begin
      if (6'h3f == s1_way_waddr_5_1_r) begin
        meta_array_63_5 <= s1_way_wdata_5_1_r;
      end else begin
        meta_array_63_5 <= _GEN_2483;
      end
    end else begin
      meta_array_63_5 <= _GEN_2483;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_63_6 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_6_1_REG) begin
      if (6'h3f == s1_way_waddr_6_1_r) begin
        meta_array_63_6 <= s1_way_wdata_6_1_r;
      end else begin
        meta_array_63_6 <= _GEN_2613;
      end
    end else begin
      meta_array_63_6 <= _GEN_2613;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[AsynchronousMetaArray.scala 156:41]
      meta_array_63_7 <= 1'h0; // @[AsynchronousMetaArray.scala 157:{55,55}]
    end else if (s1_way_wen_7_1_REG) begin
      if (6'h3f == s1_way_waddr_7_1_r) begin
        meta_array_63_7 <= s1_way_wdata_7_1_r;
      end else begin
        meta_array_63_7 <= _GEN_2743;
      end
    end else begin
      meta_array_63_7 <= _GEN_2743;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  meta_array_0_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  meta_array_0_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  meta_array_0_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  meta_array_0_3 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  meta_array_0_4 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  meta_array_0_5 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  meta_array_0_6 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  meta_array_0_7 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  meta_array_1_0 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  meta_array_1_1 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  meta_array_1_2 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  meta_array_1_3 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  meta_array_1_4 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  meta_array_1_5 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  meta_array_1_6 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  meta_array_1_7 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  meta_array_2_0 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  meta_array_2_1 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  meta_array_2_2 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  meta_array_2_3 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  meta_array_2_4 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  meta_array_2_5 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  meta_array_2_6 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  meta_array_2_7 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  meta_array_3_0 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  meta_array_3_1 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  meta_array_3_2 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  meta_array_3_3 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  meta_array_3_4 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  meta_array_3_5 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  meta_array_3_6 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  meta_array_3_7 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  meta_array_4_0 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  meta_array_4_1 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  meta_array_4_2 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  meta_array_4_3 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  meta_array_4_4 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  meta_array_4_5 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  meta_array_4_6 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  meta_array_4_7 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  meta_array_5_0 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  meta_array_5_1 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  meta_array_5_2 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  meta_array_5_3 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  meta_array_5_4 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  meta_array_5_5 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  meta_array_5_6 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  meta_array_5_7 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  meta_array_6_0 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  meta_array_6_1 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  meta_array_6_2 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  meta_array_6_3 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  meta_array_6_4 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  meta_array_6_5 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  meta_array_6_6 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  meta_array_6_7 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  meta_array_7_0 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  meta_array_7_1 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  meta_array_7_2 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  meta_array_7_3 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  meta_array_7_4 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  meta_array_7_5 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  meta_array_7_6 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  meta_array_7_7 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  meta_array_8_0 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  meta_array_8_1 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  meta_array_8_2 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  meta_array_8_3 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  meta_array_8_4 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  meta_array_8_5 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  meta_array_8_6 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  meta_array_8_7 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  meta_array_9_0 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  meta_array_9_1 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  meta_array_9_2 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  meta_array_9_3 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  meta_array_9_4 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  meta_array_9_5 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  meta_array_9_6 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  meta_array_9_7 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  meta_array_10_0 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  meta_array_10_1 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  meta_array_10_2 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  meta_array_10_3 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  meta_array_10_4 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  meta_array_10_5 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  meta_array_10_6 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  meta_array_10_7 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  meta_array_11_0 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  meta_array_11_1 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  meta_array_11_2 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  meta_array_11_3 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  meta_array_11_4 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  meta_array_11_5 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  meta_array_11_6 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  meta_array_11_7 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  meta_array_12_0 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  meta_array_12_1 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  meta_array_12_2 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  meta_array_12_3 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  meta_array_12_4 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  meta_array_12_5 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  meta_array_12_6 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  meta_array_12_7 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  meta_array_13_0 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  meta_array_13_1 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  meta_array_13_2 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  meta_array_13_3 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  meta_array_13_4 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  meta_array_13_5 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  meta_array_13_6 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  meta_array_13_7 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  meta_array_14_0 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  meta_array_14_1 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  meta_array_14_2 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  meta_array_14_3 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  meta_array_14_4 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  meta_array_14_5 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  meta_array_14_6 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  meta_array_14_7 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  meta_array_15_0 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  meta_array_15_1 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  meta_array_15_2 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  meta_array_15_3 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  meta_array_15_4 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  meta_array_15_5 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  meta_array_15_6 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  meta_array_15_7 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  meta_array_16_0 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  meta_array_16_1 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  meta_array_16_2 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  meta_array_16_3 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  meta_array_16_4 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  meta_array_16_5 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  meta_array_16_6 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  meta_array_16_7 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  meta_array_17_0 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  meta_array_17_1 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  meta_array_17_2 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  meta_array_17_3 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  meta_array_17_4 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  meta_array_17_5 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  meta_array_17_6 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  meta_array_17_7 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  meta_array_18_0 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  meta_array_18_1 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  meta_array_18_2 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  meta_array_18_3 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  meta_array_18_4 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  meta_array_18_5 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  meta_array_18_6 = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  meta_array_18_7 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  meta_array_19_0 = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  meta_array_19_1 = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  meta_array_19_2 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  meta_array_19_3 = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  meta_array_19_4 = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  meta_array_19_5 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  meta_array_19_6 = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  meta_array_19_7 = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  meta_array_20_0 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  meta_array_20_1 = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  meta_array_20_2 = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  meta_array_20_3 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  meta_array_20_4 = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  meta_array_20_5 = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  meta_array_20_6 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  meta_array_20_7 = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  meta_array_21_0 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  meta_array_21_1 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  meta_array_21_2 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  meta_array_21_3 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  meta_array_21_4 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  meta_array_21_5 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  meta_array_21_6 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  meta_array_21_7 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  meta_array_22_0 = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  meta_array_22_1 = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  meta_array_22_2 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  meta_array_22_3 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  meta_array_22_4 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  meta_array_22_5 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  meta_array_22_6 = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  meta_array_22_7 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  meta_array_23_0 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  meta_array_23_1 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  meta_array_23_2 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  meta_array_23_3 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  meta_array_23_4 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  meta_array_23_5 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  meta_array_23_6 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  meta_array_23_7 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  meta_array_24_0 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  meta_array_24_1 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  meta_array_24_2 = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  meta_array_24_3 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  meta_array_24_4 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  meta_array_24_5 = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  meta_array_24_6 = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  meta_array_24_7 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  meta_array_25_0 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  meta_array_25_1 = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  meta_array_25_2 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  meta_array_25_3 = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  meta_array_25_4 = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  meta_array_25_5 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  meta_array_25_6 = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  meta_array_25_7 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  meta_array_26_0 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  meta_array_26_1 = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  meta_array_26_2 = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  meta_array_26_3 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  meta_array_26_4 = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  meta_array_26_5 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  meta_array_26_6 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  meta_array_26_7 = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  meta_array_27_0 = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  meta_array_27_1 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  meta_array_27_2 = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  meta_array_27_3 = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  meta_array_27_4 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  meta_array_27_5 = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  meta_array_27_6 = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  meta_array_27_7 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  meta_array_28_0 = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  meta_array_28_1 = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  meta_array_28_2 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  meta_array_28_3 = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  meta_array_28_4 = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  meta_array_28_5 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  meta_array_28_6 = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  meta_array_28_7 = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  meta_array_29_0 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  meta_array_29_1 = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  meta_array_29_2 = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  meta_array_29_3 = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  meta_array_29_4 = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  meta_array_29_5 = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  meta_array_29_6 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  meta_array_29_7 = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  meta_array_30_0 = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  meta_array_30_1 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  meta_array_30_2 = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  meta_array_30_3 = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  meta_array_30_4 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  meta_array_30_5 = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  meta_array_30_6 = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  meta_array_30_7 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  meta_array_31_0 = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  meta_array_31_1 = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  meta_array_31_2 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  meta_array_31_3 = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  meta_array_31_4 = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  meta_array_31_5 = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  meta_array_31_6 = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  meta_array_31_7 = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  meta_array_32_0 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  meta_array_32_1 = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  meta_array_32_2 = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  meta_array_32_3 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  meta_array_32_4 = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  meta_array_32_5 = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  meta_array_32_6 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  meta_array_32_7 = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  meta_array_33_0 = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  meta_array_33_1 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  meta_array_33_2 = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  meta_array_33_3 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  meta_array_33_4 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  meta_array_33_5 = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  meta_array_33_6 = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  meta_array_33_7 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  meta_array_34_0 = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  meta_array_34_1 = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  meta_array_34_2 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  meta_array_34_3 = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  meta_array_34_4 = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  meta_array_34_5 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  meta_array_34_6 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  meta_array_34_7 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  meta_array_35_0 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  meta_array_35_1 = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  meta_array_35_2 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  meta_array_35_3 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  meta_array_35_4 = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  meta_array_35_5 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  meta_array_35_6 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  meta_array_35_7 = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  meta_array_36_0 = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  meta_array_36_1 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  meta_array_36_2 = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  meta_array_36_3 = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  meta_array_36_4 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  meta_array_36_5 = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  meta_array_36_6 = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  meta_array_36_7 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  meta_array_37_0 = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  meta_array_37_1 = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  meta_array_37_2 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  meta_array_37_3 = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  meta_array_37_4 = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  meta_array_37_5 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  meta_array_37_6 = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  meta_array_37_7 = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  meta_array_38_0 = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  meta_array_38_1 = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  meta_array_38_2 = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  meta_array_38_3 = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  meta_array_38_4 = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  meta_array_38_5 = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  meta_array_38_6 = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  meta_array_38_7 = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  meta_array_39_0 = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  meta_array_39_1 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  meta_array_39_2 = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  meta_array_39_3 = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  meta_array_39_4 = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  meta_array_39_5 = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  meta_array_39_6 = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  meta_array_39_7 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  meta_array_40_0 = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  meta_array_40_1 = _RAND_321[0:0];
  _RAND_322 = {1{`RANDOM}};
  meta_array_40_2 = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  meta_array_40_3 = _RAND_323[0:0];
  _RAND_324 = {1{`RANDOM}};
  meta_array_40_4 = _RAND_324[0:0];
  _RAND_325 = {1{`RANDOM}};
  meta_array_40_5 = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  meta_array_40_6 = _RAND_326[0:0];
  _RAND_327 = {1{`RANDOM}};
  meta_array_40_7 = _RAND_327[0:0];
  _RAND_328 = {1{`RANDOM}};
  meta_array_41_0 = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  meta_array_41_1 = _RAND_329[0:0];
  _RAND_330 = {1{`RANDOM}};
  meta_array_41_2 = _RAND_330[0:0];
  _RAND_331 = {1{`RANDOM}};
  meta_array_41_3 = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  meta_array_41_4 = _RAND_332[0:0];
  _RAND_333 = {1{`RANDOM}};
  meta_array_41_5 = _RAND_333[0:0];
  _RAND_334 = {1{`RANDOM}};
  meta_array_41_6 = _RAND_334[0:0];
  _RAND_335 = {1{`RANDOM}};
  meta_array_41_7 = _RAND_335[0:0];
  _RAND_336 = {1{`RANDOM}};
  meta_array_42_0 = _RAND_336[0:0];
  _RAND_337 = {1{`RANDOM}};
  meta_array_42_1 = _RAND_337[0:0];
  _RAND_338 = {1{`RANDOM}};
  meta_array_42_2 = _RAND_338[0:0];
  _RAND_339 = {1{`RANDOM}};
  meta_array_42_3 = _RAND_339[0:0];
  _RAND_340 = {1{`RANDOM}};
  meta_array_42_4 = _RAND_340[0:0];
  _RAND_341 = {1{`RANDOM}};
  meta_array_42_5 = _RAND_341[0:0];
  _RAND_342 = {1{`RANDOM}};
  meta_array_42_6 = _RAND_342[0:0];
  _RAND_343 = {1{`RANDOM}};
  meta_array_42_7 = _RAND_343[0:0];
  _RAND_344 = {1{`RANDOM}};
  meta_array_43_0 = _RAND_344[0:0];
  _RAND_345 = {1{`RANDOM}};
  meta_array_43_1 = _RAND_345[0:0];
  _RAND_346 = {1{`RANDOM}};
  meta_array_43_2 = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  meta_array_43_3 = _RAND_347[0:0];
  _RAND_348 = {1{`RANDOM}};
  meta_array_43_4 = _RAND_348[0:0];
  _RAND_349 = {1{`RANDOM}};
  meta_array_43_5 = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  meta_array_43_6 = _RAND_350[0:0];
  _RAND_351 = {1{`RANDOM}};
  meta_array_43_7 = _RAND_351[0:0];
  _RAND_352 = {1{`RANDOM}};
  meta_array_44_0 = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  meta_array_44_1 = _RAND_353[0:0];
  _RAND_354 = {1{`RANDOM}};
  meta_array_44_2 = _RAND_354[0:0];
  _RAND_355 = {1{`RANDOM}};
  meta_array_44_3 = _RAND_355[0:0];
  _RAND_356 = {1{`RANDOM}};
  meta_array_44_4 = _RAND_356[0:0];
  _RAND_357 = {1{`RANDOM}};
  meta_array_44_5 = _RAND_357[0:0];
  _RAND_358 = {1{`RANDOM}};
  meta_array_44_6 = _RAND_358[0:0];
  _RAND_359 = {1{`RANDOM}};
  meta_array_44_7 = _RAND_359[0:0];
  _RAND_360 = {1{`RANDOM}};
  meta_array_45_0 = _RAND_360[0:0];
  _RAND_361 = {1{`RANDOM}};
  meta_array_45_1 = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  meta_array_45_2 = _RAND_362[0:0];
  _RAND_363 = {1{`RANDOM}};
  meta_array_45_3 = _RAND_363[0:0];
  _RAND_364 = {1{`RANDOM}};
  meta_array_45_4 = _RAND_364[0:0];
  _RAND_365 = {1{`RANDOM}};
  meta_array_45_5 = _RAND_365[0:0];
  _RAND_366 = {1{`RANDOM}};
  meta_array_45_6 = _RAND_366[0:0];
  _RAND_367 = {1{`RANDOM}};
  meta_array_45_7 = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  meta_array_46_0 = _RAND_368[0:0];
  _RAND_369 = {1{`RANDOM}};
  meta_array_46_1 = _RAND_369[0:0];
  _RAND_370 = {1{`RANDOM}};
  meta_array_46_2 = _RAND_370[0:0];
  _RAND_371 = {1{`RANDOM}};
  meta_array_46_3 = _RAND_371[0:0];
  _RAND_372 = {1{`RANDOM}};
  meta_array_46_4 = _RAND_372[0:0];
  _RAND_373 = {1{`RANDOM}};
  meta_array_46_5 = _RAND_373[0:0];
  _RAND_374 = {1{`RANDOM}};
  meta_array_46_6 = _RAND_374[0:0];
  _RAND_375 = {1{`RANDOM}};
  meta_array_46_7 = _RAND_375[0:0];
  _RAND_376 = {1{`RANDOM}};
  meta_array_47_0 = _RAND_376[0:0];
  _RAND_377 = {1{`RANDOM}};
  meta_array_47_1 = _RAND_377[0:0];
  _RAND_378 = {1{`RANDOM}};
  meta_array_47_2 = _RAND_378[0:0];
  _RAND_379 = {1{`RANDOM}};
  meta_array_47_3 = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  meta_array_47_4 = _RAND_380[0:0];
  _RAND_381 = {1{`RANDOM}};
  meta_array_47_5 = _RAND_381[0:0];
  _RAND_382 = {1{`RANDOM}};
  meta_array_47_6 = _RAND_382[0:0];
  _RAND_383 = {1{`RANDOM}};
  meta_array_47_7 = _RAND_383[0:0];
  _RAND_384 = {1{`RANDOM}};
  meta_array_48_0 = _RAND_384[0:0];
  _RAND_385 = {1{`RANDOM}};
  meta_array_48_1 = _RAND_385[0:0];
  _RAND_386 = {1{`RANDOM}};
  meta_array_48_2 = _RAND_386[0:0];
  _RAND_387 = {1{`RANDOM}};
  meta_array_48_3 = _RAND_387[0:0];
  _RAND_388 = {1{`RANDOM}};
  meta_array_48_4 = _RAND_388[0:0];
  _RAND_389 = {1{`RANDOM}};
  meta_array_48_5 = _RAND_389[0:0];
  _RAND_390 = {1{`RANDOM}};
  meta_array_48_6 = _RAND_390[0:0];
  _RAND_391 = {1{`RANDOM}};
  meta_array_48_7 = _RAND_391[0:0];
  _RAND_392 = {1{`RANDOM}};
  meta_array_49_0 = _RAND_392[0:0];
  _RAND_393 = {1{`RANDOM}};
  meta_array_49_1 = _RAND_393[0:0];
  _RAND_394 = {1{`RANDOM}};
  meta_array_49_2 = _RAND_394[0:0];
  _RAND_395 = {1{`RANDOM}};
  meta_array_49_3 = _RAND_395[0:0];
  _RAND_396 = {1{`RANDOM}};
  meta_array_49_4 = _RAND_396[0:0];
  _RAND_397 = {1{`RANDOM}};
  meta_array_49_5 = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  meta_array_49_6 = _RAND_398[0:0];
  _RAND_399 = {1{`RANDOM}};
  meta_array_49_7 = _RAND_399[0:0];
  _RAND_400 = {1{`RANDOM}};
  meta_array_50_0 = _RAND_400[0:0];
  _RAND_401 = {1{`RANDOM}};
  meta_array_50_1 = _RAND_401[0:0];
  _RAND_402 = {1{`RANDOM}};
  meta_array_50_2 = _RAND_402[0:0];
  _RAND_403 = {1{`RANDOM}};
  meta_array_50_3 = _RAND_403[0:0];
  _RAND_404 = {1{`RANDOM}};
  meta_array_50_4 = _RAND_404[0:0];
  _RAND_405 = {1{`RANDOM}};
  meta_array_50_5 = _RAND_405[0:0];
  _RAND_406 = {1{`RANDOM}};
  meta_array_50_6 = _RAND_406[0:0];
  _RAND_407 = {1{`RANDOM}};
  meta_array_50_7 = _RAND_407[0:0];
  _RAND_408 = {1{`RANDOM}};
  meta_array_51_0 = _RAND_408[0:0];
  _RAND_409 = {1{`RANDOM}};
  meta_array_51_1 = _RAND_409[0:0];
  _RAND_410 = {1{`RANDOM}};
  meta_array_51_2 = _RAND_410[0:0];
  _RAND_411 = {1{`RANDOM}};
  meta_array_51_3 = _RAND_411[0:0];
  _RAND_412 = {1{`RANDOM}};
  meta_array_51_4 = _RAND_412[0:0];
  _RAND_413 = {1{`RANDOM}};
  meta_array_51_5 = _RAND_413[0:0];
  _RAND_414 = {1{`RANDOM}};
  meta_array_51_6 = _RAND_414[0:0];
  _RAND_415 = {1{`RANDOM}};
  meta_array_51_7 = _RAND_415[0:0];
  _RAND_416 = {1{`RANDOM}};
  meta_array_52_0 = _RAND_416[0:0];
  _RAND_417 = {1{`RANDOM}};
  meta_array_52_1 = _RAND_417[0:0];
  _RAND_418 = {1{`RANDOM}};
  meta_array_52_2 = _RAND_418[0:0];
  _RAND_419 = {1{`RANDOM}};
  meta_array_52_3 = _RAND_419[0:0];
  _RAND_420 = {1{`RANDOM}};
  meta_array_52_4 = _RAND_420[0:0];
  _RAND_421 = {1{`RANDOM}};
  meta_array_52_5 = _RAND_421[0:0];
  _RAND_422 = {1{`RANDOM}};
  meta_array_52_6 = _RAND_422[0:0];
  _RAND_423 = {1{`RANDOM}};
  meta_array_52_7 = _RAND_423[0:0];
  _RAND_424 = {1{`RANDOM}};
  meta_array_53_0 = _RAND_424[0:0];
  _RAND_425 = {1{`RANDOM}};
  meta_array_53_1 = _RAND_425[0:0];
  _RAND_426 = {1{`RANDOM}};
  meta_array_53_2 = _RAND_426[0:0];
  _RAND_427 = {1{`RANDOM}};
  meta_array_53_3 = _RAND_427[0:0];
  _RAND_428 = {1{`RANDOM}};
  meta_array_53_4 = _RAND_428[0:0];
  _RAND_429 = {1{`RANDOM}};
  meta_array_53_5 = _RAND_429[0:0];
  _RAND_430 = {1{`RANDOM}};
  meta_array_53_6 = _RAND_430[0:0];
  _RAND_431 = {1{`RANDOM}};
  meta_array_53_7 = _RAND_431[0:0];
  _RAND_432 = {1{`RANDOM}};
  meta_array_54_0 = _RAND_432[0:0];
  _RAND_433 = {1{`RANDOM}};
  meta_array_54_1 = _RAND_433[0:0];
  _RAND_434 = {1{`RANDOM}};
  meta_array_54_2 = _RAND_434[0:0];
  _RAND_435 = {1{`RANDOM}};
  meta_array_54_3 = _RAND_435[0:0];
  _RAND_436 = {1{`RANDOM}};
  meta_array_54_4 = _RAND_436[0:0];
  _RAND_437 = {1{`RANDOM}};
  meta_array_54_5 = _RAND_437[0:0];
  _RAND_438 = {1{`RANDOM}};
  meta_array_54_6 = _RAND_438[0:0];
  _RAND_439 = {1{`RANDOM}};
  meta_array_54_7 = _RAND_439[0:0];
  _RAND_440 = {1{`RANDOM}};
  meta_array_55_0 = _RAND_440[0:0];
  _RAND_441 = {1{`RANDOM}};
  meta_array_55_1 = _RAND_441[0:0];
  _RAND_442 = {1{`RANDOM}};
  meta_array_55_2 = _RAND_442[0:0];
  _RAND_443 = {1{`RANDOM}};
  meta_array_55_3 = _RAND_443[0:0];
  _RAND_444 = {1{`RANDOM}};
  meta_array_55_4 = _RAND_444[0:0];
  _RAND_445 = {1{`RANDOM}};
  meta_array_55_5 = _RAND_445[0:0];
  _RAND_446 = {1{`RANDOM}};
  meta_array_55_6 = _RAND_446[0:0];
  _RAND_447 = {1{`RANDOM}};
  meta_array_55_7 = _RAND_447[0:0];
  _RAND_448 = {1{`RANDOM}};
  meta_array_56_0 = _RAND_448[0:0];
  _RAND_449 = {1{`RANDOM}};
  meta_array_56_1 = _RAND_449[0:0];
  _RAND_450 = {1{`RANDOM}};
  meta_array_56_2 = _RAND_450[0:0];
  _RAND_451 = {1{`RANDOM}};
  meta_array_56_3 = _RAND_451[0:0];
  _RAND_452 = {1{`RANDOM}};
  meta_array_56_4 = _RAND_452[0:0];
  _RAND_453 = {1{`RANDOM}};
  meta_array_56_5 = _RAND_453[0:0];
  _RAND_454 = {1{`RANDOM}};
  meta_array_56_6 = _RAND_454[0:0];
  _RAND_455 = {1{`RANDOM}};
  meta_array_56_7 = _RAND_455[0:0];
  _RAND_456 = {1{`RANDOM}};
  meta_array_57_0 = _RAND_456[0:0];
  _RAND_457 = {1{`RANDOM}};
  meta_array_57_1 = _RAND_457[0:0];
  _RAND_458 = {1{`RANDOM}};
  meta_array_57_2 = _RAND_458[0:0];
  _RAND_459 = {1{`RANDOM}};
  meta_array_57_3 = _RAND_459[0:0];
  _RAND_460 = {1{`RANDOM}};
  meta_array_57_4 = _RAND_460[0:0];
  _RAND_461 = {1{`RANDOM}};
  meta_array_57_5 = _RAND_461[0:0];
  _RAND_462 = {1{`RANDOM}};
  meta_array_57_6 = _RAND_462[0:0];
  _RAND_463 = {1{`RANDOM}};
  meta_array_57_7 = _RAND_463[0:0];
  _RAND_464 = {1{`RANDOM}};
  meta_array_58_0 = _RAND_464[0:0];
  _RAND_465 = {1{`RANDOM}};
  meta_array_58_1 = _RAND_465[0:0];
  _RAND_466 = {1{`RANDOM}};
  meta_array_58_2 = _RAND_466[0:0];
  _RAND_467 = {1{`RANDOM}};
  meta_array_58_3 = _RAND_467[0:0];
  _RAND_468 = {1{`RANDOM}};
  meta_array_58_4 = _RAND_468[0:0];
  _RAND_469 = {1{`RANDOM}};
  meta_array_58_5 = _RAND_469[0:0];
  _RAND_470 = {1{`RANDOM}};
  meta_array_58_6 = _RAND_470[0:0];
  _RAND_471 = {1{`RANDOM}};
  meta_array_58_7 = _RAND_471[0:0];
  _RAND_472 = {1{`RANDOM}};
  meta_array_59_0 = _RAND_472[0:0];
  _RAND_473 = {1{`RANDOM}};
  meta_array_59_1 = _RAND_473[0:0];
  _RAND_474 = {1{`RANDOM}};
  meta_array_59_2 = _RAND_474[0:0];
  _RAND_475 = {1{`RANDOM}};
  meta_array_59_3 = _RAND_475[0:0];
  _RAND_476 = {1{`RANDOM}};
  meta_array_59_4 = _RAND_476[0:0];
  _RAND_477 = {1{`RANDOM}};
  meta_array_59_5 = _RAND_477[0:0];
  _RAND_478 = {1{`RANDOM}};
  meta_array_59_6 = _RAND_478[0:0];
  _RAND_479 = {1{`RANDOM}};
  meta_array_59_7 = _RAND_479[0:0];
  _RAND_480 = {1{`RANDOM}};
  meta_array_60_0 = _RAND_480[0:0];
  _RAND_481 = {1{`RANDOM}};
  meta_array_60_1 = _RAND_481[0:0];
  _RAND_482 = {1{`RANDOM}};
  meta_array_60_2 = _RAND_482[0:0];
  _RAND_483 = {1{`RANDOM}};
  meta_array_60_3 = _RAND_483[0:0];
  _RAND_484 = {1{`RANDOM}};
  meta_array_60_4 = _RAND_484[0:0];
  _RAND_485 = {1{`RANDOM}};
  meta_array_60_5 = _RAND_485[0:0];
  _RAND_486 = {1{`RANDOM}};
  meta_array_60_6 = _RAND_486[0:0];
  _RAND_487 = {1{`RANDOM}};
  meta_array_60_7 = _RAND_487[0:0];
  _RAND_488 = {1{`RANDOM}};
  meta_array_61_0 = _RAND_488[0:0];
  _RAND_489 = {1{`RANDOM}};
  meta_array_61_1 = _RAND_489[0:0];
  _RAND_490 = {1{`RANDOM}};
  meta_array_61_2 = _RAND_490[0:0];
  _RAND_491 = {1{`RANDOM}};
  meta_array_61_3 = _RAND_491[0:0];
  _RAND_492 = {1{`RANDOM}};
  meta_array_61_4 = _RAND_492[0:0];
  _RAND_493 = {1{`RANDOM}};
  meta_array_61_5 = _RAND_493[0:0];
  _RAND_494 = {1{`RANDOM}};
  meta_array_61_6 = _RAND_494[0:0];
  _RAND_495 = {1{`RANDOM}};
  meta_array_61_7 = _RAND_495[0:0];
  _RAND_496 = {1{`RANDOM}};
  meta_array_62_0 = _RAND_496[0:0];
  _RAND_497 = {1{`RANDOM}};
  meta_array_62_1 = _RAND_497[0:0];
  _RAND_498 = {1{`RANDOM}};
  meta_array_62_2 = _RAND_498[0:0];
  _RAND_499 = {1{`RANDOM}};
  meta_array_62_3 = _RAND_499[0:0];
  _RAND_500 = {1{`RANDOM}};
  meta_array_62_4 = _RAND_500[0:0];
  _RAND_501 = {1{`RANDOM}};
  meta_array_62_5 = _RAND_501[0:0];
  _RAND_502 = {1{`RANDOM}};
  meta_array_62_6 = _RAND_502[0:0];
  _RAND_503 = {1{`RANDOM}};
  meta_array_62_7 = _RAND_503[0:0];
  _RAND_504 = {1{`RANDOM}};
  meta_array_63_0 = _RAND_504[0:0];
  _RAND_505 = {1{`RANDOM}};
  meta_array_63_1 = _RAND_505[0:0];
  _RAND_506 = {1{`RANDOM}};
  meta_array_63_2 = _RAND_506[0:0];
  _RAND_507 = {1{`RANDOM}};
  meta_array_63_3 = _RAND_507[0:0];
  _RAND_508 = {1{`RANDOM}};
  meta_array_63_4 = _RAND_508[0:0];
  _RAND_509 = {1{`RANDOM}};
  meta_array_63_5 = _RAND_509[0:0];
  _RAND_510 = {1{`RANDOM}};
  meta_array_63_6 = _RAND_510[0:0];
  _RAND_511 = {1{`RANDOM}};
  meta_array_63_7 = _RAND_511[0:0];
  _RAND_512 = {1{`RANDOM}};
  s1_way_waddr_0_0_r = _RAND_512[5:0];
  _RAND_513 = {1{`RANDOM}};
  s1_way_wen_0_0_REG = _RAND_513[0:0];
  _RAND_514 = {1{`RANDOM}};
  s1_way_wdata_0_0_r = _RAND_514[0:0];
  _RAND_515 = {1{`RANDOM}};
  s1_way_waddr_0_1_r = _RAND_515[5:0];
  _RAND_516 = {1{`RANDOM}};
  s1_way_wen_0_1_REG = _RAND_516[0:0];
  _RAND_517 = {1{`RANDOM}};
  s1_way_wdata_0_1_r = _RAND_517[0:0];
  _RAND_518 = {1{`RANDOM}};
  io_resp_0_0_r = _RAND_518[0:0];
  _RAND_519 = {1{`RANDOM}};
  io_resp_0_0_r1 = _RAND_519[0:0];
  _RAND_520 = {1{`RANDOM}};
  io_resp_0_0_r2 = _RAND_520[5:0];
  _RAND_521 = {1{`RANDOM}};
  s1_way_waddr_1_0_r = _RAND_521[5:0];
  _RAND_522 = {1{`RANDOM}};
  s1_way_wen_1_0_REG = _RAND_522[0:0];
  _RAND_523 = {1{`RANDOM}};
  s1_way_wdata_1_0_r = _RAND_523[0:0];
  _RAND_524 = {1{`RANDOM}};
  s1_way_waddr_1_1_r = _RAND_524[5:0];
  _RAND_525 = {1{`RANDOM}};
  s1_way_wen_1_1_REG = _RAND_525[0:0];
  _RAND_526 = {1{`RANDOM}};
  s1_way_wdata_1_1_r = _RAND_526[0:0];
  _RAND_527 = {1{`RANDOM}};
  io_resp_0_1_r = _RAND_527[0:0];
  _RAND_528 = {1{`RANDOM}};
  io_resp_0_1_r1 = _RAND_528[0:0];
  _RAND_529 = {1{`RANDOM}};
  io_resp_0_1_r2 = _RAND_529[5:0];
  _RAND_530 = {1{`RANDOM}};
  s1_way_waddr_2_0_r = _RAND_530[5:0];
  _RAND_531 = {1{`RANDOM}};
  s1_way_wen_2_0_REG = _RAND_531[0:0];
  _RAND_532 = {1{`RANDOM}};
  s1_way_wdata_2_0_r = _RAND_532[0:0];
  _RAND_533 = {1{`RANDOM}};
  s1_way_waddr_2_1_r = _RAND_533[5:0];
  _RAND_534 = {1{`RANDOM}};
  s1_way_wen_2_1_REG = _RAND_534[0:0];
  _RAND_535 = {1{`RANDOM}};
  s1_way_wdata_2_1_r = _RAND_535[0:0];
  _RAND_536 = {1{`RANDOM}};
  io_resp_0_2_r = _RAND_536[0:0];
  _RAND_537 = {1{`RANDOM}};
  io_resp_0_2_r1 = _RAND_537[0:0];
  _RAND_538 = {1{`RANDOM}};
  io_resp_0_2_r2 = _RAND_538[5:0];
  _RAND_539 = {1{`RANDOM}};
  s1_way_waddr_3_0_r = _RAND_539[5:0];
  _RAND_540 = {1{`RANDOM}};
  s1_way_wen_3_0_REG = _RAND_540[0:0];
  _RAND_541 = {1{`RANDOM}};
  s1_way_wdata_3_0_r = _RAND_541[0:0];
  _RAND_542 = {1{`RANDOM}};
  s1_way_waddr_3_1_r = _RAND_542[5:0];
  _RAND_543 = {1{`RANDOM}};
  s1_way_wen_3_1_REG = _RAND_543[0:0];
  _RAND_544 = {1{`RANDOM}};
  s1_way_wdata_3_1_r = _RAND_544[0:0];
  _RAND_545 = {1{`RANDOM}};
  io_resp_0_3_r = _RAND_545[0:0];
  _RAND_546 = {1{`RANDOM}};
  io_resp_0_3_r1 = _RAND_546[0:0];
  _RAND_547 = {1{`RANDOM}};
  io_resp_0_3_r2 = _RAND_547[5:0];
  _RAND_548 = {1{`RANDOM}};
  s1_way_waddr_4_0_r = _RAND_548[5:0];
  _RAND_549 = {1{`RANDOM}};
  s1_way_wen_4_0_REG = _RAND_549[0:0];
  _RAND_550 = {1{`RANDOM}};
  s1_way_wdata_4_0_r = _RAND_550[0:0];
  _RAND_551 = {1{`RANDOM}};
  s1_way_waddr_4_1_r = _RAND_551[5:0];
  _RAND_552 = {1{`RANDOM}};
  s1_way_wen_4_1_REG = _RAND_552[0:0];
  _RAND_553 = {1{`RANDOM}};
  s1_way_wdata_4_1_r = _RAND_553[0:0];
  _RAND_554 = {1{`RANDOM}};
  io_resp_0_4_r = _RAND_554[0:0];
  _RAND_555 = {1{`RANDOM}};
  io_resp_0_4_r1 = _RAND_555[0:0];
  _RAND_556 = {1{`RANDOM}};
  io_resp_0_4_r2 = _RAND_556[5:0];
  _RAND_557 = {1{`RANDOM}};
  s1_way_waddr_5_0_r = _RAND_557[5:0];
  _RAND_558 = {1{`RANDOM}};
  s1_way_wen_5_0_REG = _RAND_558[0:0];
  _RAND_559 = {1{`RANDOM}};
  s1_way_wdata_5_0_r = _RAND_559[0:0];
  _RAND_560 = {1{`RANDOM}};
  s1_way_waddr_5_1_r = _RAND_560[5:0];
  _RAND_561 = {1{`RANDOM}};
  s1_way_wen_5_1_REG = _RAND_561[0:0];
  _RAND_562 = {1{`RANDOM}};
  s1_way_wdata_5_1_r = _RAND_562[0:0];
  _RAND_563 = {1{`RANDOM}};
  io_resp_0_5_r = _RAND_563[0:0];
  _RAND_564 = {1{`RANDOM}};
  io_resp_0_5_r1 = _RAND_564[0:0];
  _RAND_565 = {1{`RANDOM}};
  io_resp_0_5_r2 = _RAND_565[5:0];
  _RAND_566 = {1{`RANDOM}};
  s1_way_waddr_6_0_r = _RAND_566[5:0];
  _RAND_567 = {1{`RANDOM}};
  s1_way_wen_6_0_REG = _RAND_567[0:0];
  _RAND_568 = {1{`RANDOM}};
  s1_way_wdata_6_0_r = _RAND_568[0:0];
  _RAND_569 = {1{`RANDOM}};
  s1_way_waddr_6_1_r = _RAND_569[5:0];
  _RAND_570 = {1{`RANDOM}};
  s1_way_wen_6_1_REG = _RAND_570[0:0];
  _RAND_571 = {1{`RANDOM}};
  s1_way_wdata_6_1_r = _RAND_571[0:0];
  _RAND_572 = {1{`RANDOM}};
  io_resp_0_6_r = _RAND_572[0:0];
  _RAND_573 = {1{`RANDOM}};
  io_resp_0_6_r1 = _RAND_573[0:0];
  _RAND_574 = {1{`RANDOM}};
  io_resp_0_6_r2 = _RAND_574[5:0];
  _RAND_575 = {1{`RANDOM}};
  s1_way_waddr_7_0_r = _RAND_575[5:0];
  _RAND_576 = {1{`RANDOM}};
  s1_way_wen_7_0_REG = _RAND_576[0:0];
  _RAND_577 = {1{`RANDOM}};
  s1_way_wdata_7_0_r = _RAND_577[0:0];
  _RAND_578 = {1{`RANDOM}};
  s1_way_waddr_7_1_r = _RAND_578[5:0];
  _RAND_579 = {1{`RANDOM}};
  s1_way_wen_7_1_REG = _RAND_579[0:0];
  _RAND_580 = {1{`RANDOM}};
  s1_way_wdata_7_1_r = _RAND_580[0:0];
  _RAND_581 = {1{`RANDOM}};
  io_resp_0_7_r = _RAND_581[0:0];
  _RAND_582 = {1{`RANDOM}};
  io_resp_0_7_r1 = _RAND_582[0:0];
  _RAND_583 = {1{`RANDOM}};
  io_resp_0_7_r2 = _RAND_583[5:0];
  _RAND_584 = {1{`RANDOM}};
  io_resp_1_0_r = _RAND_584[0:0];
  _RAND_585 = {1{`RANDOM}};
  io_resp_1_0_r1 = _RAND_585[0:0];
  _RAND_586 = {1{`RANDOM}};
  io_resp_1_0_r2 = _RAND_586[5:0];
  _RAND_587 = {1{`RANDOM}};
  io_resp_1_1_r = _RAND_587[0:0];
  _RAND_588 = {1{`RANDOM}};
  io_resp_1_1_r1 = _RAND_588[0:0];
  _RAND_589 = {1{`RANDOM}};
  io_resp_1_1_r2 = _RAND_589[5:0];
  _RAND_590 = {1{`RANDOM}};
  io_resp_1_2_r = _RAND_590[0:0];
  _RAND_591 = {1{`RANDOM}};
  io_resp_1_2_r1 = _RAND_591[0:0];
  _RAND_592 = {1{`RANDOM}};
  io_resp_1_2_r2 = _RAND_592[5:0];
  _RAND_593 = {1{`RANDOM}};
  io_resp_1_3_r = _RAND_593[0:0];
  _RAND_594 = {1{`RANDOM}};
  io_resp_1_3_r1 = _RAND_594[0:0];
  _RAND_595 = {1{`RANDOM}};
  io_resp_1_3_r2 = _RAND_595[5:0];
  _RAND_596 = {1{`RANDOM}};
  io_resp_1_4_r = _RAND_596[0:0];
  _RAND_597 = {1{`RANDOM}};
  io_resp_1_4_r1 = _RAND_597[0:0];
  _RAND_598 = {1{`RANDOM}};
  io_resp_1_4_r2 = _RAND_598[5:0];
  _RAND_599 = {1{`RANDOM}};
  io_resp_1_5_r = _RAND_599[0:0];
  _RAND_600 = {1{`RANDOM}};
  io_resp_1_5_r1 = _RAND_600[0:0];
  _RAND_601 = {1{`RANDOM}};
  io_resp_1_5_r2 = _RAND_601[5:0];
  _RAND_602 = {1{`RANDOM}};
  io_resp_1_6_r = _RAND_602[0:0];
  _RAND_603 = {1{`RANDOM}};
  io_resp_1_6_r1 = _RAND_603[0:0];
  _RAND_604 = {1{`RANDOM}};
  io_resp_1_6_r2 = _RAND_604[5:0];
  _RAND_605 = {1{`RANDOM}};
  io_resp_1_7_r = _RAND_605[0:0];
  _RAND_606 = {1{`RANDOM}};
  io_resp_1_7_r1 = _RAND_606[0:0];
  _RAND_607 = {1{`RANDOM}};
  io_resp_1_7_r2 = _RAND_607[5:0];
  _RAND_608 = {1{`RANDOM}};
  io_resp_2_0_r = _RAND_608[0:0];
  _RAND_609 = {1{`RANDOM}};
  io_resp_2_0_r1 = _RAND_609[0:0];
  _RAND_610 = {1{`RANDOM}};
  io_resp_2_0_r2 = _RAND_610[5:0];
  _RAND_611 = {1{`RANDOM}};
  io_resp_2_1_r = _RAND_611[0:0];
  _RAND_612 = {1{`RANDOM}};
  io_resp_2_1_r1 = _RAND_612[0:0];
  _RAND_613 = {1{`RANDOM}};
  io_resp_2_1_r2 = _RAND_613[5:0];
  _RAND_614 = {1{`RANDOM}};
  io_resp_2_2_r = _RAND_614[0:0];
  _RAND_615 = {1{`RANDOM}};
  io_resp_2_2_r1 = _RAND_615[0:0];
  _RAND_616 = {1{`RANDOM}};
  io_resp_2_2_r2 = _RAND_616[5:0];
  _RAND_617 = {1{`RANDOM}};
  io_resp_2_3_r = _RAND_617[0:0];
  _RAND_618 = {1{`RANDOM}};
  io_resp_2_3_r1 = _RAND_618[0:0];
  _RAND_619 = {1{`RANDOM}};
  io_resp_2_3_r2 = _RAND_619[5:0];
  _RAND_620 = {1{`RANDOM}};
  io_resp_2_4_r = _RAND_620[0:0];
  _RAND_621 = {1{`RANDOM}};
  io_resp_2_4_r1 = _RAND_621[0:0];
  _RAND_622 = {1{`RANDOM}};
  io_resp_2_4_r2 = _RAND_622[5:0];
  _RAND_623 = {1{`RANDOM}};
  io_resp_2_5_r = _RAND_623[0:0];
  _RAND_624 = {1{`RANDOM}};
  io_resp_2_5_r1 = _RAND_624[0:0];
  _RAND_625 = {1{`RANDOM}};
  io_resp_2_5_r2 = _RAND_625[5:0];
  _RAND_626 = {1{`RANDOM}};
  io_resp_2_6_r = _RAND_626[0:0];
  _RAND_627 = {1{`RANDOM}};
  io_resp_2_6_r1 = _RAND_627[0:0];
  _RAND_628 = {1{`RANDOM}};
  io_resp_2_6_r2 = _RAND_628[5:0];
  _RAND_629 = {1{`RANDOM}};
  io_resp_2_7_r = _RAND_629[0:0];
  _RAND_630 = {1{`RANDOM}};
  io_resp_2_7_r1 = _RAND_630[0:0];
  _RAND_631 = {1{`RANDOM}};
  io_resp_2_7_r2 = _RAND_631[5:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    meta_array_0_0 = 1'h0;
  end
  if (reset) begin
    meta_array_0_1 = 1'h0;
  end
  if (reset) begin
    meta_array_0_2 = 1'h0;
  end
  if (reset) begin
    meta_array_0_3 = 1'h0;
  end
  if (reset) begin
    meta_array_0_4 = 1'h0;
  end
  if (reset) begin
    meta_array_0_5 = 1'h0;
  end
  if (reset) begin
    meta_array_0_6 = 1'h0;
  end
  if (reset) begin
    meta_array_0_7 = 1'h0;
  end
  if (reset) begin
    meta_array_1_0 = 1'h0;
  end
  if (reset) begin
    meta_array_1_1 = 1'h0;
  end
  if (reset) begin
    meta_array_1_2 = 1'h0;
  end
  if (reset) begin
    meta_array_1_3 = 1'h0;
  end
  if (reset) begin
    meta_array_1_4 = 1'h0;
  end
  if (reset) begin
    meta_array_1_5 = 1'h0;
  end
  if (reset) begin
    meta_array_1_6 = 1'h0;
  end
  if (reset) begin
    meta_array_1_7 = 1'h0;
  end
  if (reset) begin
    meta_array_2_0 = 1'h0;
  end
  if (reset) begin
    meta_array_2_1 = 1'h0;
  end
  if (reset) begin
    meta_array_2_2 = 1'h0;
  end
  if (reset) begin
    meta_array_2_3 = 1'h0;
  end
  if (reset) begin
    meta_array_2_4 = 1'h0;
  end
  if (reset) begin
    meta_array_2_5 = 1'h0;
  end
  if (reset) begin
    meta_array_2_6 = 1'h0;
  end
  if (reset) begin
    meta_array_2_7 = 1'h0;
  end
  if (reset) begin
    meta_array_3_0 = 1'h0;
  end
  if (reset) begin
    meta_array_3_1 = 1'h0;
  end
  if (reset) begin
    meta_array_3_2 = 1'h0;
  end
  if (reset) begin
    meta_array_3_3 = 1'h0;
  end
  if (reset) begin
    meta_array_3_4 = 1'h0;
  end
  if (reset) begin
    meta_array_3_5 = 1'h0;
  end
  if (reset) begin
    meta_array_3_6 = 1'h0;
  end
  if (reset) begin
    meta_array_3_7 = 1'h0;
  end
  if (reset) begin
    meta_array_4_0 = 1'h0;
  end
  if (reset) begin
    meta_array_4_1 = 1'h0;
  end
  if (reset) begin
    meta_array_4_2 = 1'h0;
  end
  if (reset) begin
    meta_array_4_3 = 1'h0;
  end
  if (reset) begin
    meta_array_4_4 = 1'h0;
  end
  if (reset) begin
    meta_array_4_5 = 1'h0;
  end
  if (reset) begin
    meta_array_4_6 = 1'h0;
  end
  if (reset) begin
    meta_array_4_7 = 1'h0;
  end
  if (reset) begin
    meta_array_5_0 = 1'h0;
  end
  if (reset) begin
    meta_array_5_1 = 1'h0;
  end
  if (reset) begin
    meta_array_5_2 = 1'h0;
  end
  if (reset) begin
    meta_array_5_3 = 1'h0;
  end
  if (reset) begin
    meta_array_5_4 = 1'h0;
  end
  if (reset) begin
    meta_array_5_5 = 1'h0;
  end
  if (reset) begin
    meta_array_5_6 = 1'h0;
  end
  if (reset) begin
    meta_array_5_7 = 1'h0;
  end
  if (reset) begin
    meta_array_6_0 = 1'h0;
  end
  if (reset) begin
    meta_array_6_1 = 1'h0;
  end
  if (reset) begin
    meta_array_6_2 = 1'h0;
  end
  if (reset) begin
    meta_array_6_3 = 1'h0;
  end
  if (reset) begin
    meta_array_6_4 = 1'h0;
  end
  if (reset) begin
    meta_array_6_5 = 1'h0;
  end
  if (reset) begin
    meta_array_6_6 = 1'h0;
  end
  if (reset) begin
    meta_array_6_7 = 1'h0;
  end
  if (reset) begin
    meta_array_7_0 = 1'h0;
  end
  if (reset) begin
    meta_array_7_1 = 1'h0;
  end
  if (reset) begin
    meta_array_7_2 = 1'h0;
  end
  if (reset) begin
    meta_array_7_3 = 1'h0;
  end
  if (reset) begin
    meta_array_7_4 = 1'h0;
  end
  if (reset) begin
    meta_array_7_5 = 1'h0;
  end
  if (reset) begin
    meta_array_7_6 = 1'h0;
  end
  if (reset) begin
    meta_array_7_7 = 1'h0;
  end
  if (reset) begin
    meta_array_8_0 = 1'h0;
  end
  if (reset) begin
    meta_array_8_1 = 1'h0;
  end
  if (reset) begin
    meta_array_8_2 = 1'h0;
  end
  if (reset) begin
    meta_array_8_3 = 1'h0;
  end
  if (reset) begin
    meta_array_8_4 = 1'h0;
  end
  if (reset) begin
    meta_array_8_5 = 1'h0;
  end
  if (reset) begin
    meta_array_8_6 = 1'h0;
  end
  if (reset) begin
    meta_array_8_7 = 1'h0;
  end
  if (reset) begin
    meta_array_9_0 = 1'h0;
  end
  if (reset) begin
    meta_array_9_1 = 1'h0;
  end
  if (reset) begin
    meta_array_9_2 = 1'h0;
  end
  if (reset) begin
    meta_array_9_3 = 1'h0;
  end
  if (reset) begin
    meta_array_9_4 = 1'h0;
  end
  if (reset) begin
    meta_array_9_5 = 1'h0;
  end
  if (reset) begin
    meta_array_9_6 = 1'h0;
  end
  if (reset) begin
    meta_array_9_7 = 1'h0;
  end
  if (reset) begin
    meta_array_10_0 = 1'h0;
  end
  if (reset) begin
    meta_array_10_1 = 1'h0;
  end
  if (reset) begin
    meta_array_10_2 = 1'h0;
  end
  if (reset) begin
    meta_array_10_3 = 1'h0;
  end
  if (reset) begin
    meta_array_10_4 = 1'h0;
  end
  if (reset) begin
    meta_array_10_5 = 1'h0;
  end
  if (reset) begin
    meta_array_10_6 = 1'h0;
  end
  if (reset) begin
    meta_array_10_7 = 1'h0;
  end
  if (reset) begin
    meta_array_11_0 = 1'h0;
  end
  if (reset) begin
    meta_array_11_1 = 1'h0;
  end
  if (reset) begin
    meta_array_11_2 = 1'h0;
  end
  if (reset) begin
    meta_array_11_3 = 1'h0;
  end
  if (reset) begin
    meta_array_11_4 = 1'h0;
  end
  if (reset) begin
    meta_array_11_5 = 1'h0;
  end
  if (reset) begin
    meta_array_11_6 = 1'h0;
  end
  if (reset) begin
    meta_array_11_7 = 1'h0;
  end
  if (reset) begin
    meta_array_12_0 = 1'h0;
  end
  if (reset) begin
    meta_array_12_1 = 1'h0;
  end
  if (reset) begin
    meta_array_12_2 = 1'h0;
  end
  if (reset) begin
    meta_array_12_3 = 1'h0;
  end
  if (reset) begin
    meta_array_12_4 = 1'h0;
  end
  if (reset) begin
    meta_array_12_5 = 1'h0;
  end
  if (reset) begin
    meta_array_12_6 = 1'h0;
  end
  if (reset) begin
    meta_array_12_7 = 1'h0;
  end
  if (reset) begin
    meta_array_13_0 = 1'h0;
  end
  if (reset) begin
    meta_array_13_1 = 1'h0;
  end
  if (reset) begin
    meta_array_13_2 = 1'h0;
  end
  if (reset) begin
    meta_array_13_3 = 1'h0;
  end
  if (reset) begin
    meta_array_13_4 = 1'h0;
  end
  if (reset) begin
    meta_array_13_5 = 1'h0;
  end
  if (reset) begin
    meta_array_13_6 = 1'h0;
  end
  if (reset) begin
    meta_array_13_7 = 1'h0;
  end
  if (reset) begin
    meta_array_14_0 = 1'h0;
  end
  if (reset) begin
    meta_array_14_1 = 1'h0;
  end
  if (reset) begin
    meta_array_14_2 = 1'h0;
  end
  if (reset) begin
    meta_array_14_3 = 1'h0;
  end
  if (reset) begin
    meta_array_14_4 = 1'h0;
  end
  if (reset) begin
    meta_array_14_5 = 1'h0;
  end
  if (reset) begin
    meta_array_14_6 = 1'h0;
  end
  if (reset) begin
    meta_array_14_7 = 1'h0;
  end
  if (reset) begin
    meta_array_15_0 = 1'h0;
  end
  if (reset) begin
    meta_array_15_1 = 1'h0;
  end
  if (reset) begin
    meta_array_15_2 = 1'h0;
  end
  if (reset) begin
    meta_array_15_3 = 1'h0;
  end
  if (reset) begin
    meta_array_15_4 = 1'h0;
  end
  if (reset) begin
    meta_array_15_5 = 1'h0;
  end
  if (reset) begin
    meta_array_15_6 = 1'h0;
  end
  if (reset) begin
    meta_array_15_7 = 1'h0;
  end
  if (reset) begin
    meta_array_16_0 = 1'h0;
  end
  if (reset) begin
    meta_array_16_1 = 1'h0;
  end
  if (reset) begin
    meta_array_16_2 = 1'h0;
  end
  if (reset) begin
    meta_array_16_3 = 1'h0;
  end
  if (reset) begin
    meta_array_16_4 = 1'h0;
  end
  if (reset) begin
    meta_array_16_5 = 1'h0;
  end
  if (reset) begin
    meta_array_16_6 = 1'h0;
  end
  if (reset) begin
    meta_array_16_7 = 1'h0;
  end
  if (reset) begin
    meta_array_17_0 = 1'h0;
  end
  if (reset) begin
    meta_array_17_1 = 1'h0;
  end
  if (reset) begin
    meta_array_17_2 = 1'h0;
  end
  if (reset) begin
    meta_array_17_3 = 1'h0;
  end
  if (reset) begin
    meta_array_17_4 = 1'h0;
  end
  if (reset) begin
    meta_array_17_5 = 1'h0;
  end
  if (reset) begin
    meta_array_17_6 = 1'h0;
  end
  if (reset) begin
    meta_array_17_7 = 1'h0;
  end
  if (reset) begin
    meta_array_18_0 = 1'h0;
  end
  if (reset) begin
    meta_array_18_1 = 1'h0;
  end
  if (reset) begin
    meta_array_18_2 = 1'h0;
  end
  if (reset) begin
    meta_array_18_3 = 1'h0;
  end
  if (reset) begin
    meta_array_18_4 = 1'h0;
  end
  if (reset) begin
    meta_array_18_5 = 1'h0;
  end
  if (reset) begin
    meta_array_18_6 = 1'h0;
  end
  if (reset) begin
    meta_array_18_7 = 1'h0;
  end
  if (reset) begin
    meta_array_19_0 = 1'h0;
  end
  if (reset) begin
    meta_array_19_1 = 1'h0;
  end
  if (reset) begin
    meta_array_19_2 = 1'h0;
  end
  if (reset) begin
    meta_array_19_3 = 1'h0;
  end
  if (reset) begin
    meta_array_19_4 = 1'h0;
  end
  if (reset) begin
    meta_array_19_5 = 1'h0;
  end
  if (reset) begin
    meta_array_19_6 = 1'h0;
  end
  if (reset) begin
    meta_array_19_7 = 1'h0;
  end
  if (reset) begin
    meta_array_20_0 = 1'h0;
  end
  if (reset) begin
    meta_array_20_1 = 1'h0;
  end
  if (reset) begin
    meta_array_20_2 = 1'h0;
  end
  if (reset) begin
    meta_array_20_3 = 1'h0;
  end
  if (reset) begin
    meta_array_20_4 = 1'h0;
  end
  if (reset) begin
    meta_array_20_5 = 1'h0;
  end
  if (reset) begin
    meta_array_20_6 = 1'h0;
  end
  if (reset) begin
    meta_array_20_7 = 1'h0;
  end
  if (reset) begin
    meta_array_21_0 = 1'h0;
  end
  if (reset) begin
    meta_array_21_1 = 1'h0;
  end
  if (reset) begin
    meta_array_21_2 = 1'h0;
  end
  if (reset) begin
    meta_array_21_3 = 1'h0;
  end
  if (reset) begin
    meta_array_21_4 = 1'h0;
  end
  if (reset) begin
    meta_array_21_5 = 1'h0;
  end
  if (reset) begin
    meta_array_21_6 = 1'h0;
  end
  if (reset) begin
    meta_array_21_7 = 1'h0;
  end
  if (reset) begin
    meta_array_22_0 = 1'h0;
  end
  if (reset) begin
    meta_array_22_1 = 1'h0;
  end
  if (reset) begin
    meta_array_22_2 = 1'h0;
  end
  if (reset) begin
    meta_array_22_3 = 1'h0;
  end
  if (reset) begin
    meta_array_22_4 = 1'h0;
  end
  if (reset) begin
    meta_array_22_5 = 1'h0;
  end
  if (reset) begin
    meta_array_22_6 = 1'h0;
  end
  if (reset) begin
    meta_array_22_7 = 1'h0;
  end
  if (reset) begin
    meta_array_23_0 = 1'h0;
  end
  if (reset) begin
    meta_array_23_1 = 1'h0;
  end
  if (reset) begin
    meta_array_23_2 = 1'h0;
  end
  if (reset) begin
    meta_array_23_3 = 1'h0;
  end
  if (reset) begin
    meta_array_23_4 = 1'h0;
  end
  if (reset) begin
    meta_array_23_5 = 1'h0;
  end
  if (reset) begin
    meta_array_23_6 = 1'h0;
  end
  if (reset) begin
    meta_array_23_7 = 1'h0;
  end
  if (reset) begin
    meta_array_24_0 = 1'h0;
  end
  if (reset) begin
    meta_array_24_1 = 1'h0;
  end
  if (reset) begin
    meta_array_24_2 = 1'h0;
  end
  if (reset) begin
    meta_array_24_3 = 1'h0;
  end
  if (reset) begin
    meta_array_24_4 = 1'h0;
  end
  if (reset) begin
    meta_array_24_5 = 1'h0;
  end
  if (reset) begin
    meta_array_24_6 = 1'h0;
  end
  if (reset) begin
    meta_array_24_7 = 1'h0;
  end
  if (reset) begin
    meta_array_25_0 = 1'h0;
  end
  if (reset) begin
    meta_array_25_1 = 1'h0;
  end
  if (reset) begin
    meta_array_25_2 = 1'h0;
  end
  if (reset) begin
    meta_array_25_3 = 1'h0;
  end
  if (reset) begin
    meta_array_25_4 = 1'h0;
  end
  if (reset) begin
    meta_array_25_5 = 1'h0;
  end
  if (reset) begin
    meta_array_25_6 = 1'h0;
  end
  if (reset) begin
    meta_array_25_7 = 1'h0;
  end
  if (reset) begin
    meta_array_26_0 = 1'h0;
  end
  if (reset) begin
    meta_array_26_1 = 1'h0;
  end
  if (reset) begin
    meta_array_26_2 = 1'h0;
  end
  if (reset) begin
    meta_array_26_3 = 1'h0;
  end
  if (reset) begin
    meta_array_26_4 = 1'h0;
  end
  if (reset) begin
    meta_array_26_5 = 1'h0;
  end
  if (reset) begin
    meta_array_26_6 = 1'h0;
  end
  if (reset) begin
    meta_array_26_7 = 1'h0;
  end
  if (reset) begin
    meta_array_27_0 = 1'h0;
  end
  if (reset) begin
    meta_array_27_1 = 1'h0;
  end
  if (reset) begin
    meta_array_27_2 = 1'h0;
  end
  if (reset) begin
    meta_array_27_3 = 1'h0;
  end
  if (reset) begin
    meta_array_27_4 = 1'h0;
  end
  if (reset) begin
    meta_array_27_5 = 1'h0;
  end
  if (reset) begin
    meta_array_27_6 = 1'h0;
  end
  if (reset) begin
    meta_array_27_7 = 1'h0;
  end
  if (reset) begin
    meta_array_28_0 = 1'h0;
  end
  if (reset) begin
    meta_array_28_1 = 1'h0;
  end
  if (reset) begin
    meta_array_28_2 = 1'h0;
  end
  if (reset) begin
    meta_array_28_3 = 1'h0;
  end
  if (reset) begin
    meta_array_28_4 = 1'h0;
  end
  if (reset) begin
    meta_array_28_5 = 1'h0;
  end
  if (reset) begin
    meta_array_28_6 = 1'h0;
  end
  if (reset) begin
    meta_array_28_7 = 1'h0;
  end
  if (reset) begin
    meta_array_29_0 = 1'h0;
  end
  if (reset) begin
    meta_array_29_1 = 1'h0;
  end
  if (reset) begin
    meta_array_29_2 = 1'h0;
  end
  if (reset) begin
    meta_array_29_3 = 1'h0;
  end
  if (reset) begin
    meta_array_29_4 = 1'h0;
  end
  if (reset) begin
    meta_array_29_5 = 1'h0;
  end
  if (reset) begin
    meta_array_29_6 = 1'h0;
  end
  if (reset) begin
    meta_array_29_7 = 1'h0;
  end
  if (reset) begin
    meta_array_30_0 = 1'h0;
  end
  if (reset) begin
    meta_array_30_1 = 1'h0;
  end
  if (reset) begin
    meta_array_30_2 = 1'h0;
  end
  if (reset) begin
    meta_array_30_3 = 1'h0;
  end
  if (reset) begin
    meta_array_30_4 = 1'h0;
  end
  if (reset) begin
    meta_array_30_5 = 1'h0;
  end
  if (reset) begin
    meta_array_30_6 = 1'h0;
  end
  if (reset) begin
    meta_array_30_7 = 1'h0;
  end
  if (reset) begin
    meta_array_31_0 = 1'h0;
  end
  if (reset) begin
    meta_array_31_1 = 1'h0;
  end
  if (reset) begin
    meta_array_31_2 = 1'h0;
  end
  if (reset) begin
    meta_array_31_3 = 1'h0;
  end
  if (reset) begin
    meta_array_31_4 = 1'h0;
  end
  if (reset) begin
    meta_array_31_5 = 1'h0;
  end
  if (reset) begin
    meta_array_31_6 = 1'h0;
  end
  if (reset) begin
    meta_array_31_7 = 1'h0;
  end
  if (reset) begin
    meta_array_32_0 = 1'h0;
  end
  if (reset) begin
    meta_array_32_1 = 1'h0;
  end
  if (reset) begin
    meta_array_32_2 = 1'h0;
  end
  if (reset) begin
    meta_array_32_3 = 1'h0;
  end
  if (reset) begin
    meta_array_32_4 = 1'h0;
  end
  if (reset) begin
    meta_array_32_5 = 1'h0;
  end
  if (reset) begin
    meta_array_32_6 = 1'h0;
  end
  if (reset) begin
    meta_array_32_7 = 1'h0;
  end
  if (reset) begin
    meta_array_33_0 = 1'h0;
  end
  if (reset) begin
    meta_array_33_1 = 1'h0;
  end
  if (reset) begin
    meta_array_33_2 = 1'h0;
  end
  if (reset) begin
    meta_array_33_3 = 1'h0;
  end
  if (reset) begin
    meta_array_33_4 = 1'h0;
  end
  if (reset) begin
    meta_array_33_5 = 1'h0;
  end
  if (reset) begin
    meta_array_33_6 = 1'h0;
  end
  if (reset) begin
    meta_array_33_7 = 1'h0;
  end
  if (reset) begin
    meta_array_34_0 = 1'h0;
  end
  if (reset) begin
    meta_array_34_1 = 1'h0;
  end
  if (reset) begin
    meta_array_34_2 = 1'h0;
  end
  if (reset) begin
    meta_array_34_3 = 1'h0;
  end
  if (reset) begin
    meta_array_34_4 = 1'h0;
  end
  if (reset) begin
    meta_array_34_5 = 1'h0;
  end
  if (reset) begin
    meta_array_34_6 = 1'h0;
  end
  if (reset) begin
    meta_array_34_7 = 1'h0;
  end
  if (reset) begin
    meta_array_35_0 = 1'h0;
  end
  if (reset) begin
    meta_array_35_1 = 1'h0;
  end
  if (reset) begin
    meta_array_35_2 = 1'h0;
  end
  if (reset) begin
    meta_array_35_3 = 1'h0;
  end
  if (reset) begin
    meta_array_35_4 = 1'h0;
  end
  if (reset) begin
    meta_array_35_5 = 1'h0;
  end
  if (reset) begin
    meta_array_35_6 = 1'h0;
  end
  if (reset) begin
    meta_array_35_7 = 1'h0;
  end
  if (reset) begin
    meta_array_36_0 = 1'h0;
  end
  if (reset) begin
    meta_array_36_1 = 1'h0;
  end
  if (reset) begin
    meta_array_36_2 = 1'h0;
  end
  if (reset) begin
    meta_array_36_3 = 1'h0;
  end
  if (reset) begin
    meta_array_36_4 = 1'h0;
  end
  if (reset) begin
    meta_array_36_5 = 1'h0;
  end
  if (reset) begin
    meta_array_36_6 = 1'h0;
  end
  if (reset) begin
    meta_array_36_7 = 1'h0;
  end
  if (reset) begin
    meta_array_37_0 = 1'h0;
  end
  if (reset) begin
    meta_array_37_1 = 1'h0;
  end
  if (reset) begin
    meta_array_37_2 = 1'h0;
  end
  if (reset) begin
    meta_array_37_3 = 1'h0;
  end
  if (reset) begin
    meta_array_37_4 = 1'h0;
  end
  if (reset) begin
    meta_array_37_5 = 1'h0;
  end
  if (reset) begin
    meta_array_37_6 = 1'h0;
  end
  if (reset) begin
    meta_array_37_7 = 1'h0;
  end
  if (reset) begin
    meta_array_38_0 = 1'h0;
  end
  if (reset) begin
    meta_array_38_1 = 1'h0;
  end
  if (reset) begin
    meta_array_38_2 = 1'h0;
  end
  if (reset) begin
    meta_array_38_3 = 1'h0;
  end
  if (reset) begin
    meta_array_38_4 = 1'h0;
  end
  if (reset) begin
    meta_array_38_5 = 1'h0;
  end
  if (reset) begin
    meta_array_38_6 = 1'h0;
  end
  if (reset) begin
    meta_array_38_7 = 1'h0;
  end
  if (reset) begin
    meta_array_39_0 = 1'h0;
  end
  if (reset) begin
    meta_array_39_1 = 1'h0;
  end
  if (reset) begin
    meta_array_39_2 = 1'h0;
  end
  if (reset) begin
    meta_array_39_3 = 1'h0;
  end
  if (reset) begin
    meta_array_39_4 = 1'h0;
  end
  if (reset) begin
    meta_array_39_5 = 1'h0;
  end
  if (reset) begin
    meta_array_39_6 = 1'h0;
  end
  if (reset) begin
    meta_array_39_7 = 1'h0;
  end
  if (reset) begin
    meta_array_40_0 = 1'h0;
  end
  if (reset) begin
    meta_array_40_1 = 1'h0;
  end
  if (reset) begin
    meta_array_40_2 = 1'h0;
  end
  if (reset) begin
    meta_array_40_3 = 1'h0;
  end
  if (reset) begin
    meta_array_40_4 = 1'h0;
  end
  if (reset) begin
    meta_array_40_5 = 1'h0;
  end
  if (reset) begin
    meta_array_40_6 = 1'h0;
  end
  if (reset) begin
    meta_array_40_7 = 1'h0;
  end
  if (reset) begin
    meta_array_41_0 = 1'h0;
  end
  if (reset) begin
    meta_array_41_1 = 1'h0;
  end
  if (reset) begin
    meta_array_41_2 = 1'h0;
  end
  if (reset) begin
    meta_array_41_3 = 1'h0;
  end
  if (reset) begin
    meta_array_41_4 = 1'h0;
  end
  if (reset) begin
    meta_array_41_5 = 1'h0;
  end
  if (reset) begin
    meta_array_41_6 = 1'h0;
  end
  if (reset) begin
    meta_array_41_7 = 1'h0;
  end
  if (reset) begin
    meta_array_42_0 = 1'h0;
  end
  if (reset) begin
    meta_array_42_1 = 1'h0;
  end
  if (reset) begin
    meta_array_42_2 = 1'h0;
  end
  if (reset) begin
    meta_array_42_3 = 1'h0;
  end
  if (reset) begin
    meta_array_42_4 = 1'h0;
  end
  if (reset) begin
    meta_array_42_5 = 1'h0;
  end
  if (reset) begin
    meta_array_42_6 = 1'h0;
  end
  if (reset) begin
    meta_array_42_7 = 1'h0;
  end
  if (reset) begin
    meta_array_43_0 = 1'h0;
  end
  if (reset) begin
    meta_array_43_1 = 1'h0;
  end
  if (reset) begin
    meta_array_43_2 = 1'h0;
  end
  if (reset) begin
    meta_array_43_3 = 1'h0;
  end
  if (reset) begin
    meta_array_43_4 = 1'h0;
  end
  if (reset) begin
    meta_array_43_5 = 1'h0;
  end
  if (reset) begin
    meta_array_43_6 = 1'h0;
  end
  if (reset) begin
    meta_array_43_7 = 1'h0;
  end
  if (reset) begin
    meta_array_44_0 = 1'h0;
  end
  if (reset) begin
    meta_array_44_1 = 1'h0;
  end
  if (reset) begin
    meta_array_44_2 = 1'h0;
  end
  if (reset) begin
    meta_array_44_3 = 1'h0;
  end
  if (reset) begin
    meta_array_44_4 = 1'h0;
  end
  if (reset) begin
    meta_array_44_5 = 1'h0;
  end
  if (reset) begin
    meta_array_44_6 = 1'h0;
  end
  if (reset) begin
    meta_array_44_7 = 1'h0;
  end
  if (reset) begin
    meta_array_45_0 = 1'h0;
  end
  if (reset) begin
    meta_array_45_1 = 1'h0;
  end
  if (reset) begin
    meta_array_45_2 = 1'h0;
  end
  if (reset) begin
    meta_array_45_3 = 1'h0;
  end
  if (reset) begin
    meta_array_45_4 = 1'h0;
  end
  if (reset) begin
    meta_array_45_5 = 1'h0;
  end
  if (reset) begin
    meta_array_45_6 = 1'h0;
  end
  if (reset) begin
    meta_array_45_7 = 1'h0;
  end
  if (reset) begin
    meta_array_46_0 = 1'h0;
  end
  if (reset) begin
    meta_array_46_1 = 1'h0;
  end
  if (reset) begin
    meta_array_46_2 = 1'h0;
  end
  if (reset) begin
    meta_array_46_3 = 1'h0;
  end
  if (reset) begin
    meta_array_46_4 = 1'h0;
  end
  if (reset) begin
    meta_array_46_5 = 1'h0;
  end
  if (reset) begin
    meta_array_46_6 = 1'h0;
  end
  if (reset) begin
    meta_array_46_7 = 1'h0;
  end
  if (reset) begin
    meta_array_47_0 = 1'h0;
  end
  if (reset) begin
    meta_array_47_1 = 1'h0;
  end
  if (reset) begin
    meta_array_47_2 = 1'h0;
  end
  if (reset) begin
    meta_array_47_3 = 1'h0;
  end
  if (reset) begin
    meta_array_47_4 = 1'h0;
  end
  if (reset) begin
    meta_array_47_5 = 1'h0;
  end
  if (reset) begin
    meta_array_47_6 = 1'h0;
  end
  if (reset) begin
    meta_array_47_7 = 1'h0;
  end
  if (reset) begin
    meta_array_48_0 = 1'h0;
  end
  if (reset) begin
    meta_array_48_1 = 1'h0;
  end
  if (reset) begin
    meta_array_48_2 = 1'h0;
  end
  if (reset) begin
    meta_array_48_3 = 1'h0;
  end
  if (reset) begin
    meta_array_48_4 = 1'h0;
  end
  if (reset) begin
    meta_array_48_5 = 1'h0;
  end
  if (reset) begin
    meta_array_48_6 = 1'h0;
  end
  if (reset) begin
    meta_array_48_7 = 1'h0;
  end
  if (reset) begin
    meta_array_49_0 = 1'h0;
  end
  if (reset) begin
    meta_array_49_1 = 1'h0;
  end
  if (reset) begin
    meta_array_49_2 = 1'h0;
  end
  if (reset) begin
    meta_array_49_3 = 1'h0;
  end
  if (reset) begin
    meta_array_49_4 = 1'h0;
  end
  if (reset) begin
    meta_array_49_5 = 1'h0;
  end
  if (reset) begin
    meta_array_49_6 = 1'h0;
  end
  if (reset) begin
    meta_array_49_7 = 1'h0;
  end
  if (reset) begin
    meta_array_50_0 = 1'h0;
  end
  if (reset) begin
    meta_array_50_1 = 1'h0;
  end
  if (reset) begin
    meta_array_50_2 = 1'h0;
  end
  if (reset) begin
    meta_array_50_3 = 1'h0;
  end
  if (reset) begin
    meta_array_50_4 = 1'h0;
  end
  if (reset) begin
    meta_array_50_5 = 1'h0;
  end
  if (reset) begin
    meta_array_50_6 = 1'h0;
  end
  if (reset) begin
    meta_array_50_7 = 1'h0;
  end
  if (reset) begin
    meta_array_51_0 = 1'h0;
  end
  if (reset) begin
    meta_array_51_1 = 1'h0;
  end
  if (reset) begin
    meta_array_51_2 = 1'h0;
  end
  if (reset) begin
    meta_array_51_3 = 1'h0;
  end
  if (reset) begin
    meta_array_51_4 = 1'h0;
  end
  if (reset) begin
    meta_array_51_5 = 1'h0;
  end
  if (reset) begin
    meta_array_51_6 = 1'h0;
  end
  if (reset) begin
    meta_array_51_7 = 1'h0;
  end
  if (reset) begin
    meta_array_52_0 = 1'h0;
  end
  if (reset) begin
    meta_array_52_1 = 1'h0;
  end
  if (reset) begin
    meta_array_52_2 = 1'h0;
  end
  if (reset) begin
    meta_array_52_3 = 1'h0;
  end
  if (reset) begin
    meta_array_52_4 = 1'h0;
  end
  if (reset) begin
    meta_array_52_5 = 1'h0;
  end
  if (reset) begin
    meta_array_52_6 = 1'h0;
  end
  if (reset) begin
    meta_array_52_7 = 1'h0;
  end
  if (reset) begin
    meta_array_53_0 = 1'h0;
  end
  if (reset) begin
    meta_array_53_1 = 1'h0;
  end
  if (reset) begin
    meta_array_53_2 = 1'h0;
  end
  if (reset) begin
    meta_array_53_3 = 1'h0;
  end
  if (reset) begin
    meta_array_53_4 = 1'h0;
  end
  if (reset) begin
    meta_array_53_5 = 1'h0;
  end
  if (reset) begin
    meta_array_53_6 = 1'h0;
  end
  if (reset) begin
    meta_array_53_7 = 1'h0;
  end
  if (reset) begin
    meta_array_54_0 = 1'h0;
  end
  if (reset) begin
    meta_array_54_1 = 1'h0;
  end
  if (reset) begin
    meta_array_54_2 = 1'h0;
  end
  if (reset) begin
    meta_array_54_3 = 1'h0;
  end
  if (reset) begin
    meta_array_54_4 = 1'h0;
  end
  if (reset) begin
    meta_array_54_5 = 1'h0;
  end
  if (reset) begin
    meta_array_54_6 = 1'h0;
  end
  if (reset) begin
    meta_array_54_7 = 1'h0;
  end
  if (reset) begin
    meta_array_55_0 = 1'h0;
  end
  if (reset) begin
    meta_array_55_1 = 1'h0;
  end
  if (reset) begin
    meta_array_55_2 = 1'h0;
  end
  if (reset) begin
    meta_array_55_3 = 1'h0;
  end
  if (reset) begin
    meta_array_55_4 = 1'h0;
  end
  if (reset) begin
    meta_array_55_5 = 1'h0;
  end
  if (reset) begin
    meta_array_55_6 = 1'h0;
  end
  if (reset) begin
    meta_array_55_7 = 1'h0;
  end
  if (reset) begin
    meta_array_56_0 = 1'h0;
  end
  if (reset) begin
    meta_array_56_1 = 1'h0;
  end
  if (reset) begin
    meta_array_56_2 = 1'h0;
  end
  if (reset) begin
    meta_array_56_3 = 1'h0;
  end
  if (reset) begin
    meta_array_56_4 = 1'h0;
  end
  if (reset) begin
    meta_array_56_5 = 1'h0;
  end
  if (reset) begin
    meta_array_56_6 = 1'h0;
  end
  if (reset) begin
    meta_array_56_7 = 1'h0;
  end
  if (reset) begin
    meta_array_57_0 = 1'h0;
  end
  if (reset) begin
    meta_array_57_1 = 1'h0;
  end
  if (reset) begin
    meta_array_57_2 = 1'h0;
  end
  if (reset) begin
    meta_array_57_3 = 1'h0;
  end
  if (reset) begin
    meta_array_57_4 = 1'h0;
  end
  if (reset) begin
    meta_array_57_5 = 1'h0;
  end
  if (reset) begin
    meta_array_57_6 = 1'h0;
  end
  if (reset) begin
    meta_array_57_7 = 1'h0;
  end
  if (reset) begin
    meta_array_58_0 = 1'h0;
  end
  if (reset) begin
    meta_array_58_1 = 1'h0;
  end
  if (reset) begin
    meta_array_58_2 = 1'h0;
  end
  if (reset) begin
    meta_array_58_3 = 1'h0;
  end
  if (reset) begin
    meta_array_58_4 = 1'h0;
  end
  if (reset) begin
    meta_array_58_5 = 1'h0;
  end
  if (reset) begin
    meta_array_58_6 = 1'h0;
  end
  if (reset) begin
    meta_array_58_7 = 1'h0;
  end
  if (reset) begin
    meta_array_59_0 = 1'h0;
  end
  if (reset) begin
    meta_array_59_1 = 1'h0;
  end
  if (reset) begin
    meta_array_59_2 = 1'h0;
  end
  if (reset) begin
    meta_array_59_3 = 1'h0;
  end
  if (reset) begin
    meta_array_59_4 = 1'h0;
  end
  if (reset) begin
    meta_array_59_5 = 1'h0;
  end
  if (reset) begin
    meta_array_59_6 = 1'h0;
  end
  if (reset) begin
    meta_array_59_7 = 1'h0;
  end
  if (reset) begin
    meta_array_60_0 = 1'h0;
  end
  if (reset) begin
    meta_array_60_1 = 1'h0;
  end
  if (reset) begin
    meta_array_60_2 = 1'h0;
  end
  if (reset) begin
    meta_array_60_3 = 1'h0;
  end
  if (reset) begin
    meta_array_60_4 = 1'h0;
  end
  if (reset) begin
    meta_array_60_5 = 1'h0;
  end
  if (reset) begin
    meta_array_60_6 = 1'h0;
  end
  if (reset) begin
    meta_array_60_7 = 1'h0;
  end
  if (reset) begin
    meta_array_61_0 = 1'h0;
  end
  if (reset) begin
    meta_array_61_1 = 1'h0;
  end
  if (reset) begin
    meta_array_61_2 = 1'h0;
  end
  if (reset) begin
    meta_array_61_3 = 1'h0;
  end
  if (reset) begin
    meta_array_61_4 = 1'h0;
  end
  if (reset) begin
    meta_array_61_5 = 1'h0;
  end
  if (reset) begin
    meta_array_61_6 = 1'h0;
  end
  if (reset) begin
    meta_array_61_7 = 1'h0;
  end
  if (reset) begin
    meta_array_62_0 = 1'h0;
  end
  if (reset) begin
    meta_array_62_1 = 1'h0;
  end
  if (reset) begin
    meta_array_62_2 = 1'h0;
  end
  if (reset) begin
    meta_array_62_3 = 1'h0;
  end
  if (reset) begin
    meta_array_62_4 = 1'h0;
  end
  if (reset) begin
    meta_array_62_5 = 1'h0;
  end
  if (reset) begin
    meta_array_62_6 = 1'h0;
  end
  if (reset) begin
    meta_array_62_7 = 1'h0;
  end
  if (reset) begin
    meta_array_63_0 = 1'h0;
  end
  if (reset) begin
    meta_array_63_1 = 1'h0;
  end
  if (reset) begin
    meta_array_63_2 = 1'h0;
  end
  if (reset) begin
    meta_array_63_3 = 1'h0;
  end
  if (reset) begin
    meta_array_63_4 = 1'h0;
  end
  if (reset) begin
    meta_array_63_5 = 1'h0;
  end
  if (reset) begin
    meta_array_63_6 = 1'h0;
  end
  if (reset) begin
    meta_array_63_7 = 1'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule

