module ImmExtractor(
  input  [63:0] io_data_in_0,
  output [63:0] io_data_out_0
);
  assign io_data_out_0 = io_data_in_0; // @[DataArray.scala 110:15]
endmodule

