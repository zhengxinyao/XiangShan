module PLICFanIn(
  input  [2:0]  io_prio_0,
  input  [2:0]  io_prio_1,
  input  [2:0]  io_prio_2,
  input  [2:0]  io_prio_3,
  input  [2:0]  io_prio_4,
  input  [2:0]  io_prio_5,
  input  [2:0]  io_prio_6,
  input  [2:0]  io_prio_7,
  input  [2:0]  io_prio_8,
  input  [2:0]  io_prio_9,
  input  [2:0]  io_prio_10,
  input  [2:0]  io_prio_11,
  input  [2:0]  io_prio_12,
  input  [2:0]  io_prio_13,
  input  [2:0]  io_prio_14,
  input  [2:0]  io_prio_15,
  input  [2:0]  io_prio_16,
  input  [2:0]  io_prio_17,
  input  [2:0]  io_prio_18,
  input  [2:0]  io_prio_19,
  input  [2:0]  io_prio_20,
  input  [2:0]  io_prio_21,
  input  [2:0]  io_prio_22,
  input  [2:0]  io_prio_23,
  input  [2:0]  io_prio_24,
  input  [2:0]  io_prio_25,
  input  [2:0]  io_prio_26,
  input  [2:0]  io_prio_27,
  input  [2:0]  io_prio_28,
  input  [2:0]  io_prio_29,
  input  [2:0]  io_prio_30,
  input  [2:0]  io_prio_31,
  input  [2:0]  io_prio_32,
  input  [2:0]  io_prio_33,
  input  [2:0]  io_prio_34,
  input  [2:0]  io_prio_35,
  input  [2:0]  io_prio_36,
  input  [2:0]  io_prio_37,
  input  [2:0]  io_prio_38,
  input  [2:0]  io_prio_39,
  input  [2:0]  io_prio_40,
  input  [2:0]  io_prio_41,
  input  [2:0]  io_prio_42,
  input  [2:0]  io_prio_43,
  input  [2:0]  io_prio_44,
  input  [2:0]  io_prio_45,
  input  [2:0]  io_prio_46,
  input  [2:0]  io_prio_47,
  input  [2:0]  io_prio_48,
  input  [2:0]  io_prio_49,
  input  [2:0]  io_prio_50,
  input  [2:0]  io_prio_51,
  input  [2:0]  io_prio_52,
  input  [2:0]  io_prio_53,
  input  [2:0]  io_prio_54,
  input  [2:0]  io_prio_55,
  input  [2:0]  io_prio_56,
  input  [2:0]  io_prio_57,
  input  [2:0]  io_prio_58,
  input  [2:0]  io_prio_59,
  input  [2:0]  io_prio_60,
  input  [2:0]  io_prio_61,
  input  [2:0]  io_prio_62,
  input  [2:0]  io_prio_63,
  input  [2:0]  io_prio_64,
  input  [64:0] io_ip,
  output [6:0]  io_dev,
  output [2:0]  io_max
);
  wire [3:0] effectivePriority_1 = {io_ip[0],io_prio_0}; // @[Cat.scala 31:58]
  wire [3:0] effectivePriority_2 = {io_ip[1],io_prio_1}; // @[Cat.scala 31:58]
  wire [3:0] effectivePriority_3 = {io_ip[2],io_prio_2}; // @[Cat.scala 31:58]
  wire [3:0] effectivePriority_4 = {io_ip[3],io_prio_3}; // @[Cat.scala 31:58]
  wire [3:0] effectivePriority_5 = {io_ip[4],io_prio_4}; // @[Cat.scala 31:58]
  wire [3:0] effectivePriority_6 = {io_ip[5],io_prio_5}; // @[Cat.scala 31:58]
  wire [3:0] effectivePriority_7 = {io_ip[6],io_prio_6}; // @[Cat.scala 31:58]
  wire [3:0] effectivePriority_8 = {io_ip[7],io_prio_7}; // @[Cat.scala 31:58]
  wire [3:0] effectivePriority_9 = {io_ip[8],io_prio_8}; // @[Cat.scala 31:58]
  wire [3:0] effectivePriority_10 = {io_ip[9],io_prio_9}; // @[Cat.scala 31:58]
  wire [3:0] effectivePriority_11 = {io_ip[10],io_prio_10}; // @[Cat.scala 31:58]
  wire [3:0] effectivePriority_12 = {io_ip[11],io_prio_11}; // @[Cat.scala 31:58]
  wire [3:0] effectivePriority_13 = {io_ip[12],io_prio_12}; // @[Cat.scala 31:58]
  wire [3:0] effectivePriority_14 = {io_ip[13],io_prio_13}; // @[Cat.scala 31:58]
  wire [3:0] effectivePriority_15 = {io_ip[14],io_prio_14}; // @[Cat.scala 31:58]
  wire [3:0] effectivePriority_16 = {io_ip[15],io_prio_15}; // @[Cat.scala 31:58]
  wire [3:0] effectivePriority_17 = {io_ip[16],io_prio_16}; // @[Cat.scala 31:58]
  wire [3:0] effectivePriority_18 = {io_ip[17],io_prio_17}; // @[Cat.scala 31:58]
  wire [3:0] effectivePriority_19 = {io_ip[18],io_prio_18}; // @[Cat.scala 31:58]
  wire [3:0] effectivePriority_20 = {io_ip[19],io_prio_19}; // @[Cat.scala 31:58]
  wire [3:0] effectivePriority_21 = {io_ip[20],io_prio_20}; // @[Cat.scala 31:58]
  wire [3:0] effectivePriority_22 = {io_ip[21],io_prio_21}; // @[Cat.scala 31:58]
  wire [3:0] effectivePriority_23 = {io_ip[22],io_prio_22}; // @[Cat.scala 31:58]
  wire [3:0] effectivePriority_24 = {io_ip[23],io_prio_23}; // @[Cat.scala 31:58]
  wire [3:0] effectivePriority_25 = {io_ip[24],io_prio_24}; // @[Cat.scala 31:58]
  wire [3:0] effectivePriority_26 = {io_ip[25],io_prio_25}; // @[Cat.scala 31:58]
  wire [3:0] effectivePriority_27 = {io_ip[26],io_prio_26}; // @[Cat.scala 31:58]
  wire [3:0] effectivePriority_28 = {io_ip[27],io_prio_27}; // @[Cat.scala 31:58]
  wire [3:0] effectivePriority_29 = {io_ip[28],io_prio_28}; // @[Cat.scala 31:58]
  wire [3:0] effectivePriority_30 = {io_ip[29],io_prio_29}; // @[Cat.scala 31:58]
  wire [3:0] effectivePriority_31 = {io_ip[30],io_prio_30}; // @[Cat.scala 31:58]
  wire [3:0] effectivePriority_32 = {io_ip[31],io_prio_31}; // @[Cat.scala 31:58]
  wire [3:0] effectivePriority_33 = {io_ip[32],io_prio_32}; // @[Cat.scala 31:58]
  wire [3:0] effectivePriority_34 = {io_ip[33],io_prio_33}; // @[Cat.scala 31:58]
  wire [3:0] effectivePriority_35 = {io_ip[34],io_prio_34}; // @[Cat.scala 31:58]
  wire [3:0] effectivePriority_36 = {io_ip[35],io_prio_35}; // @[Cat.scala 31:58]
  wire [3:0] effectivePriority_37 = {io_ip[36],io_prio_36}; // @[Cat.scala 31:58]
  wire [3:0] effectivePriority_38 = {io_ip[37],io_prio_37}; // @[Cat.scala 31:58]
  wire [3:0] effectivePriority_39 = {io_ip[38],io_prio_38}; // @[Cat.scala 31:58]
  wire [3:0] effectivePriority_40 = {io_ip[39],io_prio_39}; // @[Cat.scala 31:58]
  wire [3:0] effectivePriority_41 = {io_ip[40],io_prio_40}; // @[Cat.scala 31:58]
  wire [3:0] effectivePriority_42 = {io_ip[41],io_prio_41}; // @[Cat.scala 31:58]
  wire [3:0] effectivePriority_43 = {io_ip[42],io_prio_42}; // @[Cat.scala 31:58]
  wire [3:0] effectivePriority_44 = {io_ip[43],io_prio_43}; // @[Cat.scala 31:58]
  wire [3:0] effectivePriority_45 = {io_ip[44],io_prio_44}; // @[Cat.scala 31:58]
  wire [3:0] effectivePriority_46 = {io_ip[45],io_prio_45}; // @[Cat.scala 31:58]
  wire [3:0] effectivePriority_47 = {io_ip[46],io_prio_46}; // @[Cat.scala 31:58]
  wire [3:0] effectivePriority_48 = {io_ip[47],io_prio_47}; // @[Cat.scala 31:58]
  wire [3:0] effectivePriority_49 = {io_ip[48],io_prio_48}; // @[Cat.scala 31:58]
  wire [3:0] effectivePriority_50 = {io_ip[49],io_prio_49}; // @[Cat.scala 31:58]
  wire [3:0] effectivePriority_51 = {io_ip[50],io_prio_50}; // @[Cat.scala 31:58]
  wire [3:0] effectivePriority_52 = {io_ip[51],io_prio_51}; // @[Cat.scala 31:58]
  wire [3:0] effectivePriority_53 = {io_ip[52],io_prio_52}; // @[Cat.scala 31:58]
  wire [3:0] effectivePriority_54 = {io_ip[53],io_prio_53}; // @[Cat.scala 31:58]
  wire [3:0] effectivePriority_55 = {io_ip[54],io_prio_54}; // @[Cat.scala 31:58]
  wire [3:0] effectivePriority_56 = {io_ip[55],io_prio_55}; // @[Cat.scala 31:58]
  wire [3:0] effectivePriority_57 = {io_ip[56],io_prio_56}; // @[Cat.scala 31:58]
  wire [3:0] effectivePriority_58 = {io_ip[57],io_prio_57}; // @[Cat.scala 31:58]
  wire [3:0] effectivePriority_59 = {io_ip[58],io_prio_58}; // @[Cat.scala 31:58]
  wire [3:0] effectivePriority_60 = {io_ip[59],io_prio_59}; // @[Cat.scala 31:58]
  wire [3:0] effectivePriority_61 = {io_ip[60],io_prio_60}; // @[Cat.scala 31:58]
  wire [3:0] effectivePriority_62 = {io_ip[61],io_prio_61}; // @[Cat.scala 31:58]
  wire [3:0] effectivePriority_63 = {io_ip[62],io_prio_62}; // @[Cat.scala 31:58]
  wire [3:0] effectivePriority_64 = {io_ip[63],io_prio_63}; // @[Cat.scala 31:58]
  wire [3:0] effectivePriority_65 = {io_ip[64],io_prio_64}; // @[Cat.scala 31:58]
  wire  _T = 4'h8 >= effectivePriority_1; // @[Plic.scala 344:20]
  wire [3:0] _T_2 = _T ? 4'h8 : effectivePriority_1; // @[Misc.scala 34:9]
  wire  _T_3 = _T ? 1'h0 : 1'h1; // @[Misc.scala 34:36]
  wire  _T_4 = effectivePriority_2 >= effectivePriority_3; // @[Plic.scala 344:20]
  wire [3:0] _T_6 = _T_4 ? effectivePriority_2 : effectivePriority_3; // @[Misc.scala 34:9]
  wire  _T_7 = _T_4 ? 1'h0 : 1'h1; // @[Misc.scala 34:36]
  wire  _T_8 = _T_2 >= _T_6; // @[Plic.scala 344:20]
  wire [1:0] _GEN_0 = {{1'd0}, _T_7}; // @[Plic.scala 344:61]
  wire [1:0] _T_9 = 2'h2 | _GEN_0; // @[Plic.scala 344:61]
  wire [3:0] _T_10 = _T_8 ? _T_2 : _T_6; // @[Misc.scala 34:9]
  wire [1:0] _T_11 = _T_8 ? {{1'd0}, _T_3} : _T_9; // @[Misc.scala 34:36]
  wire  _T_12 = effectivePriority_4 >= effectivePriority_5; // @[Plic.scala 344:20]
  wire [3:0] _T_14 = _T_12 ? effectivePriority_4 : effectivePriority_5; // @[Misc.scala 34:9]
  wire  _T_15 = _T_12 ? 1'h0 : 1'h1; // @[Misc.scala 34:36]
  wire  _T_16 = effectivePriority_6 >= effectivePriority_7; // @[Plic.scala 344:20]
  wire [3:0] _T_18 = _T_16 ? effectivePriority_6 : effectivePriority_7; // @[Misc.scala 34:9]
  wire  _T_19 = _T_16 ? 1'h0 : 1'h1; // @[Misc.scala 34:36]
  wire  _T_20 = _T_14 >= _T_18; // @[Plic.scala 344:20]
  wire [1:0] _GEN_1 = {{1'd0}, _T_19}; // @[Plic.scala 344:61]
  wire [1:0] _T_21 = 2'h2 | _GEN_1; // @[Plic.scala 344:61]
  wire [3:0] _T_22 = _T_20 ? _T_14 : _T_18; // @[Misc.scala 34:9]
  wire [1:0] _T_23 = _T_20 ? {{1'd0}, _T_15} : _T_21; // @[Misc.scala 34:36]
  wire  _T_24 = _T_10 >= _T_22; // @[Plic.scala 344:20]
  wire [2:0] _GEN_2 = {{1'd0}, _T_23}; // @[Plic.scala 344:61]
  wire [2:0] _T_25 = 3'h4 | _GEN_2; // @[Plic.scala 344:61]
  wire [3:0] _T_26 = _T_24 ? _T_10 : _T_22; // @[Misc.scala 34:9]
  wire [2:0] _T_27 = _T_24 ? {{1'd0}, _T_11} : _T_25; // @[Misc.scala 34:36]
  wire  _T_28 = effectivePriority_8 >= effectivePriority_9; // @[Plic.scala 344:20]
  wire [3:0] _T_30 = _T_28 ? effectivePriority_8 : effectivePriority_9; // @[Misc.scala 34:9]
  wire  _T_31 = _T_28 ? 1'h0 : 1'h1; // @[Misc.scala 34:36]
  wire  _T_32 = effectivePriority_10 >= effectivePriority_11; // @[Plic.scala 344:20]
  wire [3:0] _T_34 = _T_32 ? effectivePriority_10 : effectivePriority_11; // @[Misc.scala 34:9]
  wire  _T_35 = _T_32 ? 1'h0 : 1'h1; // @[Misc.scala 34:36]
  wire  _T_36 = _T_30 >= _T_34; // @[Plic.scala 344:20]
  wire [1:0] _GEN_3 = {{1'd0}, _T_35}; // @[Plic.scala 344:61]
  wire [1:0] _T_37 = 2'h2 | _GEN_3; // @[Plic.scala 344:61]
  wire [3:0] _T_38 = _T_36 ? _T_30 : _T_34; // @[Misc.scala 34:9]
  wire [1:0] _T_39 = _T_36 ? {{1'd0}, _T_31} : _T_37; // @[Misc.scala 34:36]
  wire  _T_40 = effectivePriority_12 >= effectivePriority_13; // @[Plic.scala 344:20]
  wire [3:0] _T_42 = _T_40 ? effectivePriority_12 : effectivePriority_13; // @[Misc.scala 34:9]
  wire  _T_43 = _T_40 ? 1'h0 : 1'h1; // @[Misc.scala 34:36]
  wire  _T_44 = effectivePriority_14 >= effectivePriority_15; // @[Plic.scala 344:20]
  wire [3:0] _T_46 = _T_44 ? effectivePriority_14 : effectivePriority_15; // @[Misc.scala 34:9]
  wire  _T_47 = _T_44 ? 1'h0 : 1'h1; // @[Misc.scala 34:36]
  wire  _T_48 = _T_42 >= _T_46; // @[Plic.scala 344:20]
  wire [1:0] _GEN_4 = {{1'd0}, _T_47}; // @[Plic.scala 344:61]
  wire [1:0] _T_49 = 2'h2 | _GEN_4; // @[Plic.scala 344:61]
  wire [3:0] _T_50 = _T_48 ? _T_42 : _T_46; // @[Misc.scala 34:9]
  wire [1:0] _T_51 = _T_48 ? {{1'd0}, _T_43} : _T_49; // @[Misc.scala 34:36]
  wire  _T_52 = _T_38 >= _T_50; // @[Plic.scala 344:20]
  wire [2:0] _GEN_5 = {{1'd0}, _T_51}; // @[Plic.scala 344:61]
  wire [2:0] _T_53 = 3'h4 | _GEN_5; // @[Plic.scala 344:61]
  wire [3:0] _T_54 = _T_52 ? _T_38 : _T_50; // @[Misc.scala 34:9]
  wire [2:0] _T_55 = _T_52 ? {{1'd0}, _T_39} : _T_53; // @[Misc.scala 34:36]
  wire  _T_56 = _T_26 >= _T_54; // @[Plic.scala 344:20]
  wire [3:0] _GEN_6 = {{1'd0}, _T_55}; // @[Plic.scala 344:61]
  wire [3:0] _T_57 = 4'h8 | _GEN_6; // @[Plic.scala 344:61]
  wire [3:0] _T_58 = _T_56 ? _T_26 : _T_54; // @[Misc.scala 34:9]
  wire [3:0] _T_59 = _T_56 ? {{1'd0}, _T_27} : _T_57; // @[Misc.scala 34:36]
  wire  _T_60 = effectivePriority_16 >= effectivePriority_17; // @[Plic.scala 344:20]
  wire [3:0] _T_62 = _T_60 ? effectivePriority_16 : effectivePriority_17; // @[Misc.scala 34:9]
  wire  _T_63 = _T_60 ? 1'h0 : 1'h1; // @[Misc.scala 34:36]
  wire  _T_64 = effectivePriority_18 >= effectivePriority_19; // @[Plic.scala 344:20]
  wire [3:0] _T_66 = _T_64 ? effectivePriority_18 : effectivePriority_19; // @[Misc.scala 34:9]
  wire  _T_67 = _T_64 ? 1'h0 : 1'h1; // @[Misc.scala 34:36]
  wire  _T_68 = _T_62 >= _T_66; // @[Plic.scala 344:20]
  wire [1:0] _GEN_7 = {{1'd0}, _T_67}; // @[Plic.scala 344:61]
  wire [1:0] _T_69 = 2'h2 | _GEN_7; // @[Plic.scala 344:61]
  wire [3:0] _T_70 = _T_68 ? _T_62 : _T_66; // @[Misc.scala 34:9]
  wire [1:0] _T_71 = _T_68 ? {{1'd0}, _T_63} : _T_69; // @[Misc.scala 34:36]
  wire  _T_72 = effectivePriority_20 >= effectivePriority_21; // @[Plic.scala 344:20]
  wire [3:0] _T_74 = _T_72 ? effectivePriority_20 : effectivePriority_21; // @[Misc.scala 34:9]
  wire  _T_75 = _T_72 ? 1'h0 : 1'h1; // @[Misc.scala 34:36]
  wire  _T_76 = effectivePriority_22 >= effectivePriority_23; // @[Plic.scala 344:20]
  wire [3:0] _T_78 = _T_76 ? effectivePriority_22 : effectivePriority_23; // @[Misc.scala 34:9]
  wire  _T_79 = _T_76 ? 1'h0 : 1'h1; // @[Misc.scala 34:36]
  wire  _T_80 = _T_74 >= _T_78; // @[Plic.scala 344:20]
  wire [1:0] _GEN_8 = {{1'd0}, _T_79}; // @[Plic.scala 344:61]
  wire [1:0] _T_81 = 2'h2 | _GEN_8; // @[Plic.scala 344:61]
  wire [3:0] _T_82 = _T_80 ? _T_74 : _T_78; // @[Misc.scala 34:9]
  wire [1:0] _T_83 = _T_80 ? {{1'd0}, _T_75} : _T_81; // @[Misc.scala 34:36]
  wire  _T_84 = _T_70 >= _T_82; // @[Plic.scala 344:20]
  wire [2:0] _GEN_9 = {{1'd0}, _T_83}; // @[Plic.scala 344:61]
  wire [2:0] _T_85 = 3'h4 | _GEN_9; // @[Plic.scala 344:61]
  wire [3:0] _T_86 = _T_84 ? _T_70 : _T_82; // @[Misc.scala 34:9]
  wire [2:0] _T_87 = _T_84 ? {{1'd0}, _T_71} : _T_85; // @[Misc.scala 34:36]
  wire  _T_88 = effectivePriority_24 >= effectivePriority_25; // @[Plic.scala 344:20]
  wire [3:0] _T_90 = _T_88 ? effectivePriority_24 : effectivePriority_25; // @[Misc.scala 34:9]
  wire  _T_91 = _T_88 ? 1'h0 : 1'h1; // @[Misc.scala 34:36]
  wire  _T_92 = effectivePriority_26 >= effectivePriority_27; // @[Plic.scala 344:20]
  wire [3:0] _T_94 = _T_92 ? effectivePriority_26 : effectivePriority_27; // @[Misc.scala 34:9]
  wire  _T_95 = _T_92 ? 1'h0 : 1'h1; // @[Misc.scala 34:36]
  wire  _T_96 = _T_90 >= _T_94; // @[Plic.scala 344:20]
  wire [1:0] _GEN_10 = {{1'd0}, _T_95}; // @[Plic.scala 344:61]
  wire [1:0] _T_97 = 2'h2 | _GEN_10; // @[Plic.scala 344:61]
  wire [3:0] _T_98 = _T_96 ? _T_90 : _T_94; // @[Misc.scala 34:9]
  wire [1:0] _T_99 = _T_96 ? {{1'd0}, _T_91} : _T_97; // @[Misc.scala 34:36]
  wire  _T_100 = effectivePriority_28 >= effectivePriority_29; // @[Plic.scala 344:20]
  wire [3:0] _T_102 = _T_100 ? effectivePriority_28 : effectivePriority_29; // @[Misc.scala 34:9]
  wire  _T_103 = _T_100 ? 1'h0 : 1'h1; // @[Misc.scala 34:36]
  wire  _T_104 = effectivePriority_30 >= effectivePriority_31; // @[Plic.scala 344:20]
  wire [3:0] _T_106 = _T_104 ? effectivePriority_30 : effectivePriority_31; // @[Misc.scala 34:9]
  wire  _T_107 = _T_104 ? 1'h0 : 1'h1; // @[Misc.scala 34:36]
  wire  _T_108 = _T_102 >= _T_106; // @[Plic.scala 344:20]
  wire [1:0] _GEN_11 = {{1'd0}, _T_107}; // @[Plic.scala 344:61]
  wire [1:0] _T_109 = 2'h2 | _GEN_11; // @[Plic.scala 344:61]
  wire [3:0] _T_110 = _T_108 ? _T_102 : _T_106; // @[Misc.scala 34:9]
  wire [1:0] _T_111 = _T_108 ? {{1'd0}, _T_103} : _T_109; // @[Misc.scala 34:36]
  wire  _T_112 = _T_98 >= _T_110; // @[Plic.scala 344:20]
  wire [2:0] _GEN_12 = {{1'd0}, _T_111}; // @[Plic.scala 344:61]
  wire [2:0] _T_113 = 3'h4 | _GEN_12; // @[Plic.scala 344:61]
  wire [3:0] _T_114 = _T_112 ? _T_98 : _T_110; // @[Misc.scala 34:9]
  wire [2:0] _T_115 = _T_112 ? {{1'd0}, _T_99} : _T_113; // @[Misc.scala 34:36]
  wire  _T_116 = _T_86 >= _T_114; // @[Plic.scala 344:20]
  wire [3:0] _GEN_13 = {{1'd0}, _T_115}; // @[Plic.scala 344:61]
  wire [3:0] _T_117 = 4'h8 | _GEN_13; // @[Plic.scala 344:61]
  wire [3:0] _T_118 = _T_116 ? _T_86 : _T_114; // @[Misc.scala 34:9]
  wire [3:0] _T_119 = _T_116 ? {{1'd0}, _T_87} : _T_117; // @[Misc.scala 34:36]
  wire  _T_120 = _T_58 >= _T_118; // @[Plic.scala 344:20]
  wire [4:0] _GEN_14 = {{1'd0}, _T_119}; // @[Plic.scala 344:61]
  wire [4:0] _T_121 = 5'h10 | _GEN_14; // @[Plic.scala 344:61]
  wire [3:0] _T_122 = _T_120 ? _T_58 : _T_118; // @[Misc.scala 34:9]
  wire [4:0] _T_123 = _T_120 ? {{1'd0}, _T_59} : _T_121; // @[Misc.scala 34:36]
  wire  _T_124 = effectivePriority_32 >= effectivePriority_33; // @[Plic.scala 344:20]
  wire [3:0] _T_126 = _T_124 ? effectivePriority_32 : effectivePriority_33; // @[Misc.scala 34:9]
  wire  _T_127 = _T_124 ? 1'h0 : 1'h1; // @[Misc.scala 34:36]
  wire  _T_128 = effectivePriority_34 >= effectivePriority_35; // @[Plic.scala 344:20]
  wire [3:0] _T_130 = _T_128 ? effectivePriority_34 : effectivePriority_35; // @[Misc.scala 34:9]
  wire  _T_131 = _T_128 ? 1'h0 : 1'h1; // @[Misc.scala 34:36]
  wire  _T_132 = _T_126 >= _T_130; // @[Plic.scala 344:20]
  wire [1:0] _GEN_15 = {{1'd0}, _T_131}; // @[Plic.scala 344:61]
  wire [1:0] _T_133 = 2'h2 | _GEN_15; // @[Plic.scala 344:61]
  wire [3:0] _T_134 = _T_132 ? _T_126 : _T_130; // @[Misc.scala 34:9]
  wire [1:0] _T_135 = _T_132 ? {{1'd0}, _T_127} : _T_133; // @[Misc.scala 34:36]
  wire  _T_136 = effectivePriority_36 >= effectivePriority_37; // @[Plic.scala 344:20]
  wire [3:0] _T_138 = _T_136 ? effectivePriority_36 : effectivePriority_37; // @[Misc.scala 34:9]
  wire  _T_139 = _T_136 ? 1'h0 : 1'h1; // @[Misc.scala 34:36]
  wire  _T_140 = effectivePriority_38 >= effectivePriority_39; // @[Plic.scala 344:20]
  wire [3:0] _T_142 = _T_140 ? effectivePriority_38 : effectivePriority_39; // @[Misc.scala 34:9]
  wire  _T_143 = _T_140 ? 1'h0 : 1'h1; // @[Misc.scala 34:36]
  wire  _T_144 = _T_138 >= _T_142; // @[Plic.scala 344:20]
  wire [1:0] _GEN_16 = {{1'd0}, _T_143}; // @[Plic.scala 344:61]
  wire [1:0] _T_145 = 2'h2 | _GEN_16; // @[Plic.scala 344:61]
  wire [3:0] _T_146 = _T_144 ? _T_138 : _T_142; // @[Misc.scala 34:9]
  wire [1:0] _T_147 = _T_144 ? {{1'd0}, _T_139} : _T_145; // @[Misc.scala 34:36]
  wire  _T_148 = _T_134 >= _T_146; // @[Plic.scala 344:20]
  wire [2:0] _GEN_17 = {{1'd0}, _T_147}; // @[Plic.scala 344:61]
  wire [2:0] _T_149 = 3'h4 | _GEN_17; // @[Plic.scala 344:61]
  wire [3:0] _T_150 = _T_148 ? _T_134 : _T_146; // @[Misc.scala 34:9]
  wire [2:0] _T_151 = _T_148 ? {{1'd0}, _T_135} : _T_149; // @[Misc.scala 34:36]
  wire  _T_152 = effectivePriority_40 >= effectivePriority_41; // @[Plic.scala 344:20]
  wire [3:0] _T_154 = _T_152 ? effectivePriority_40 : effectivePriority_41; // @[Misc.scala 34:9]
  wire  _T_155 = _T_152 ? 1'h0 : 1'h1; // @[Misc.scala 34:36]
  wire  _T_156 = effectivePriority_42 >= effectivePriority_43; // @[Plic.scala 344:20]
  wire [3:0] _T_158 = _T_156 ? effectivePriority_42 : effectivePriority_43; // @[Misc.scala 34:9]
  wire  _T_159 = _T_156 ? 1'h0 : 1'h1; // @[Misc.scala 34:36]
  wire  _T_160 = _T_154 >= _T_158; // @[Plic.scala 344:20]
  wire [1:0] _GEN_18 = {{1'd0}, _T_159}; // @[Plic.scala 344:61]
  wire [1:0] _T_161 = 2'h2 | _GEN_18; // @[Plic.scala 344:61]
  wire [3:0] _T_162 = _T_160 ? _T_154 : _T_158; // @[Misc.scala 34:9]
  wire [1:0] _T_163 = _T_160 ? {{1'd0}, _T_155} : _T_161; // @[Misc.scala 34:36]
  wire  _T_164 = effectivePriority_44 >= effectivePriority_45; // @[Plic.scala 344:20]
  wire [3:0] _T_166 = _T_164 ? effectivePriority_44 : effectivePriority_45; // @[Misc.scala 34:9]
  wire  _T_167 = _T_164 ? 1'h0 : 1'h1; // @[Misc.scala 34:36]
  wire  _T_168 = effectivePriority_46 >= effectivePriority_47; // @[Plic.scala 344:20]
  wire [3:0] _T_170 = _T_168 ? effectivePriority_46 : effectivePriority_47; // @[Misc.scala 34:9]
  wire  _T_171 = _T_168 ? 1'h0 : 1'h1; // @[Misc.scala 34:36]
  wire  _T_172 = _T_166 >= _T_170; // @[Plic.scala 344:20]
  wire [1:0] _GEN_19 = {{1'd0}, _T_171}; // @[Plic.scala 344:61]
  wire [1:0] _T_173 = 2'h2 | _GEN_19; // @[Plic.scala 344:61]
  wire [3:0] _T_174 = _T_172 ? _T_166 : _T_170; // @[Misc.scala 34:9]
  wire [1:0] _T_175 = _T_172 ? {{1'd0}, _T_167} : _T_173; // @[Misc.scala 34:36]
  wire  _T_176 = _T_162 >= _T_174; // @[Plic.scala 344:20]
  wire [2:0] _GEN_20 = {{1'd0}, _T_175}; // @[Plic.scala 344:61]
  wire [2:0] _T_177 = 3'h4 | _GEN_20; // @[Plic.scala 344:61]
  wire [3:0] _T_178 = _T_176 ? _T_162 : _T_174; // @[Misc.scala 34:9]
  wire [2:0] _T_179 = _T_176 ? {{1'd0}, _T_163} : _T_177; // @[Misc.scala 34:36]
  wire  _T_180 = _T_150 >= _T_178; // @[Plic.scala 344:20]
  wire [3:0] _GEN_21 = {{1'd0}, _T_179}; // @[Plic.scala 344:61]
  wire [3:0] _T_181 = 4'h8 | _GEN_21; // @[Plic.scala 344:61]
  wire [3:0] _T_182 = _T_180 ? _T_150 : _T_178; // @[Misc.scala 34:9]
  wire [3:0] _T_183 = _T_180 ? {{1'd0}, _T_151} : _T_181; // @[Misc.scala 34:36]
  wire  _T_184 = effectivePriority_48 >= effectivePriority_49; // @[Plic.scala 344:20]
  wire [3:0] _T_186 = _T_184 ? effectivePriority_48 : effectivePriority_49; // @[Misc.scala 34:9]
  wire  _T_187 = _T_184 ? 1'h0 : 1'h1; // @[Misc.scala 34:36]
  wire  _T_188 = effectivePriority_50 >= effectivePriority_51; // @[Plic.scala 344:20]
  wire [3:0] _T_190 = _T_188 ? effectivePriority_50 : effectivePriority_51; // @[Misc.scala 34:9]
  wire  _T_191 = _T_188 ? 1'h0 : 1'h1; // @[Misc.scala 34:36]
  wire  _T_192 = _T_186 >= _T_190; // @[Plic.scala 344:20]
  wire [1:0] _GEN_22 = {{1'd0}, _T_191}; // @[Plic.scala 344:61]
  wire [1:0] _T_193 = 2'h2 | _GEN_22; // @[Plic.scala 344:61]
  wire [3:0] _T_194 = _T_192 ? _T_186 : _T_190; // @[Misc.scala 34:9]
  wire [1:0] _T_195 = _T_192 ? {{1'd0}, _T_187} : _T_193; // @[Misc.scala 34:36]
  wire  _T_196 = effectivePriority_52 >= effectivePriority_53; // @[Plic.scala 344:20]
  wire [3:0] _T_198 = _T_196 ? effectivePriority_52 : effectivePriority_53; // @[Misc.scala 34:9]
  wire  _T_199 = _T_196 ? 1'h0 : 1'h1; // @[Misc.scala 34:36]
  wire  _T_200 = effectivePriority_54 >= effectivePriority_55; // @[Plic.scala 344:20]
  wire [3:0] _T_202 = _T_200 ? effectivePriority_54 : effectivePriority_55; // @[Misc.scala 34:9]
  wire  _T_203 = _T_200 ? 1'h0 : 1'h1; // @[Misc.scala 34:36]
  wire  _T_204 = _T_198 >= _T_202; // @[Plic.scala 344:20]
  wire [1:0] _GEN_23 = {{1'd0}, _T_203}; // @[Plic.scala 344:61]
  wire [1:0] _T_205 = 2'h2 | _GEN_23; // @[Plic.scala 344:61]
  wire [3:0] _T_206 = _T_204 ? _T_198 : _T_202; // @[Misc.scala 34:9]
  wire [1:0] _T_207 = _T_204 ? {{1'd0}, _T_199} : _T_205; // @[Misc.scala 34:36]
  wire  _T_208 = _T_194 >= _T_206; // @[Plic.scala 344:20]
  wire [2:0] _GEN_24 = {{1'd0}, _T_207}; // @[Plic.scala 344:61]
  wire [2:0] _T_209 = 3'h4 | _GEN_24; // @[Plic.scala 344:61]
  wire [3:0] _T_210 = _T_208 ? _T_194 : _T_206; // @[Misc.scala 34:9]
  wire [2:0] _T_211 = _T_208 ? {{1'd0}, _T_195} : _T_209; // @[Misc.scala 34:36]
  wire  _T_212 = effectivePriority_56 >= effectivePriority_57; // @[Plic.scala 344:20]
  wire [3:0] _T_214 = _T_212 ? effectivePriority_56 : effectivePriority_57; // @[Misc.scala 34:9]
  wire  _T_215 = _T_212 ? 1'h0 : 1'h1; // @[Misc.scala 34:36]
  wire  _T_216 = effectivePriority_58 >= effectivePriority_59; // @[Plic.scala 344:20]
  wire [3:0] _T_218 = _T_216 ? effectivePriority_58 : effectivePriority_59; // @[Misc.scala 34:9]
  wire  _T_219 = _T_216 ? 1'h0 : 1'h1; // @[Misc.scala 34:36]
  wire  _T_220 = _T_214 >= _T_218; // @[Plic.scala 344:20]
  wire [1:0] _GEN_25 = {{1'd0}, _T_219}; // @[Plic.scala 344:61]
  wire [1:0] _T_221 = 2'h2 | _GEN_25; // @[Plic.scala 344:61]
  wire [3:0] _T_222 = _T_220 ? _T_214 : _T_218; // @[Misc.scala 34:9]
  wire [1:0] _T_223 = _T_220 ? {{1'd0}, _T_215} : _T_221; // @[Misc.scala 34:36]
  wire  _T_224 = effectivePriority_60 >= effectivePriority_61; // @[Plic.scala 344:20]
  wire [3:0] _T_226 = _T_224 ? effectivePriority_60 : effectivePriority_61; // @[Misc.scala 34:9]
  wire  _T_227 = _T_224 ? 1'h0 : 1'h1; // @[Misc.scala 34:36]
  wire  _T_228 = effectivePriority_62 >= effectivePriority_63; // @[Plic.scala 344:20]
  wire [3:0] _T_230 = _T_228 ? effectivePriority_62 : effectivePriority_63; // @[Misc.scala 34:9]
  wire  _T_231 = _T_228 ? 1'h0 : 1'h1; // @[Misc.scala 34:36]
  wire  _T_232 = _T_226 >= _T_230; // @[Plic.scala 344:20]
  wire [1:0] _GEN_26 = {{1'd0}, _T_231}; // @[Plic.scala 344:61]
  wire [1:0] _T_233 = 2'h2 | _GEN_26; // @[Plic.scala 344:61]
  wire [3:0] _T_234 = _T_232 ? _T_226 : _T_230; // @[Misc.scala 34:9]
  wire [1:0] _T_235 = _T_232 ? {{1'd0}, _T_227} : _T_233; // @[Misc.scala 34:36]
  wire  _T_236 = _T_222 >= _T_234; // @[Plic.scala 344:20]
  wire [2:0] _GEN_27 = {{1'd0}, _T_235}; // @[Plic.scala 344:61]
  wire [2:0] _T_237 = 3'h4 | _GEN_27; // @[Plic.scala 344:61]
  wire [3:0] _T_238 = _T_236 ? _T_222 : _T_234; // @[Misc.scala 34:9]
  wire [2:0] _T_239 = _T_236 ? {{1'd0}, _T_223} : _T_237; // @[Misc.scala 34:36]
  wire  _T_240 = _T_210 >= _T_238; // @[Plic.scala 344:20]
  wire [3:0] _GEN_28 = {{1'd0}, _T_239}; // @[Plic.scala 344:61]
  wire [3:0] _T_241 = 4'h8 | _GEN_28; // @[Plic.scala 344:61]
  wire [3:0] _T_242 = _T_240 ? _T_210 : _T_238; // @[Misc.scala 34:9]
  wire [3:0] _T_243 = _T_240 ? {{1'd0}, _T_211} : _T_241; // @[Misc.scala 34:36]
  wire  _T_244 = _T_182 >= _T_242; // @[Plic.scala 344:20]
  wire [4:0] _GEN_29 = {{1'd0}, _T_243}; // @[Plic.scala 344:61]
  wire [4:0] _T_245 = 5'h10 | _GEN_29; // @[Plic.scala 344:61]
  wire [3:0] _T_246 = _T_244 ? _T_182 : _T_242; // @[Misc.scala 34:9]
  wire [4:0] _T_247 = _T_244 ? {{1'd0}, _T_183} : _T_245; // @[Misc.scala 34:36]
  wire  _T_248 = _T_122 >= _T_246; // @[Plic.scala 344:20]
  wire [5:0] _GEN_30 = {{1'd0}, _T_247}; // @[Plic.scala 344:61]
  wire [5:0] _T_249 = 6'h20 | _GEN_30; // @[Plic.scala 344:61]
  wire [3:0] _T_250 = _T_248 ? _T_122 : _T_246; // @[Misc.scala 34:9]
  wire [5:0] _T_251 = _T_248 ? {{1'd0}, _T_123} : _T_249; // @[Misc.scala 34:36]
  wire  _T_252 = effectivePriority_64 >= effectivePriority_65; // @[Plic.scala 344:20]
  wire [3:0] _T_254 = _T_252 ? effectivePriority_64 : effectivePriority_65; // @[Misc.scala 34:9]
  wire  _T_255 = _T_252 ? 1'h0 : 1'h1; // @[Misc.scala 34:36]
  wire  _T_256 = _T_250 >= _T_254; // @[Plic.scala 344:20]
  wire [6:0] _GEN_31 = {{6'd0}, _T_255}; // @[Plic.scala 344:61]
  wire [6:0] _T_257 = 7'h40 | _GEN_31; // @[Plic.scala 344:61]
  wire [3:0] maxPri = _T_256 ? _T_250 : _T_254; // @[Misc.scala 34:9]
  assign io_dev = _T_256 ? {{1'd0}, _T_251} : _T_257; // @[Misc.scala 34:36]
  assign io_max = maxPri[2:0]; // @[Plic.scala 350:10]
endmodule

