module bosc_Frontend(
  input          clock,
  input          reset,
  input          auto_icache_client_out_a_ready,
  output         auto_icache_client_out_a_valid,
  output [2:0]   auto_icache_client_out_a_bits_opcode,
  output [2:0]   auto_icache_client_out_a_bits_size,
  output [1:0]   auto_icache_client_out_a_bits_source,
  output [35:0]  auto_icache_client_out_a_bits_address,
  output [31:0]  auto_icache_client_out_a_bits_mask,
  output         auto_icache_client_out_bready,
  input          auto_icache_client_out_bvalid,
  input  [1:0]   auto_icache_client_out_bparam,
  input  [35:0]  auto_icache_client_out_baddress,
  input  [255:0] auto_icache_client_out_bdata,
  input          auto_icache_client_out_c_ready,
  output         auto_icache_client_out_c_valid,
  output [2:0]   auto_icache_client_out_c_bits_opcode,
  output [2:0]   auto_icache_client_out_c_bits_param,
  output [35:0]  auto_icache_client_out_c_bits_address,
  output         auto_icache_client_out_c_bits_echo_blockisdirty,
  output [255:0] auto_icache_client_out_c_bits_data,
  output         auto_icache_client_out_d_ready,
  input          auto_icache_client_out_d_valid,
  input  [2:0]   auto_icache_client_out_d_bits_opcode,
  input  [1:0]   auto_icache_client_out_d_bits_param,
  input  [1:0]   auto_icache_client_out_d_bits_source,
  input  [3:0]   auto_icache_client_out_d_bits_sink,
  input          auto_icache_client_out_d_bits_echo_blockisdirty,
  input  [255:0] auto_icache_client_out_d_bits_data,
  input          auto_icache_client_out_d_bits_corrupt,
  input          auto_icache_client_out_e_ready,
  output         auto_icache_client_out_e_valid,
  output [3:0]   auto_icache_client_out_e_bits_sink,
  input          auto_instrUncache_client_out_a_ready,
  output         auto_instrUncache_client_out_a_valid,
  output [35:0]  auto_instrUncache_client_out_a_bits_address,
  output         auto_instrUncache_client_out_d_ready,
  input          auto_instrUncache_client_out_d_valid,
  input          auto_instrUncache_client_out_d_bits_source,
  input  [63:0]  auto_instrUncache_client_out_d_bits_data,
  input  [35:0]  io_reset_vector,
  input          io_ptw_req_0_ready,
  output         io_ptw_req_0_valid,
  output [26:0]  io_ptw_req_0_bits_vpn,
  input          io_ptw_req_1_ready,
  output         io_ptw_req_1_valid,
  output [26:0]  io_ptw_req_1_bits_vpn,
  input          io_ptw_req_3_ready,
  output         io_ptw_req_3_valid,
  output [26:0]  io_ptw_req_3_bits_vpn,
  input          io_ptw_resp_valid,
  input  [26:0]  io_ptw_resp_bits_data_entry_tag,
  input  [15:0]  io_ptw_resp_bits_data_entry_asid,
  input  [23:0]  io_ptw_resp_bits_data_entry_ppn,
  input          io_ptw_resp_bits_data_entry_perm_d,
  input          io_ptw_resp_bits_data_entry_perm_a,
  input          io_ptw_resp_bits_data_entry_perm_g,
  input          io_ptw_resp_bits_data_entry_perm_u,
  input          io_ptw_resp_bits_data_entry_perm_x,
  input          io_ptw_resp_bits_data_entry_perm_w,
  input          io_ptw_resp_bits_data_entry_perm_r,
  input  [1:0]   io_ptw_resp_bits_data_entry_level,
  input          io_ptw_resp_bits_data_pf,
  input          io_ptw_resp_bits_data_af,
  input          io_backend_cfVec_0_ready,
  output         io_backend_cfVec_0_valid,
  output [31:0]  io_backend_cfVec_0_bits_instr,
  output [9:0]   io_backend_cfVec_0_bits_foldpc,
  output         io_backend_cfVec_0_bits_exceptionVec_1,
  output         io_backend_cfVec_0_bits_exceptionVec_12,
  output         io_backend_cfVec_0_bits_trigger_frontendHit_0,
  output         io_backend_cfVec_0_bits_trigger_frontendHit_1,
  output         io_backend_cfVec_0_bits_trigger_frontendHit_2,
  output         io_backend_cfVec_0_bits_trigger_frontendHit_3,
  output         io_backend_cfVec_0_bits_trigger_backendEn_0,
  output         io_backend_cfVec_0_bits_trigger_backendEn_1,
  output         io_backend_cfVec_0_bits_pd_isRVC,
  output [1:0]   io_backend_cfVec_0_bits_pd_brType,
  output         io_backend_cfVec_0_bits_pd_isCall,
  output         io_backend_cfVec_0_bits_pd_isRet,
  output         io_backend_cfVec_0_bits_pred_taken,
  output         io_backend_cfVec_0_bits_crossPageIPFFix,
  output         io_backend_cfVec_0_bits_ftqPtr_flag,
  output [2:0]   io_backend_cfVec_0_bits_ftqPtr_value,
  output [2:0]   io_backend_cfVec_0_bits_ftqOffset,
  input          io_backend_cfVec_1_ready,
  output         io_backend_cfVec_1_valid,
  output [31:0]  io_backend_cfVec_1_bits_instr,
  output [9:0]   io_backend_cfVec_1_bits_foldpc,
  output         io_backend_cfVec_1_bits_exceptionVec_1,
  output         io_backend_cfVec_1_bits_exceptionVec_12,
  output         io_backend_cfVec_1_bits_trigger_frontendHit_0,
  output         io_backend_cfVec_1_bits_trigger_frontendHit_1,
  output         io_backend_cfVec_1_bits_trigger_frontendHit_2,
  output         io_backend_cfVec_1_bits_trigger_frontendHit_3,
  output         io_backend_cfVec_1_bits_trigger_backendEn_0,
  output         io_backend_cfVec_1_bits_trigger_backendEn_1,
  output         io_backend_cfVec_1_bits_pd_isRVC,
  output [1:0]   io_backend_cfVec_1_bits_pd_brType,
  output         io_backend_cfVec_1_bits_pd_isCall,
  output         io_backend_cfVec_1_bits_pd_isRet,
  output         io_backend_cfVec_1_bits_pred_taken,
  output         io_backend_cfVec_1_bits_crossPageIPFFix,
  output         io_backend_cfVec_1_bits_ftqPtr_flag,
  output [2:0]   io_backend_cfVec_1_bits_ftqPtr_value,
  output [2:0]   io_backend_cfVec_1_bits_ftqOffset,
  output         io_backend_fromFtq_pc_mem_wen,
  output [2:0]   io_backend_fromFtq_pc_mem_waddr,
  output [38:0]  io_backend_fromFtq_pc_mem_wdata_startAddr,
  output [38:0]  io_backend_fromFtq_pc_mem_wdata_nextLineAddr,
  output         io_backend_fromFtq_pc_mem_wdata_isNextMask_0,
  output         io_backend_fromFtq_pc_mem_wdata_isNextMask_1,
  output         io_backend_fromFtq_pc_mem_wdata_isNextMask_2,
  output         io_backend_fromFtq_pc_mem_wdata_isNextMask_3,
  output         io_backend_fromFtq_pc_mem_wdata_isNextMask_4,
  output         io_backend_fromFtq_pc_mem_wdata_isNextMask_5,
  output         io_backend_fromFtq_pc_mem_wdata_isNextMask_6,
  output         io_backend_fromFtq_pc_mem_wdata_isNextMask_7,
  output [38:0]  io_backend_fromFtq_newest_entry_target,
  output         io_backend_fromFtq_newest_entry_ptr_flag,
  output [2:0]   io_backend_fromFtq_newest_entry_ptr_value,
  input          io_backend_toFtq_rob_commits_0_valid,
  input  [2:0]   io_backend_toFtq_rob_commits_0_bits_commitType,
  input          io_backend_toFtq_rob_commits_0_bits_ftqIdx_flag,
  input  [2:0]   io_backend_toFtq_rob_commits_0_bits_ftqIdx_value,
  input  [2:0]   io_backend_toFtq_rob_commits_0_bits_ftqOffset,
  input          io_backend_toFtq_rob_commits_1_valid,
  input  [2:0]   io_backend_toFtq_rob_commits_1_bits_commitType,
  input          io_backend_toFtq_rob_commits_1_bits_ftqIdx_flag,
  input  [2:0]   io_backend_toFtq_rob_commits_1_bits_ftqIdx_value,
  input  [2:0]   io_backend_toFtq_rob_commits_1_bits_ftqOffset,
  input          io_backend_toFtq_redirect_valid,
  input          io_backend_toFtq_redirect_bits_ftqIdx_flag,
  input  [2:0]   io_backend_toFtq_redirect_bits_ftqIdx_value,
  input  [2:0]   io_backend_toFtq_redirect_bits_ftqOffset,
  input          io_backend_toFtq_redirect_bits_level,
  input  [38:0]  io_backend_toFtq_redirect_bits_cfiUpdate_pc,
  input          io_backend_toFtq_redirect_bits_cfiUpdate_pd_isRVC,
  input  [1:0]   io_backend_toFtq_redirect_bits_cfiUpdate_pd_brType,
  input          io_backend_toFtq_redirect_bits_cfiUpdate_pd_isCall,
  input          io_backend_toFtq_redirect_bits_cfiUpdate_pd_isRet,
  input  [38:0]  io_backend_toFtq_redirect_bits_cfiUpdate_target,
  input          io_backend_toFtq_redirect_bits_cfiUpdate_taken,
  input          io_backend_toFtq_redirect_bits_cfiUpdate_isMisPred,
  input          io_sfence_valid,
  input          io_sfence_bits_rs1,
  input          io_sfence_bits_rs2,
  input  [38:0]  io_sfence_bits_addr,
  input  [15:0]  io_sfence_bits_asid,
  input  [3:0]   io_tlbCsr_satp_mode,
  input  [15:0]  io_tlbCsr_satp_asid,
  input  [43:0]  io_tlbCsr_satp_ppn,
  input          io_tlbCsr_satp_changed,
  input          io_tlbCsr_priv_mxr,
  input          io_tlbCsr_priv_sum,
  input  [1:0]   io_tlbCsr_priv_imode,
  input  [1:0]   io_tlbCsr_priv_dmode,
  input          io_csrCtrl_icache_parity_enable,
  input          io_csrCtrl_lvpred_disable,
  input          io_csrCtrl_no_spec_load,
  input          io_csrCtrl_storeset_wait_store,
  input  [4:0]   io_csrCtrl_lvpred_timeout,
  input          io_csrCtrl_bp_ctrl_ubtb_enable,
  input          io_csrCtrl_bp_ctrl_btb_enable,
  input          io_csrCtrl_bp_ctrl_tage_enable,
  input          io_csrCtrl_bp_ctrl_sc_enable,
  input          io_csrCtrl_bp_ctrl_ras_enable,
  input  [3:0]   io_csrCtrl_sbuffer_threshold,
  input          io_csrCtrl_ldld_vio_check_enable,
  input          io_csrCtrl_cache_error_enable,
  input          io_csrCtrl_uncache_write_outstanding_enable,
  input          io_csrCtrl_fusion_enable,
  input          io_csrCtrl_wfi_enable,
  input          io_csrCtrl_svinval_enable,
  input          io_csrCtrl_distribute_csr_wvalid,
  input  [11:0]  io_csrCtrl_distribute_csr_waddr,
  input  [63:0]  io_csrCtrl_distribute_csr_wdata,
  input          io_csrCtrl_singlestep,
  input          io_csrCtrl_frontend_trigger_t_valid,
  input  [1:0]   io_csrCtrl_frontend_trigger_t_bits_addr,
  input  [1:0]   io_csrCtrl_frontend_trigger_t_bits_tdata_matchType,
  input          io_csrCtrl_frontend_trigger_t_bits_tdata_select,
  input          io_csrCtrl_frontend_trigger_t_bits_tdata_timing,
  input          io_csrCtrl_frontend_trigger_t_bits_tdata_chain,
  input  [63:0]  io_csrCtrl_frontend_trigger_t_bits_tdata_tdata2,
  input          io_csrCtrl_mem_trigger_t_valid,
  input  [2:0]   io_csrCtrl_mem_trigger_t_bits_addr,
  input  [1:0]   io_csrCtrl_mem_trigger_t_bits_tdata_matchType,
  input          io_csrCtrl_mem_trigger_t_bits_tdata_select,
  input          io_csrCtrl_mem_trigger_t_bits_tdata_chain,
  input  [63:0]  io_csrCtrl_mem_trigger_t_bits_tdata_tdata2,
  input          io_csrCtrl_trigger_enable_0,
  input          io_csrCtrl_trigger_enable_1,
  input          io_csrCtrl_trigger_enable_2,
  input          io_csrCtrl_trigger_enable_3,
  input          io_csrCtrl_trigger_enable_4,
  input          io_csrCtrl_trigger_enable_5,
  input          io_csrCtrl_trigger_enable_6,
  input          io_csrCtrl_trigger_enable_7,
  input          io_csrCtrl_trigger_enable_8,
  input          io_csrCtrl_trigger_enable_9,
  output         io_csrUpdate_wvalid,
  output [11:0]  io_csrUpdate_waddr,
  output [63:0]  io_csrUpdate_wdata,
  output [35:0]  io_error_paddr,
  output         io_error_report_to_beu,
  output [5:0]   io_perf_0_value,
  output [5:0]   io_perf_1_value,
  output [5:0]   io_perf_2_value,
  output [5:0]   io_perf_3_value,
  output [5:0]   io_perf_4_value,
  output [5:0]   io_perf_5_value,
  output [5:0]   io_perf_6_value,
  output [5:0]   io_perf_7_value
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
`endif // RANDOMIZE_REG_INIT
  wire  instrUncache_clock; // @[Frontend.scala 32:33]
  wire  instrUncache_reset; // @[Frontend.scala 32:33]
  wire  instrUncache_auto_client_out_a_ready; // @[Frontend.scala 32:33]
  wire  instrUncache_auto_client_out_a_valid; // @[Frontend.scala 32:33]
  wire [35:0] instrUncache_auto_client_out_a_bits_address; // @[Frontend.scala 32:33]
  wire  instrUncache_auto_client_out_d_ready; // @[Frontend.scala 32:33]
  wire  instrUncache_auto_client_out_d_valid; // @[Frontend.scala 32:33]
  wire  instrUncache_auto_client_out_d_bits_source; // @[Frontend.scala 32:33]
  wire [63:0] instrUncache_auto_client_out_d_bits_data; // @[Frontend.scala 32:33]
  wire  instrUncache_io_req_ready; // @[Frontend.scala 32:33]
  wire  instrUncache_io_req_valid; // @[Frontend.scala 32:33]
  wire [35:0] instrUncache_io_req_bits_addr; // @[Frontend.scala 32:33]
  wire  instrUncache_io_resp_valid; // @[Frontend.scala 32:33]
  wire [31:0] instrUncache_io_resp_bits_data; // @[Frontend.scala 32:33]
  wire  icache_clock; // @[Frontend.scala 33:33]
  wire  icache_reset; // @[Frontend.scala 33:33]
  wire  icache_auto_client_out_a_ready; // @[Frontend.scala 33:33]
  wire  icache_auto_client_out_a_valid; // @[Frontend.scala 33:33]
  wire [2:0] icache_auto_client_out_a_bits_opcode; // @[Frontend.scala 33:33]
  wire [2:0] icache_auto_client_out_a_bits_size; // @[Frontend.scala 33:33]
  wire [1:0] icache_auto_client_out_a_bits_source; // @[Frontend.scala 33:33]
  wire [35:0] icache_auto_client_out_a_bits_address; // @[Frontend.scala 33:33]
  wire [31:0] icache_auto_client_out_a_bits_mask; // @[Frontend.scala 33:33]
  wire  icache_auto_client_out_bready; // @[Frontend.scala 33:33]
  wire  icache_auto_client_out_bvalid; // @[Frontend.scala 33:33]
  wire [1:0] icache_auto_client_out_bparam; // @[Frontend.scala 33:33]
  wire [35:0] icache_auto_client_out_baddress; // @[Frontend.scala 33:33]
  wire [255:0] icache_auto_client_out_bdata; // @[Frontend.scala 33:33]
  wire  icache_auto_client_out_c_ready; // @[Frontend.scala 33:33]
  wire  icache_auto_client_out_c_valid; // @[Frontend.scala 33:33]
  wire [2:0] icache_auto_client_out_c_bits_opcode; // @[Frontend.scala 33:33]
  wire [2:0] icache_auto_client_out_c_bits_param; // @[Frontend.scala 33:33]
  wire [35:0] icache_auto_client_out_c_bits_address; // @[Frontend.scala 33:33]
  wire  icache_auto_client_out_c_bits_echo_blockisdirty; // @[Frontend.scala 33:33]
  wire [255:0] icache_auto_client_out_c_bits_data; // @[Frontend.scala 33:33]
  wire  icache_auto_client_out_d_ready; // @[Frontend.scala 33:33]
  wire  icache_auto_client_out_d_valid; // @[Frontend.scala 33:33]
  wire [2:0] icache_auto_client_out_d_bits_opcode; // @[Frontend.scala 33:33]
  wire [1:0] icache_auto_client_out_d_bits_param; // @[Frontend.scala 33:33]
  wire [1:0] icache_auto_client_out_d_bits_source; // @[Frontend.scala 33:33]
  wire [3:0] icache_auto_client_out_d_bits_sink; // @[Frontend.scala 33:33]
  wire  icache_auto_client_out_d_bits_echo_blockisdirty; // @[Frontend.scala 33:33]
  wire [255:0] icache_auto_client_out_d_bits_data; // @[Frontend.scala 33:33]
  wire  icache_auto_client_out_d_bits_corrupt; // @[Frontend.scala 33:33]
  wire  icache_auto_client_out_e_ready; // @[Frontend.scala 33:33]
  wire  icache_auto_client_out_e_valid; // @[Frontend.scala 33:33]
  wire [3:0] icache_auto_client_out_e_bits_sink; // @[Frontend.scala 33:33]
  wire  icache_io_stop; // @[Frontend.scala 33:33]
  wire  icache_io_fetch_req_ready; // @[Frontend.scala 33:33]
  wire  icache_io_fetch_req_valid; // @[Frontend.scala 33:33]
  wire [38:0] icache_io_fetch_req_bits_pcMemRead_0_startAddr; // @[Frontend.scala 33:33]
  wire [38:0] icache_io_fetch_req_bits_pcMemRead_0_nextlineStart; // @[Frontend.scala 33:33]
  wire [38:0] icache_io_fetch_req_bits_pcMemRead_1_startAddr; // @[Frontend.scala 33:33]
  wire [38:0] icache_io_fetch_req_bits_pcMemRead_1_nextlineStart; // @[Frontend.scala 33:33]
  wire [38:0] icache_io_fetch_req_bits_pcMemRead_2_startAddr; // @[Frontend.scala 33:33]
  wire [38:0] icache_io_fetch_req_bits_pcMemRead_2_nextlineStart; // @[Frontend.scala 33:33]
  wire [38:0] icache_io_fetch_req_bits_pcMemRead_3_startAddr; // @[Frontend.scala 33:33]
  wire [38:0] icache_io_fetch_req_bits_pcMemRead_3_nextlineStart; // @[Frontend.scala 33:33]
  wire [38:0] icache_io_fetch_req_bits_pcMemRead_4_startAddr; // @[Frontend.scala 33:33]
  wire [38:0] icache_io_fetch_req_bits_pcMemRead_4_nextlineStart; // @[Frontend.scala 33:33]
  wire  icache_io_fetch_req_bits_readValid_0; // @[Frontend.scala 33:33]
  wire  icache_io_fetch_req_bits_readValid_1; // @[Frontend.scala 33:33]
  wire  icache_io_fetch_req_bits_readValid_2; // @[Frontend.scala 33:33]
  wire  icache_io_fetch_req_bits_readValid_3; // @[Frontend.scala 33:33]
  wire  icache_io_fetch_req_bits_readValid_4; // @[Frontend.scala 33:33]
  wire  icache_io_fetch_resp_0_valid; // @[Frontend.scala 33:33]
  wire [38:0] icache_io_fetch_resp_0_bits_vaddr; // @[Frontend.scala 33:33]
  wire [511:0] icache_io_fetch_resp_0_bits_registerData; // @[Frontend.scala 33:33]
  wire [511:0] icache_io_fetch_resp_0_bits_sramData; // @[Frontend.scala 33:33]
  wire  icache_io_fetch_resp_0_bits_select; // @[Frontend.scala 33:33]
  wire [35:0] icache_io_fetch_resp_0_bits_paddr; // @[Frontend.scala 33:33]
  wire  icache_io_fetch_resp_0_bits_tlbExcp_pageFault; // @[Frontend.scala 33:33]
  wire  icache_io_fetch_resp_0_bits_tlbExcp_accessFault; // @[Frontend.scala 33:33]
  wire  icache_io_fetch_resp_0_bits_tlbExcp_mmio; // @[Frontend.scala 33:33]
  wire  icache_io_fetch_resp_1_valid; // @[Frontend.scala 33:33]
  wire [38:0] icache_io_fetch_resp_1_bits_vaddr; // @[Frontend.scala 33:33]
  wire [511:0] icache_io_fetch_resp_1_bits_registerData; // @[Frontend.scala 33:33]
  wire [511:0] icache_io_fetch_resp_1_bits_sramData; // @[Frontend.scala 33:33]
  wire  icache_io_fetch_resp_1_bits_select; // @[Frontend.scala 33:33]
  wire  icache_io_fetch_resp_1_bits_tlbExcp_pageFault; // @[Frontend.scala 33:33]
  wire  icache_io_fetch_resp_1_bits_tlbExcp_accessFault; // @[Frontend.scala 33:33]
  wire  icache_io_toIFU; // @[Frontend.scala 33:33]
  wire [35:0] icache_io_pmp_0_req_bits_addr; // @[Frontend.scala 33:33]
  wire  icache_io_pmp_0_resp_instr; // @[Frontend.scala 33:33]
  wire  icache_io_pmp_0_resp_mmio; // @[Frontend.scala 33:33]
  wire [35:0] icache_io_pmp_1_req_bits_addr; // @[Frontend.scala 33:33]
  wire  icache_io_pmp_1_resp_instr; // @[Frontend.scala 33:33]
  wire  icache_io_itlb_0_req_ready; // @[Frontend.scala 33:33]
  wire  icache_io_itlb_0_req_valid; // @[Frontend.scala 33:33]
  wire [38:0] icache_io_itlb_0_req_bits_vaddr; // @[Frontend.scala 33:33]
  wire  icache_io_itlb_0_req_bits_kill; // @[Frontend.scala 33:33]
  wire  icache_io_itlb_0_resp_ready; // @[Frontend.scala 33:33]
  wire  icache_io_itlb_0_resp_valid; // @[Frontend.scala 33:33]
  wire [35:0] icache_io_itlb_0_resp_bits_paddr_0; // @[Frontend.scala 33:33]
  wire  icache_io_itlb_0_resp_bits_excp_0_pf_instr; // @[Frontend.scala 33:33]
  wire  icache_io_itlb_0_resp_bits_excp_0_af_instr; // @[Frontend.scala 33:33]
  wire  icache_io_itlb_1_req_ready; // @[Frontend.scala 33:33]
  wire  icache_io_itlb_1_req_valid; // @[Frontend.scala 33:33]
  wire [38:0] icache_io_itlb_1_req_bits_vaddr; // @[Frontend.scala 33:33]
  wire  icache_io_itlb_1_req_bits_kill; // @[Frontend.scala 33:33]
  wire  icache_io_itlb_1_resp_ready; // @[Frontend.scala 33:33]
  wire  icache_io_itlb_1_resp_valid; // @[Frontend.scala 33:33]
  wire [35:0] icache_io_itlb_1_resp_bits_paddr_0; // @[Frontend.scala 33:33]
  wire  icache_io_itlb_1_resp_bits_excp_0_pf_instr; // @[Frontend.scala 33:33]
  wire  icache_io_itlb_1_resp_bits_excp_0_af_instr; // @[Frontend.scala 33:33]
  wire  icache_io_perfInfo_only_0_hit; // @[Frontend.scala 33:33]
  wire  icache_io_perfInfo_only_0_miss; // @[Frontend.scala 33:33]
  wire  icache_io_perfInfo_hit_0_hit_1; // @[Frontend.scala 33:33]
  wire  icache_io_perfInfo_hit_0_miss_1; // @[Frontend.scala 33:33]
  wire  icache_io_perfInfo_miss_0_hit_1; // @[Frontend.scala 33:33]
  wire  icache_io_perfInfo_miss_0_miss_1; // @[Frontend.scala 33:33]
  wire  icache_io_perfInfo_hit_0_except_1; // @[Frontend.scala 33:33]
  wire  icache_io_perfInfo_miss_0_except_1; // @[Frontend.scala 33:33]
  wire  icache_io_perfInfo_except_0; // @[Frontend.scala 33:33]
  wire  icache_io_perfInfo_bank_hit_1; // @[Frontend.scala 33:33]
  wire  icache_io_perfInfo_hit; // @[Frontend.scala 33:33]
  wire  icache_io_error_source_tag; // @[Frontend.scala 33:33]
  wire  icache_io_error_source_data; // @[Frontend.scala 33:33]
  wire  icache_io_error_source_l2; // @[Frontend.scala 33:33]
  wire  icache_io_error_opType_fetch; // @[Frontend.scala 33:33]
  wire  icache_io_error_opType_load; // @[Frontend.scala 33:33]
  wire  icache_io_error_opType_store; // @[Frontend.scala 33:33]
  wire  icache_io_error_opType_probe; // @[Frontend.scala 33:33]
  wire  icache_io_error_opType_release; // @[Frontend.scala 33:33]
  wire  icache_io_error_opType_atom; // @[Frontend.scala 33:33]
  wire [35:0] icache_io_error_paddr; // @[Frontend.scala 33:33]
  wire  icache_io_error_report_to_beu; // @[Frontend.scala 33:33]
  wire  icache_io_error_valid; // @[Frontend.scala 33:33]
  wire  icache_io_csr_distribute_csr_wvalid; // @[Frontend.scala 33:33]
  wire [11:0] icache_io_csr_distribute_csr_waddr; // @[Frontend.scala 33:33]
  wire [63:0] icache_io_csr_distribute_csr_wdata; // @[Frontend.scala 33:33]
  wire  icache_io_csr_update_wvalid; // @[Frontend.scala 33:33]
  wire [11:0] icache_io_csr_update_waddr; // @[Frontend.scala 33:33]
  wire [63:0] icache_io_csr_update_wdata; // @[Frontend.scala 33:33]
  wire  icache_io_csr_parity_enable; // @[Frontend.scala 33:33]
  wire  bpu_clock; // @[Frontend.scala 66:23]
  wire  bpu_reset; // @[Frontend.scala 66:23]
  wire  bpu_io_bpu_to_ftq_resp_ready; // @[Frontend.scala 66:23]
  wire  bpu_io_bpu_to_ftq_resp_valid; // @[Frontend.scala 66:23]
  wire [38:0] bpu_io_bpu_to_ftq_resp_bits_s1_pc; // @[Frontend.scala 66:23]
  wire  bpu_io_bpu_to_ftq_resp_bits_s1_full_pred_br_taken_mask_0; // @[Frontend.scala 66:23]
  wire  bpu_io_bpu_to_ftq_resp_bits_s1_full_pred_br_taken_mask_1; // @[Frontend.scala 66:23]
  wire  bpu_io_bpu_to_ftq_resp_bits_s1_full_pred_slot_valids_0; // @[Frontend.scala 66:23]
  wire  bpu_io_bpu_to_ftq_resp_bits_s1_full_pred_slot_valids_1; // @[Frontend.scala 66:23]
  wire [38:0] bpu_io_bpu_to_ftq_resp_bits_s1_full_pred_targets_0; // @[Frontend.scala 66:23]
  wire [38:0] bpu_io_bpu_to_ftq_resp_bits_s1_full_pred_targets_1; // @[Frontend.scala 66:23]
  wire [2:0] bpu_io_bpu_to_ftq_resp_bits_s1_full_pred_offsets_0; // @[Frontend.scala 66:23]
  wire [2:0] bpu_io_bpu_to_ftq_resp_bits_s1_full_pred_offsets_1; // @[Frontend.scala 66:23]
  wire [38:0] bpu_io_bpu_to_ftq_resp_bits_s1_full_pred_fallThroughAddr; // @[Frontend.scala 66:23]
  wire  bpu_io_bpu_to_ftq_resp_bits_s1_full_pred_fallThroughErr; // @[Frontend.scala 66:23]
  wire  bpu_io_bpu_to_ftq_resp_bits_s1_full_pred_is_br_sharing; // @[Frontend.scala 66:23]
  wire  bpu_io_bpu_to_ftq_resp_bits_s1_full_pred_hit; // @[Frontend.scala 66:23]
  wire [38:0] bpu_io_bpu_to_ftq_resp_bits_s2_pc; // @[Frontend.scala 66:23]
  wire  bpu_io_bpu_to_ftq_resp_bits_s2_valid; // @[Frontend.scala 66:23]
  wire  bpu_io_bpu_to_ftq_resp_bits_s2_hasRedirect; // @[Frontend.scala 66:23]
  wire  bpu_io_bpu_to_ftq_resp_bits_s2_ftq_idx_flag; // @[Frontend.scala 66:23]
  wire [2:0] bpu_io_bpu_to_ftq_resp_bits_s2_ftq_idx_value; // @[Frontend.scala 66:23]
  wire  bpu_io_bpu_to_ftq_resp_bits_s2_full_pred_br_taken_mask_0; // @[Frontend.scala 66:23]
  wire  bpu_io_bpu_to_ftq_resp_bits_s2_full_pred_br_taken_mask_1; // @[Frontend.scala 66:23]
  wire  bpu_io_bpu_to_ftq_resp_bits_s2_full_pred_slot_valids_0; // @[Frontend.scala 66:23]
  wire  bpu_io_bpu_to_ftq_resp_bits_s2_full_pred_slot_valids_1; // @[Frontend.scala 66:23]
  wire [38:0] bpu_io_bpu_to_ftq_resp_bits_s2_full_pred_targets_0; // @[Frontend.scala 66:23]
  wire [38:0] bpu_io_bpu_to_ftq_resp_bits_s2_full_pred_targets_1; // @[Frontend.scala 66:23]
  wire [2:0] bpu_io_bpu_to_ftq_resp_bits_s2_full_pred_offsets_0; // @[Frontend.scala 66:23]
  wire [2:0] bpu_io_bpu_to_ftq_resp_bits_s2_full_pred_offsets_1; // @[Frontend.scala 66:23]
  wire [38:0] bpu_io_bpu_to_ftq_resp_bits_s2_full_pred_fallThroughAddr; // @[Frontend.scala 66:23]
  wire  bpu_io_bpu_to_ftq_resp_bits_s2_full_pred_fallThroughErr; // @[Frontend.scala 66:23]
  wire  bpu_io_bpu_to_ftq_resp_bits_s2_full_pred_is_br_sharing; // @[Frontend.scala 66:23]
  wire  bpu_io_bpu_to_ftq_resp_bits_s2_full_pred_hit; // @[Frontend.scala 66:23]
  wire [38:0] bpu_io_bpu_to_ftq_resp_bits_s3_pc; // @[Frontend.scala 66:23]
  wire  bpu_io_bpu_to_ftq_resp_bits_s3_valid; // @[Frontend.scala 66:23]
  wire  bpu_io_bpu_to_ftq_resp_bits_s3_hasRedirect; // @[Frontend.scala 66:23]
  wire  bpu_io_bpu_to_ftq_resp_bits_s3_ftq_idx_flag; // @[Frontend.scala 66:23]
  wire [2:0] bpu_io_bpu_to_ftq_resp_bits_s3_ftq_idx_value; // @[Frontend.scala 66:23]
  wire  bpu_io_bpu_to_ftq_resp_bits_s3_full_pred_br_taken_mask_0; // @[Frontend.scala 66:23]
  wire  bpu_io_bpu_to_ftq_resp_bits_s3_full_pred_br_taken_mask_1; // @[Frontend.scala 66:23]
  wire  bpu_io_bpu_to_ftq_resp_bits_s3_full_pred_slot_valids_0; // @[Frontend.scala 66:23]
  wire  bpu_io_bpu_to_ftq_resp_bits_s3_full_pred_slot_valids_1; // @[Frontend.scala 66:23]
  wire [38:0] bpu_io_bpu_to_ftq_resp_bits_s3_full_pred_targets_0; // @[Frontend.scala 66:23]
  wire [38:0] bpu_io_bpu_to_ftq_resp_bits_s3_full_pred_targets_1; // @[Frontend.scala 66:23]
  wire [2:0] bpu_io_bpu_to_ftq_resp_bits_s3_full_pred_offsets_0; // @[Frontend.scala 66:23]
  wire [2:0] bpu_io_bpu_to_ftq_resp_bits_s3_full_pred_offsets_1; // @[Frontend.scala 66:23]
  wire [38:0] bpu_io_bpu_to_ftq_resp_bits_s3_full_pred_fallThroughAddr; // @[Frontend.scala 66:23]
  wire  bpu_io_bpu_to_ftq_resp_bits_s3_full_pred_fallThroughErr; // @[Frontend.scala 66:23]
  wire  bpu_io_bpu_to_ftq_resp_bits_s3_full_pred_is_br_sharing; // @[Frontend.scala 66:23]
  wire  bpu_io_bpu_to_ftq_resp_bits_s3_full_pred_hit; // @[Frontend.scala 66:23]
  wire [255:0] bpu_io_bpu_to_ftq_resp_bits_last_stage_meta; // @[Frontend.scala 66:23]
  wire [7:0] bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_17_folded_hist; // @[Frontend.scala 66:23]
  wire [7:0] bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_16_folded_hist; // @[Frontend.scala 66:23]
  wire [10:0] bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_15_folded_hist; // @[Frontend.scala 66:23]
  wire [6:0] bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_14_folded_hist; // @[Frontend.scala 66:23]
  wire [6:0] bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_13_folded_hist; // @[Frontend.scala 66:23]
  wire [6:0] bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_12_folded_hist; // @[Frontend.scala 66:23]
  wire [7:0] bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_11_folded_hist; // @[Frontend.scala 66:23]
  wire [8:0] bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_10_folded_hist; // @[Frontend.scala 66:23]
  wire [6:0] bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_9_folded_hist; // @[Frontend.scala 66:23]
  wire [7:0] bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_8_folded_hist; // @[Frontend.scala 66:23]
  wire [8:0] bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_7_folded_hist; // @[Frontend.scala 66:23]
  wire [8:0] bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_6_folded_hist; // @[Frontend.scala 66:23]
  wire [10:0] bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_5_folded_hist; // @[Frontend.scala 66:23]
  wire [3:0] bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_4_folded_hist; // @[Frontend.scala 66:23]
  wire [10:0] bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_3_folded_hist; // @[Frontend.scala 66:23]
  wire [7:0] bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_2_folded_hist; // @[Frontend.scala 66:23]
  wire [7:0] bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_1_folded_hist; // @[Frontend.scala 66:23]
  wire [7:0] bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_0_folded_hist; // @[Frontend.scala 66:23]
  wire  bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_5_bits_0; // @[Frontend.scala 66:23]
  wire  bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_5_bits_1; // @[Frontend.scala 66:23]
  wire  bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_5_bits_2; // @[Frontend.scala 66:23]
  wire  bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_5_bits_3; // @[Frontend.scala 66:23]
  wire  bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_4_bits_0; // @[Frontend.scala 66:23]
  wire  bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_4_bits_1; // @[Frontend.scala 66:23]
  wire  bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_4_bits_2; // @[Frontend.scala 66:23]
  wire  bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_4_bits_3; // @[Frontend.scala 66:23]
  wire  bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_3_bits_0; // @[Frontend.scala 66:23]
  wire  bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_3_bits_1; // @[Frontend.scala 66:23]
  wire  bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_3_bits_2; // @[Frontend.scala 66:23]
  wire  bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_3_bits_3; // @[Frontend.scala 66:23]
  wire  bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_2_bits_0; // @[Frontend.scala 66:23]
  wire  bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_2_bits_1; // @[Frontend.scala 66:23]
  wire  bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_2_bits_2; // @[Frontend.scala 66:23]
  wire  bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_2_bits_3; // @[Frontend.scala 66:23]
  wire  bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_1_bits_0; // @[Frontend.scala 66:23]
  wire  bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_1_bits_1; // @[Frontend.scala 66:23]
  wire  bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_1_bits_2; // @[Frontend.scala 66:23]
  wire  bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_1_bits_3; // @[Frontend.scala 66:23]
  wire  bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_0_bits_0; // @[Frontend.scala 66:23]
  wire  bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_0_bits_1; // @[Frontend.scala 66:23]
  wire  bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_0_bits_2; // @[Frontend.scala 66:23]
  wire  bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_0_bits_3; // @[Frontend.scala 66:23]
  wire [2:0] bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_lastBrNumOH; // @[Frontend.scala 66:23]
  wire  bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_histPtr_flag; // @[Frontend.scala 66:23]
  wire [7:0] bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_histPtr_value; // @[Frontend.scala 66:23]
  wire [4:0] bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_rasSp; // @[Frontend.scala 66:23]
  wire [38:0] bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_rasTop_retAddr; // @[Frontend.scala 66:23]
  wire [7:0] bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_rasTop_ctr; // @[Frontend.scala 66:23]
  wire  bpu_io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_valid; // @[Frontend.scala 66:23]
  wire [2:0] bpu_io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_brSlots_0_offset; // @[Frontend.scala 66:23]
  wire [11:0] bpu_io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_brSlots_0_lower; // @[Frontend.scala 66:23]
  wire [1:0] bpu_io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_brSlots_0_tarStat; // @[Frontend.scala 66:23]
  wire  bpu_io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_brSlots_0_sharing; // @[Frontend.scala 66:23]
  wire  bpu_io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_brSlots_0_valid; // @[Frontend.scala 66:23]
  wire [2:0] bpu_io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_tailSlot_offset; // @[Frontend.scala 66:23]
  wire [19:0] bpu_io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_tailSlot_lower; // @[Frontend.scala 66:23]
  wire [1:0] bpu_io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_tailSlot_tarStat; // @[Frontend.scala 66:23]
  wire  bpu_io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_tailSlot_sharing; // @[Frontend.scala 66:23]
  wire  bpu_io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_tailSlot_valid; // @[Frontend.scala 66:23]
  wire [2:0] bpu_io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_pftAddr; // @[Frontend.scala 66:23]
  wire  bpu_io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_carry; // @[Frontend.scala 66:23]
  wire  bpu_io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_isCall; // @[Frontend.scala 66:23]
  wire  bpu_io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_isRet; // @[Frontend.scala 66:23]
  wire  bpu_io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_isJalr; // @[Frontend.scala 66:23]
  wire  bpu_io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_last_may_be_rvi_call; // @[Frontend.scala 66:23]
  wire  bpu_io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_always_taken_0; // @[Frontend.scala 66:23]
  wire  bpu_io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_always_taken_1; // @[Frontend.scala 66:23]
  wire  bpu_io_ftq_to_bpu_redirect_valid; // @[Frontend.scala 66:23]
  wire  bpu_io_ftq_to_bpu_redirect_bits_level; // @[Frontend.scala 66:23]
  wire [38:0] bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_pc; // @[Frontend.scala 66:23]
  wire  bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_pd_isRVC; // @[Frontend.scala 66:23]
  wire  bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_pd_isCall; // @[Frontend.scala 66:23]
  wire  bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_pd_isRet; // @[Frontend.scala 66:23]
  wire [4:0] bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_rasSp; // @[Frontend.scala 66:23]
  wire [38:0] bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_rasEntry_retAddr; // @[Frontend.scala 66:23]
  wire [7:0] bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_rasEntry_ctr; // @[Frontend.scala 66:23]
  wire [7:0] bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_17_folded_hist; // @[Frontend.scala 66:23]
  wire [7:0] bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_16_folded_hist; // @[Frontend.scala 66:23]
  wire [10:0] bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_15_folded_hist; // @[Frontend.scala 66:23]
  wire [6:0] bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_14_folded_hist; // @[Frontend.scala 66:23]
  wire [6:0] bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_13_folded_hist; // @[Frontend.scala 66:23]
  wire [6:0] bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_12_folded_hist; // @[Frontend.scala 66:23]
  wire [7:0] bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_11_folded_hist; // @[Frontend.scala 66:23]
  wire [8:0] bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_10_folded_hist; // @[Frontend.scala 66:23]
  wire [6:0] bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_9_folded_hist; // @[Frontend.scala 66:23]
  wire [7:0] bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_8_folded_hist; // @[Frontend.scala 66:23]
  wire [8:0] bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_7_folded_hist; // @[Frontend.scala 66:23]
  wire [8:0] bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_6_folded_hist; // @[Frontend.scala 66:23]
  wire [10:0] bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_5_folded_hist; // @[Frontend.scala 66:23]
  wire [3:0] bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_4_folded_hist; // @[Frontend.scala 66:23]
  wire [10:0] bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_3_folded_hist; // @[Frontend.scala 66:23]
  wire [7:0] bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_2_folded_hist; // @[Frontend.scala 66:23]
  wire [7:0] bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_1_folded_hist; // @[Frontend.scala 66:23]
  wire [7:0] bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_0_folded_hist; // @[Frontend.scala 66:23]
  wire  bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_5_bits_0; // @[Frontend.scala 66:23]
  wire  bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_5_bits_1; // @[Frontend.scala 66:23]
  wire  bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_5_bits_2; // @[Frontend.scala 66:23]
  wire  bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_5_bits_3; // @[Frontend.scala 66:23]
  wire  bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_4_bits_0; // @[Frontend.scala 66:23]
  wire  bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_4_bits_1; // @[Frontend.scala 66:23]
  wire  bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_4_bits_2; // @[Frontend.scala 66:23]
  wire  bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_3_bits_0; // @[Frontend.scala 66:23]
  wire  bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_3_bits_1; // @[Frontend.scala 66:23]
  wire  bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_3_bits_2; // @[Frontend.scala 66:23]
  wire  bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_3_bits_3; // @[Frontend.scala 66:23]
  wire  bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_2_bits_0; // @[Frontend.scala 66:23]
  wire  bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_2_bits_1; // @[Frontend.scala 66:23]
  wire  bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_2_bits_2; // @[Frontend.scala 66:23]
  wire  bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_2_bits_3; // @[Frontend.scala 66:23]
  wire  bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_1_bits_0; // @[Frontend.scala 66:23]
  wire  bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_1_bits_1; // @[Frontend.scala 66:23]
  wire  bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_1_bits_2; // @[Frontend.scala 66:23]
  wire  bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_1_bits_3; // @[Frontend.scala 66:23]
  wire  bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_0_bits_0; // @[Frontend.scala 66:23]
  wire  bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_0_bits_1; // @[Frontend.scala 66:23]
  wire  bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_0_bits_2; // @[Frontend.scala 66:23]
  wire  bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_0_bits_3; // @[Frontend.scala 66:23]
  wire [2:0] bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_lastBrNumOH; // @[Frontend.scala 66:23]
  wire  bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_histPtr_flag; // @[Frontend.scala 66:23]
  wire [7:0] bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_histPtr_value; // @[Frontend.scala 66:23]
  wire [38:0] bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_target; // @[Frontend.scala 66:23]
  wire  bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_taken; // @[Frontend.scala 66:23]
  wire [1:0] bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_shift; // @[Frontend.scala 66:23]
  wire  bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_addIntoHist; // @[Frontend.scala 66:23]
  wire  bpu_io_ftq_to_bpu_update_valid; // @[Frontend.scala 66:23]
  wire [38:0] bpu_io_ftq_to_bpu_update_bits_pc; // @[Frontend.scala 66:23]
  wire [7:0] bpu_io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_17_folded_hist; // @[Frontend.scala 66:23]
  wire [7:0] bpu_io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_16_folded_hist; // @[Frontend.scala 66:23]
  wire [10:0] bpu_io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_15_folded_hist; // @[Frontend.scala 66:23]
  wire [6:0] bpu_io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_14_folded_hist; // @[Frontend.scala 66:23]
  wire [6:0] bpu_io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_13_folded_hist; // @[Frontend.scala 66:23]
  wire [6:0] bpu_io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_12_folded_hist; // @[Frontend.scala 66:23]
  wire [8:0] bpu_io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_10_folded_hist; // @[Frontend.scala 66:23]
  wire [6:0] bpu_io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_9_folded_hist; // @[Frontend.scala 66:23]
  wire [7:0] bpu_io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_8_folded_hist; // @[Frontend.scala 66:23]
  wire [8:0] bpu_io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_7_folded_hist; // @[Frontend.scala 66:23]
  wire [8:0] bpu_io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_6_folded_hist; // @[Frontend.scala 66:23]
  wire [10:0] bpu_io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_5_folded_hist; // @[Frontend.scala 66:23]
  wire [3:0] bpu_io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_4_folded_hist; // @[Frontend.scala 66:23]
  wire [10:0] bpu_io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_3_folded_hist; // @[Frontend.scala 66:23]
  wire [7:0] bpu_io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_2_folded_hist; // @[Frontend.scala 66:23]
  wire [7:0] bpu_io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_1_folded_hist; // @[Frontend.scala 66:23]
  wire [7:0] bpu_io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_0_folded_hist; // @[Frontend.scala 66:23]
  wire  bpu_io_ftq_to_bpu_update_bits_ftb_entry_valid; // @[Frontend.scala 66:23]
  wire [2:0] bpu_io_ftq_to_bpu_update_bits_ftb_entry_brSlots_0_offset; // @[Frontend.scala 66:23]
  wire [11:0] bpu_io_ftq_to_bpu_update_bits_ftb_entry_brSlots_0_lower; // @[Frontend.scala 66:23]
  wire [1:0] bpu_io_ftq_to_bpu_update_bits_ftb_entry_brSlots_0_tarStat; // @[Frontend.scala 66:23]
  wire  bpu_io_ftq_to_bpu_update_bits_ftb_entry_brSlots_0_sharing; // @[Frontend.scala 66:23]
  wire  bpu_io_ftq_to_bpu_update_bits_ftb_entry_brSlots_0_valid; // @[Frontend.scala 66:23]
  wire [2:0] bpu_io_ftq_to_bpu_update_bits_ftb_entry_tailSlot_offset; // @[Frontend.scala 66:23]
  wire [19:0] bpu_io_ftq_to_bpu_update_bits_ftb_entry_tailSlot_lower; // @[Frontend.scala 66:23]
  wire [1:0] bpu_io_ftq_to_bpu_update_bits_ftb_entry_tailSlot_tarStat; // @[Frontend.scala 66:23]
  wire  bpu_io_ftq_to_bpu_update_bits_ftb_entry_tailSlot_sharing; // @[Frontend.scala 66:23]
  wire  bpu_io_ftq_to_bpu_update_bits_ftb_entry_tailSlot_valid; // @[Frontend.scala 66:23]
  wire [2:0] bpu_io_ftq_to_bpu_update_bits_ftb_entry_pftAddr; // @[Frontend.scala 66:23]
  wire  bpu_io_ftq_to_bpu_update_bits_ftb_entry_carry; // @[Frontend.scala 66:23]
  wire  bpu_io_ftq_to_bpu_update_bits_ftb_entry_isCall; // @[Frontend.scala 66:23]
  wire  bpu_io_ftq_to_bpu_update_bits_ftb_entry_isRet; // @[Frontend.scala 66:23]
  wire  bpu_io_ftq_to_bpu_update_bits_ftb_entry_isJalr; // @[Frontend.scala 66:23]
  wire  bpu_io_ftq_to_bpu_update_bits_ftb_entry_last_may_be_rvi_call; // @[Frontend.scala 66:23]
  wire  bpu_io_ftq_to_bpu_update_bits_ftb_entry_always_taken_0; // @[Frontend.scala 66:23]
  wire  bpu_io_ftq_to_bpu_update_bits_ftb_entry_always_taken_1; // @[Frontend.scala 66:23]
  wire  bpu_io_ftq_to_bpu_update_bits_br_taken_mask_0; // @[Frontend.scala 66:23]
  wire  bpu_io_ftq_to_bpu_update_bits_br_taken_mask_1; // @[Frontend.scala 66:23]
  wire  bpu_io_ftq_to_bpu_update_bits_jmp_taken; // @[Frontend.scala 66:23]
  wire  bpu_io_ftq_to_bpu_update_bits_mispred_mask_0; // @[Frontend.scala 66:23]
  wire  bpu_io_ftq_to_bpu_update_bits_mispred_mask_1; // @[Frontend.scala 66:23]
  wire  bpu_io_ftq_to_bpu_update_bits_mispred_mask_2; // @[Frontend.scala 66:23]
  wire  bpu_io_ftq_to_bpu_update_bits_old_entry; // @[Frontend.scala 66:23]
  wire [255:0] bpu_io_ftq_to_bpu_update_bits_meta; // @[Frontend.scala 66:23]
  wire [38:0] bpu_io_ftq_to_bpu_update_bits_full_target; // @[Frontend.scala 66:23]
  wire  bpu_io_ftq_to_bpu_enq_ptr_flag; // @[Frontend.scala 66:23]
  wire [2:0] bpu_io_ftq_to_bpu_enq_ptr_value; // @[Frontend.scala 66:23]
  wire  bpu_io_ctrl_ubtb_enable; // @[Frontend.scala 66:23]
  wire  bpu_io_ctrl_btb_enable; // @[Frontend.scala 66:23]
  wire  bpu_io_ctrl_tage_enable; // @[Frontend.scala 66:23]
  wire  bpu_io_ctrl_sc_enable; // @[Frontend.scala 66:23]
  wire  bpu_io_ctrl_ras_enable; // @[Frontend.scala 66:23]
  wire [35:0] bpu_io_reset_vector; // @[Frontend.scala 66:23]
  wire [5:0] bpu_io_perf_0_value; // @[Frontend.scala 66:23]
  wire [5:0] bpu_io_perf_1_value; // @[Frontend.scala 66:23]
  wire [5:0] bpu_io_perf_2_value; // @[Frontend.scala 66:23]
  wire [5:0] bpu_io_perf_3_value; // @[Frontend.scala 66:23]
  wire [5:0] bpu_io_perf_4_value; // @[Frontend.scala 66:23]
  wire [5:0] bpu_io_perf_5_value; // @[Frontend.scala 66:23]
  wire [5:0] bpu_io_perf_6_value; // @[Frontend.scala 66:23]
  wire  ifu_clock; // @[Frontend.scala 67:23]
  wire  ifu_reset; // @[Frontend.scala 67:23]
  wire  ifu_io_ftqInter_fromFtq_req_ready; // @[Frontend.scala 67:23]
  wire  ifu_io_ftqInter_fromFtq_req_valid; // @[Frontend.scala 67:23]
  wire [38:0] ifu_io_ftqInter_fromFtq_req_bits_startAddr; // @[Frontend.scala 67:23]
  wire [38:0] ifu_io_ftqInter_fromFtq_req_bits_nextlineStart; // @[Frontend.scala 67:23]
  wire [38:0] ifu_io_ftqInter_fromFtq_req_bits_nextStartAddr; // @[Frontend.scala 67:23]
  wire  ifu_io_ftqInter_fromFtq_req_bits_ftqIdx_flag; // @[Frontend.scala 67:23]
  wire [2:0] ifu_io_ftqInter_fromFtq_req_bits_ftqIdx_value; // @[Frontend.scala 67:23]
  wire  ifu_io_ftqInter_fromFtq_req_bits_ftqOffset_valid; // @[Frontend.scala 67:23]
  wire [2:0] ifu_io_ftqInter_fromFtq_req_bits_ftqOffset_bits; // @[Frontend.scala 67:23]
  wire  ifu_io_ftqInter_fromFtq_redirect_valid; // @[Frontend.scala 67:23]
  wire  ifu_io_ftqInter_fromFtq_redirect_bits_ftqIdx_flag; // @[Frontend.scala 67:23]
  wire [2:0] ifu_io_ftqInter_fromFtq_redirect_bits_ftqIdx_value; // @[Frontend.scala 67:23]
  wire [2:0] ifu_io_ftqInter_fromFtq_redirect_bits_ftqOffset; // @[Frontend.scala 67:23]
  wire  ifu_io_ftqInter_fromFtq_redirect_bits_level; // @[Frontend.scala 67:23]
  wire  ifu_io_ftqInter_fromFtq_flushFromBpu_s2_valid; // @[Frontend.scala 67:23]
  wire  ifu_io_ftqInter_fromFtq_flushFromBpu_s2_bits_flag; // @[Frontend.scala 67:23]
  wire [2:0] ifu_io_ftqInter_fromFtq_flushFromBpu_s2_bits_value; // @[Frontend.scala 67:23]
  wire  ifu_io_ftqInter_fromFtq_flushFromBpu_s3_valid; // @[Frontend.scala 67:23]
  wire  ifu_io_ftqInter_fromFtq_flushFromBpu_s3_bits_flag; // @[Frontend.scala 67:23]
  wire [2:0] ifu_io_ftqInter_fromFtq_flushFromBpu_s3_bits_value; // @[Frontend.scala 67:23]
  wire  ifu_io_ftqInter_toFtq_pdWb_valid; // @[Frontend.scala 67:23]
  wire [38:0] ifu_io_ftqInter_toFtq_pdWb_bits_pc_0; // @[Frontend.scala 67:23]
  wire [38:0] ifu_io_ftqInter_toFtq_pdWb_bits_pc_1; // @[Frontend.scala 67:23]
  wire [38:0] ifu_io_ftqInter_toFtq_pdWb_bits_pc_2; // @[Frontend.scala 67:23]
  wire [38:0] ifu_io_ftqInter_toFtq_pdWb_bits_pc_3; // @[Frontend.scala 67:23]
  wire [38:0] ifu_io_ftqInter_toFtq_pdWb_bits_pc_4; // @[Frontend.scala 67:23]
  wire [38:0] ifu_io_ftqInter_toFtq_pdWb_bits_pc_5; // @[Frontend.scala 67:23]
  wire [38:0] ifu_io_ftqInter_toFtq_pdWb_bits_pc_6; // @[Frontend.scala 67:23]
  wire [38:0] ifu_io_ftqInter_toFtq_pdWb_bits_pc_7; // @[Frontend.scala 67:23]
  wire  ifu_io_ftqInter_toFtq_pdWb_bits_pd_0_valid; // @[Frontend.scala 67:23]
  wire  ifu_io_ftqInter_toFtq_pdWb_bits_pd_0_isRVC; // @[Frontend.scala 67:23]
  wire [1:0] ifu_io_ftqInter_toFtq_pdWb_bits_pd_0_brType; // @[Frontend.scala 67:23]
  wire  ifu_io_ftqInter_toFtq_pdWb_bits_pd_0_isCall; // @[Frontend.scala 67:23]
  wire  ifu_io_ftqInter_toFtq_pdWb_bits_pd_0_isRet; // @[Frontend.scala 67:23]
  wire  ifu_io_ftqInter_toFtq_pdWb_bits_pd_1_valid; // @[Frontend.scala 67:23]
  wire  ifu_io_ftqInter_toFtq_pdWb_bits_pd_1_isRVC; // @[Frontend.scala 67:23]
  wire [1:0] ifu_io_ftqInter_toFtq_pdWb_bits_pd_1_brType; // @[Frontend.scala 67:23]
  wire  ifu_io_ftqInter_toFtq_pdWb_bits_pd_1_isCall; // @[Frontend.scala 67:23]
  wire  ifu_io_ftqInter_toFtq_pdWb_bits_pd_1_isRet; // @[Frontend.scala 67:23]
  wire  ifu_io_ftqInter_toFtq_pdWb_bits_pd_2_valid; // @[Frontend.scala 67:23]
  wire  ifu_io_ftqInter_toFtq_pdWb_bits_pd_2_isRVC; // @[Frontend.scala 67:23]
  wire [1:0] ifu_io_ftqInter_toFtq_pdWb_bits_pd_2_brType; // @[Frontend.scala 67:23]
  wire  ifu_io_ftqInter_toFtq_pdWb_bits_pd_2_isCall; // @[Frontend.scala 67:23]
  wire  ifu_io_ftqInter_toFtq_pdWb_bits_pd_2_isRet; // @[Frontend.scala 67:23]
  wire  ifu_io_ftqInter_toFtq_pdWb_bits_pd_3_valid; // @[Frontend.scala 67:23]
  wire  ifu_io_ftqInter_toFtq_pdWb_bits_pd_3_isRVC; // @[Frontend.scala 67:23]
  wire [1:0] ifu_io_ftqInter_toFtq_pdWb_bits_pd_3_brType; // @[Frontend.scala 67:23]
  wire  ifu_io_ftqInter_toFtq_pdWb_bits_pd_3_isCall; // @[Frontend.scala 67:23]
  wire  ifu_io_ftqInter_toFtq_pdWb_bits_pd_3_isRet; // @[Frontend.scala 67:23]
  wire  ifu_io_ftqInter_toFtq_pdWb_bits_pd_4_valid; // @[Frontend.scala 67:23]
  wire  ifu_io_ftqInter_toFtq_pdWb_bits_pd_4_isRVC; // @[Frontend.scala 67:23]
  wire [1:0] ifu_io_ftqInter_toFtq_pdWb_bits_pd_4_brType; // @[Frontend.scala 67:23]
  wire  ifu_io_ftqInter_toFtq_pdWb_bits_pd_4_isCall; // @[Frontend.scala 67:23]
  wire  ifu_io_ftqInter_toFtq_pdWb_bits_pd_4_isRet; // @[Frontend.scala 67:23]
  wire  ifu_io_ftqInter_toFtq_pdWb_bits_pd_5_valid; // @[Frontend.scala 67:23]
  wire  ifu_io_ftqInter_toFtq_pdWb_bits_pd_5_isRVC; // @[Frontend.scala 67:23]
  wire [1:0] ifu_io_ftqInter_toFtq_pdWb_bits_pd_5_brType; // @[Frontend.scala 67:23]
  wire  ifu_io_ftqInter_toFtq_pdWb_bits_pd_5_isCall; // @[Frontend.scala 67:23]
  wire  ifu_io_ftqInter_toFtq_pdWb_bits_pd_5_isRet; // @[Frontend.scala 67:23]
  wire  ifu_io_ftqInter_toFtq_pdWb_bits_pd_6_valid; // @[Frontend.scala 67:23]
  wire  ifu_io_ftqInter_toFtq_pdWb_bits_pd_6_isRVC; // @[Frontend.scala 67:23]
  wire [1:0] ifu_io_ftqInter_toFtq_pdWb_bits_pd_6_brType; // @[Frontend.scala 67:23]
  wire  ifu_io_ftqInter_toFtq_pdWb_bits_pd_6_isCall; // @[Frontend.scala 67:23]
  wire  ifu_io_ftqInter_toFtq_pdWb_bits_pd_6_isRet; // @[Frontend.scala 67:23]
  wire  ifu_io_ftqInter_toFtq_pdWb_bits_pd_7_valid; // @[Frontend.scala 67:23]
  wire  ifu_io_ftqInter_toFtq_pdWb_bits_pd_7_isRVC; // @[Frontend.scala 67:23]
  wire [1:0] ifu_io_ftqInter_toFtq_pdWb_bits_pd_7_brType; // @[Frontend.scala 67:23]
  wire  ifu_io_ftqInter_toFtq_pdWb_bits_pd_7_isCall; // @[Frontend.scala 67:23]
  wire  ifu_io_ftqInter_toFtq_pdWb_bits_pd_7_isRet; // @[Frontend.scala 67:23]
  wire  ifu_io_ftqInter_toFtq_pdWb_bits_ftqIdx_flag; // @[Frontend.scala 67:23]
  wire [2:0] ifu_io_ftqInter_toFtq_pdWb_bits_ftqIdx_value; // @[Frontend.scala 67:23]
  wire  ifu_io_ftqInter_toFtq_pdWb_bits_misOffset_valid; // @[Frontend.scala 67:23]
  wire [2:0] ifu_io_ftqInter_toFtq_pdWb_bits_misOffset_bits; // @[Frontend.scala 67:23]
  wire  ifu_io_ftqInter_toFtq_pdWb_bits_cfiOffset_valid; // @[Frontend.scala 67:23]
  wire [38:0] ifu_io_ftqInter_toFtq_pdWb_bits_target; // @[Frontend.scala 67:23]
  wire [38:0] ifu_io_ftqInter_toFtq_pdWb_bits_jalTarget; // @[Frontend.scala 67:23]
  wire  ifu_io_ftqInter_toFtq_pdWb_bits_instrRange_0; // @[Frontend.scala 67:23]
  wire  ifu_io_ftqInter_toFtq_pdWb_bits_instrRange_1; // @[Frontend.scala 67:23]
  wire  ifu_io_ftqInter_toFtq_pdWb_bits_instrRange_2; // @[Frontend.scala 67:23]
  wire  ifu_io_ftqInter_toFtq_pdWb_bits_instrRange_3; // @[Frontend.scala 67:23]
  wire  ifu_io_ftqInter_toFtq_pdWb_bits_instrRange_4; // @[Frontend.scala 67:23]
  wire  ifu_io_ftqInter_toFtq_pdWb_bits_instrRange_5; // @[Frontend.scala 67:23]
  wire  ifu_io_ftqInter_toFtq_pdWb_bits_instrRange_6; // @[Frontend.scala 67:23]
  wire  ifu_io_ftqInter_toFtq_pdWb_bits_instrRange_7; // @[Frontend.scala 67:23]
  wire  ifu_io_icacheInter_icacheReady; // @[Frontend.scala 67:23]
  wire  ifu_io_icacheInter_resp_0_valid; // @[Frontend.scala 67:23]
  wire [38:0] ifu_io_icacheInter_resp_0_bits_vaddr; // @[Frontend.scala 67:23]
  wire [511:0] ifu_io_icacheInter_resp_0_bits_registerData; // @[Frontend.scala 67:23]
  wire [511:0] ifu_io_icacheInter_resp_0_bits_sramData; // @[Frontend.scala 67:23]
  wire  ifu_io_icacheInter_resp_0_bits_select; // @[Frontend.scala 67:23]
  wire [35:0] ifu_io_icacheInter_resp_0_bits_paddr; // @[Frontend.scala 67:23]
  wire  ifu_io_icacheInter_resp_0_bits_tlbExcp_pageFault; // @[Frontend.scala 67:23]
  wire  ifu_io_icacheInter_resp_0_bits_tlbExcp_accessFault; // @[Frontend.scala 67:23]
  wire  ifu_io_icacheInter_resp_0_bits_tlbExcp_mmio; // @[Frontend.scala 67:23]
  wire  ifu_io_icacheInter_resp_1_valid; // @[Frontend.scala 67:23]
  wire [38:0] ifu_io_icacheInter_resp_1_bits_vaddr; // @[Frontend.scala 67:23]
  wire [511:0] ifu_io_icacheInter_resp_1_bits_registerData; // @[Frontend.scala 67:23]
  wire [511:0] ifu_io_icacheInter_resp_1_bits_sramData; // @[Frontend.scala 67:23]
  wire  ifu_io_icacheInter_resp_1_bits_select; // @[Frontend.scala 67:23]
  wire  ifu_io_icacheInter_resp_1_bits_tlbExcp_pageFault; // @[Frontend.scala 67:23]
  wire  ifu_io_icacheInter_resp_1_bits_tlbExcp_accessFault; // @[Frontend.scala 67:23]
  wire  ifu_io_icacheStop; // @[Frontend.scala 67:23]
  wire  ifu_io_icachePerfInfo_only_0_hit; // @[Frontend.scala 67:23]
  wire  ifu_io_icachePerfInfo_only_0_miss; // @[Frontend.scala 67:23]
  wire  ifu_io_icachePerfInfo_hit_0_hit_1; // @[Frontend.scala 67:23]
  wire  ifu_io_icachePerfInfo_hit_0_miss_1; // @[Frontend.scala 67:23]
  wire  ifu_io_icachePerfInfo_miss_0_hit_1; // @[Frontend.scala 67:23]
  wire  ifu_io_icachePerfInfo_miss_0_miss_1; // @[Frontend.scala 67:23]
  wire  ifu_io_icachePerfInfo_hit_0_except_1; // @[Frontend.scala 67:23]
  wire  ifu_io_icachePerfInfo_miss_0_except_1; // @[Frontend.scala 67:23]
  wire  ifu_io_icachePerfInfo_except_0; // @[Frontend.scala 67:23]
  wire  ifu_io_icachePerfInfo_bank_hit_1; // @[Frontend.scala 67:23]
  wire  ifu_io_icachePerfInfo_hit; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_ready; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_valid; // @[Frontend.scala 67:23]
  wire [31:0] ifu_io_toIbuffer_bits_instrs_0; // @[Frontend.scala 67:23]
  wire [31:0] ifu_io_toIbuffer_bits_instrs_1; // @[Frontend.scala 67:23]
  wire [31:0] ifu_io_toIbuffer_bits_instrs_2; // @[Frontend.scala 67:23]
  wire [31:0] ifu_io_toIbuffer_bits_instrs_3; // @[Frontend.scala 67:23]
  wire [31:0] ifu_io_toIbuffer_bits_instrs_4; // @[Frontend.scala 67:23]
  wire [31:0] ifu_io_toIbuffer_bits_instrs_5; // @[Frontend.scala 67:23]
  wire [31:0] ifu_io_toIbuffer_bits_instrs_6; // @[Frontend.scala 67:23]
  wire [31:0] ifu_io_toIbuffer_bits_instrs_7; // @[Frontend.scala 67:23]
  wire [7:0] ifu_io_toIbuffer_bits_valid; // @[Frontend.scala 67:23]
  wire [7:0] ifu_io_toIbuffer_bits_enqEnable; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_pd_0_isRVC; // @[Frontend.scala 67:23]
  wire [1:0] ifu_io_toIbuffer_bits_pd_0_brType; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_pd_0_isCall; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_pd_0_isRet; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_pd_1_isRVC; // @[Frontend.scala 67:23]
  wire [1:0] ifu_io_toIbuffer_bits_pd_1_brType; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_pd_1_isCall; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_pd_1_isRet; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_pd_2_isRVC; // @[Frontend.scala 67:23]
  wire [1:0] ifu_io_toIbuffer_bits_pd_2_brType; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_pd_2_isCall; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_pd_2_isRet; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_pd_3_isRVC; // @[Frontend.scala 67:23]
  wire [1:0] ifu_io_toIbuffer_bits_pd_3_brType; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_pd_3_isCall; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_pd_3_isRet; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_pd_4_isRVC; // @[Frontend.scala 67:23]
  wire [1:0] ifu_io_toIbuffer_bits_pd_4_brType; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_pd_4_isCall; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_pd_4_isRet; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_pd_5_isRVC; // @[Frontend.scala 67:23]
  wire [1:0] ifu_io_toIbuffer_bits_pd_5_brType; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_pd_5_isCall; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_pd_5_isRet; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_pd_6_isRVC; // @[Frontend.scala 67:23]
  wire [1:0] ifu_io_toIbuffer_bits_pd_6_brType; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_pd_6_isCall; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_pd_6_isRet; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_pd_7_isRVC; // @[Frontend.scala 67:23]
  wire [1:0] ifu_io_toIbuffer_bits_pd_7_brType; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_pd_7_isCall; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_pd_7_isRet; // @[Frontend.scala 67:23]
  wire [9:0] ifu_io_toIbuffer_bits_foldpc_0; // @[Frontend.scala 67:23]
  wire [9:0] ifu_io_toIbuffer_bits_foldpc_1; // @[Frontend.scala 67:23]
  wire [9:0] ifu_io_toIbuffer_bits_foldpc_2; // @[Frontend.scala 67:23]
  wire [9:0] ifu_io_toIbuffer_bits_foldpc_3; // @[Frontend.scala 67:23]
  wire [9:0] ifu_io_toIbuffer_bits_foldpc_4; // @[Frontend.scala 67:23]
  wire [9:0] ifu_io_toIbuffer_bits_foldpc_5; // @[Frontend.scala 67:23]
  wire [9:0] ifu_io_toIbuffer_bits_foldpc_6; // @[Frontend.scala 67:23]
  wire [9:0] ifu_io_toIbuffer_bits_foldpc_7; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_ftqPtr_flag; // @[Frontend.scala 67:23]
  wire [2:0] ifu_io_toIbuffer_bits_ftqPtr_value; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_ftqOffset_0_valid; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_ftqOffset_1_valid; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_ftqOffset_2_valid; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_ftqOffset_3_valid; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_ftqOffset_4_valid; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_ftqOffset_5_valid; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_ftqOffset_6_valid; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_ftqOffset_7_valid; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_ipf_0; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_ipf_1; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_ipf_2; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_ipf_3; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_ipf_4; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_ipf_5; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_ipf_6; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_ipf_7; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_acf_0; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_acf_1; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_acf_2; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_acf_3; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_acf_4; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_acf_5; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_acf_6; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_acf_7; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_crossPageIPFFix_0; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_crossPageIPFFix_1; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_crossPageIPFFix_2; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_crossPageIPFFix_3; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_crossPageIPFFix_4; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_crossPageIPFFix_5; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_crossPageIPFFix_6; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_crossPageIPFFix_7; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_triggered_0_frontendHit_0; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_triggered_0_frontendHit_1; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_triggered_0_frontendHit_2; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_triggered_0_frontendHit_3; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_triggered_0_backendEn_0; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_triggered_0_backendEn_1; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_triggered_1_frontendHit_0; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_triggered_1_frontendHit_1; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_triggered_1_frontendHit_2; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_triggered_1_frontendHit_3; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_triggered_1_backendEn_0; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_triggered_1_backendEn_1; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_triggered_2_frontendHit_0; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_triggered_2_frontendHit_1; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_triggered_2_frontendHit_2; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_triggered_2_frontendHit_3; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_triggered_2_backendEn_0; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_triggered_2_backendEn_1; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_triggered_3_frontendHit_0; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_triggered_3_frontendHit_1; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_triggered_3_frontendHit_2; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_triggered_3_frontendHit_3; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_triggered_3_backendEn_0; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_triggered_3_backendEn_1; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_triggered_4_frontendHit_0; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_triggered_4_frontendHit_1; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_triggered_4_frontendHit_2; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_triggered_4_frontendHit_3; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_triggered_4_backendEn_0; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_triggered_4_backendEn_1; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_triggered_5_frontendHit_0; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_triggered_5_frontendHit_1; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_triggered_5_frontendHit_2; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_triggered_5_frontendHit_3; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_triggered_5_backendEn_0; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_triggered_5_backendEn_1; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_triggered_6_frontendHit_0; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_triggered_6_frontendHit_1; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_triggered_6_frontendHit_2; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_triggered_6_frontendHit_3; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_triggered_6_backendEn_0; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_triggered_6_backendEn_1; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_triggered_7_frontendHit_0; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_triggered_7_frontendHit_1; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_triggered_7_frontendHit_2; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_triggered_7_frontendHit_3; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_triggered_7_backendEn_0; // @[Frontend.scala 67:23]
  wire  ifu_io_toIbuffer_bits_triggered_7_backendEn_1; // @[Frontend.scala 67:23]
  wire  ifu_io_uncacheInter_fromUncache_ready; // @[Frontend.scala 67:23]
  wire  ifu_io_uncacheInter_fromUncache_valid; // @[Frontend.scala 67:23]
  wire [31:0] ifu_io_uncacheInter_fromUncache_bits_data; // @[Frontend.scala 67:23]
  wire  ifu_io_uncacheInter_toUncache_ready; // @[Frontend.scala 67:23]
  wire  ifu_io_uncacheInter_toUncache_valid; // @[Frontend.scala 67:23]
  wire [35:0] ifu_io_uncacheInter_toUncache_bits_addr; // @[Frontend.scala 67:23]
  wire  ifu_io_frontendTrigger_t_valid; // @[Frontend.scala 67:23]
  wire [1:0] ifu_io_frontendTrigger_t_bits_addr; // @[Frontend.scala 67:23]
  wire [1:0] ifu_io_frontendTrigger_t_bits_tdata_matchType; // @[Frontend.scala 67:23]
  wire  ifu_io_frontendTrigger_t_bits_tdata_select; // @[Frontend.scala 67:23]
  wire  ifu_io_frontendTrigger_t_bits_tdata_timing; // @[Frontend.scala 67:23]
  wire  ifu_io_frontendTrigger_t_bits_tdata_chain; // @[Frontend.scala 67:23]
  wire [63:0] ifu_io_frontendTrigger_t_bits_tdata_tdata2; // @[Frontend.scala 67:23]
  wire  ifu_io_csrTriggerEnable_0; // @[Frontend.scala 67:23]
  wire  ifu_io_csrTriggerEnable_1; // @[Frontend.scala 67:23]
  wire  ifu_io_csrTriggerEnable_2; // @[Frontend.scala 67:23]
  wire  ifu_io_csrTriggerEnable_3; // @[Frontend.scala 67:23]
  wire  ifu_io_rob_commits_0_valid; // @[Frontend.scala 67:23]
  wire  ifu_io_rob_commits_0_bits_ftqIdx_flag; // @[Frontend.scala 67:23]
  wire [2:0] ifu_io_rob_commits_0_bits_ftqIdx_value; // @[Frontend.scala 67:23]
  wire [2:0] ifu_io_rob_commits_0_bits_ftqOffset; // @[Frontend.scala 67:23]
  wire  ifu_io_rob_commits_1_valid; // @[Frontend.scala 67:23]
  wire  ifu_io_rob_commits_1_bits_ftqIdx_flag; // @[Frontend.scala 67:23]
  wire [2:0] ifu_io_rob_commits_1_bits_ftqIdx_value; // @[Frontend.scala 67:23]
  wire [2:0] ifu_io_rob_commits_1_bits_ftqOffset; // @[Frontend.scala 67:23]
  wire  ifu_io_iTLBInter_req_valid; // @[Frontend.scala 67:23]
  wire [38:0] ifu_io_iTLBInter_req_bits_vaddr; // @[Frontend.scala 67:23]
  wire [35:0] ifu_io_iTLBInter_resp_bits_paddr_0; // @[Frontend.scala 67:23]
  wire  ifu_io_iTLBInter_resp_bits_miss; // @[Frontend.scala 67:23]
  wire  ifu_io_iTLBInter_resp_bits_excp_0_pf_instr; // @[Frontend.scala 67:23]
  wire  ifu_io_iTLBInter_resp_bits_excp_0_af_instr; // @[Frontend.scala 67:23]
  wire [35:0] ifu_io_pmp_req_bits_addr; // @[Frontend.scala 67:23]
  wire  ifu_io_pmp_resp_instr; // @[Frontend.scala 67:23]
  wire  ifu_io_pmp_resp_mmio; // @[Frontend.scala 67:23]
  wire  ifu_io_mmioCommitRead_mmioFtqPtr_flag; // @[Frontend.scala 67:23]
  wire [2:0] ifu_io_mmioCommitRead_mmioFtqPtr_value; // @[Frontend.scala 67:23]
  wire  ifu_io_mmioCommitRead_mmioLastCommit; // @[Frontend.scala 67:23]
  wire [5:0] ifu_io_perf_0_value; // @[Frontend.scala 67:23]
  wire [5:0] ifu_io_perf_1_value; // @[Frontend.scala 67:23]
  wire [5:0] ifu_io_perf_2_value; // @[Frontend.scala 67:23]
  wire [5:0] ifu_io_perf_3_value; // @[Frontend.scala 67:23]
  wire [5:0] ifu_io_perf_4_value; // @[Frontend.scala 67:23]
  wire [5:0] ifu_io_perf_5_value; // @[Frontend.scala 67:23]
  wire [5:0] ifu_io_perf_6_value; // @[Frontend.scala 67:23]
  wire [5:0] ifu_io_perf_7_value; // @[Frontend.scala 67:23]
  wire [5:0] ifu_io_perf_8_value; // @[Frontend.scala 67:23]
  wire [5:0] ifu_io_perf_9_value; // @[Frontend.scala 67:23]
  wire [5:0] ifu_io_perf_10_value; // @[Frontend.scala 67:23]
  wire [5:0] ifu_io_perf_11_value; // @[Frontend.scala 67:23]
  wire [5:0] ifu_io_perf_12_value; // @[Frontend.scala 67:23]
  wire  ibuffer_clock; // @[Frontend.scala 68:24]
  wire  ibuffer_reset; // @[Frontend.scala 68:24]
  wire  ibuffer_io_flush; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_ready; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_valid; // @[Frontend.scala 68:24]
  wire [31:0] ibuffer_io_in_bits_instrs_0; // @[Frontend.scala 68:24]
  wire [31:0] ibuffer_io_in_bits_instrs_1; // @[Frontend.scala 68:24]
  wire [31:0] ibuffer_io_in_bits_instrs_2; // @[Frontend.scala 68:24]
  wire [31:0] ibuffer_io_in_bits_instrs_3; // @[Frontend.scala 68:24]
  wire [31:0] ibuffer_io_in_bits_instrs_4; // @[Frontend.scala 68:24]
  wire [31:0] ibuffer_io_in_bits_instrs_5; // @[Frontend.scala 68:24]
  wire [31:0] ibuffer_io_in_bits_instrs_6; // @[Frontend.scala 68:24]
  wire [31:0] ibuffer_io_in_bits_instrs_7; // @[Frontend.scala 68:24]
  wire [7:0] ibuffer_io_in_bits_valid; // @[Frontend.scala 68:24]
  wire [7:0] ibuffer_io_in_bits_enqEnable; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_pd_0_isRVC; // @[Frontend.scala 68:24]
  wire [1:0] ibuffer_io_in_bits_pd_0_brType; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_pd_0_isCall; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_pd_0_isRet; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_pd_1_isRVC; // @[Frontend.scala 68:24]
  wire [1:0] ibuffer_io_in_bits_pd_1_brType; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_pd_1_isCall; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_pd_1_isRet; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_pd_2_isRVC; // @[Frontend.scala 68:24]
  wire [1:0] ibuffer_io_in_bits_pd_2_brType; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_pd_2_isCall; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_pd_2_isRet; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_pd_3_isRVC; // @[Frontend.scala 68:24]
  wire [1:0] ibuffer_io_in_bits_pd_3_brType; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_pd_3_isCall; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_pd_3_isRet; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_pd_4_isRVC; // @[Frontend.scala 68:24]
  wire [1:0] ibuffer_io_in_bits_pd_4_brType; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_pd_4_isCall; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_pd_4_isRet; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_pd_5_isRVC; // @[Frontend.scala 68:24]
  wire [1:0] ibuffer_io_in_bits_pd_5_brType; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_pd_5_isCall; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_pd_5_isRet; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_pd_6_isRVC; // @[Frontend.scala 68:24]
  wire [1:0] ibuffer_io_in_bits_pd_6_brType; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_pd_6_isCall; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_pd_6_isRet; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_pd_7_isRVC; // @[Frontend.scala 68:24]
  wire [1:0] ibuffer_io_in_bits_pd_7_brType; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_pd_7_isCall; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_pd_7_isRet; // @[Frontend.scala 68:24]
  wire [9:0] ibuffer_io_in_bits_foldpc_0; // @[Frontend.scala 68:24]
  wire [9:0] ibuffer_io_in_bits_foldpc_1; // @[Frontend.scala 68:24]
  wire [9:0] ibuffer_io_in_bits_foldpc_2; // @[Frontend.scala 68:24]
  wire [9:0] ibuffer_io_in_bits_foldpc_3; // @[Frontend.scala 68:24]
  wire [9:0] ibuffer_io_in_bits_foldpc_4; // @[Frontend.scala 68:24]
  wire [9:0] ibuffer_io_in_bits_foldpc_5; // @[Frontend.scala 68:24]
  wire [9:0] ibuffer_io_in_bits_foldpc_6; // @[Frontend.scala 68:24]
  wire [9:0] ibuffer_io_in_bits_foldpc_7; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_ftqPtr_flag; // @[Frontend.scala 68:24]
  wire [2:0] ibuffer_io_in_bits_ftqPtr_value; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_ftqOffset_0_valid; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_ftqOffset_1_valid; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_ftqOffset_2_valid; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_ftqOffset_3_valid; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_ftqOffset_4_valid; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_ftqOffset_5_valid; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_ftqOffset_6_valid; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_ftqOffset_7_valid; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_ipf_0; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_ipf_1; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_ipf_2; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_ipf_3; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_ipf_4; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_ipf_5; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_ipf_6; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_ipf_7; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_acf_0; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_acf_1; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_acf_2; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_acf_3; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_acf_4; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_acf_5; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_acf_6; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_acf_7; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_crossPageIPFFix_0; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_crossPageIPFFix_1; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_crossPageIPFFix_2; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_crossPageIPFFix_3; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_crossPageIPFFix_4; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_crossPageIPFFix_5; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_crossPageIPFFix_6; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_crossPageIPFFix_7; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_triggered_0_frontendHit_0; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_triggered_0_frontendHit_1; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_triggered_0_frontendHit_2; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_triggered_0_frontendHit_3; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_triggered_0_backendEn_0; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_triggered_0_backendEn_1; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_triggered_1_frontendHit_0; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_triggered_1_frontendHit_1; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_triggered_1_frontendHit_2; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_triggered_1_frontendHit_3; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_triggered_1_backendEn_0; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_triggered_1_backendEn_1; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_triggered_2_frontendHit_0; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_triggered_2_frontendHit_1; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_triggered_2_frontendHit_2; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_triggered_2_frontendHit_3; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_triggered_2_backendEn_0; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_triggered_2_backendEn_1; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_triggered_3_frontendHit_0; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_triggered_3_frontendHit_1; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_triggered_3_frontendHit_2; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_triggered_3_frontendHit_3; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_triggered_3_backendEn_0; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_triggered_3_backendEn_1; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_triggered_4_frontendHit_0; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_triggered_4_frontendHit_1; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_triggered_4_frontendHit_2; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_triggered_4_frontendHit_3; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_triggered_4_backendEn_0; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_triggered_4_backendEn_1; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_triggered_5_frontendHit_0; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_triggered_5_frontendHit_1; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_triggered_5_frontendHit_2; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_triggered_5_frontendHit_3; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_triggered_5_backendEn_0; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_triggered_5_backendEn_1; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_triggered_6_frontendHit_0; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_triggered_6_frontendHit_1; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_triggered_6_frontendHit_2; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_triggered_6_frontendHit_3; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_triggered_6_backendEn_0; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_triggered_6_backendEn_1; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_triggered_7_frontendHit_0; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_triggered_7_frontendHit_1; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_triggered_7_frontendHit_2; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_triggered_7_frontendHit_3; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_triggered_7_backendEn_0; // @[Frontend.scala 68:24]
  wire  ibuffer_io_in_bits_triggered_7_backendEn_1; // @[Frontend.scala 68:24]
  wire  ibuffer_io_out_0_ready; // @[Frontend.scala 68:24]
  wire  ibuffer_io_out_0_valid; // @[Frontend.scala 68:24]
  wire [31:0] ibuffer_io_out_0_bits_instr; // @[Frontend.scala 68:24]
  wire [9:0] ibuffer_io_out_0_bits_foldpc; // @[Frontend.scala 68:24]
  wire  ibuffer_io_out_0_bits_exceptionVec_1; // @[Frontend.scala 68:24]
  wire  ibuffer_io_out_0_bits_exceptionVec_12; // @[Frontend.scala 68:24]
  wire  ibuffer_io_out_0_bits_trigger_frontendHit_0; // @[Frontend.scala 68:24]
  wire  ibuffer_io_out_0_bits_trigger_frontendHit_1; // @[Frontend.scala 68:24]
  wire  ibuffer_io_out_0_bits_trigger_frontendHit_2; // @[Frontend.scala 68:24]
  wire  ibuffer_io_out_0_bits_trigger_frontendHit_3; // @[Frontend.scala 68:24]
  wire  ibuffer_io_out_0_bits_trigger_backendEn_0; // @[Frontend.scala 68:24]
  wire  ibuffer_io_out_0_bits_trigger_backendEn_1; // @[Frontend.scala 68:24]
  wire  ibuffer_io_out_0_bits_pd_isRVC; // @[Frontend.scala 68:24]
  wire [1:0] ibuffer_io_out_0_bits_pd_brType; // @[Frontend.scala 68:24]
  wire  ibuffer_io_out_0_bits_pd_isCall; // @[Frontend.scala 68:24]
  wire  ibuffer_io_out_0_bits_pd_isRet; // @[Frontend.scala 68:24]
  wire  ibuffer_io_out_0_bits_pred_taken; // @[Frontend.scala 68:24]
  wire  ibuffer_io_out_0_bits_crossPageIPFFix; // @[Frontend.scala 68:24]
  wire  ibuffer_io_out_0_bits_ftqPtr_flag; // @[Frontend.scala 68:24]
  wire [2:0] ibuffer_io_out_0_bits_ftqPtr_value; // @[Frontend.scala 68:24]
  wire [2:0] ibuffer_io_out_0_bits_ftqOffset; // @[Frontend.scala 68:24]
  wire  ibuffer_io_out_1_ready; // @[Frontend.scala 68:24]
  wire  ibuffer_io_out_1_valid; // @[Frontend.scala 68:24]
  wire [31:0] ibuffer_io_out_1_bits_instr; // @[Frontend.scala 68:24]
  wire [9:0] ibuffer_io_out_1_bits_foldpc; // @[Frontend.scala 68:24]
  wire  ibuffer_io_out_1_bits_exceptionVec_1; // @[Frontend.scala 68:24]
  wire  ibuffer_io_out_1_bits_exceptionVec_12; // @[Frontend.scala 68:24]
  wire  ibuffer_io_out_1_bits_trigger_frontendHit_0; // @[Frontend.scala 68:24]
  wire  ibuffer_io_out_1_bits_trigger_frontendHit_1; // @[Frontend.scala 68:24]
  wire  ibuffer_io_out_1_bits_trigger_frontendHit_2; // @[Frontend.scala 68:24]
  wire  ibuffer_io_out_1_bits_trigger_frontendHit_3; // @[Frontend.scala 68:24]
  wire  ibuffer_io_out_1_bits_trigger_backendEn_0; // @[Frontend.scala 68:24]
  wire  ibuffer_io_out_1_bits_trigger_backendEn_1; // @[Frontend.scala 68:24]
  wire  ibuffer_io_out_1_bits_pd_isRVC; // @[Frontend.scala 68:24]
  wire [1:0] ibuffer_io_out_1_bits_pd_brType; // @[Frontend.scala 68:24]
  wire  ibuffer_io_out_1_bits_pd_isCall; // @[Frontend.scala 68:24]
  wire  ibuffer_io_out_1_bits_pd_isRet; // @[Frontend.scala 68:24]
  wire  ibuffer_io_out_1_bits_pred_taken; // @[Frontend.scala 68:24]
  wire  ibuffer_io_out_1_bits_crossPageIPFFix; // @[Frontend.scala 68:24]
  wire  ibuffer_io_out_1_bits_ftqPtr_flag; // @[Frontend.scala 68:24]
  wire [2:0] ibuffer_io_out_1_bits_ftqPtr_value; // @[Frontend.scala 68:24]
  wire [2:0] ibuffer_io_out_1_bits_ftqOffset; // @[Frontend.scala 68:24]
  wire [5:0] ibuffer_io_perf_0_value; // @[Frontend.scala 68:24]
  wire [5:0] ibuffer_io_perf_1_value; // @[Frontend.scala 68:24]
  wire [5:0] ibuffer_io_perf_2_value; // @[Frontend.scala 68:24]
  wire [5:0] ibuffer_io_perf_3_value; // @[Frontend.scala 68:24]
  wire [5:0] ibuffer_io_perf_4_value; // @[Frontend.scala 68:24]
  wire [5:0] ibuffer_io_perf_5_value; // @[Frontend.scala 68:24]
  wire [5:0] ibuffer_io_perf_6_value; // @[Frontend.scala 68:24]
  wire [5:0] ibuffer_io_perf_7_value; // @[Frontend.scala 68:24]
  wire  ftq_clock; // @[Frontend.scala 69:19]
  wire  ftq_reset; // @[Frontend.scala 69:19]
  wire  ftq_io_fromBpu_resp_ready; // @[Frontend.scala 69:19]
  wire  ftq_io_fromBpu_resp_valid; // @[Frontend.scala 69:19]
  wire [38:0] ftq_io_fromBpu_resp_bits_s1_pc; // @[Frontend.scala 69:19]
  wire  ftq_io_fromBpu_resp_bits_s1_full_pred_br_taken_mask_0; // @[Frontend.scala 69:19]
  wire  ftq_io_fromBpu_resp_bits_s1_full_pred_br_taken_mask_1; // @[Frontend.scala 69:19]
  wire  ftq_io_fromBpu_resp_bits_s1_full_pred_slot_valids_0; // @[Frontend.scala 69:19]
  wire  ftq_io_fromBpu_resp_bits_s1_full_pred_slot_valids_1; // @[Frontend.scala 69:19]
  wire [38:0] ftq_io_fromBpu_resp_bits_s1_full_pred_targets_0; // @[Frontend.scala 69:19]
  wire [38:0] ftq_io_fromBpu_resp_bits_s1_full_pred_targets_1; // @[Frontend.scala 69:19]
  wire [2:0] ftq_io_fromBpu_resp_bits_s1_full_pred_offsets_0; // @[Frontend.scala 69:19]
  wire [2:0] ftq_io_fromBpu_resp_bits_s1_full_pred_offsets_1; // @[Frontend.scala 69:19]
  wire [38:0] ftq_io_fromBpu_resp_bits_s1_full_pred_fallThroughAddr; // @[Frontend.scala 69:19]
  wire  ftq_io_fromBpu_resp_bits_s1_full_pred_fallThroughErr; // @[Frontend.scala 69:19]
  wire  ftq_io_fromBpu_resp_bits_s1_full_pred_is_br_sharing; // @[Frontend.scala 69:19]
  wire  ftq_io_fromBpu_resp_bits_s1_full_pred_hit; // @[Frontend.scala 69:19]
  wire [38:0] ftq_io_fromBpu_resp_bits_s2_pc; // @[Frontend.scala 69:19]
  wire  ftq_io_fromBpu_resp_bits_s2_valid; // @[Frontend.scala 69:19]
  wire  ftq_io_fromBpu_resp_bits_s2_hasRedirect; // @[Frontend.scala 69:19]
  wire  ftq_io_fromBpu_resp_bits_s2_ftq_idx_flag; // @[Frontend.scala 69:19]
  wire [2:0] ftq_io_fromBpu_resp_bits_s2_ftq_idx_value; // @[Frontend.scala 69:19]
  wire  ftq_io_fromBpu_resp_bits_s2_full_pred_br_taken_mask_0; // @[Frontend.scala 69:19]
  wire  ftq_io_fromBpu_resp_bits_s2_full_pred_br_taken_mask_1; // @[Frontend.scala 69:19]
  wire  ftq_io_fromBpu_resp_bits_s2_full_pred_slot_valids_0; // @[Frontend.scala 69:19]
  wire  ftq_io_fromBpu_resp_bits_s2_full_pred_slot_valids_1; // @[Frontend.scala 69:19]
  wire [38:0] ftq_io_fromBpu_resp_bits_s2_full_pred_targets_0; // @[Frontend.scala 69:19]
  wire [38:0] ftq_io_fromBpu_resp_bits_s2_full_pred_targets_1; // @[Frontend.scala 69:19]
  wire [2:0] ftq_io_fromBpu_resp_bits_s2_full_pred_offsets_0; // @[Frontend.scala 69:19]
  wire [2:0] ftq_io_fromBpu_resp_bits_s2_full_pred_offsets_1; // @[Frontend.scala 69:19]
  wire [38:0] ftq_io_fromBpu_resp_bits_s2_full_pred_fallThroughAddr; // @[Frontend.scala 69:19]
  wire  ftq_io_fromBpu_resp_bits_s2_full_pred_fallThroughErr; // @[Frontend.scala 69:19]
  wire  ftq_io_fromBpu_resp_bits_s2_full_pred_is_br_sharing; // @[Frontend.scala 69:19]
  wire  ftq_io_fromBpu_resp_bits_s2_full_pred_hit; // @[Frontend.scala 69:19]
  wire [38:0] ftq_io_fromBpu_resp_bits_s3_pc; // @[Frontend.scala 69:19]
  wire  ftq_io_fromBpu_resp_bits_s3_valid; // @[Frontend.scala 69:19]
  wire  ftq_io_fromBpu_resp_bits_s3_hasRedirect; // @[Frontend.scala 69:19]
  wire  ftq_io_fromBpu_resp_bits_s3_ftq_idx_flag; // @[Frontend.scala 69:19]
  wire [2:0] ftq_io_fromBpu_resp_bits_s3_ftq_idx_value; // @[Frontend.scala 69:19]
  wire  ftq_io_fromBpu_resp_bits_s3_full_pred_br_taken_mask_0; // @[Frontend.scala 69:19]
  wire  ftq_io_fromBpu_resp_bits_s3_full_pred_br_taken_mask_1; // @[Frontend.scala 69:19]
  wire  ftq_io_fromBpu_resp_bits_s3_full_pred_slot_valids_0; // @[Frontend.scala 69:19]
  wire  ftq_io_fromBpu_resp_bits_s3_full_pred_slot_valids_1; // @[Frontend.scala 69:19]
  wire [38:0] ftq_io_fromBpu_resp_bits_s3_full_pred_targets_0; // @[Frontend.scala 69:19]
  wire [38:0] ftq_io_fromBpu_resp_bits_s3_full_pred_targets_1; // @[Frontend.scala 69:19]
  wire [2:0] ftq_io_fromBpu_resp_bits_s3_full_pred_offsets_0; // @[Frontend.scala 69:19]
  wire [2:0] ftq_io_fromBpu_resp_bits_s3_full_pred_offsets_1; // @[Frontend.scala 69:19]
  wire [38:0] ftq_io_fromBpu_resp_bits_s3_full_pred_fallThroughAddr; // @[Frontend.scala 69:19]
  wire  ftq_io_fromBpu_resp_bits_s3_full_pred_fallThroughErr; // @[Frontend.scala 69:19]
  wire  ftq_io_fromBpu_resp_bits_s3_full_pred_is_br_sharing; // @[Frontend.scala 69:19]
  wire  ftq_io_fromBpu_resp_bits_s3_full_pred_hit; // @[Frontend.scala 69:19]
  wire [255:0] ftq_io_fromBpu_resp_bits_last_stage_meta; // @[Frontend.scala 69:19]
  wire [7:0] ftq_io_fromBpu_resp_bits_last_stage_spec_info_folded_hist_hist_17_folded_hist; // @[Frontend.scala 69:19]
  wire [7:0] ftq_io_fromBpu_resp_bits_last_stage_spec_info_folded_hist_hist_16_folded_hist; // @[Frontend.scala 69:19]
  wire [10:0] ftq_io_fromBpu_resp_bits_last_stage_spec_info_folded_hist_hist_15_folded_hist; // @[Frontend.scala 69:19]
  wire [6:0] ftq_io_fromBpu_resp_bits_last_stage_spec_info_folded_hist_hist_14_folded_hist; // @[Frontend.scala 69:19]
  wire [6:0] ftq_io_fromBpu_resp_bits_last_stage_spec_info_folded_hist_hist_13_folded_hist; // @[Frontend.scala 69:19]
  wire [6:0] ftq_io_fromBpu_resp_bits_last_stage_spec_info_folded_hist_hist_12_folded_hist; // @[Frontend.scala 69:19]
  wire [7:0] ftq_io_fromBpu_resp_bits_last_stage_spec_info_folded_hist_hist_11_folded_hist; // @[Frontend.scala 69:19]
  wire [8:0] ftq_io_fromBpu_resp_bits_last_stage_spec_info_folded_hist_hist_10_folded_hist; // @[Frontend.scala 69:19]
  wire [6:0] ftq_io_fromBpu_resp_bits_last_stage_spec_info_folded_hist_hist_9_folded_hist; // @[Frontend.scala 69:19]
  wire [7:0] ftq_io_fromBpu_resp_bits_last_stage_spec_info_folded_hist_hist_8_folded_hist; // @[Frontend.scala 69:19]
  wire [8:0] ftq_io_fromBpu_resp_bits_last_stage_spec_info_folded_hist_hist_7_folded_hist; // @[Frontend.scala 69:19]
  wire [8:0] ftq_io_fromBpu_resp_bits_last_stage_spec_info_folded_hist_hist_6_folded_hist; // @[Frontend.scala 69:19]
  wire [10:0] ftq_io_fromBpu_resp_bits_last_stage_spec_info_folded_hist_hist_5_folded_hist; // @[Frontend.scala 69:19]
  wire [3:0] ftq_io_fromBpu_resp_bits_last_stage_spec_info_folded_hist_hist_4_folded_hist; // @[Frontend.scala 69:19]
  wire [10:0] ftq_io_fromBpu_resp_bits_last_stage_spec_info_folded_hist_hist_3_folded_hist; // @[Frontend.scala 69:19]
  wire [7:0] ftq_io_fromBpu_resp_bits_last_stage_spec_info_folded_hist_hist_2_folded_hist; // @[Frontend.scala 69:19]
  wire [7:0] ftq_io_fromBpu_resp_bits_last_stage_spec_info_folded_hist_hist_1_folded_hist; // @[Frontend.scala 69:19]
  wire [7:0] ftq_io_fromBpu_resp_bits_last_stage_spec_info_folded_hist_hist_0_folded_hist; // @[Frontend.scala 69:19]
  wire  ftq_io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_5_bits_0; // @[Frontend.scala 69:19]
  wire  ftq_io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_5_bits_1; // @[Frontend.scala 69:19]
  wire  ftq_io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_5_bits_2; // @[Frontend.scala 69:19]
  wire  ftq_io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_5_bits_3; // @[Frontend.scala 69:19]
  wire  ftq_io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_4_bits_0; // @[Frontend.scala 69:19]
  wire  ftq_io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_4_bits_1; // @[Frontend.scala 69:19]
  wire  ftq_io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_4_bits_2; // @[Frontend.scala 69:19]
  wire  ftq_io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_4_bits_3; // @[Frontend.scala 69:19]
  wire  ftq_io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_3_bits_0; // @[Frontend.scala 69:19]
  wire  ftq_io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_3_bits_1; // @[Frontend.scala 69:19]
  wire  ftq_io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_3_bits_2; // @[Frontend.scala 69:19]
  wire  ftq_io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_3_bits_3; // @[Frontend.scala 69:19]
  wire  ftq_io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_2_bits_0; // @[Frontend.scala 69:19]
  wire  ftq_io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_2_bits_1; // @[Frontend.scala 69:19]
  wire  ftq_io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_2_bits_2; // @[Frontend.scala 69:19]
  wire  ftq_io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_2_bits_3; // @[Frontend.scala 69:19]
  wire  ftq_io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_1_bits_0; // @[Frontend.scala 69:19]
  wire  ftq_io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_1_bits_1; // @[Frontend.scala 69:19]
  wire  ftq_io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_1_bits_2; // @[Frontend.scala 69:19]
  wire  ftq_io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_1_bits_3; // @[Frontend.scala 69:19]
  wire  ftq_io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_0_bits_0; // @[Frontend.scala 69:19]
  wire  ftq_io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_0_bits_1; // @[Frontend.scala 69:19]
  wire  ftq_io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_0_bits_2; // @[Frontend.scala 69:19]
  wire  ftq_io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_0_bits_3; // @[Frontend.scala 69:19]
  wire [2:0] ftq_io_fromBpu_resp_bits_last_stage_spec_info_lastBrNumOH; // @[Frontend.scala 69:19]
  wire  ftq_io_fromBpu_resp_bits_last_stage_spec_info_histPtr_flag; // @[Frontend.scala 69:19]
  wire [7:0] ftq_io_fromBpu_resp_bits_last_stage_spec_info_histPtr_value; // @[Frontend.scala 69:19]
  wire [4:0] ftq_io_fromBpu_resp_bits_last_stage_spec_info_rasSp; // @[Frontend.scala 69:19]
  wire [38:0] ftq_io_fromBpu_resp_bits_last_stage_spec_info_rasTop_retAddr; // @[Frontend.scala 69:19]
  wire [7:0] ftq_io_fromBpu_resp_bits_last_stage_spec_info_rasTop_ctr; // @[Frontend.scala 69:19]
  wire  ftq_io_fromBpu_resp_bits_last_stage_ftb_entry_valid; // @[Frontend.scala 69:19]
  wire [2:0] ftq_io_fromBpu_resp_bits_last_stage_ftb_entry_brSlots_0_offset; // @[Frontend.scala 69:19]
  wire [11:0] ftq_io_fromBpu_resp_bits_last_stage_ftb_entry_brSlots_0_lower; // @[Frontend.scala 69:19]
  wire [1:0] ftq_io_fromBpu_resp_bits_last_stage_ftb_entry_brSlots_0_tarStat; // @[Frontend.scala 69:19]
  wire  ftq_io_fromBpu_resp_bits_last_stage_ftb_entry_brSlots_0_sharing; // @[Frontend.scala 69:19]
  wire  ftq_io_fromBpu_resp_bits_last_stage_ftb_entry_brSlots_0_valid; // @[Frontend.scala 69:19]
  wire [2:0] ftq_io_fromBpu_resp_bits_last_stage_ftb_entry_tailSlot_offset; // @[Frontend.scala 69:19]
  wire [19:0] ftq_io_fromBpu_resp_bits_last_stage_ftb_entry_tailSlot_lower; // @[Frontend.scala 69:19]
  wire [1:0] ftq_io_fromBpu_resp_bits_last_stage_ftb_entry_tailSlot_tarStat; // @[Frontend.scala 69:19]
  wire  ftq_io_fromBpu_resp_bits_last_stage_ftb_entry_tailSlot_sharing; // @[Frontend.scala 69:19]
  wire  ftq_io_fromBpu_resp_bits_last_stage_ftb_entry_tailSlot_valid; // @[Frontend.scala 69:19]
  wire [2:0] ftq_io_fromBpu_resp_bits_last_stage_ftb_entry_pftAddr; // @[Frontend.scala 69:19]
  wire  ftq_io_fromBpu_resp_bits_last_stage_ftb_entry_carry; // @[Frontend.scala 69:19]
  wire  ftq_io_fromBpu_resp_bits_last_stage_ftb_entry_isCall; // @[Frontend.scala 69:19]
  wire  ftq_io_fromBpu_resp_bits_last_stage_ftb_entry_isRet; // @[Frontend.scala 69:19]
  wire  ftq_io_fromBpu_resp_bits_last_stage_ftb_entry_isJalr; // @[Frontend.scala 69:19]
  wire  ftq_io_fromBpu_resp_bits_last_stage_ftb_entry_last_may_be_rvi_call; // @[Frontend.scala 69:19]
  wire  ftq_io_fromBpu_resp_bits_last_stage_ftb_entry_always_taken_0; // @[Frontend.scala 69:19]
  wire  ftq_io_fromBpu_resp_bits_last_stage_ftb_entry_always_taken_1; // @[Frontend.scala 69:19]
  wire  ftq_io_fromIfu_pdWb_valid; // @[Frontend.scala 69:19]
  wire [38:0] ftq_io_fromIfu_pdWb_bits_pc_0; // @[Frontend.scala 69:19]
  wire [38:0] ftq_io_fromIfu_pdWb_bits_pc_1; // @[Frontend.scala 69:19]
  wire [38:0] ftq_io_fromIfu_pdWb_bits_pc_2; // @[Frontend.scala 69:19]
  wire [38:0] ftq_io_fromIfu_pdWb_bits_pc_3; // @[Frontend.scala 69:19]
  wire [38:0] ftq_io_fromIfu_pdWb_bits_pc_4; // @[Frontend.scala 69:19]
  wire [38:0] ftq_io_fromIfu_pdWb_bits_pc_5; // @[Frontend.scala 69:19]
  wire [38:0] ftq_io_fromIfu_pdWb_bits_pc_6; // @[Frontend.scala 69:19]
  wire [38:0] ftq_io_fromIfu_pdWb_bits_pc_7; // @[Frontend.scala 69:19]
  wire  ftq_io_fromIfu_pdWb_bits_pd_0_valid; // @[Frontend.scala 69:19]
  wire  ftq_io_fromIfu_pdWb_bits_pd_0_isRVC; // @[Frontend.scala 69:19]
  wire [1:0] ftq_io_fromIfu_pdWb_bits_pd_0_brType; // @[Frontend.scala 69:19]
  wire  ftq_io_fromIfu_pdWb_bits_pd_0_isCall; // @[Frontend.scala 69:19]
  wire  ftq_io_fromIfu_pdWb_bits_pd_0_isRet; // @[Frontend.scala 69:19]
  wire  ftq_io_fromIfu_pdWb_bits_pd_1_valid; // @[Frontend.scala 69:19]
  wire  ftq_io_fromIfu_pdWb_bits_pd_1_isRVC; // @[Frontend.scala 69:19]
  wire [1:0] ftq_io_fromIfu_pdWb_bits_pd_1_brType; // @[Frontend.scala 69:19]
  wire  ftq_io_fromIfu_pdWb_bits_pd_1_isCall; // @[Frontend.scala 69:19]
  wire  ftq_io_fromIfu_pdWb_bits_pd_1_isRet; // @[Frontend.scala 69:19]
  wire  ftq_io_fromIfu_pdWb_bits_pd_2_valid; // @[Frontend.scala 69:19]
  wire  ftq_io_fromIfu_pdWb_bits_pd_2_isRVC; // @[Frontend.scala 69:19]
  wire [1:0] ftq_io_fromIfu_pdWb_bits_pd_2_brType; // @[Frontend.scala 69:19]
  wire  ftq_io_fromIfu_pdWb_bits_pd_2_isCall; // @[Frontend.scala 69:19]
  wire  ftq_io_fromIfu_pdWb_bits_pd_2_isRet; // @[Frontend.scala 69:19]
  wire  ftq_io_fromIfu_pdWb_bits_pd_3_valid; // @[Frontend.scala 69:19]
  wire  ftq_io_fromIfu_pdWb_bits_pd_3_isRVC; // @[Frontend.scala 69:19]
  wire [1:0] ftq_io_fromIfu_pdWb_bits_pd_3_brType; // @[Frontend.scala 69:19]
  wire  ftq_io_fromIfu_pdWb_bits_pd_3_isCall; // @[Frontend.scala 69:19]
  wire  ftq_io_fromIfu_pdWb_bits_pd_3_isRet; // @[Frontend.scala 69:19]
  wire  ftq_io_fromIfu_pdWb_bits_pd_4_valid; // @[Frontend.scala 69:19]
  wire  ftq_io_fromIfu_pdWb_bits_pd_4_isRVC; // @[Frontend.scala 69:19]
  wire [1:0] ftq_io_fromIfu_pdWb_bits_pd_4_brType; // @[Frontend.scala 69:19]
  wire  ftq_io_fromIfu_pdWb_bits_pd_4_isCall; // @[Frontend.scala 69:19]
  wire  ftq_io_fromIfu_pdWb_bits_pd_4_isRet; // @[Frontend.scala 69:19]
  wire  ftq_io_fromIfu_pdWb_bits_pd_5_valid; // @[Frontend.scala 69:19]
  wire  ftq_io_fromIfu_pdWb_bits_pd_5_isRVC; // @[Frontend.scala 69:19]
  wire [1:0] ftq_io_fromIfu_pdWb_bits_pd_5_brType; // @[Frontend.scala 69:19]
  wire  ftq_io_fromIfu_pdWb_bits_pd_5_isCall; // @[Frontend.scala 69:19]
  wire  ftq_io_fromIfu_pdWb_bits_pd_5_isRet; // @[Frontend.scala 69:19]
  wire  ftq_io_fromIfu_pdWb_bits_pd_6_valid; // @[Frontend.scala 69:19]
  wire  ftq_io_fromIfu_pdWb_bits_pd_6_isRVC; // @[Frontend.scala 69:19]
  wire [1:0] ftq_io_fromIfu_pdWb_bits_pd_6_brType; // @[Frontend.scala 69:19]
  wire  ftq_io_fromIfu_pdWb_bits_pd_6_isCall; // @[Frontend.scala 69:19]
  wire  ftq_io_fromIfu_pdWb_bits_pd_6_isRet; // @[Frontend.scala 69:19]
  wire  ftq_io_fromIfu_pdWb_bits_pd_7_valid; // @[Frontend.scala 69:19]
  wire  ftq_io_fromIfu_pdWb_bits_pd_7_isRVC; // @[Frontend.scala 69:19]
  wire [1:0] ftq_io_fromIfu_pdWb_bits_pd_7_brType; // @[Frontend.scala 69:19]
  wire  ftq_io_fromIfu_pdWb_bits_pd_7_isCall; // @[Frontend.scala 69:19]
  wire  ftq_io_fromIfu_pdWb_bits_pd_7_isRet; // @[Frontend.scala 69:19]
  wire  ftq_io_fromIfu_pdWb_bits_ftqIdx_flag; // @[Frontend.scala 69:19]
  wire [2:0] ftq_io_fromIfu_pdWb_bits_ftqIdx_value; // @[Frontend.scala 69:19]
  wire  ftq_io_fromIfu_pdWb_bits_misOffset_valid; // @[Frontend.scala 69:19]
  wire [2:0] ftq_io_fromIfu_pdWb_bits_misOffset_bits; // @[Frontend.scala 69:19]
  wire  ftq_io_fromIfu_pdWb_bits_cfiOffset_valid; // @[Frontend.scala 69:19]
  wire [38:0] ftq_io_fromIfu_pdWb_bits_target; // @[Frontend.scala 69:19]
  wire [38:0] ftq_io_fromIfu_pdWb_bits_jalTarget; // @[Frontend.scala 69:19]
  wire  ftq_io_fromIfu_pdWb_bits_instrRange_0; // @[Frontend.scala 69:19]
  wire  ftq_io_fromIfu_pdWb_bits_instrRange_1; // @[Frontend.scala 69:19]
  wire  ftq_io_fromIfu_pdWb_bits_instrRange_2; // @[Frontend.scala 69:19]
  wire  ftq_io_fromIfu_pdWb_bits_instrRange_3; // @[Frontend.scala 69:19]
  wire  ftq_io_fromIfu_pdWb_bits_instrRange_4; // @[Frontend.scala 69:19]
  wire  ftq_io_fromIfu_pdWb_bits_instrRange_5; // @[Frontend.scala 69:19]
  wire  ftq_io_fromIfu_pdWb_bits_instrRange_6; // @[Frontend.scala 69:19]
  wire  ftq_io_fromIfu_pdWb_bits_instrRange_7; // @[Frontend.scala 69:19]
  wire  ftq_io_fromBackend_rob_commits_0_valid; // @[Frontend.scala 69:19]
  wire [2:0] ftq_io_fromBackend_rob_commits_0_bits_commitType; // @[Frontend.scala 69:19]
  wire  ftq_io_fromBackend_rob_commits_0_bits_ftqIdx_flag; // @[Frontend.scala 69:19]
  wire [2:0] ftq_io_fromBackend_rob_commits_0_bits_ftqIdx_value; // @[Frontend.scala 69:19]
  wire [2:0] ftq_io_fromBackend_rob_commits_0_bits_ftqOffset; // @[Frontend.scala 69:19]
  wire  ftq_io_fromBackend_rob_commits_1_valid; // @[Frontend.scala 69:19]
  wire [2:0] ftq_io_fromBackend_rob_commits_1_bits_commitType; // @[Frontend.scala 69:19]
  wire  ftq_io_fromBackend_rob_commits_1_bits_ftqIdx_flag; // @[Frontend.scala 69:19]
  wire [2:0] ftq_io_fromBackend_rob_commits_1_bits_ftqIdx_value; // @[Frontend.scala 69:19]
  wire [2:0] ftq_io_fromBackend_rob_commits_1_bits_ftqOffset; // @[Frontend.scala 69:19]
  wire  ftq_io_fromBackend_redirect_valid; // @[Frontend.scala 69:19]
  wire  ftq_io_fromBackend_redirect_bits_ftqIdx_flag; // @[Frontend.scala 69:19]
  wire [2:0] ftq_io_fromBackend_redirect_bits_ftqIdx_value; // @[Frontend.scala 69:19]
  wire [2:0] ftq_io_fromBackend_redirect_bits_ftqOffset; // @[Frontend.scala 69:19]
  wire  ftq_io_fromBackend_redirect_bits_level; // @[Frontend.scala 69:19]
  wire [38:0] ftq_io_fromBackend_redirect_bits_cfiUpdate_pc; // @[Frontend.scala 69:19]
  wire  ftq_io_fromBackend_redirect_bits_cfiUpdate_pd_isRVC; // @[Frontend.scala 69:19]
  wire [1:0] ftq_io_fromBackend_redirect_bits_cfiUpdate_pd_brType; // @[Frontend.scala 69:19]
  wire  ftq_io_fromBackend_redirect_bits_cfiUpdate_pd_isCall; // @[Frontend.scala 69:19]
  wire  ftq_io_fromBackend_redirect_bits_cfiUpdate_pd_isRet; // @[Frontend.scala 69:19]
  wire [38:0] ftq_io_fromBackend_redirect_bits_cfiUpdate_target; // @[Frontend.scala 69:19]
  wire  ftq_io_fromBackend_redirect_bits_cfiUpdate_taken; // @[Frontend.scala 69:19]
  wire  ftq_io_fromBackend_redirect_bits_cfiUpdate_isMisPred; // @[Frontend.scala 69:19]
  wire  ftq_io_toBpu_redirect_valid; // @[Frontend.scala 69:19]
  wire  ftq_io_toBpu_redirect_bits_level; // @[Frontend.scala 69:19]
  wire [38:0] ftq_io_toBpu_redirect_bits_cfiUpdate_pc; // @[Frontend.scala 69:19]
  wire  ftq_io_toBpu_redirect_bits_cfiUpdate_pd_isRVC; // @[Frontend.scala 69:19]
  wire  ftq_io_toBpu_redirect_bits_cfiUpdate_pd_isCall; // @[Frontend.scala 69:19]
  wire  ftq_io_toBpu_redirect_bits_cfiUpdate_pd_isRet; // @[Frontend.scala 69:19]
  wire [4:0] ftq_io_toBpu_redirect_bits_cfiUpdate_rasSp; // @[Frontend.scala 69:19]
  wire [38:0] ftq_io_toBpu_redirect_bits_cfiUpdate_rasEntry_retAddr; // @[Frontend.scala 69:19]
  wire [7:0] ftq_io_toBpu_redirect_bits_cfiUpdate_rasEntry_ctr; // @[Frontend.scala 69:19]
  wire [7:0] ftq_io_toBpu_redirect_bits_cfiUpdate_folded_hist_hist_17_folded_hist; // @[Frontend.scala 69:19]
  wire [7:0] ftq_io_toBpu_redirect_bits_cfiUpdate_folded_hist_hist_16_folded_hist; // @[Frontend.scala 69:19]
  wire [10:0] ftq_io_toBpu_redirect_bits_cfiUpdate_folded_hist_hist_15_folded_hist; // @[Frontend.scala 69:19]
  wire [6:0] ftq_io_toBpu_redirect_bits_cfiUpdate_folded_hist_hist_14_folded_hist; // @[Frontend.scala 69:19]
  wire [6:0] ftq_io_toBpu_redirect_bits_cfiUpdate_folded_hist_hist_13_folded_hist; // @[Frontend.scala 69:19]
  wire [6:0] ftq_io_toBpu_redirect_bits_cfiUpdate_folded_hist_hist_12_folded_hist; // @[Frontend.scala 69:19]
  wire [7:0] ftq_io_toBpu_redirect_bits_cfiUpdate_folded_hist_hist_11_folded_hist; // @[Frontend.scala 69:19]
  wire [8:0] ftq_io_toBpu_redirect_bits_cfiUpdate_folded_hist_hist_10_folded_hist; // @[Frontend.scala 69:19]
  wire [6:0] ftq_io_toBpu_redirect_bits_cfiUpdate_folded_hist_hist_9_folded_hist; // @[Frontend.scala 69:19]
  wire [7:0] ftq_io_toBpu_redirect_bits_cfiUpdate_folded_hist_hist_8_folded_hist; // @[Frontend.scala 69:19]
  wire [8:0] ftq_io_toBpu_redirect_bits_cfiUpdate_folded_hist_hist_7_folded_hist; // @[Frontend.scala 69:19]
  wire [8:0] ftq_io_toBpu_redirect_bits_cfiUpdate_folded_hist_hist_6_folded_hist; // @[Frontend.scala 69:19]
  wire [10:0] ftq_io_toBpu_redirect_bits_cfiUpdate_folded_hist_hist_5_folded_hist; // @[Frontend.scala 69:19]
  wire [3:0] ftq_io_toBpu_redirect_bits_cfiUpdate_folded_hist_hist_4_folded_hist; // @[Frontend.scala 69:19]
  wire [10:0] ftq_io_toBpu_redirect_bits_cfiUpdate_folded_hist_hist_3_folded_hist; // @[Frontend.scala 69:19]
  wire [7:0] ftq_io_toBpu_redirect_bits_cfiUpdate_folded_hist_hist_2_folded_hist; // @[Frontend.scala 69:19]
  wire [7:0] ftq_io_toBpu_redirect_bits_cfiUpdate_folded_hist_hist_1_folded_hist; // @[Frontend.scala 69:19]
  wire [7:0] ftq_io_toBpu_redirect_bits_cfiUpdate_folded_hist_hist_0_folded_hist; // @[Frontend.scala 69:19]
  wire  ftq_io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_5_bits_0; // @[Frontend.scala 69:19]
  wire  ftq_io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_5_bits_1; // @[Frontend.scala 69:19]
  wire  ftq_io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_5_bits_2; // @[Frontend.scala 69:19]
  wire  ftq_io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_5_bits_3; // @[Frontend.scala 69:19]
  wire  ftq_io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_4_bits_0; // @[Frontend.scala 69:19]
  wire  ftq_io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_4_bits_1; // @[Frontend.scala 69:19]
  wire  ftq_io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_4_bits_2; // @[Frontend.scala 69:19]
  wire  ftq_io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_3_bits_0; // @[Frontend.scala 69:19]
  wire  ftq_io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_3_bits_1; // @[Frontend.scala 69:19]
  wire  ftq_io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_3_bits_2; // @[Frontend.scala 69:19]
  wire  ftq_io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_3_bits_3; // @[Frontend.scala 69:19]
  wire  ftq_io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_2_bits_0; // @[Frontend.scala 69:19]
  wire  ftq_io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_2_bits_1; // @[Frontend.scala 69:19]
  wire  ftq_io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_2_bits_2; // @[Frontend.scala 69:19]
  wire  ftq_io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_2_bits_3; // @[Frontend.scala 69:19]
  wire  ftq_io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_1_bits_0; // @[Frontend.scala 69:19]
  wire  ftq_io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_1_bits_1; // @[Frontend.scala 69:19]
  wire  ftq_io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_1_bits_2; // @[Frontend.scala 69:19]
  wire  ftq_io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_1_bits_3; // @[Frontend.scala 69:19]
  wire  ftq_io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_0_bits_0; // @[Frontend.scala 69:19]
  wire  ftq_io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_0_bits_1; // @[Frontend.scala 69:19]
  wire  ftq_io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_0_bits_2; // @[Frontend.scala 69:19]
  wire  ftq_io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_0_bits_3; // @[Frontend.scala 69:19]
  wire [2:0] ftq_io_toBpu_redirect_bits_cfiUpdate_lastBrNumOH; // @[Frontend.scala 69:19]
  wire  ftq_io_toBpu_redirect_bits_cfiUpdate_histPtr_flag; // @[Frontend.scala 69:19]
  wire [7:0] ftq_io_toBpu_redirect_bits_cfiUpdate_histPtr_value; // @[Frontend.scala 69:19]
  wire [38:0] ftq_io_toBpu_redirect_bits_cfiUpdate_target; // @[Frontend.scala 69:19]
  wire  ftq_io_toBpu_redirect_bits_cfiUpdate_taken; // @[Frontend.scala 69:19]
  wire [1:0] ftq_io_toBpu_redirect_bits_cfiUpdate_shift; // @[Frontend.scala 69:19]
  wire  ftq_io_toBpu_redirect_bits_cfiUpdate_addIntoHist; // @[Frontend.scala 69:19]
  wire  ftq_io_toBpu_update_valid; // @[Frontend.scala 69:19]
  wire [38:0] ftq_io_toBpu_update_bits_pc; // @[Frontend.scala 69:19]
  wire [7:0] ftq_io_toBpu_update_bits_spec_info_folded_hist_hist_17_folded_hist; // @[Frontend.scala 69:19]
  wire [7:0] ftq_io_toBpu_update_bits_spec_info_folded_hist_hist_16_folded_hist; // @[Frontend.scala 69:19]
  wire [10:0] ftq_io_toBpu_update_bits_spec_info_folded_hist_hist_15_folded_hist; // @[Frontend.scala 69:19]
  wire [6:0] ftq_io_toBpu_update_bits_spec_info_folded_hist_hist_14_folded_hist; // @[Frontend.scala 69:19]
  wire [6:0] ftq_io_toBpu_update_bits_spec_info_folded_hist_hist_13_folded_hist; // @[Frontend.scala 69:19]
  wire [6:0] ftq_io_toBpu_update_bits_spec_info_folded_hist_hist_12_folded_hist; // @[Frontend.scala 69:19]
  wire [8:0] ftq_io_toBpu_update_bits_spec_info_folded_hist_hist_10_folded_hist; // @[Frontend.scala 69:19]
  wire [6:0] ftq_io_toBpu_update_bits_spec_info_folded_hist_hist_9_folded_hist; // @[Frontend.scala 69:19]
  wire [7:0] ftq_io_toBpu_update_bits_spec_info_folded_hist_hist_8_folded_hist; // @[Frontend.scala 69:19]
  wire [8:0] ftq_io_toBpu_update_bits_spec_info_folded_hist_hist_7_folded_hist; // @[Frontend.scala 69:19]
  wire [8:0] ftq_io_toBpu_update_bits_spec_info_folded_hist_hist_6_folded_hist; // @[Frontend.scala 69:19]
  wire [10:0] ftq_io_toBpu_update_bits_spec_info_folded_hist_hist_5_folded_hist; // @[Frontend.scala 69:19]
  wire [3:0] ftq_io_toBpu_update_bits_spec_info_folded_hist_hist_4_folded_hist; // @[Frontend.scala 69:19]
  wire [10:0] ftq_io_toBpu_update_bits_spec_info_folded_hist_hist_3_folded_hist; // @[Frontend.scala 69:19]
  wire [7:0] ftq_io_toBpu_update_bits_spec_info_folded_hist_hist_2_folded_hist; // @[Frontend.scala 69:19]
  wire [7:0] ftq_io_toBpu_update_bits_spec_info_folded_hist_hist_1_folded_hist; // @[Frontend.scala 69:19]
  wire [7:0] ftq_io_toBpu_update_bits_spec_info_folded_hist_hist_0_folded_hist; // @[Frontend.scala 69:19]
  wire  ftq_io_toBpu_update_bits_ftb_entry_valid; // @[Frontend.scala 69:19]
  wire [2:0] ftq_io_toBpu_update_bits_ftb_entry_brSlots_0_offset; // @[Frontend.scala 69:19]
  wire [11:0] ftq_io_toBpu_update_bits_ftb_entry_brSlots_0_lower; // @[Frontend.scala 69:19]
  wire [1:0] ftq_io_toBpu_update_bits_ftb_entry_brSlots_0_tarStat; // @[Frontend.scala 69:19]
  wire  ftq_io_toBpu_update_bits_ftb_entry_brSlots_0_sharing; // @[Frontend.scala 69:19]
  wire  ftq_io_toBpu_update_bits_ftb_entry_brSlots_0_valid; // @[Frontend.scala 69:19]
  wire [2:0] ftq_io_toBpu_update_bits_ftb_entry_tailSlot_offset; // @[Frontend.scala 69:19]
  wire [19:0] ftq_io_toBpu_update_bits_ftb_entry_tailSlot_lower; // @[Frontend.scala 69:19]
  wire [1:0] ftq_io_toBpu_update_bits_ftb_entry_tailSlot_tarStat; // @[Frontend.scala 69:19]
  wire  ftq_io_toBpu_update_bits_ftb_entry_tailSlot_sharing; // @[Frontend.scala 69:19]
  wire  ftq_io_toBpu_update_bits_ftb_entry_tailSlot_valid; // @[Frontend.scala 69:19]
  wire [2:0] ftq_io_toBpu_update_bits_ftb_entry_pftAddr; // @[Frontend.scala 69:19]
  wire  ftq_io_toBpu_update_bits_ftb_entry_carry; // @[Frontend.scala 69:19]
  wire  ftq_io_toBpu_update_bits_ftb_entry_isCall; // @[Frontend.scala 69:19]
  wire  ftq_io_toBpu_update_bits_ftb_entry_isRet; // @[Frontend.scala 69:19]
  wire  ftq_io_toBpu_update_bits_ftb_entry_isJalr; // @[Frontend.scala 69:19]
  wire  ftq_io_toBpu_update_bits_ftb_entry_last_may_be_rvi_call; // @[Frontend.scala 69:19]
  wire  ftq_io_toBpu_update_bits_ftb_entry_always_taken_0; // @[Frontend.scala 69:19]
  wire  ftq_io_toBpu_update_bits_ftb_entry_always_taken_1; // @[Frontend.scala 69:19]
  wire  ftq_io_toBpu_update_bits_br_taken_mask_0; // @[Frontend.scala 69:19]
  wire  ftq_io_toBpu_update_bits_br_taken_mask_1; // @[Frontend.scala 69:19]
  wire  ftq_io_toBpu_update_bits_jmp_taken; // @[Frontend.scala 69:19]
  wire  ftq_io_toBpu_update_bits_mispred_mask_0; // @[Frontend.scala 69:19]
  wire  ftq_io_toBpu_update_bits_mispred_mask_1; // @[Frontend.scala 69:19]
  wire  ftq_io_toBpu_update_bits_mispred_mask_2; // @[Frontend.scala 69:19]
  wire  ftq_io_toBpu_update_bits_false_hit; // @[Frontend.scala 69:19]
  wire  ftq_io_toBpu_update_bits_old_entry; // @[Frontend.scala 69:19]
  wire [255:0] ftq_io_toBpu_update_bits_meta; // @[Frontend.scala 69:19]
  wire [38:0] ftq_io_toBpu_update_bits_full_target; // @[Frontend.scala 69:19]
  wire  ftq_io_toBpu_enq_ptr_flag; // @[Frontend.scala 69:19]
  wire [2:0] ftq_io_toBpu_enq_ptr_value; // @[Frontend.scala 69:19]
  wire  ftq_io_toIfu_req_ready; // @[Frontend.scala 69:19]
  wire  ftq_io_toIfu_req_valid; // @[Frontend.scala 69:19]
  wire [38:0] ftq_io_toIfu_req_bits_startAddr; // @[Frontend.scala 69:19]
  wire [38:0] ftq_io_toIfu_req_bits_nextlineStart; // @[Frontend.scala 69:19]
  wire [38:0] ftq_io_toIfu_req_bits_nextStartAddr; // @[Frontend.scala 69:19]
  wire  ftq_io_toIfu_req_bits_ftqIdx_flag; // @[Frontend.scala 69:19]
  wire [2:0] ftq_io_toIfu_req_bits_ftqIdx_value; // @[Frontend.scala 69:19]
  wire  ftq_io_toIfu_req_bits_ftqOffset_valid; // @[Frontend.scala 69:19]
  wire [2:0] ftq_io_toIfu_req_bits_ftqOffset_bits; // @[Frontend.scala 69:19]
  wire  ftq_io_toIfu_redirect_valid; // @[Frontend.scala 69:19]
  wire  ftq_io_toIfu_redirect_bits_ftqIdx_flag; // @[Frontend.scala 69:19]
  wire [2:0] ftq_io_toIfu_redirect_bits_ftqIdx_value; // @[Frontend.scala 69:19]
  wire [2:0] ftq_io_toIfu_redirect_bits_ftqOffset; // @[Frontend.scala 69:19]
  wire  ftq_io_toIfu_redirect_bits_level; // @[Frontend.scala 69:19]
  wire  ftq_io_toIfu_flushFromBpu_s2_valid; // @[Frontend.scala 69:19]
  wire  ftq_io_toIfu_flushFromBpu_s2_bits_flag; // @[Frontend.scala 69:19]
  wire [2:0] ftq_io_toIfu_flushFromBpu_s2_bits_value; // @[Frontend.scala 69:19]
  wire  ftq_io_toIfu_flushFromBpu_s3_valid; // @[Frontend.scala 69:19]
  wire  ftq_io_toIfu_flushFromBpu_s3_bits_flag; // @[Frontend.scala 69:19]
  wire [2:0] ftq_io_toIfu_flushFromBpu_s3_bits_value; // @[Frontend.scala 69:19]
  wire  ftq_io_toICache_req_valid; // @[Frontend.scala 69:19]
  wire [38:0] ftq_io_toICache_req_bits_pcMemRead_0_startAddr; // @[Frontend.scala 69:19]
  wire [38:0] ftq_io_toICache_req_bits_pcMemRead_0_nextlineStart; // @[Frontend.scala 69:19]
  wire [38:0] ftq_io_toICache_req_bits_pcMemRead_1_startAddr; // @[Frontend.scala 69:19]
  wire [38:0] ftq_io_toICache_req_bits_pcMemRead_1_nextlineStart; // @[Frontend.scala 69:19]
  wire [38:0] ftq_io_toICache_req_bits_pcMemRead_2_startAddr; // @[Frontend.scala 69:19]
  wire [38:0] ftq_io_toICache_req_bits_pcMemRead_2_nextlineStart; // @[Frontend.scala 69:19]
  wire [38:0] ftq_io_toICache_req_bits_pcMemRead_3_startAddr; // @[Frontend.scala 69:19]
  wire [38:0] ftq_io_toICache_req_bits_pcMemRead_3_nextlineStart; // @[Frontend.scala 69:19]
  wire [38:0] ftq_io_toICache_req_bits_pcMemRead_4_startAddr; // @[Frontend.scala 69:19]
  wire [38:0] ftq_io_toICache_req_bits_pcMemRead_4_nextlineStart; // @[Frontend.scala 69:19]
  wire  ftq_io_toICache_req_bits_readValid_0; // @[Frontend.scala 69:19]
  wire  ftq_io_toICache_req_bits_readValid_1; // @[Frontend.scala 69:19]
  wire  ftq_io_toICache_req_bits_readValid_2; // @[Frontend.scala 69:19]
  wire  ftq_io_toICache_req_bits_readValid_3; // @[Frontend.scala 69:19]
  wire  ftq_io_toICache_req_bits_readValid_4; // @[Frontend.scala 69:19]
  wire  ftq_io_toBackend_pc_mem_wen; // @[Frontend.scala 69:19]
  wire [2:0] ftq_io_toBackend_pc_mem_waddr; // @[Frontend.scala 69:19]
  wire [38:0] ftq_io_toBackend_pc_mem_wdata_startAddr; // @[Frontend.scala 69:19]
  wire [38:0] ftq_io_toBackend_pc_mem_wdata_nextLineAddr; // @[Frontend.scala 69:19]
  wire  ftq_io_toBackend_pc_mem_wdata_isNextMask_0; // @[Frontend.scala 69:19]
  wire  ftq_io_toBackend_pc_mem_wdata_isNextMask_1; // @[Frontend.scala 69:19]
  wire  ftq_io_toBackend_pc_mem_wdata_isNextMask_2; // @[Frontend.scala 69:19]
  wire  ftq_io_toBackend_pc_mem_wdata_isNextMask_3; // @[Frontend.scala 69:19]
  wire  ftq_io_toBackend_pc_mem_wdata_isNextMask_4; // @[Frontend.scala 69:19]
  wire  ftq_io_toBackend_pc_mem_wdata_isNextMask_5; // @[Frontend.scala 69:19]
  wire  ftq_io_toBackend_pc_mem_wdata_isNextMask_6; // @[Frontend.scala 69:19]
  wire  ftq_io_toBackend_pc_mem_wdata_isNextMask_7; // @[Frontend.scala 69:19]
  wire [38:0] ftq_io_toBackend_newest_entry_target; // @[Frontend.scala 69:19]
  wire  ftq_io_toBackend_newest_entry_ptr_flag; // @[Frontend.scala 69:19]
  wire [2:0] ftq_io_toBackend_newest_entry_ptr_value; // @[Frontend.scala 69:19]
  wire  ftq_io_mmioCommitRead_mmioFtqPtr_flag; // @[Frontend.scala 69:19]
  wire [2:0] ftq_io_mmioCommitRead_mmioFtqPtr_value; // @[Frontend.scala 69:19]
  wire  ftq_io_mmioCommitRead_mmioLastCommit; // @[Frontend.scala 69:19]
  wire [5:0] ftq_io_perf_0_value; // @[Frontend.scala 69:19]
  wire [5:0] ftq_io_perf_1_value; // @[Frontend.scala 69:19]
  wire [5:0] ftq_io_perf_2_value; // @[Frontend.scala 69:19]
  wire [5:0] ftq_io_perf_3_value; // @[Frontend.scala 69:19]
  wire [5:0] ftq_io_perf_4_value; // @[Frontend.scala 69:19]
  wire [5:0] ftq_io_perf_5_value; // @[Frontend.scala 69:19]
  wire [5:0] ftq_io_perf_6_value; // @[Frontend.scala 69:19]
  wire [5:0] ftq_io_perf_7_value; // @[Frontend.scala 69:19]
  wire [5:0] ftq_io_perf_8_value; // @[Frontend.scala 69:19]
  wire [5:0] ftq_io_perf_9_value; // @[Frontend.scala 69:19]
  wire [5:0] ftq_io_perf_10_value; // @[Frontend.scala 69:19]
  wire [5:0] ftq_io_perf_11_value; // @[Frontend.scala 69:19]
  wire [5:0] ftq_io_perf_12_value; // @[Frontend.scala 69:19]
  wire [5:0] ftq_io_perf_13_value; // @[Frontend.scala 69:19]
  wire [5:0] ftq_io_perf_14_value; // @[Frontend.scala 69:19]
  wire [5:0] ftq_io_perf_15_value; // @[Frontend.scala 69:19]
  wire [5:0] ftq_io_perf_16_value; // @[Frontend.scala 69:19]
  wire [5:0] ftq_io_perf_17_value; // @[Frontend.scala 69:19]
  wire [5:0] ftq_io_perf_18_value; // @[Frontend.scala 69:19]
  wire [5:0] ftq_io_perf_19_value; // @[Frontend.scala 69:19]
  wire [5:0] ftq_io_perf_20_value; // @[Frontend.scala 69:19]
  wire [5:0] ftq_io_perf_21_value; // @[Frontend.scala 69:19]
  wire [5:0] ftq_io_perf_22_value; // @[Frontend.scala 69:19]
  wire [5:0] ftq_io_perf_23_value; // @[Frontend.scala 69:19]
  wire  tlbCsr_delay_clock; // @[Hold.scala 97:23]
  wire [3:0] tlbCsr_delay_io_in_satp_mode; // @[Hold.scala 97:23]
  wire [15:0] tlbCsr_delay_io_in_satp_asid; // @[Hold.scala 97:23]
  wire [43:0] tlbCsr_delay_io_in_satp_ppn; // @[Hold.scala 97:23]
  wire  tlbCsr_delay_io_in_satp_changed; // @[Hold.scala 97:23]
  wire  tlbCsr_delay_io_in_priv_mxr; // @[Hold.scala 97:23]
  wire  tlbCsr_delay_io_in_priv_sum; // @[Hold.scala 97:23]
  wire [1:0] tlbCsr_delay_io_in_priv_imode; // @[Hold.scala 97:23]
  wire [1:0] tlbCsr_delay_io_in_priv_dmode; // @[Hold.scala 97:23]
  wire [3:0] tlbCsr_delay_io_out_satp_mode; // @[Hold.scala 97:23]
  wire [15:0] tlbCsr_delay_io_out_satp_asid; // @[Hold.scala 97:23]
  wire [43:0] tlbCsr_delay_io_out_satp_ppn; // @[Hold.scala 97:23]
  wire  tlbCsr_delay_io_out_satp_changed; // @[Hold.scala 97:23]
  wire  tlbCsr_delay_io_out_priv_mxr; // @[Hold.scala 97:23]
  wire  tlbCsr_delay_io_out_priv_sum; // @[Hold.scala 97:23]
  wire [1:0] tlbCsr_delay_io_out_priv_imode; // @[Hold.scala 97:23]
  wire [1:0] tlbCsr_delay_io_out_priv_dmode; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_clock; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_in_icache_parity_enable; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_in_lvpred_disable; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_in_no_spec_load; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_in_storeset_wait_store; // @[Hold.scala 97:23]
  wire [4:0] csrCtrl_delay_io_in_lvpred_timeout; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_in_bp_ctrl_ubtb_enable; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_in_bp_ctrl_btb_enable; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_in_bp_ctrl_tage_enable; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_in_bp_ctrl_sc_enable; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_in_bp_ctrl_ras_enable; // @[Hold.scala 97:23]
  wire [3:0] csrCtrl_delay_io_in_sbuffer_threshold; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_in_ldld_vio_check_enable; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_in_cache_error_enable; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_in_uncache_write_outstanding_enable; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_in_fusion_enable; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_in_wfi_enable; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_in_svinval_enable; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_in_distribute_csr_wvalid; // @[Hold.scala 97:23]
  wire [11:0] csrCtrl_delay_io_in_distribute_csr_waddr; // @[Hold.scala 97:23]
  wire [63:0] csrCtrl_delay_io_in_distribute_csr_wdata; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_in_singlestep; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_in_frontend_trigger_t_valid; // @[Hold.scala 97:23]
  wire [1:0] csrCtrl_delay_io_in_frontend_trigger_t_bits_addr; // @[Hold.scala 97:23]
  wire [1:0] csrCtrl_delay_io_in_frontend_trigger_t_bits_tdata_matchType; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_in_frontend_trigger_t_bits_tdata_select; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_in_frontend_trigger_t_bits_tdata_timing; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_in_frontend_trigger_t_bits_tdata_chain; // @[Hold.scala 97:23]
  wire [63:0] csrCtrl_delay_io_in_frontend_trigger_t_bits_tdata_tdata2; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_in_mem_trigger_t_valid; // @[Hold.scala 97:23]
  wire [2:0] csrCtrl_delay_io_in_mem_trigger_t_bits_addr; // @[Hold.scala 97:23]
  wire [1:0] csrCtrl_delay_io_in_mem_trigger_t_bits_tdata_matchType; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_in_mem_trigger_t_bits_tdata_select; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_in_mem_trigger_t_bits_tdata_chain; // @[Hold.scala 97:23]
  wire [63:0] csrCtrl_delay_io_in_mem_trigger_t_bits_tdata_tdata2; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_in_trigger_enable_0; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_in_trigger_enable_1; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_in_trigger_enable_2; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_in_trigger_enable_3; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_in_trigger_enable_4; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_in_trigger_enable_5; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_in_trigger_enable_6; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_in_trigger_enable_7; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_in_trigger_enable_8; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_in_trigger_enable_9; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_out_icache_parity_enable; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_out_lvpred_disable; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_out_no_spec_load; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_out_storeset_wait_store; // @[Hold.scala 97:23]
  wire [4:0] csrCtrl_delay_io_out_lvpred_timeout; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_out_bp_ctrl_ubtb_enable; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_out_bp_ctrl_btb_enable; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_out_bp_ctrl_tage_enable; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_out_bp_ctrl_sc_enable; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_out_bp_ctrl_ras_enable; // @[Hold.scala 97:23]
  wire [3:0] csrCtrl_delay_io_out_sbuffer_threshold; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_out_ldld_vio_check_enable; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_out_cache_error_enable; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_out_uncache_write_outstanding_enable; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_out_fusion_enable; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_out_wfi_enable; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_out_svinval_enable; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_out_distribute_csr_wvalid; // @[Hold.scala 97:23]
  wire [11:0] csrCtrl_delay_io_out_distribute_csr_waddr; // @[Hold.scala 97:23]
  wire [63:0] csrCtrl_delay_io_out_distribute_csr_wdata; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_out_singlestep; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_out_frontend_trigger_t_valid; // @[Hold.scala 97:23]
  wire [1:0] csrCtrl_delay_io_out_frontend_trigger_t_bits_addr; // @[Hold.scala 97:23]
  wire [1:0] csrCtrl_delay_io_out_frontend_trigger_t_bits_tdata_matchType; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_out_frontend_trigger_t_bits_tdata_select; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_out_frontend_trigger_t_bits_tdata_timing; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_out_frontend_trigger_t_bits_tdata_chain; // @[Hold.scala 97:23]
  wire [63:0] csrCtrl_delay_io_out_frontend_trigger_t_bits_tdata_tdata2; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_out_mem_trigger_t_valid; // @[Hold.scala 97:23]
  wire [2:0] csrCtrl_delay_io_out_mem_trigger_t_bits_addr; // @[Hold.scala 97:23]
  wire [1:0] csrCtrl_delay_io_out_mem_trigger_t_bits_tdata_matchType; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_out_mem_trigger_t_bits_tdata_select; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_out_mem_trigger_t_bits_tdata_chain; // @[Hold.scala 97:23]
  wire [63:0] csrCtrl_delay_io_out_mem_trigger_t_bits_tdata_tdata2; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_out_trigger_enable_0; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_out_trigger_enable_1; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_out_trigger_enable_2; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_out_trigger_enable_3; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_out_trigger_enable_4; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_out_trigger_enable_5; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_out_trigger_enable_6; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_out_trigger_enable_7; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_out_trigger_enable_8; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_out_trigger_enable_9; // @[Hold.scala 97:23]
  wire  pmp_clock; // @[Frontend.scala 87:19]
  wire  pmp_reset; // @[Frontend.scala 87:19]
  wire  pmp_io_distribute_csr_wvalid; // @[Frontend.scala 87:19]
  wire [11:0] pmp_io_distribute_csr_waddr; // @[Frontend.scala 87:19]
  wire [63:0] pmp_io_distribute_csr_wdata; // @[Frontend.scala 87:19]
  wire  pmp_io_pmp_0_cfg_l; // @[Frontend.scala 87:19]
  wire [1:0] pmp_io_pmp_0_cfg_a; // @[Frontend.scala 87:19]
  wire  pmp_io_pmp_0_cfg_x; // @[Frontend.scala 87:19]
  wire  pmp_io_pmp_0_cfg_w; // @[Frontend.scala 87:19]
  wire  pmp_io_pmp_0_cfg_r; // @[Frontend.scala 87:19]
  wire [33:0] pmp_io_pmp_0_addr; // @[Frontend.scala 87:19]
  wire [35:0] pmp_io_pmp_0_mask; // @[Frontend.scala 87:19]
  wire  pmp_io_pmp_1_cfg_l; // @[Frontend.scala 87:19]
  wire [1:0] pmp_io_pmp_1_cfg_a; // @[Frontend.scala 87:19]
  wire  pmp_io_pmp_1_cfg_x; // @[Frontend.scala 87:19]
  wire  pmp_io_pmp_1_cfg_w; // @[Frontend.scala 87:19]
  wire  pmp_io_pmp_1_cfg_r; // @[Frontend.scala 87:19]
  wire [33:0] pmp_io_pmp_1_addr; // @[Frontend.scala 87:19]
  wire [35:0] pmp_io_pmp_1_mask; // @[Frontend.scala 87:19]
  wire  pmp_io_pmp_2_cfg_l; // @[Frontend.scala 87:19]
  wire [1:0] pmp_io_pmp_2_cfg_a; // @[Frontend.scala 87:19]
  wire  pmp_io_pmp_2_cfg_x; // @[Frontend.scala 87:19]
  wire  pmp_io_pmp_2_cfg_w; // @[Frontend.scala 87:19]
  wire  pmp_io_pmp_2_cfg_r; // @[Frontend.scala 87:19]
  wire [33:0] pmp_io_pmp_2_addr; // @[Frontend.scala 87:19]
  wire [35:0] pmp_io_pmp_2_mask; // @[Frontend.scala 87:19]
  wire  pmp_io_pmp_3_cfg_l; // @[Frontend.scala 87:19]
  wire [1:0] pmp_io_pmp_3_cfg_a; // @[Frontend.scala 87:19]
  wire  pmp_io_pmp_3_cfg_x; // @[Frontend.scala 87:19]
  wire  pmp_io_pmp_3_cfg_w; // @[Frontend.scala 87:19]
  wire  pmp_io_pmp_3_cfg_r; // @[Frontend.scala 87:19]
  wire [33:0] pmp_io_pmp_3_addr; // @[Frontend.scala 87:19]
  wire [35:0] pmp_io_pmp_3_mask; // @[Frontend.scala 87:19]
  wire  pmp_io_pmp_4_cfg_l; // @[Frontend.scala 87:19]
  wire [1:0] pmp_io_pmp_4_cfg_a; // @[Frontend.scala 87:19]
  wire  pmp_io_pmp_4_cfg_x; // @[Frontend.scala 87:19]
  wire  pmp_io_pmp_4_cfg_w; // @[Frontend.scala 87:19]
  wire  pmp_io_pmp_4_cfg_r; // @[Frontend.scala 87:19]
  wire [33:0] pmp_io_pmp_4_addr; // @[Frontend.scala 87:19]
  wire [35:0] pmp_io_pmp_4_mask; // @[Frontend.scala 87:19]
  wire  pmp_io_pmp_5_cfg_l; // @[Frontend.scala 87:19]
  wire [1:0] pmp_io_pmp_5_cfg_a; // @[Frontend.scala 87:19]
  wire  pmp_io_pmp_5_cfg_x; // @[Frontend.scala 87:19]
  wire  pmp_io_pmp_5_cfg_w; // @[Frontend.scala 87:19]
  wire  pmp_io_pmp_5_cfg_r; // @[Frontend.scala 87:19]
  wire [33:0] pmp_io_pmp_5_addr; // @[Frontend.scala 87:19]
  wire [35:0] pmp_io_pmp_5_mask; // @[Frontend.scala 87:19]
  wire  pmp_io_pmp_6_cfg_l; // @[Frontend.scala 87:19]
  wire [1:0] pmp_io_pmp_6_cfg_a; // @[Frontend.scala 87:19]
  wire  pmp_io_pmp_6_cfg_x; // @[Frontend.scala 87:19]
  wire  pmp_io_pmp_6_cfg_w; // @[Frontend.scala 87:19]
  wire  pmp_io_pmp_6_cfg_r; // @[Frontend.scala 87:19]
  wire [33:0] pmp_io_pmp_6_addr; // @[Frontend.scala 87:19]
  wire [35:0] pmp_io_pmp_6_mask; // @[Frontend.scala 87:19]
  wire  pmp_io_pmp_7_cfg_l; // @[Frontend.scala 87:19]
  wire [1:0] pmp_io_pmp_7_cfg_a; // @[Frontend.scala 87:19]
  wire  pmp_io_pmp_7_cfg_x; // @[Frontend.scala 87:19]
  wire  pmp_io_pmp_7_cfg_w; // @[Frontend.scala 87:19]
  wire  pmp_io_pmp_7_cfg_r; // @[Frontend.scala 87:19]
  wire [33:0] pmp_io_pmp_7_addr; // @[Frontend.scala 87:19]
  wire [35:0] pmp_io_pmp_7_mask; // @[Frontend.scala 87:19]
  wire  pmp_io_pmp_8_cfg_l; // @[Frontend.scala 87:19]
  wire [1:0] pmp_io_pmp_8_cfg_a; // @[Frontend.scala 87:19]
  wire  pmp_io_pmp_8_cfg_x; // @[Frontend.scala 87:19]
  wire  pmp_io_pmp_8_cfg_w; // @[Frontend.scala 87:19]
  wire  pmp_io_pmp_8_cfg_r; // @[Frontend.scala 87:19]
  wire [33:0] pmp_io_pmp_8_addr; // @[Frontend.scala 87:19]
  wire [35:0] pmp_io_pmp_8_mask; // @[Frontend.scala 87:19]
  wire  pmp_io_pmp_9_cfg_l; // @[Frontend.scala 87:19]
  wire [1:0] pmp_io_pmp_9_cfg_a; // @[Frontend.scala 87:19]
  wire  pmp_io_pmp_9_cfg_x; // @[Frontend.scala 87:19]
  wire  pmp_io_pmp_9_cfg_w; // @[Frontend.scala 87:19]
  wire  pmp_io_pmp_9_cfg_r; // @[Frontend.scala 87:19]
  wire [33:0] pmp_io_pmp_9_addr; // @[Frontend.scala 87:19]
  wire [35:0] pmp_io_pmp_9_mask; // @[Frontend.scala 87:19]
  wire  pmp_io_pmp_10_cfg_l; // @[Frontend.scala 87:19]
  wire [1:0] pmp_io_pmp_10_cfg_a; // @[Frontend.scala 87:19]
  wire  pmp_io_pmp_10_cfg_x; // @[Frontend.scala 87:19]
  wire  pmp_io_pmp_10_cfg_w; // @[Frontend.scala 87:19]
  wire  pmp_io_pmp_10_cfg_r; // @[Frontend.scala 87:19]
  wire [33:0] pmp_io_pmp_10_addr; // @[Frontend.scala 87:19]
  wire [35:0] pmp_io_pmp_10_mask; // @[Frontend.scala 87:19]
  wire  pmp_io_pmp_11_cfg_l; // @[Frontend.scala 87:19]
  wire [1:0] pmp_io_pmp_11_cfg_a; // @[Frontend.scala 87:19]
  wire  pmp_io_pmp_11_cfg_x; // @[Frontend.scala 87:19]
  wire  pmp_io_pmp_11_cfg_w; // @[Frontend.scala 87:19]
  wire  pmp_io_pmp_11_cfg_r; // @[Frontend.scala 87:19]
  wire [33:0] pmp_io_pmp_11_addr; // @[Frontend.scala 87:19]
  wire [35:0] pmp_io_pmp_11_mask; // @[Frontend.scala 87:19]
  wire  pmp_io_pmp_12_cfg_l; // @[Frontend.scala 87:19]
  wire [1:0] pmp_io_pmp_12_cfg_a; // @[Frontend.scala 87:19]
  wire  pmp_io_pmp_12_cfg_x; // @[Frontend.scala 87:19]
  wire  pmp_io_pmp_12_cfg_w; // @[Frontend.scala 87:19]
  wire  pmp_io_pmp_12_cfg_r; // @[Frontend.scala 87:19]
  wire [33:0] pmp_io_pmp_12_addr; // @[Frontend.scala 87:19]
  wire [35:0] pmp_io_pmp_12_mask; // @[Frontend.scala 87:19]
  wire  pmp_io_pmp_13_cfg_l; // @[Frontend.scala 87:19]
  wire [1:0] pmp_io_pmp_13_cfg_a; // @[Frontend.scala 87:19]
  wire  pmp_io_pmp_13_cfg_x; // @[Frontend.scala 87:19]
  wire  pmp_io_pmp_13_cfg_w; // @[Frontend.scala 87:19]
  wire  pmp_io_pmp_13_cfg_r; // @[Frontend.scala 87:19]
  wire [33:0] pmp_io_pmp_13_addr; // @[Frontend.scala 87:19]
  wire [35:0] pmp_io_pmp_13_mask; // @[Frontend.scala 87:19]
  wire  pmp_io_pmp_14_cfg_l; // @[Frontend.scala 87:19]
  wire [1:0] pmp_io_pmp_14_cfg_a; // @[Frontend.scala 87:19]
  wire  pmp_io_pmp_14_cfg_x; // @[Frontend.scala 87:19]
  wire  pmp_io_pmp_14_cfg_w; // @[Frontend.scala 87:19]
  wire  pmp_io_pmp_14_cfg_r; // @[Frontend.scala 87:19]
  wire [33:0] pmp_io_pmp_14_addr; // @[Frontend.scala 87:19]
  wire [35:0] pmp_io_pmp_14_mask; // @[Frontend.scala 87:19]
  wire  pmp_io_pmp_15_cfg_l; // @[Frontend.scala 87:19]
  wire [1:0] pmp_io_pmp_15_cfg_a; // @[Frontend.scala 87:19]
  wire  pmp_io_pmp_15_cfg_x; // @[Frontend.scala 87:19]
  wire  pmp_io_pmp_15_cfg_w; // @[Frontend.scala 87:19]
  wire  pmp_io_pmp_15_cfg_r; // @[Frontend.scala 87:19]
  wire [33:0] pmp_io_pmp_15_addr; // @[Frontend.scala 87:19]
  wire [35:0] pmp_io_pmp_15_mask; // @[Frontend.scala 87:19]
  wire  pmp_io_pma_0_cfg_c; // @[Frontend.scala 87:19]
  wire  pmp_io_pma_0_cfg_atomic; // @[Frontend.scala 87:19]
  wire [1:0] pmp_io_pma_0_cfg_a; // @[Frontend.scala 87:19]
  wire  pmp_io_pma_0_cfg_x; // @[Frontend.scala 87:19]
  wire  pmp_io_pma_0_cfg_w; // @[Frontend.scala 87:19]
  wire  pmp_io_pma_0_cfg_r; // @[Frontend.scala 87:19]
  wire [33:0] pmp_io_pma_0_addr; // @[Frontend.scala 87:19]
  wire [35:0] pmp_io_pma_0_mask; // @[Frontend.scala 87:19]
  wire  pmp_io_pma_1_cfg_c; // @[Frontend.scala 87:19]
  wire  pmp_io_pma_1_cfg_atomic; // @[Frontend.scala 87:19]
  wire [1:0] pmp_io_pma_1_cfg_a; // @[Frontend.scala 87:19]
  wire  pmp_io_pma_1_cfg_x; // @[Frontend.scala 87:19]
  wire  pmp_io_pma_1_cfg_w; // @[Frontend.scala 87:19]
  wire  pmp_io_pma_1_cfg_r; // @[Frontend.scala 87:19]
  wire [33:0] pmp_io_pma_1_addr; // @[Frontend.scala 87:19]
  wire [35:0] pmp_io_pma_1_mask; // @[Frontend.scala 87:19]
  wire  pmp_io_pma_2_cfg_c; // @[Frontend.scala 87:19]
  wire  pmp_io_pma_2_cfg_atomic; // @[Frontend.scala 87:19]
  wire [1:0] pmp_io_pma_2_cfg_a; // @[Frontend.scala 87:19]
  wire  pmp_io_pma_2_cfg_x; // @[Frontend.scala 87:19]
  wire  pmp_io_pma_2_cfg_w; // @[Frontend.scala 87:19]
  wire  pmp_io_pma_2_cfg_r; // @[Frontend.scala 87:19]
  wire [33:0] pmp_io_pma_2_addr; // @[Frontend.scala 87:19]
  wire [35:0] pmp_io_pma_2_mask; // @[Frontend.scala 87:19]
  wire  pmp_io_pma_3_cfg_c; // @[Frontend.scala 87:19]
  wire  pmp_io_pma_3_cfg_atomic; // @[Frontend.scala 87:19]
  wire [1:0] pmp_io_pma_3_cfg_a; // @[Frontend.scala 87:19]
  wire  pmp_io_pma_3_cfg_x; // @[Frontend.scala 87:19]
  wire  pmp_io_pma_3_cfg_w; // @[Frontend.scala 87:19]
  wire  pmp_io_pma_3_cfg_r; // @[Frontend.scala 87:19]
  wire [33:0] pmp_io_pma_3_addr; // @[Frontend.scala 87:19]
  wire [35:0] pmp_io_pma_3_mask; // @[Frontend.scala 87:19]
  wire  pmp_io_pma_4_cfg_c; // @[Frontend.scala 87:19]
  wire  pmp_io_pma_4_cfg_atomic; // @[Frontend.scala 87:19]
  wire [1:0] pmp_io_pma_4_cfg_a; // @[Frontend.scala 87:19]
  wire  pmp_io_pma_4_cfg_x; // @[Frontend.scala 87:19]
  wire  pmp_io_pma_4_cfg_w; // @[Frontend.scala 87:19]
  wire  pmp_io_pma_4_cfg_r; // @[Frontend.scala 87:19]
  wire [33:0] pmp_io_pma_4_addr; // @[Frontend.scala 87:19]
  wire [35:0] pmp_io_pma_4_mask; // @[Frontend.scala 87:19]
  wire  pmp_io_pma_5_cfg_c; // @[Frontend.scala 87:19]
  wire  pmp_io_pma_5_cfg_atomic; // @[Frontend.scala 87:19]
  wire [1:0] pmp_io_pma_5_cfg_a; // @[Frontend.scala 87:19]
  wire  pmp_io_pma_5_cfg_x; // @[Frontend.scala 87:19]
  wire  pmp_io_pma_5_cfg_w; // @[Frontend.scala 87:19]
  wire  pmp_io_pma_5_cfg_r; // @[Frontend.scala 87:19]
  wire [33:0] pmp_io_pma_5_addr; // @[Frontend.scala 87:19]
  wire [35:0] pmp_io_pma_5_mask; // @[Frontend.scala 87:19]
  wire  pmp_io_pma_6_cfg_c; // @[Frontend.scala 87:19]
  wire  pmp_io_pma_6_cfg_atomic; // @[Frontend.scala 87:19]
  wire [1:0] pmp_io_pma_6_cfg_a; // @[Frontend.scala 87:19]
  wire  pmp_io_pma_6_cfg_x; // @[Frontend.scala 87:19]
  wire  pmp_io_pma_6_cfg_w; // @[Frontend.scala 87:19]
  wire  pmp_io_pma_6_cfg_r; // @[Frontend.scala 87:19]
  wire [33:0] pmp_io_pma_6_addr; // @[Frontend.scala 87:19]
  wire [35:0] pmp_io_pma_6_mask; // @[Frontend.scala 87:19]
  wire  pmp_io_pma_7_cfg_c; // @[Frontend.scala 87:19]
  wire  pmp_io_pma_7_cfg_atomic; // @[Frontend.scala 87:19]
  wire [1:0] pmp_io_pma_7_cfg_a; // @[Frontend.scala 87:19]
  wire  pmp_io_pma_7_cfg_x; // @[Frontend.scala 87:19]
  wire  pmp_io_pma_7_cfg_w; // @[Frontend.scala 87:19]
  wire  pmp_io_pma_7_cfg_r; // @[Frontend.scala 87:19]
  wire [33:0] pmp_io_pma_7_addr; // @[Frontend.scala 87:19]
  wire [35:0] pmp_io_pma_7_mask; // @[Frontend.scala 87:19]
  wire  pmp_io_pma_8_cfg_c; // @[Frontend.scala 87:19]
  wire  pmp_io_pma_8_cfg_atomic; // @[Frontend.scala 87:19]
  wire [1:0] pmp_io_pma_8_cfg_a; // @[Frontend.scala 87:19]
  wire  pmp_io_pma_8_cfg_x; // @[Frontend.scala 87:19]
  wire  pmp_io_pma_8_cfg_w; // @[Frontend.scala 87:19]
  wire  pmp_io_pma_8_cfg_r; // @[Frontend.scala 87:19]
  wire [33:0] pmp_io_pma_8_addr; // @[Frontend.scala 87:19]
  wire [35:0] pmp_io_pma_8_mask; // @[Frontend.scala 87:19]
  wire  pmp_io_pma_9_cfg_c; // @[Frontend.scala 87:19]
  wire  pmp_io_pma_9_cfg_atomic; // @[Frontend.scala 87:19]
  wire [1:0] pmp_io_pma_9_cfg_a; // @[Frontend.scala 87:19]
  wire  pmp_io_pma_9_cfg_x; // @[Frontend.scala 87:19]
  wire  pmp_io_pma_9_cfg_w; // @[Frontend.scala 87:19]
  wire  pmp_io_pma_9_cfg_r; // @[Frontend.scala 87:19]
  wire [33:0] pmp_io_pma_9_addr; // @[Frontend.scala 87:19]
  wire [35:0] pmp_io_pma_9_mask; // @[Frontend.scala 87:19]
  wire  pmp_io_pma_10_cfg_c; // @[Frontend.scala 87:19]
  wire  pmp_io_pma_10_cfg_atomic; // @[Frontend.scala 87:19]
  wire [1:0] pmp_io_pma_10_cfg_a; // @[Frontend.scala 87:19]
  wire  pmp_io_pma_10_cfg_x; // @[Frontend.scala 87:19]
  wire  pmp_io_pma_10_cfg_w; // @[Frontend.scala 87:19]
  wire  pmp_io_pma_10_cfg_r; // @[Frontend.scala 87:19]
  wire [33:0] pmp_io_pma_10_addr; // @[Frontend.scala 87:19]
  wire [35:0] pmp_io_pma_10_mask; // @[Frontend.scala 87:19]
  wire  pmp_io_pma_11_cfg_c; // @[Frontend.scala 87:19]
  wire  pmp_io_pma_11_cfg_atomic; // @[Frontend.scala 87:19]
  wire [1:0] pmp_io_pma_11_cfg_a; // @[Frontend.scala 87:19]
  wire  pmp_io_pma_11_cfg_x; // @[Frontend.scala 87:19]
  wire  pmp_io_pma_11_cfg_w; // @[Frontend.scala 87:19]
  wire  pmp_io_pma_11_cfg_r; // @[Frontend.scala 87:19]
  wire [33:0] pmp_io_pma_11_addr; // @[Frontend.scala 87:19]
  wire [35:0] pmp_io_pma_11_mask; // @[Frontend.scala 87:19]
  wire  pmp_io_pma_12_cfg_c; // @[Frontend.scala 87:19]
  wire  pmp_io_pma_12_cfg_atomic; // @[Frontend.scala 87:19]
  wire [1:0] pmp_io_pma_12_cfg_a; // @[Frontend.scala 87:19]
  wire  pmp_io_pma_12_cfg_x; // @[Frontend.scala 87:19]
  wire  pmp_io_pma_12_cfg_w; // @[Frontend.scala 87:19]
  wire  pmp_io_pma_12_cfg_r; // @[Frontend.scala 87:19]
  wire [33:0] pmp_io_pma_12_addr; // @[Frontend.scala 87:19]
  wire [35:0] pmp_io_pma_12_mask; // @[Frontend.scala 87:19]
  wire  pmp_io_pma_13_cfg_c; // @[Frontend.scala 87:19]
  wire  pmp_io_pma_13_cfg_atomic; // @[Frontend.scala 87:19]
  wire [1:0] pmp_io_pma_13_cfg_a; // @[Frontend.scala 87:19]
  wire  pmp_io_pma_13_cfg_x; // @[Frontend.scala 87:19]
  wire  pmp_io_pma_13_cfg_w; // @[Frontend.scala 87:19]
  wire  pmp_io_pma_13_cfg_r; // @[Frontend.scala 87:19]
  wire [33:0] pmp_io_pma_13_addr; // @[Frontend.scala 87:19]
  wire [35:0] pmp_io_pma_13_mask; // @[Frontend.scala 87:19]
  wire  pmp_io_pma_14_cfg_c; // @[Frontend.scala 87:19]
  wire  pmp_io_pma_14_cfg_atomic; // @[Frontend.scala 87:19]
  wire [1:0] pmp_io_pma_14_cfg_a; // @[Frontend.scala 87:19]
  wire  pmp_io_pma_14_cfg_x; // @[Frontend.scala 87:19]
  wire  pmp_io_pma_14_cfg_w; // @[Frontend.scala 87:19]
  wire  pmp_io_pma_14_cfg_r; // @[Frontend.scala 87:19]
  wire [33:0] pmp_io_pma_14_addr; // @[Frontend.scala 87:19]
  wire [35:0] pmp_io_pma_14_mask; // @[Frontend.scala 87:19]
  wire  pmp_io_pma_15_cfg_c; // @[Frontend.scala 87:19]
  wire  pmp_io_pma_15_cfg_atomic; // @[Frontend.scala 87:19]
  wire [1:0] pmp_io_pma_15_cfg_a; // @[Frontend.scala 87:19]
  wire  pmp_io_pma_15_cfg_x; // @[Frontend.scala 87:19]
  wire  pmp_io_pma_15_cfg_w; // @[Frontend.scala 87:19]
  wire  pmp_io_pma_15_cfg_r; // @[Frontend.scala 87:19]
  wire [33:0] pmp_io_pma_15_addr; // @[Frontend.scala 87:19]
  wire [35:0] pmp_io_pma_15_mask; // @[Frontend.scala 87:19]
  wire [1:0] PMPChecker_io_check_env_mode; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pmp_0_cfg_l; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_io_check_env_pmp_0_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pmp_0_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pmp_0_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pmp_0_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_io_check_env_pmp_0_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_io_check_env_pmp_0_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pmp_1_cfg_l; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_io_check_env_pmp_1_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pmp_1_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pmp_1_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pmp_1_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_io_check_env_pmp_1_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_io_check_env_pmp_1_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pmp_2_cfg_l; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_io_check_env_pmp_2_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pmp_2_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pmp_2_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pmp_2_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_io_check_env_pmp_2_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_io_check_env_pmp_2_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pmp_3_cfg_l; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_io_check_env_pmp_3_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pmp_3_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pmp_3_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pmp_3_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_io_check_env_pmp_3_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_io_check_env_pmp_3_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pmp_4_cfg_l; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_io_check_env_pmp_4_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pmp_4_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pmp_4_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pmp_4_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_io_check_env_pmp_4_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_io_check_env_pmp_4_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pmp_5_cfg_l; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_io_check_env_pmp_5_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pmp_5_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pmp_5_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pmp_5_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_io_check_env_pmp_5_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_io_check_env_pmp_5_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pmp_6_cfg_l; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_io_check_env_pmp_6_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pmp_6_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pmp_6_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pmp_6_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_io_check_env_pmp_6_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_io_check_env_pmp_6_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pmp_7_cfg_l; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_io_check_env_pmp_7_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pmp_7_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pmp_7_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pmp_7_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_io_check_env_pmp_7_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_io_check_env_pmp_7_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pmp_8_cfg_l; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_io_check_env_pmp_8_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pmp_8_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pmp_8_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pmp_8_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_io_check_env_pmp_8_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_io_check_env_pmp_8_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pmp_9_cfg_l; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_io_check_env_pmp_9_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pmp_9_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pmp_9_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pmp_9_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_io_check_env_pmp_9_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_io_check_env_pmp_9_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pmp_10_cfg_l; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_io_check_env_pmp_10_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pmp_10_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pmp_10_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pmp_10_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_io_check_env_pmp_10_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_io_check_env_pmp_10_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pmp_11_cfg_l; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_io_check_env_pmp_11_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pmp_11_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pmp_11_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pmp_11_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_io_check_env_pmp_11_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_io_check_env_pmp_11_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pmp_12_cfg_l; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_io_check_env_pmp_12_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pmp_12_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pmp_12_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pmp_12_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_io_check_env_pmp_12_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_io_check_env_pmp_12_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pmp_13_cfg_l; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_io_check_env_pmp_13_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pmp_13_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pmp_13_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pmp_13_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_io_check_env_pmp_13_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_io_check_env_pmp_13_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pmp_14_cfg_l; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_io_check_env_pmp_14_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pmp_14_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pmp_14_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pmp_14_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_io_check_env_pmp_14_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_io_check_env_pmp_14_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pmp_15_cfg_l; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_io_check_env_pmp_15_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pmp_15_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pmp_15_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pmp_15_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_io_check_env_pmp_15_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_io_check_env_pmp_15_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pma_0_cfg_c; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pma_0_cfg_atomic; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_io_check_env_pma_0_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pma_0_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pma_0_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pma_0_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_io_check_env_pma_0_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_io_check_env_pma_0_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pma_1_cfg_c; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pma_1_cfg_atomic; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_io_check_env_pma_1_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pma_1_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pma_1_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pma_1_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_io_check_env_pma_1_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_io_check_env_pma_1_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pma_2_cfg_c; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pma_2_cfg_atomic; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_io_check_env_pma_2_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pma_2_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pma_2_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pma_2_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_io_check_env_pma_2_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_io_check_env_pma_2_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pma_3_cfg_c; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pma_3_cfg_atomic; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_io_check_env_pma_3_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pma_3_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pma_3_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pma_3_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_io_check_env_pma_3_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_io_check_env_pma_3_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pma_4_cfg_c; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pma_4_cfg_atomic; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_io_check_env_pma_4_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pma_4_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pma_4_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pma_4_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_io_check_env_pma_4_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_io_check_env_pma_4_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pma_5_cfg_c; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pma_5_cfg_atomic; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_io_check_env_pma_5_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pma_5_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pma_5_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pma_5_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_io_check_env_pma_5_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_io_check_env_pma_5_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pma_6_cfg_c; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pma_6_cfg_atomic; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_io_check_env_pma_6_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pma_6_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pma_6_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pma_6_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_io_check_env_pma_6_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_io_check_env_pma_6_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pma_7_cfg_c; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pma_7_cfg_atomic; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_io_check_env_pma_7_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pma_7_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pma_7_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pma_7_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_io_check_env_pma_7_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_io_check_env_pma_7_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pma_8_cfg_c; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pma_8_cfg_atomic; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_io_check_env_pma_8_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pma_8_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pma_8_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pma_8_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_io_check_env_pma_8_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_io_check_env_pma_8_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pma_9_cfg_c; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pma_9_cfg_atomic; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_io_check_env_pma_9_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pma_9_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pma_9_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pma_9_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_io_check_env_pma_9_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_io_check_env_pma_9_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pma_10_cfg_c; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pma_10_cfg_atomic; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_io_check_env_pma_10_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pma_10_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pma_10_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pma_10_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_io_check_env_pma_10_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_io_check_env_pma_10_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pma_11_cfg_c; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pma_11_cfg_atomic; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_io_check_env_pma_11_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pma_11_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pma_11_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pma_11_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_io_check_env_pma_11_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_io_check_env_pma_11_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pma_12_cfg_c; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pma_12_cfg_atomic; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_io_check_env_pma_12_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pma_12_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pma_12_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pma_12_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_io_check_env_pma_12_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_io_check_env_pma_12_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pma_13_cfg_c; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pma_13_cfg_atomic; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_io_check_env_pma_13_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pma_13_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pma_13_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pma_13_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_io_check_env_pma_13_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_io_check_env_pma_13_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pma_14_cfg_c; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pma_14_cfg_atomic; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_io_check_env_pma_14_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pma_14_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pma_14_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pma_14_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_io_check_env_pma_14_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_io_check_env_pma_14_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pma_15_cfg_c; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pma_15_cfg_atomic; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_io_check_env_pma_15_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pma_15_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pma_15_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_check_env_pma_15_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_io_check_env_pma_15_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_io_check_env_pma_15_mask; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_io_req_bits_addr; // @[Frontend.scala 88:45]
  wire [2:0] PMPChecker_io_req_bits_cmd; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_resp_ld; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_resp_st; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_resp_instr; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_resp_mmio; // @[Frontend.scala 88:45]
  wire  PMPChecker_io_resp_atomic; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_1_io_check_env_mode; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pmp_0_cfg_l; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_1_io_check_env_pmp_0_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pmp_0_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pmp_0_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pmp_0_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_1_io_check_env_pmp_0_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_1_io_check_env_pmp_0_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pmp_1_cfg_l; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_1_io_check_env_pmp_1_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pmp_1_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pmp_1_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pmp_1_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_1_io_check_env_pmp_1_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_1_io_check_env_pmp_1_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pmp_2_cfg_l; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_1_io_check_env_pmp_2_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pmp_2_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pmp_2_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pmp_2_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_1_io_check_env_pmp_2_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_1_io_check_env_pmp_2_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pmp_3_cfg_l; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_1_io_check_env_pmp_3_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pmp_3_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pmp_3_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pmp_3_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_1_io_check_env_pmp_3_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_1_io_check_env_pmp_3_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pmp_4_cfg_l; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_1_io_check_env_pmp_4_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pmp_4_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pmp_4_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pmp_4_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_1_io_check_env_pmp_4_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_1_io_check_env_pmp_4_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pmp_5_cfg_l; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_1_io_check_env_pmp_5_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pmp_5_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pmp_5_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pmp_5_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_1_io_check_env_pmp_5_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_1_io_check_env_pmp_5_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pmp_6_cfg_l; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_1_io_check_env_pmp_6_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pmp_6_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pmp_6_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pmp_6_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_1_io_check_env_pmp_6_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_1_io_check_env_pmp_6_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pmp_7_cfg_l; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_1_io_check_env_pmp_7_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pmp_7_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pmp_7_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pmp_7_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_1_io_check_env_pmp_7_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_1_io_check_env_pmp_7_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pmp_8_cfg_l; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_1_io_check_env_pmp_8_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pmp_8_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pmp_8_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pmp_8_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_1_io_check_env_pmp_8_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_1_io_check_env_pmp_8_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pmp_9_cfg_l; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_1_io_check_env_pmp_9_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pmp_9_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pmp_9_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pmp_9_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_1_io_check_env_pmp_9_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_1_io_check_env_pmp_9_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pmp_10_cfg_l; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_1_io_check_env_pmp_10_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pmp_10_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pmp_10_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pmp_10_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_1_io_check_env_pmp_10_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_1_io_check_env_pmp_10_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pmp_11_cfg_l; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_1_io_check_env_pmp_11_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pmp_11_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pmp_11_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pmp_11_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_1_io_check_env_pmp_11_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_1_io_check_env_pmp_11_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pmp_12_cfg_l; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_1_io_check_env_pmp_12_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pmp_12_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pmp_12_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pmp_12_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_1_io_check_env_pmp_12_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_1_io_check_env_pmp_12_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pmp_13_cfg_l; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_1_io_check_env_pmp_13_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pmp_13_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pmp_13_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pmp_13_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_1_io_check_env_pmp_13_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_1_io_check_env_pmp_13_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pmp_14_cfg_l; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_1_io_check_env_pmp_14_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pmp_14_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pmp_14_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pmp_14_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_1_io_check_env_pmp_14_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_1_io_check_env_pmp_14_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pmp_15_cfg_l; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_1_io_check_env_pmp_15_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pmp_15_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pmp_15_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pmp_15_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_1_io_check_env_pmp_15_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_1_io_check_env_pmp_15_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pma_0_cfg_c; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pma_0_cfg_atomic; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_1_io_check_env_pma_0_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pma_0_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pma_0_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pma_0_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_1_io_check_env_pma_0_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_1_io_check_env_pma_0_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pma_1_cfg_c; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pma_1_cfg_atomic; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_1_io_check_env_pma_1_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pma_1_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pma_1_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pma_1_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_1_io_check_env_pma_1_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_1_io_check_env_pma_1_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pma_2_cfg_c; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pma_2_cfg_atomic; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_1_io_check_env_pma_2_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pma_2_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pma_2_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pma_2_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_1_io_check_env_pma_2_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_1_io_check_env_pma_2_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pma_3_cfg_c; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pma_3_cfg_atomic; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_1_io_check_env_pma_3_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pma_3_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pma_3_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pma_3_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_1_io_check_env_pma_3_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_1_io_check_env_pma_3_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pma_4_cfg_c; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pma_4_cfg_atomic; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_1_io_check_env_pma_4_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pma_4_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pma_4_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pma_4_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_1_io_check_env_pma_4_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_1_io_check_env_pma_4_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pma_5_cfg_c; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pma_5_cfg_atomic; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_1_io_check_env_pma_5_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pma_5_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pma_5_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pma_5_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_1_io_check_env_pma_5_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_1_io_check_env_pma_5_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pma_6_cfg_c; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pma_6_cfg_atomic; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_1_io_check_env_pma_6_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pma_6_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pma_6_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pma_6_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_1_io_check_env_pma_6_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_1_io_check_env_pma_6_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pma_7_cfg_c; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pma_7_cfg_atomic; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_1_io_check_env_pma_7_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pma_7_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pma_7_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pma_7_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_1_io_check_env_pma_7_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_1_io_check_env_pma_7_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pma_8_cfg_c; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pma_8_cfg_atomic; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_1_io_check_env_pma_8_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pma_8_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pma_8_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pma_8_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_1_io_check_env_pma_8_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_1_io_check_env_pma_8_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pma_9_cfg_c; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pma_9_cfg_atomic; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_1_io_check_env_pma_9_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pma_9_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pma_9_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pma_9_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_1_io_check_env_pma_9_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_1_io_check_env_pma_9_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pma_10_cfg_c; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pma_10_cfg_atomic; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_1_io_check_env_pma_10_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pma_10_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pma_10_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pma_10_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_1_io_check_env_pma_10_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_1_io_check_env_pma_10_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pma_11_cfg_c; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pma_11_cfg_atomic; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_1_io_check_env_pma_11_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pma_11_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pma_11_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pma_11_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_1_io_check_env_pma_11_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_1_io_check_env_pma_11_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pma_12_cfg_c; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pma_12_cfg_atomic; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_1_io_check_env_pma_12_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pma_12_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pma_12_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pma_12_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_1_io_check_env_pma_12_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_1_io_check_env_pma_12_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pma_13_cfg_c; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pma_13_cfg_atomic; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_1_io_check_env_pma_13_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pma_13_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pma_13_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pma_13_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_1_io_check_env_pma_13_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_1_io_check_env_pma_13_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pma_14_cfg_c; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pma_14_cfg_atomic; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_1_io_check_env_pma_14_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pma_14_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pma_14_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pma_14_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_1_io_check_env_pma_14_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_1_io_check_env_pma_14_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pma_15_cfg_c; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pma_15_cfg_atomic; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_1_io_check_env_pma_15_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pma_15_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pma_15_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_check_env_pma_15_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_1_io_check_env_pma_15_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_1_io_check_env_pma_15_mask; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_1_io_req_bits_addr; // @[Frontend.scala 88:45]
  wire [2:0] PMPChecker_1_io_req_bits_cmd; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_resp_ld; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_resp_st; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_resp_instr; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_resp_mmio; // @[Frontend.scala 88:45]
  wire  PMPChecker_1_io_resp_atomic; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_2_io_check_env_mode; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pmp_0_cfg_l; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_2_io_check_env_pmp_0_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pmp_0_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pmp_0_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pmp_0_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_2_io_check_env_pmp_0_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_2_io_check_env_pmp_0_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pmp_1_cfg_l; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_2_io_check_env_pmp_1_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pmp_1_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pmp_1_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pmp_1_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_2_io_check_env_pmp_1_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_2_io_check_env_pmp_1_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pmp_2_cfg_l; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_2_io_check_env_pmp_2_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pmp_2_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pmp_2_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pmp_2_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_2_io_check_env_pmp_2_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_2_io_check_env_pmp_2_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pmp_3_cfg_l; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_2_io_check_env_pmp_3_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pmp_3_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pmp_3_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pmp_3_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_2_io_check_env_pmp_3_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_2_io_check_env_pmp_3_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pmp_4_cfg_l; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_2_io_check_env_pmp_4_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pmp_4_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pmp_4_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pmp_4_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_2_io_check_env_pmp_4_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_2_io_check_env_pmp_4_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pmp_5_cfg_l; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_2_io_check_env_pmp_5_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pmp_5_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pmp_5_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pmp_5_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_2_io_check_env_pmp_5_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_2_io_check_env_pmp_5_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pmp_6_cfg_l; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_2_io_check_env_pmp_6_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pmp_6_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pmp_6_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pmp_6_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_2_io_check_env_pmp_6_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_2_io_check_env_pmp_6_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pmp_7_cfg_l; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_2_io_check_env_pmp_7_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pmp_7_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pmp_7_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pmp_7_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_2_io_check_env_pmp_7_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_2_io_check_env_pmp_7_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pmp_8_cfg_l; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_2_io_check_env_pmp_8_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pmp_8_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pmp_8_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pmp_8_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_2_io_check_env_pmp_8_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_2_io_check_env_pmp_8_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pmp_9_cfg_l; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_2_io_check_env_pmp_9_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pmp_9_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pmp_9_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pmp_9_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_2_io_check_env_pmp_9_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_2_io_check_env_pmp_9_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pmp_10_cfg_l; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_2_io_check_env_pmp_10_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pmp_10_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pmp_10_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pmp_10_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_2_io_check_env_pmp_10_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_2_io_check_env_pmp_10_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pmp_11_cfg_l; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_2_io_check_env_pmp_11_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pmp_11_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pmp_11_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pmp_11_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_2_io_check_env_pmp_11_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_2_io_check_env_pmp_11_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pmp_12_cfg_l; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_2_io_check_env_pmp_12_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pmp_12_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pmp_12_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pmp_12_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_2_io_check_env_pmp_12_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_2_io_check_env_pmp_12_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pmp_13_cfg_l; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_2_io_check_env_pmp_13_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pmp_13_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pmp_13_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pmp_13_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_2_io_check_env_pmp_13_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_2_io_check_env_pmp_13_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pmp_14_cfg_l; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_2_io_check_env_pmp_14_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pmp_14_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pmp_14_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pmp_14_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_2_io_check_env_pmp_14_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_2_io_check_env_pmp_14_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pmp_15_cfg_l; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_2_io_check_env_pmp_15_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pmp_15_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pmp_15_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pmp_15_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_2_io_check_env_pmp_15_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_2_io_check_env_pmp_15_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pma_0_cfg_c; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pma_0_cfg_atomic; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_2_io_check_env_pma_0_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pma_0_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pma_0_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pma_0_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_2_io_check_env_pma_0_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_2_io_check_env_pma_0_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pma_1_cfg_c; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pma_1_cfg_atomic; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_2_io_check_env_pma_1_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pma_1_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pma_1_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pma_1_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_2_io_check_env_pma_1_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_2_io_check_env_pma_1_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pma_2_cfg_c; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pma_2_cfg_atomic; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_2_io_check_env_pma_2_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pma_2_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pma_2_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pma_2_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_2_io_check_env_pma_2_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_2_io_check_env_pma_2_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pma_3_cfg_c; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pma_3_cfg_atomic; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_2_io_check_env_pma_3_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pma_3_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pma_3_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pma_3_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_2_io_check_env_pma_3_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_2_io_check_env_pma_3_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pma_4_cfg_c; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pma_4_cfg_atomic; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_2_io_check_env_pma_4_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pma_4_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pma_4_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pma_4_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_2_io_check_env_pma_4_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_2_io_check_env_pma_4_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pma_5_cfg_c; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pma_5_cfg_atomic; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_2_io_check_env_pma_5_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pma_5_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pma_5_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pma_5_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_2_io_check_env_pma_5_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_2_io_check_env_pma_5_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pma_6_cfg_c; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pma_6_cfg_atomic; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_2_io_check_env_pma_6_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pma_6_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pma_6_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pma_6_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_2_io_check_env_pma_6_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_2_io_check_env_pma_6_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pma_7_cfg_c; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pma_7_cfg_atomic; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_2_io_check_env_pma_7_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pma_7_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pma_7_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pma_7_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_2_io_check_env_pma_7_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_2_io_check_env_pma_7_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pma_8_cfg_c; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pma_8_cfg_atomic; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_2_io_check_env_pma_8_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pma_8_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pma_8_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pma_8_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_2_io_check_env_pma_8_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_2_io_check_env_pma_8_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pma_9_cfg_c; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pma_9_cfg_atomic; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_2_io_check_env_pma_9_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pma_9_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pma_9_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pma_9_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_2_io_check_env_pma_9_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_2_io_check_env_pma_9_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pma_10_cfg_c; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pma_10_cfg_atomic; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_2_io_check_env_pma_10_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pma_10_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pma_10_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pma_10_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_2_io_check_env_pma_10_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_2_io_check_env_pma_10_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pma_11_cfg_c; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pma_11_cfg_atomic; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_2_io_check_env_pma_11_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pma_11_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pma_11_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pma_11_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_2_io_check_env_pma_11_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_2_io_check_env_pma_11_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pma_12_cfg_c; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pma_12_cfg_atomic; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_2_io_check_env_pma_12_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pma_12_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pma_12_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pma_12_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_2_io_check_env_pma_12_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_2_io_check_env_pma_12_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pma_13_cfg_c; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pma_13_cfg_atomic; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_2_io_check_env_pma_13_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pma_13_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pma_13_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pma_13_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_2_io_check_env_pma_13_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_2_io_check_env_pma_13_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pma_14_cfg_c; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pma_14_cfg_atomic; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_2_io_check_env_pma_14_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pma_14_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pma_14_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pma_14_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_2_io_check_env_pma_14_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_2_io_check_env_pma_14_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pma_15_cfg_c; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pma_15_cfg_atomic; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_2_io_check_env_pma_15_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pma_15_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pma_15_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_check_env_pma_15_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_2_io_check_env_pma_15_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_2_io_check_env_pma_15_mask; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_2_io_req_bits_addr; // @[Frontend.scala 88:45]
  wire [2:0] PMPChecker_2_io_req_bits_cmd; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_resp_ld; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_resp_st; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_resp_instr; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_resp_mmio; // @[Frontend.scala 88:45]
  wire  PMPChecker_2_io_resp_atomic; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_3_io_check_env_mode; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pmp_0_cfg_l; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_3_io_check_env_pmp_0_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pmp_0_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pmp_0_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pmp_0_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_3_io_check_env_pmp_0_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_3_io_check_env_pmp_0_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pmp_1_cfg_l; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_3_io_check_env_pmp_1_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pmp_1_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pmp_1_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pmp_1_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_3_io_check_env_pmp_1_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_3_io_check_env_pmp_1_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pmp_2_cfg_l; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_3_io_check_env_pmp_2_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pmp_2_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pmp_2_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pmp_2_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_3_io_check_env_pmp_2_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_3_io_check_env_pmp_2_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pmp_3_cfg_l; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_3_io_check_env_pmp_3_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pmp_3_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pmp_3_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pmp_3_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_3_io_check_env_pmp_3_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_3_io_check_env_pmp_3_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pmp_4_cfg_l; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_3_io_check_env_pmp_4_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pmp_4_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pmp_4_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pmp_4_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_3_io_check_env_pmp_4_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_3_io_check_env_pmp_4_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pmp_5_cfg_l; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_3_io_check_env_pmp_5_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pmp_5_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pmp_5_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pmp_5_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_3_io_check_env_pmp_5_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_3_io_check_env_pmp_5_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pmp_6_cfg_l; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_3_io_check_env_pmp_6_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pmp_6_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pmp_6_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pmp_6_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_3_io_check_env_pmp_6_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_3_io_check_env_pmp_6_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pmp_7_cfg_l; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_3_io_check_env_pmp_7_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pmp_7_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pmp_7_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pmp_7_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_3_io_check_env_pmp_7_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_3_io_check_env_pmp_7_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pmp_8_cfg_l; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_3_io_check_env_pmp_8_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pmp_8_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pmp_8_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pmp_8_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_3_io_check_env_pmp_8_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_3_io_check_env_pmp_8_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pmp_9_cfg_l; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_3_io_check_env_pmp_9_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pmp_9_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pmp_9_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pmp_9_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_3_io_check_env_pmp_9_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_3_io_check_env_pmp_9_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pmp_10_cfg_l; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_3_io_check_env_pmp_10_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pmp_10_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pmp_10_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pmp_10_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_3_io_check_env_pmp_10_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_3_io_check_env_pmp_10_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pmp_11_cfg_l; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_3_io_check_env_pmp_11_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pmp_11_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pmp_11_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pmp_11_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_3_io_check_env_pmp_11_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_3_io_check_env_pmp_11_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pmp_12_cfg_l; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_3_io_check_env_pmp_12_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pmp_12_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pmp_12_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pmp_12_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_3_io_check_env_pmp_12_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_3_io_check_env_pmp_12_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pmp_13_cfg_l; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_3_io_check_env_pmp_13_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pmp_13_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pmp_13_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pmp_13_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_3_io_check_env_pmp_13_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_3_io_check_env_pmp_13_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pmp_14_cfg_l; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_3_io_check_env_pmp_14_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pmp_14_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pmp_14_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pmp_14_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_3_io_check_env_pmp_14_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_3_io_check_env_pmp_14_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pmp_15_cfg_l; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_3_io_check_env_pmp_15_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pmp_15_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pmp_15_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pmp_15_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_3_io_check_env_pmp_15_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_3_io_check_env_pmp_15_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pma_0_cfg_c; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pma_0_cfg_atomic; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_3_io_check_env_pma_0_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pma_0_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pma_0_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pma_0_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_3_io_check_env_pma_0_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_3_io_check_env_pma_0_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pma_1_cfg_c; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pma_1_cfg_atomic; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_3_io_check_env_pma_1_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pma_1_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pma_1_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pma_1_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_3_io_check_env_pma_1_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_3_io_check_env_pma_1_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pma_2_cfg_c; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pma_2_cfg_atomic; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_3_io_check_env_pma_2_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pma_2_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pma_2_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pma_2_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_3_io_check_env_pma_2_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_3_io_check_env_pma_2_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pma_3_cfg_c; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pma_3_cfg_atomic; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_3_io_check_env_pma_3_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pma_3_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pma_3_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pma_3_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_3_io_check_env_pma_3_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_3_io_check_env_pma_3_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pma_4_cfg_c; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pma_4_cfg_atomic; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_3_io_check_env_pma_4_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pma_4_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pma_4_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pma_4_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_3_io_check_env_pma_4_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_3_io_check_env_pma_4_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pma_5_cfg_c; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pma_5_cfg_atomic; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_3_io_check_env_pma_5_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pma_5_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pma_5_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pma_5_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_3_io_check_env_pma_5_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_3_io_check_env_pma_5_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pma_6_cfg_c; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pma_6_cfg_atomic; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_3_io_check_env_pma_6_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pma_6_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pma_6_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pma_6_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_3_io_check_env_pma_6_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_3_io_check_env_pma_6_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pma_7_cfg_c; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pma_7_cfg_atomic; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_3_io_check_env_pma_7_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pma_7_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pma_7_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pma_7_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_3_io_check_env_pma_7_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_3_io_check_env_pma_7_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pma_8_cfg_c; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pma_8_cfg_atomic; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_3_io_check_env_pma_8_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pma_8_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pma_8_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pma_8_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_3_io_check_env_pma_8_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_3_io_check_env_pma_8_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pma_9_cfg_c; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pma_9_cfg_atomic; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_3_io_check_env_pma_9_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pma_9_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pma_9_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pma_9_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_3_io_check_env_pma_9_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_3_io_check_env_pma_9_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pma_10_cfg_c; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pma_10_cfg_atomic; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_3_io_check_env_pma_10_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pma_10_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pma_10_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pma_10_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_3_io_check_env_pma_10_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_3_io_check_env_pma_10_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pma_11_cfg_c; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pma_11_cfg_atomic; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_3_io_check_env_pma_11_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pma_11_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pma_11_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pma_11_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_3_io_check_env_pma_11_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_3_io_check_env_pma_11_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pma_12_cfg_c; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pma_12_cfg_atomic; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_3_io_check_env_pma_12_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pma_12_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pma_12_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pma_12_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_3_io_check_env_pma_12_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_3_io_check_env_pma_12_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pma_13_cfg_c; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pma_13_cfg_atomic; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_3_io_check_env_pma_13_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pma_13_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pma_13_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pma_13_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_3_io_check_env_pma_13_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_3_io_check_env_pma_13_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pma_14_cfg_c; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pma_14_cfg_atomic; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_3_io_check_env_pma_14_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pma_14_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pma_14_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pma_14_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_3_io_check_env_pma_14_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_3_io_check_env_pma_14_mask; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pma_15_cfg_c; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pma_15_cfg_atomic; // @[Frontend.scala 88:45]
  wire [1:0] PMPChecker_3_io_check_env_pma_15_cfg_a; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pma_15_cfg_x; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pma_15_cfg_w; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_check_env_pma_15_cfg_r; // @[Frontend.scala 88:45]
  wire [33:0] PMPChecker_3_io_check_env_pma_15_addr; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_3_io_check_env_pma_15_mask; // @[Frontend.scala 88:45]
  wire [35:0] PMPChecker_3_io_req_bits_addr; // @[Frontend.scala 88:45]
  wire [2:0] PMPChecker_3_io_req_bits_cmd; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_resp_ld; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_resp_st; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_resp_instr; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_resp_mmio; // @[Frontend.scala 88:45]
  wire  PMPChecker_3_io_resp_atomic; // @[Frontend.scala 88:45]
  wire  itlb_clock; // @[Frontend.scala 104:20]
  wire  itlb_reset; // @[Frontend.scala 104:20]
  wire  itlb_io_sfence_valid; // @[Frontend.scala 104:20]
  wire  itlb_io_sfence_bits_rs1; // @[Frontend.scala 104:20]
  wire  itlb_io_sfence_bits_rs2; // @[Frontend.scala 104:20]
  wire [38:0] itlb_io_sfence_bits_addr; // @[Frontend.scala 104:20]
  wire [15:0] itlb_io_sfence_bits_asid; // @[Frontend.scala 104:20]
  wire [3:0] itlb_io_csr_satp_mode; // @[Frontend.scala 104:20]
  wire [15:0] itlb_io_csr_satp_asid; // @[Frontend.scala 104:20]
  wire  itlb_io_csr_satp_changed; // @[Frontend.scala 104:20]
  wire [1:0] itlb_io_csr_priv_imode; // @[Frontend.scala 104:20]
  wire  itlb_io_requestor_0_req_ready; // @[Frontend.scala 104:20]
  wire  itlb_io_requestor_0_req_valid; // @[Frontend.scala 104:20]
  wire [38:0] itlb_io_requestor_0_req_bits_vaddr; // @[Frontend.scala 104:20]
  wire  itlb_io_requestor_0_req_bits_kill; // @[Frontend.scala 104:20]
  wire  itlb_io_requestor_0_resp_ready; // @[Frontend.scala 104:20]
  wire  itlb_io_requestor_0_resp_valid; // @[Frontend.scala 104:20]
  wire [35:0] itlb_io_requestor_0_resp_bits_paddr_0; // @[Frontend.scala 104:20]
  wire  itlb_io_requestor_0_resp_bits_excp_0_pf_instr; // @[Frontend.scala 104:20]
  wire  itlb_io_requestor_0_resp_bits_excp_0_af_instr; // @[Frontend.scala 104:20]
  wire  itlb_io_requestor_1_req_ready; // @[Frontend.scala 104:20]
  wire  itlb_io_requestor_1_req_valid; // @[Frontend.scala 104:20]
  wire [38:0] itlb_io_requestor_1_req_bits_vaddr; // @[Frontend.scala 104:20]
  wire  itlb_io_requestor_1_req_bits_kill; // @[Frontend.scala 104:20]
  wire  itlb_io_requestor_1_resp_ready; // @[Frontend.scala 104:20]
  wire  itlb_io_requestor_1_resp_valid; // @[Frontend.scala 104:20]
  wire [35:0] itlb_io_requestor_1_resp_bits_paddr_0; // @[Frontend.scala 104:20]
  wire  itlb_io_requestor_1_resp_bits_excp_0_pf_instr; // @[Frontend.scala 104:20]
  wire  itlb_io_requestor_1_resp_bits_excp_0_af_instr; // @[Frontend.scala 104:20]
  wire  itlb_io_requestor_3_req_ready; // @[Frontend.scala 104:20]
  wire  itlb_io_requestor_3_req_valid; // @[Frontend.scala 104:20]
  wire [38:0] itlb_io_requestor_3_req_bits_vaddr; // @[Frontend.scala 104:20]
  wire  itlb_io_requestor_3_resp_valid; // @[Frontend.scala 104:20]
  wire [35:0] itlb_io_requestor_3_resp_bits_paddr_0; // @[Frontend.scala 104:20]
  wire  itlb_io_requestor_3_resp_bits_miss; // @[Frontend.scala 104:20]
  wire  itlb_io_requestor_3_resp_bits_excp_0_pf_instr; // @[Frontend.scala 104:20]
  wire  itlb_io_requestor_3_resp_bits_excp_0_af_instr; // @[Frontend.scala 104:20]
  wire  itlb_io_flushPipe_0; // @[Frontend.scala 104:20]
  wire  itlb_io_flushPipe_1; // @[Frontend.scala 104:20]
  wire  itlb_io_flushPipe_3; // @[Frontend.scala 104:20]
  wire  itlb_io_ptw_req_0_ready; // @[Frontend.scala 104:20]
  wire  itlb_io_ptw_req_0_valid; // @[Frontend.scala 104:20]
  wire [26:0] itlb_io_ptw_req_0_bits_vpn; // @[Frontend.scala 104:20]
  wire  itlb_io_ptw_req_1_ready; // @[Frontend.scala 104:20]
  wire  itlb_io_ptw_req_1_valid; // @[Frontend.scala 104:20]
  wire [26:0] itlb_io_ptw_req_1_bits_vpn; // @[Frontend.scala 104:20]
  wire  itlb_io_ptw_req_3_ready; // @[Frontend.scala 104:20]
  wire  itlb_io_ptw_req_3_valid; // @[Frontend.scala 104:20]
  wire [26:0] itlb_io_ptw_req_3_bits_vpn; // @[Frontend.scala 104:20]
  wire  itlb_io_ptw_resp_ready; // @[Frontend.scala 104:20]
  wire  itlb_io_ptw_resp_valid; // @[Frontend.scala 104:20]
  wire [26:0] itlb_io_ptw_resp_bits_entry_tag; // @[Frontend.scala 104:20]
  wire [15:0] itlb_io_ptw_resp_bits_entry_asid; // @[Frontend.scala 104:20]
  wire [23:0] itlb_io_ptw_resp_bits_entry_ppn; // @[Frontend.scala 104:20]
  wire  itlb_io_ptw_resp_bits_entry_perm_d; // @[Frontend.scala 104:20]
  wire  itlb_io_ptw_resp_bits_entry_perm_a; // @[Frontend.scala 104:20]
  wire  itlb_io_ptw_resp_bits_entry_perm_g; // @[Frontend.scala 104:20]
  wire  itlb_io_ptw_resp_bits_entry_perm_u; // @[Frontend.scala 104:20]
  wire  itlb_io_ptw_resp_bits_entry_perm_x; // @[Frontend.scala 104:20]
  wire  itlb_io_ptw_resp_bits_entry_perm_w; // @[Frontend.scala 104:20]
  wire  itlb_io_ptw_resp_bits_entry_perm_r; // @[Frontend.scala 104:20]
  wire [1:0] itlb_io_ptw_resp_bits_entry_level; // @[Frontend.scala 104:20]
  wire  itlb_io_ptw_resp_bits_pf; // @[Frontend.scala 104:20]
  wire  itlb_io_ptw_resp_bits_af; // @[Frontend.scala 104:20]
  wire  pfevent_clock; // @[Frontend.scala 165:23]
  wire  pfevent_reset; // @[Frontend.scala 165:23]
  wire  pfevent_io_distribute_csr_wvalid; // @[Frontend.scala 165:23]
  wire [11:0] pfevent_io_distribute_csr_waddr; // @[Frontend.scala 165:23]
  wire [63:0] pfevent_io_distribute_csr_wdata; // @[Frontend.scala 165:23]
  wire [63:0] pfevent_io_hpmevent_0; // @[Frontend.scala 165:23]
  wire [63:0] pfevent_io_hpmevent_1; // @[Frontend.scala 165:23]
  wire [63:0] pfevent_io_hpmevent_2; // @[Frontend.scala 165:23]
  wire [63:0] pfevent_io_hpmevent_3; // @[Frontend.scala 165:23]
  wire [63:0] pfevent_io_hpmevent_4; // @[Frontend.scala 165:23]
  wire [63:0] pfevent_io_hpmevent_5; // @[Frontend.scala 165:23]
  wire [63:0] pfevent_io_hpmevent_6; // @[Frontend.scala 165:23]
  wire [63:0] pfevent_io_hpmevent_7; // @[Frontend.scala 165:23]
  wire [63:0] pfevent_io_hpmevent_8; // @[Frontend.scala 165:23]
  wire [63:0] pfevent_io_hpmevent_9; // @[Frontend.scala 165:23]
  wire [63:0] pfevent_io_hpmevent_10; // @[Frontend.scala 165:23]
  wire [63:0] pfevent_io_hpmevent_11; // @[Frontend.scala 165:23]
  wire [63:0] pfevent_io_hpmevent_12; // @[Frontend.scala 165:23]
  wire [63:0] pfevent_io_hpmevent_13; // @[Frontend.scala 165:23]
  wire [63:0] pfevent_io_hpmevent_14; // @[Frontend.scala 165:23]
  wire [63:0] pfevent_io_hpmevent_15; // @[Frontend.scala 165:23]
  wire [63:0] pfevent_io_hpmevent_16; // @[Frontend.scala 165:23]
  wire [63:0] pfevent_io_hpmevent_17; // @[Frontend.scala 165:23]
  wire [63:0] pfevent_io_hpmevent_18; // @[Frontend.scala 165:23]
  wire [63:0] pfevent_io_hpmevent_19; // @[Frontend.scala 165:23]
  wire [63:0] pfevent_io_hpmevent_20; // @[Frontend.scala 165:23]
  wire [63:0] pfevent_io_hpmevent_21; // @[Frontend.scala 165:23]
  wire [63:0] pfevent_io_hpmevent_22; // @[Frontend.scala 165:23]
  wire [63:0] pfevent_io_hpmevent_23; // @[Frontend.scala 165:23]
  wire  hpm_clock; // @[PerfCounterUtils.scala 255:21]
  wire [63:0] hpm_io_hpm_event_0; // @[PerfCounterUtils.scala 255:21]
  wire [63:0] hpm_io_hpm_event_1; // @[PerfCounterUtils.scala 255:21]
  wire [63:0] hpm_io_hpm_event_2; // @[PerfCounterUtils.scala 255:21]
  wire [63:0] hpm_io_hpm_event_3; // @[PerfCounterUtils.scala 255:21]
  wire [63:0] hpm_io_hpm_event_4; // @[PerfCounterUtils.scala 255:21]
  wire [63:0] hpm_io_hpm_event_5; // @[PerfCounterUtils.scala 255:21]
  wire [63:0] hpm_io_hpm_event_6; // @[PerfCounterUtils.scala 255:21]
  wire [63:0] hpm_io_hpm_event_7; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_0_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_1_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_2_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_3_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_4_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_5_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_6_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_7_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_8_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_9_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_10_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_11_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_12_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_13_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_14_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_15_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_16_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_17_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_18_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_19_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_20_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_23_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_24_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_25_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_26_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_27_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_28_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_29_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_30_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_31_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_32_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_33_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_34_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_35_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_36_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_37_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_38_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_39_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_40_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_41_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_42_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_43_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_44_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_45_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_46_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_47_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_48_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_49_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_50_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_51_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_52_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_53_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_perf_0_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_perf_1_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_perf_2_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_perf_3_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_perf_4_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_perf_5_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_perf_6_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_perf_7_value; // @[PerfCounterUtils.scala 255:21]
  reg  needFlush; // @[Frontend.scala 71:26]
  reg  io_csrUpdate_REG_wvalid; // @[Frontend.scala 136:26]
  reg [11:0] io_csrUpdate_REG_waddr; // @[Frontend.scala 136:26]
  reg [63:0] io_csrUpdate_REG_wdata; // @[Frontend.scala 136:26]
  reg  icache_io_csr_parity_enable_REG; // @[Frontend.scala 139:41]
  reg [35:0] io_error_REG_paddr; // @[Frontend.scala 156:30]
  reg  io_error_REG_report_to_beu; // @[Frontend.scala 156:30]
  reg [35:0] io_error_REG_1_paddr; // @[Frontend.scala 156:22]
  reg  io_error_REG_1_report_to_beu; // @[Frontend.scala 156:22]
  reg [5:0] io_perf_0_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg [5:0] io_perf_0_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  reg [5:0] io_perf_1_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg [5:0] io_perf_1_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  reg [5:0] io_perf_2_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg [5:0] io_perf_2_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  reg [5:0] io_perf_3_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg [5:0] io_perf_3_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  reg [5:0] io_perf_4_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg [5:0] io_perf_4_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  reg [5:0] io_perf_5_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg [5:0] io_perf_5_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  reg [5:0] io_perf_6_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg [5:0] io_perf_6_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  reg [5:0] io_perf_7_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg [5:0] io_perf_7_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  InstrUncache instrUncache ( // @[Frontend.scala 32:33]
    .clock(instrUncache_clock),
    .reset(instrUncache_reset),
    .auto_client_out_a_ready(instrUncache_auto_client_out_a_ready),
    .auto_client_out_a_valid(instrUncache_auto_client_out_a_valid),
    .auto_client_out_a_bits_address(instrUncache_auto_client_out_a_bits_address),
    .auto_client_out_d_ready(instrUncache_auto_client_out_d_ready),
    .auto_client_out_d_valid(instrUncache_auto_client_out_d_valid),
    .auto_client_out_d_bits_source(instrUncache_auto_client_out_d_bits_source),
    .auto_client_out_d_bits_data(instrUncache_auto_client_out_d_bits_data),
    .io_req_ready(instrUncache_io_req_ready),
    .io_req_valid(instrUncache_io_req_valid),
    .io_req_bits_addr(instrUncache_io_req_bits_addr),
    .io_resp_valid(instrUncache_io_resp_valid),
    .io_resp_bits_data(instrUncache_io_resp_bits_data)
  );
  ICache icache ( // @[Frontend.scala 33:33]
    .clock(icache_clock),
    .reset(icache_reset),
    .auto_client_out_a_ready(icache_auto_client_out_a_ready),
    .auto_client_out_a_valid(icache_auto_client_out_a_valid),
    .auto_client_out_a_bits_opcode(icache_auto_client_out_a_bits_opcode),
    .auto_client_out_a_bits_size(icache_auto_client_out_a_bits_size),
    .auto_client_out_a_bits_source(icache_auto_client_out_a_bits_source),
    .auto_client_out_a_bits_address(icache_auto_client_out_a_bits_address),
    .auto_client_out_a_bits_mask(icache_auto_client_out_a_bits_mask),
    .auto_client_out_bready(icache_auto_client_out_bready),
    .auto_client_out_bvalid(icache_auto_client_out_bvalid),
    .auto_client_out_bparam(icache_auto_client_out_bparam),
    .auto_client_out_baddress(icache_auto_client_out_baddress),
    .auto_client_out_bdata(icache_auto_client_out_bdata),
    .auto_client_out_c_ready(icache_auto_client_out_c_ready),
    .auto_client_out_c_valid(icache_auto_client_out_c_valid),
    .auto_client_out_c_bits_opcode(icache_auto_client_out_c_bits_opcode),
    .auto_client_out_c_bits_param(icache_auto_client_out_c_bits_param),
    .auto_client_out_c_bits_address(icache_auto_client_out_c_bits_address),
    .auto_client_out_c_bits_echo_blockisdirty(icache_auto_client_out_c_bits_echo_blockisdirty),
    .auto_client_out_c_bits_data(icache_auto_client_out_c_bits_data),
    .auto_client_out_d_ready(icache_auto_client_out_d_ready),
    .auto_client_out_d_valid(icache_auto_client_out_d_valid),
    .auto_client_out_d_bits_opcode(icache_auto_client_out_d_bits_opcode),
    .auto_client_out_d_bits_param(icache_auto_client_out_d_bits_param),
    .auto_client_out_d_bits_source(icache_auto_client_out_d_bits_source),
    .auto_client_out_d_bits_sink(icache_auto_client_out_d_bits_sink),
    .auto_client_out_d_bits_echo_blockisdirty(icache_auto_client_out_d_bits_echo_blockisdirty),
    .auto_client_out_d_bits_data(icache_auto_client_out_d_bits_data),
    .auto_client_out_d_bits_corrupt(icache_auto_client_out_d_bits_corrupt),
    .auto_client_out_e_ready(icache_auto_client_out_e_ready),
    .auto_client_out_e_valid(icache_auto_client_out_e_valid),
    .auto_client_out_e_bits_sink(icache_auto_client_out_e_bits_sink),
    .io_stop(icache_io_stop),
    .io_fetch_req_ready(icache_io_fetch_req_ready),
    .io_fetch_req_valid(icache_io_fetch_req_valid),
    .io_fetch_req_bits_pcMemRead_0_startAddr(icache_io_fetch_req_bits_pcMemRead_0_startAddr),
    .io_fetch_req_bits_pcMemRead_0_nextlineStart(icache_io_fetch_req_bits_pcMemRead_0_nextlineStart),
    .io_fetch_req_bits_pcMemRead_1_startAddr(icache_io_fetch_req_bits_pcMemRead_1_startAddr),
    .io_fetch_req_bits_pcMemRead_1_nextlineStart(icache_io_fetch_req_bits_pcMemRead_1_nextlineStart),
    .io_fetch_req_bits_pcMemRead_2_startAddr(icache_io_fetch_req_bits_pcMemRead_2_startAddr),
    .io_fetch_req_bits_pcMemRead_2_nextlineStart(icache_io_fetch_req_bits_pcMemRead_2_nextlineStart),
    .io_fetch_req_bits_pcMemRead_3_startAddr(icache_io_fetch_req_bits_pcMemRead_3_startAddr),
    .io_fetch_req_bits_pcMemRead_3_nextlineStart(icache_io_fetch_req_bits_pcMemRead_3_nextlineStart),
    .io_fetch_req_bits_pcMemRead_4_startAddr(icache_io_fetch_req_bits_pcMemRead_4_startAddr),
    .io_fetch_req_bits_pcMemRead_4_nextlineStart(icache_io_fetch_req_bits_pcMemRead_4_nextlineStart),
    .io_fetch_req_bits_readValid_0(icache_io_fetch_req_bits_readValid_0),
    .io_fetch_req_bits_readValid_1(icache_io_fetch_req_bits_readValid_1),
    .io_fetch_req_bits_readValid_2(icache_io_fetch_req_bits_readValid_2),
    .io_fetch_req_bits_readValid_3(icache_io_fetch_req_bits_readValid_3),
    .io_fetch_req_bits_readValid_4(icache_io_fetch_req_bits_readValid_4),
    .io_fetch_resp_0_valid(icache_io_fetch_resp_0_valid),
    .io_fetch_resp_0_bits_vaddr(icache_io_fetch_resp_0_bits_vaddr),
    .io_fetch_resp_0_bits_registerData(icache_io_fetch_resp_0_bits_registerData),
    .io_fetch_resp_0_bits_sramData(icache_io_fetch_resp_0_bits_sramData),
    .io_fetch_resp_0_bits_select(icache_io_fetch_resp_0_bits_select),
    .io_fetch_resp_0_bits_paddr(icache_io_fetch_resp_0_bits_paddr),
    .io_fetch_resp_0_bits_tlbExcp_pageFault(icache_io_fetch_resp_0_bits_tlbExcp_pageFault),
    .io_fetch_resp_0_bits_tlbExcp_accessFault(icache_io_fetch_resp_0_bits_tlbExcp_accessFault),
    .io_fetch_resp_0_bits_tlbExcp_mmio(icache_io_fetch_resp_0_bits_tlbExcp_mmio),
    .io_fetch_resp_1_valid(icache_io_fetch_resp_1_valid),
    .io_fetch_resp_1_bits_vaddr(icache_io_fetch_resp_1_bits_vaddr),
    .io_fetch_resp_1_bits_registerData(icache_io_fetch_resp_1_bits_registerData),
    .io_fetch_resp_1_bits_sramData(icache_io_fetch_resp_1_bits_sramData),
    .io_fetch_resp_1_bits_select(icache_io_fetch_resp_1_bits_select),
    .io_fetch_resp_1_bits_tlbExcp_pageFault(icache_io_fetch_resp_1_bits_tlbExcp_pageFault),
    .io_fetch_resp_1_bits_tlbExcp_accessFault(icache_io_fetch_resp_1_bits_tlbExcp_accessFault),
    .io_toIFU(icache_io_toIFU),
    .io_pmp_0_req_bits_addr(icache_io_pmp_0_req_bits_addr),
    .io_pmp_0_resp_instr(icache_io_pmp_0_resp_instr),
    .io_pmp_0_resp_mmio(icache_io_pmp_0_resp_mmio),
    .io_pmp_1_req_bits_addr(icache_io_pmp_1_req_bits_addr),
    .io_pmp_1_resp_instr(icache_io_pmp_1_resp_instr),
    .io_itlb_0_req_ready(icache_io_itlb_0_req_ready),
    .io_itlb_0_req_valid(icache_io_itlb_0_req_valid),
    .io_itlb_0_req_bits_vaddr(icache_io_itlb_0_req_bits_vaddr),
    .io_itlb_0_req_bits_kill(icache_io_itlb_0_req_bits_kill),
    .io_itlb_0_resp_ready(icache_io_itlb_0_resp_ready),
    .io_itlb_0_resp_valid(icache_io_itlb_0_resp_valid),
    .io_itlb_0_resp_bits_paddr_0(icache_io_itlb_0_resp_bits_paddr_0),
    .io_itlb_0_resp_bits_excp_0_pf_instr(icache_io_itlb_0_resp_bits_excp_0_pf_instr),
    .io_itlb_0_resp_bits_excp_0_af_instr(icache_io_itlb_0_resp_bits_excp_0_af_instr),
    .io_itlb_1_req_ready(icache_io_itlb_1_req_ready),
    .io_itlb_1_req_valid(icache_io_itlb_1_req_valid),
    .io_itlb_1_req_bits_vaddr(icache_io_itlb_1_req_bits_vaddr),
    .io_itlb_1_req_bits_kill(icache_io_itlb_1_req_bits_kill),
    .io_itlb_1_resp_ready(icache_io_itlb_1_resp_ready),
    .io_itlb_1_resp_valid(icache_io_itlb_1_resp_valid),
    .io_itlb_1_resp_bits_paddr_0(icache_io_itlb_1_resp_bits_paddr_0),
    .io_itlb_1_resp_bits_excp_0_pf_instr(icache_io_itlb_1_resp_bits_excp_0_pf_instr),
    .io_itlb_1_resp_bits_excp_0_af_instr(icache_io_itlb_1_resp_bits_excp_0_af_instr),
    .io_perfInfo_only_0_hit(icache_io_perfInfo_only_0_hit),
    .io_perfInfo_only_0_miss(icache_io_perfInfo_only_0_miss),
    .io_perfInfo_hit_0_hit_1(icache_io_perfInfo_hit_0_hit_1),
    .io_perfInfo_hit_0_miss_1(icache_io_perfInfo_hit_0_miss_1),
    .io_perfInfo_miss_0_hit_1(icache_io_perfInfo_miss_0_hit_1),
    .io_perfInfo_miss_0_miss_1(icache_io_perfInfo_miss_0_miss_1),
    .io_perfInfo_hit_0_except_1(icache_io_perfInfo_hit_0_except_1),
    .io_perfInfo_miss_0_except_1(icache_io_perfInfo_miss_0_except_1),
    .io_perfInfo_except_0(icache_io_perfInfo_except_0),
    .io_perfInfo_bank_hit_1(icache_io_perfInfo_bank_hit_1),
    .io_perfInfo_hit(icache_io_perfInfo_hit),
    .io_error_source_tag(icache_io_error_source_tag),
    .io_error_source_data(icache_io_error_source_data),
    .io_error_source_l2(icache_io_error_source_l2),
    .io_error_opType_fetch(icache_io_error_opType_fetch),
    .io_error_opType_load(icache_io_error_opType_load),
    .io_error_opType_store(icache_io_error_opType_store),
    .io_error_opType_probe(icache_io_error_opType_probe),
    .io_error_opType_release(icache_io_error_opType_release),
    .io_error_opType_atom(icache_io_error_opType_atom),
    .io_error_paddr(icache_io_error_paddr),
    .io_error_report_to_beu(icache_io_error_report_to_beu),
    .io_error_valid(icache_io_error_valid),
    .io_csr_distribute_csr_wvalid(icache_io_csr_distribute_csr_wvalid),
    .io_csr_distribute_csr_waddr(icache_io_csr_distribute_csr_waddr),
    .io_csr_distribute_csr_wdata(icache_io_csr_distribute_csr_wdata),
    .io_csr_update_wvalid(icache_io_csr_update_wvalid),
    .io_csr_update_waddr(icache_io_csr_update_waddr),
    .io_csr_update_wdata(icache_io_csr_update_wdata),
    .io_csr_parity_enable(icache_io_csr_parity_enable)
  );
  Predictor bpu ( // @[Frontend.scala 66:23]
    .clock(bpu_clock),
    .reset(bpu_reset),
    .io_bpu_to_ftq_resp_ready(bpu_io_bpu_to_ftq_resp_ready),
    .io_bpu_to_ftq_resp_valid(bpu_io_bpu_to_ftq_resp_valid),
    .io_bpu_to_ftq_resp_bits_s1_pc(bpu_io_bpu_to_ftq_resp_bits_s1_pc),
    .io_bpu_to_ftq_resp_bits_s1_full_pred_br_taken_mask_0(bpu_io_bpu_to_ftq_resp_bits_s1_full_pred_br_taken_mask_0),
    .io_bpu_to_ftq_resp_bits_s1_full_pred_br_taken_mask_1(bpu_io_bpu_to_ftq_resp_bits_s1_full_pred_br_taken_mask_1),
    .io_bpu_to_ftq_resp_bits_s1_full_pred_slot_valids_0(bpu_io_bpu_to_ftq_resp_bits_s1_full_pred_slot_valids_0),
    .io_bpu_to_ftq_resp_bits_s1_full_pred_slot_valids_1(bpu_io_bpu_to_ftq_resp_bits_s1_full_pred_slot_valids_1),
    .io_bpu_to_ftq_resp_bits_s1_full_pred_targets_0(bpu_io_bpu_to_ftq_resp_bits_s1_full_pred_targets_0),
    .io_bpu_to_ftq_resp_bits_s1_full_pred_targets_1(bpu_io_bpu_to_ftq_resp_bits_s1_full_pred_targets_1),
    .io_bpu_to_ftq_resp_bits_s1_full_pred_offsets_0(bpu_io_bpu_to_ftq_resp_bits_s1_full_pred_offsets_0),
    .io_bpu_to_ftq_resp_bits_s1_full_pred_offsets_1(bpu_io_bpu_to_ftq_resp_bits_s1_full_pred_offsets_1),
    .io_bpu_to_ftq_resp_bits_s1_full_pred_fallThroughAddr(bpu_io_bpu_to_ftq_resp_bits_s1_full_pred_fallThroughAddr),
    .io_bpu_to_ftq_resp_bits_s1_full_pred_fallThroughErr(bpu_io_bpu_to_ftq_resp_bits_s1_full_pred_fallThroughErr),
    .io_bpu_to_ftq_resp_bits_s1_full_pred_is_br_sharing(bpu_io_bpu_to_ftq_resp_bits_s1_full_pred_is_br_sharing),
    .io_bpu_to_ftq_resp_bits_s1_full_pred_hit(bpu_io_bpu_to_ftq_resp_bits_s1_full_pred_hit),
    .io_bpu_to_ftq_resp_bits_s2_pc(bpu_io_bpu_to_ftq_resp_bits_s2_pc),
    .io_bpu_to_ftq_resp_bits_s2_valid(bpu_io_bpu_to_ftq_resp_bits_s2_valid),
    .io_bpu_to_ftq_resp_bits_s2_hasRedirect(bpu_io_bpu_to_ftq_resp_bits_s2_hasRedirect),
    .io_bpu_to_ftq_resp_bits_s2_ftq_idx_flag(bpu_io_bpu_to_ftq_resp_bits_s2_ftq_idx_flag),
    .io_bpu_to_ftq_resp_bits_s2_ftq_idx_value(bpu_io_bpu_to_ftq_resp_bits_s2_ftq_idx_value),
    .io_bpu_to_ftq_resp_bits_s2_full_pred_br_taken_mask_0(bpu_io_bpu_to_ftq_resp_bits_s2_full_pred_br_taken_mask_0),
    .io_bpu_to_ftq_resp_bits_s2_full_pred_br_taken_mask_1(bpu_io_bpu_to_ftq_resp_bits_s2_full_pred_br_taken_mask_1),
    .io_bpu_to_ftq_resp_bits_s2_full_pred_slot_valids_0(bpu_io_bpu_to_ftq_resp_bits_s2_full_pred_slot_valids_0),
    .io_bpu_to_ftq_resp_bits_s2_full_pred_slot_valids_1(bpu_io_bpu_to_ftq_resp_bits_s2_full_pred_slot_valids_1),
    .io_bpu_to_ftq_resp_bits_s2_full_pred_targets_0(bpu_io_bpu_to_ftq_resp_bits_s2_full_pred_targets_0),
    .io_bpu_to_ftq_resp_bits_s2_full_pred_targets_1(bpu_io_bpu_to_ftq_resp_bits_s2_full_pred_targets_1),
    .io_bpu_to_ftq_resp_bits_s2_full_pred_offsets_0(bpu_io_bpu_to_ftq_resp_bits_s2_full_pred_offsets_0),
    .io_bpu_to_ftq_resp_bits_s2_full_pred_offsets_1(bpu_io_bpu_to_ftq_resp_bits_s2_full_pred_offsets_1),
    .io_bpu_to_ftq_resp_bits_s2_full_pred_fallThroughAddr(bpu_io_bpu_to_ftq_resp_bits_s2_full_pred_fallThroughAddr),
    .io_bpu_to_ftq_resp_bits_s2_full_pred_fallThroughErr(bpu_io_bpu_to_ftq_resp_bits_s2_full_pred_fallThroughErr),
    .io_bpu_to_ftq_resp_bits_s2_full_pred_is_br_sharing(bpu_io_bpu_to_ftq_resp_bits_s2_full_pred_is_br_sharing),
    .io_bpu_to_ftq_resp_bits_s2_full_pred_hit(bpu_io_bpu_to_ftq_resp_bits_s2_full_pred_hit),
    .io_bpu_to_ftq_resp_bits_s3_pc(bpu_io_bpu_to_ftq_resp_bits_s3_pc),
    .io_bpu_to_ftq_resp_bits_s3_valid(bpu_io_bpu_to_ftq_resp_bits_s3_valid),
    .io_bpu_to_ftq_resp_bits_s3_hasRedirect(bpu_io_bpu_to_ftq_resp_bits_s3_hasRedirect),
    .io_bpu_to_ftq_resp_bits_s3_ftq_idx_flag(bpu_io_bpu_to_ftq_resp_bits_s3_ftq_idx_flag),
    .io_bpu_to_ftq_resp_bits_s3_ftq_idx_value(bpu_io_bpu_to_ftq_resp_bits_s3_ftq_idx_value),
    .io_bpu_to_ftq_resp_bits_s3_full_pred_br_taken_mask_0(bpu_io_bpu_to_ftq_resp_bits_s3_full_pred_br_taken_mask_0),
    .io_bpu_to_ftq_resp_bits_s3_full_pred_br_taken_mask_1(bpu_io_bpu_to_ftq_resp_bits_s3_full_pred_br_taken_mask_1),
    .io_bpu_to_ftq_resp_bits_s3_full_pred_slot_valids_0(bpu_io_bpu_to_ftq_resp_bits_s3_full_pred_slot_valids_0),
    .io_bpu_to_ftq_resp_bits_s3_full_pred_slot_valids_1(bpu_io_bpu_to_ftq_resp_bits_s3_full_pred_slot_valids_1),
    .io_bpu_to_ftq_resp_bits_s3_full_pred_targets_0(bpu_io_bpu_to_ftq_resp_bits_s3_full_pred_targets_0),
    .io_bpu_to_ftq_resp_bits_s3_full_pred_targets_1(bpu_io_bpu_to_ftq_resp_bits_s3_full_pred_targets_1),
    .io_bpu_to_ftq_resp_bits_s3_full_pred_offsets_0(bpu_io_bpu_to_ftq_resp_bits_s3_full_pred_offsets_0),
    .io_bpu_to_ftq_resp_bits_s3_full_pred_offsets_1(bpu_io_bpu_to_ftq_resp_bits_s3_full_pred_offsets_1),
    .io_bpu_to_ftq_resp_bits_s3_full_pred_fallThroughAddr(bpu_io_bpu_to_ftq_resp_bits_s3_full_pred_fallThroughAddr),
    .io_bpu_to_ftq_resp_bits_s3_full_pred_fallThroughErr(bpu_io_bpu_to_ftq_resp_bits_s3_full_pred_fallThroughErr),
    .io_bpu_to_ftq_resp_bits_s3_full_pred_is_br_sharing(bpu_io_bpu_to_ftq_resp_bits_s3_full_pred_is_br_sharing),
    .io_bpu_to_ftq_resp_bits_s3_full_pred_hit(bpu_io_bpu_to_ftq_resp_bits_s3_full_pred_hit),
    .io_bpu_to_ftq_resp_bits_last_stage_meta(bpu_io_bpu_to_ftq_resp_bits_last_stage_meta),
    .io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_17_folded_hist(
      bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_17_folded_hist),
    .io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_16_folded_hist(
      bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_16_folded_hist),
    .io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_15_folded_hist(
      bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_15_folded_hist),
    .io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_14_folded_hist(
      bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_14_folded_hist),
    .io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_13_folded_hist(
      bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_13_folded_hist),
    .io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_12_folded_hist(
      bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_12_folded_hist),
    .io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_11_folded_hist(
      bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_11_folded_hist),
    .io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_10_folded_hist(
      bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_10_folded_hist),
    .io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_9_folded_hist(
      bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_9_folded_hist),
    .io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_8_folded_hist(
      bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_8_folded_hist),
    .io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_7_folded_hist(
      bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_7_folded_hist),
    .io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_6_folded_hist(
      bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_6_folded_hist),
    .io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_5_folded_hist(
      bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_5_folded_hist),
    .io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_4_folded_hist(
      bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_4_folded_hist),
    .io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_3_folded_hist(
      bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_3_folded_hist),
    .io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_2_folded_hist(
      bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_2_folded_hist),
    .io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_1_folded_hist(
      bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_1_folded_hist),
    .io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_0_folded_hist(
      bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_0_folded_hist),
    .io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_5_bits_0(
      bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_5_bits_0),
    .io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_5_bits_1(
      bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_5_bits_1),
    .io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_5_bits_2(
      bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_5_bits_2),
    .io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_5_bits_3(
      bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_5_bits_3),
    .io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_4_bits_0(
      bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_4_bits_0),
    .io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_4_bits_1(
      bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_4_bits_1),
    .io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_4_bits_2(
      bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_4_bits_2),
    .io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_4_bits_3(
      bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_4_bits_3),
    .io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_3_bits_0(
      bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_3_bits_0),
    .io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_3_bits_1(
      bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_3_bits_1),
    .io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_3_bits_2(
      bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_3_bits_2),
    .io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_3_bits_3(
      bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_3_bits_3),
    .io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_2_bits_0(
      bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_2_bits_0),
    .io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_2_bits_1(
      bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_2_bits_1),
    .io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_2_bits_2(
      bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_2_bits_2),
    .io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_2_bits_3(
      bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_2_bits_3),
    .io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_1_bits_0(
      bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_1_bits_0),
    .io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_1_bits_1(
      bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_1_bits_1),
    .io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_1_bits_2(
      bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_1_bits_2),
    .io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_1_bits_3(
      bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_1_bits_3),
    .io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_0_bits_0(
      bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_0_bits_0),
    .io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_0_bits_1(
      bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_0_bits_1),
    .io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_0_bits_2(
      bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_0_bits_2),
    .io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_0_bits_3(
      bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_0_bits_3),
    .io_bpu_to_ftq_resp_bits_last_stage_spec_info_lastBrNumOH(
      bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_lastBrNumOH),
    .io_bpu_to_ftq_resp_bits_last_stage_spec_info_histPtr_flag(
      bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_histPtr_flag),
    .io_bpu_to_ftq_resp_bits_last_stage_spec_info_histPtr_value(
      bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_histPtr_value),
    .io_bpu_to_ftq_resp_bits_last_stage_spec_info_rasSp(bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_rasSp),
    .io_bpu_to_ftq_resp_bits_last_stage_spec_info_rasTop_retAddr(
      bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_rasTop_retAddr),
    .io_bpu_to_ftq_resp_bits_last_stage_spec_info_rasTop_ctr(bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_rasTop_ctr
      ),
    .io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_valid(bpu_io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_valid),
    .io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_brSlots_0_offset(
      bpu_io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_brSlots_0_offset),
    .io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_brSlots_0_lower(
      bpu_io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_brSlots_0_lower),
    .io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_brSlots_0_tarStat(
      bpu_io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_brSlots_0_tarStat),
    .io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_brSlots_0_sharing(
      bpu_io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_brSlots_0_sharing),
    .io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_brSlots_0_valid(
      bpu_io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_brSlots_0_valid),
    .io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_tailSlot_offset(
      bpu_io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_tailSlot_offset),
    .io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_tailSlot_lower(
      bpu_io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_tailSlot_lower),
    .io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_tailSlot_tarStat(
      bpu_io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_tailSlot_tarStat),
    .io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_tailSlot_sharing(
      bpu_io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_tailSlot_sharing),
    .io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_tailSlot_valid(
      bpu_io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_tailSlot_valid),
    .io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_pftAddr(bpu_io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_pftAddr),
    .io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_carry(bpu_io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_carry),
    .io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_isCall(bpu_io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_isCall),
    .io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_isRet(bpu_io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_isRet),
    .io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_isJalr(bpu_io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_isJalr),
    .io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_last_may_be_rvi_call(
      bpu_io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_last_may_be_rvi_call),
    .io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_always_taken_0(
      bpu_io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_always_taken_0),
    .io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_always_taken_1(
      bpu_io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_always_taken_1),
    .io_ftq_to_bpu_redirect_valid(bpu_io_ftq_to_bpu_redirect_valid),
    .io_ftq_to_bpu_redirect_bits_level(bpu_io_ftq_to_bpu_redirect_bits_level),
    .io_ftq_to_bpu_redirect_bits_cfiUpdate_pc(bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_pc),
    .io_ftq_to_bpu_redirect_bits_cfiUpdate_pd_isRVC(bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_pd_isRVC),
    .io_ftq_to_bpu_redirect_bits_cfiUpdate_pd_isCall(bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_pd_isCall),
    .io_ftq_to_bpu_redirect_bits_cfiUpdate_pd_isRet(bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_pd_isRet),
    .io_ftq_to_bpu_redirect_bits_cfiUpdate_rasSp(bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_rasSp),
    .io_ftq_to_bpu_redirect_bits_cfiUpdate_rasEntry_retAddr(bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_rasEntry_retAddr),
    .io_ftq_to_bpu_redirect_bits_cfiUpdate_rasEntry_ctr(bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_rasEntry_ctr),
    .io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_17_folded_hist(
      bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_17_folded_hist),
    .io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_16_folded_hist(
      bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_16_folded_hist),
    .io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_15_folded_hist(
      bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_15_folded_hist),
    .io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_14_folded_hist(
      bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_14_folded_hist),
    .io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_13_folded_hist(
      bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_13_folded_hist),
    .io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_12_folded_hist(
      bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_12_folded_hist),
    .io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_11_folded_hist(
      bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_11_folded_hist),
    .io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_10_folded_hist(
      bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_10_folded_hist),
    .io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_9_folded_hist(
      bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_9_folded_hist),
    .io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_8_folded_hist(
      bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_8_folded_hist),
    .io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_7_folded_hist(
      bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_7_folded_hist),
    .io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_6_folded_hist(
      bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_6_folded_hist),
    .io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_5_folded_hist(
      bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_5_folded_hist),
    .io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_4_folded_hist(
      bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_4_folded_hist),
    .io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_3_folded_hist(
      bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_3_folded_hist),
    .io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_2_folded_hist(
      bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_2_folded_hist),
    .io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_1_folded_hist(
      bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_1_folded_hist),
    .io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_0_folded_hist(
      bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_0_folded_hist),
    .io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_5_bits_0(
      bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_5_bits_0),
    .io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_5_bits_1(
      bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_5_bits_1),
    .io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_5_bits_2(
      bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_5_bits_2),
    .io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_5_bits_3(
      bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_5_bits_3),
    .io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_4_bits_0(
      bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_4_bits_0),
    .io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_4_bits_1(
      bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_4_bits_1),
    .io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_4_bits_2(
      bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_4_bits_2),
    .io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_3_bits_0(
      bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_3_bits_0),
    .io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_3_bits_1(
      bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_3_bits_1),
    .io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_3_bits_2(
      bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_3_bits_2),
    .io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_3_bits_3(
      bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_3_bits_3),
    .io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_2_bits_0(
      bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_2_bits_0),
    .io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_2_bits_1(
      bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_2_bits_1),
    .io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_2_bits_2(
      bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_2_bits_2),
    .io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_2_bits_3(
      bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_2_bits_3),
    .io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_1_bits_0(
      bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_1_bits_0),
    .io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_1_bits_1(
      bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_1_bits_1),
    .io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_1_bits_2(
      bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_1_bits_2),
    .io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_1_bits_3(
      bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_1_bits_3),
    .io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_0_bits_0(
      bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_0_bits_0),
    .io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_0_bits_1(
      bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_0_bits_1),
    .io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_0_bits_2(
      bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_0_bits_2),
    .io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_0_bits_3(
      bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_0_bits_3),
    .io_ftq_to_bpu_redirect_bits_cfiUpdate_lastBrNumOH(bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_lastBrNumOH),
    .io_ftq_to_bpu_redirect_bits_cfiUpdate_histPtr_flag(bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_histPtr_flag),
    .io_ftq_to_bpu_redirect_bits_cfiUpdate_histPtr_value(bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_histPtr_value),
    .io_ftq_to_bpu_redirect_bits_cfiUpdate_target(bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_target),
    .io_ftq_to_bpu_redirect_bits_cfiUpdate_taken(bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_taken),
    .io_ftq_to_bpu_redirect_bits_cfiUpdate_shift(bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_shift),
    .io_ftq_to_bpu_redirect_bits_cfiUpdate_addIntoHist(bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_addIntoHist),
    .io_ftq_to_bpu_update_valid(bpu_io_ftq_to_bpu_update_valid),
    .io_ftq_to_bpu_update_bits_pc(bpu_io_ftq_to_bpu_update_bits_pc),
    .io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_17_folded_hist(
      bpu_io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_17_folded_hist),
    .io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_16_folded_hist(
      bpu_io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_16_folded_hist),
    .io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_15_folded_hist(
      bpu_io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_15_folded_hist),
    .io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_14_folded_hist(
      bpu_io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_14_folded_hist),
    .io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_13_folded_hist(
      bpu_io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_13_folded_hist),
    .io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_12_folded_hist(
      bpu_io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_12_folded_hist),
    .io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_10_folded_hist(
      bpu_io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_10_folded_hist),
    .io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_9_folded_hist(
      bpu_io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_9_folded_hist),
    .io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_8_folded_hist(
      bpu_io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_8_folded_hist),
    .io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_7_folded_hist(
      bpu_io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_7_folded_hist),
    .io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_6_folded_hist(
      bpu_io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_6_folded_hist),
    .io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_5_folded_hist(
      bpu_io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_5_folded_hist),
    .io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_4_folded_hist(
      bpu_io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_4_folded_hist),
    .io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_3_folded_hist(
      bpu_io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_3_folded_hist),
    .io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_2_folded_hist(
      bpu_io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_2_folded_hist),
    .io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_1_folded_hist(
      bpu_io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_1_folded_hist),
    .io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_0_folded_hist(
      bpu_io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_0_folded_hist),
    .io_ftq_to_bpu_update_bits_ftb_entry_valid(bpu_io_ftq_to_bpu_update_bits_ftb_entry_valid),
    .io_ftq_to_bpu_update_bits_ftb_entry_brSlots_0_offset(bpu_io_ftq_to_bpu_update_bits_ftb_entry_brSlots_0_offset),
    .io_ftq_to_bpu_update_bits_ftb_entry_brSlots_0_lower(bpu_io_ftq_to_bpu_update_bits_ftb_entry_brSlots_0_lower),
    .io_ftq_to_bpu_update_bits_ftb_entry_brSlots_0_tarStat(bpu_io_ftq_to_bpu_update_bits_ftb_entry_brSlots_0_tarStat),
    .io_ftq_to_bpu_update_bits_ftb_entry_brSlots_0_sharing(bpu_io_ftq_to_bpu_update_bits_ftb_entry_brSlots_0_sharing),
    .io_ftq_to_bpu_update_bits_ftb_entry_brSlots_0_valid(bpu_io_ftq_to_bpu_update_bits_ftb_entry_brSlots_0_valid),
    .io_ftq_to_bpu_update_bits_ftb_entry_tailSlot_offset(bpu_io_ftq_to_bpu_update_bits_ftb_entry_tailSlot_offset),
    .io_ftq_to_bpu_update_bits_ftb_entry_tailSlot_lower(bpu_io_ftq_to_bpu_update_bits_ftb_entry_tailSlot_lower),
    .io_ftq_to_bpu_update_bits_ftb_entry_tailSlot_tarStat(bpu_io_ftq_to_bpu_update_bits_ftb_entry_tailSlot_tarStat),
    .io_ftq_to_bpu_update_bits_ftb_entry_tailSlot_sharing(bpu_io_ftq_to_bpu_update_bits_ftb_entry_tailSlot_sharing),
    .io_ftq_to_bpu_update_bits_ftb_entry_tailSlot_valid(bpu_io_ftq_to_bpu_update_bits_ftb_entry_tailSlot_valid),
    .io_ftq_to_bpu_update_bits_ftb_entry_pftAddr(bpu_io_ftq_to_bpu_update_bits_ftb_entry_pftAddr),
    .io_ftq_to_bpu_update_bits_ftb_entry_carry(bpu_io_ftq_to_bpu_update_bits_ftb_entry_carry),
    .io_ftq_to_bpu_update_bits_ftb_entry_isCall(bpu_io_ftq_to_bpu_update_bits_ftb_entry_isCall),
    .io_ftq_to_bpu_update_bits_ftb_entry_isRet(bpu_io_ftq_to_bpu_update_bits_ftb_entry_isRet),
    .io_ftq_to_bpu_update_bits_ftb_entry_isJalr(bpu_io_ftq_to_bpu_update_bits_ftb_entry_isJalr),
    .io_ftq_to_bpu_update_bits_ftb_entry_last_may_be_rvi_call(
      bpu_io_ftq_to_bpu_update_bits_ftb_entry_last_may_be_rvi_call),
    .io_ftq_to_bpu_update_bits_ftb_entry_always_taken_0(bpu_io_ftq_to_bpu_update_bits_ftb_entry_always_taken_0),
    .io_ftq_to_bpu_update_bits_ftb_entry_always_taken_1(bpu_io_ftq_to_bpu_update_bits_ftb_entry_always_taken_1),
    .io_ftq_to_bpu_update_bits_br_taken_mask_0(bpu_io_ftq_to_bpu_update_bits_br_taken_mask_0),
    .io_ftq_to_bpu_update_bits_br_taken_mask_1(bpu_io_ftq_to_bpu_update_bits_br_taken_mask_1),
    .io_ftq_to_bpu_update_bits_jmp_taken(bpu_io_ftq_to_bpu_update_bits_jmp_taken),
    .io_ftq_to_bpu_update_bits_mispred_mask_0(bpu_io_ftq_to_bpu_update_bits_mispred_mask_0),
    .io_ftq_to_bpu_update_bits_mispred_mask_1(bpu_io_ftq_to_bpu_update_bits_mispred_mask_1),
    .io_ftq_to_bpu_update_bits_mispred_mask_2(bpu_io_ftq_to_bpu_update_bits_mispred_mask_2),
    .io_ftq_to_bpu_update_bits_old_entry(bpu_io_ftq_to_bpu_update_bits_old_entry),
    .io_ftq_to_bpu_update_bits_meta(bpu_io_ftq_to_bpu_update_bits_meta),
    .io_ftq_to_bpu_update_bits_full_target(bpu_io_ftq_to_bpu_update_bits_full_target),
    .io_ftq_to_bpu_enq_ptr_flag(bpu_io_ftq_to_bpu_enq_ptr_flag),
    .io_ftq_to_bpu_enq_ptr_value(bpu_io_ftq_to_bpu_enq_ptr_value),
    .io_ctrl_ubtb_enable(bpu_io_ctrl_ubtb_enable),
    .io_ctrl_btb_enable(bpu_io_ctrl_btb_enable),
    .io_ctrl_tage_enable(bpu_io_ctrl_tage_enable),
    .io_ctrl_sc_enable(bpu_io_ctrl_sc_enable),
    .io_ctrl_ras_enable(bpu_io_ctrl_ras_enable),
    .io_reset_vector(bpu_io_reset_vector),
    .io_perf_0_value(bpu_io_perf_0_value),
    .io_perf_1_value(bpu_io_perf_1_value),
    .io_perf_2_value(bpu_io_perf_2_value),
    .io_perf_3_value(bpu_io_perf_3_value),
    .io_perf_4_value(bpu_io_perf_4_value),
    .io_perf_5_value(bpu_io_perf_5_value),
    .io_perf_6_value(bpu_io_perf_6_value)
  );
  NewIFU ifu ( // @[Frontend.scala 67:23]
    .clock(ifu_clock),
    .reset(ifu_reset),
    .io_ftqInter_fromFtq_req_ready(ifu_io_ftqInter_fromFtq_req_ready),
    .io_ftqInter_fromFtq_req_valid(ifu_io_ftqInter_fromFtq_req_valid),
    .io_ftqInter_fromFtq_req_bits_startAddr(ifu_io_ftqInter_fromFtq_req_bits_startAddr),
    .io_ftqInter_fromFtq_req_bits_nextlineStart(ifu_io_ftqInter_fromFtq_req_bits_nextlineStart),
    .io_ftqInter_fromFtq_req_bits_nextStartAddr(ifu_io_ftqInter_fromFtq_req_bits_nextStartAddr),
    .io_ftqInter_fromFtq_req_bits_ftqIdx_flag(ifu_io_ftqInter_fromFtq_req_bits_ftqIdx_flag),
    .io_ftqInter_fromFtq_req_bits_ftqIdx_value(ifu_io_ftqInter_fromFtq_req_bits_ftqIdx_value),
    .io_ftqInter_fromFtq_req_bits_ftqOffset_valid(ifu_io_ftqInter_fromFtq_req_bits_ftqOffset_valid),
    .io_ftqInter_fromFtq_req_bits_ftqOffset_bits(ifu_io_ftqInter_fromFtq_req_bits_ftqOffset_bits),
    .io_ftqInter_fromFtq_redirect_valid(ifu_io_ftqInter_fromFtq_redirect_valid),
    .io_ftqInter_fromFtq_redirect_bits_ftqIdx_flag(ifu_io_ftqInter_fromFtq_redirect_bits_ftqIdx_flag),
    .io_ftqInter_fromFtq_redirect_bits_ftqIdx_value(ifu_io_ftqInter_fromFtq_redirect_bits_ftqIdx_value),
    .io_ftqInter_fromFtq_redirect_bits_ftqOffset(ifu_io_ftqInter_fromFtq_redirect_bits_ftqOffset),
    .io_ftqInter_fromFtq_redirect_bits_level(ifu_io_ftqInter_fromFtq_redirect_bits_level),
    .io_ftqInter_fromFtq_flushFromBpu_s2_valid(ifu_io_ftqInter_fromFtq_flushFromBpu_s2_valid),
    .io_ftqInter_fromFtq_flushFromBpu_s2_bits_flag(ifu_io_ftqInter_fromFtq_flushFromBpu_s2_bits_flag),
    .io_ftqInter_fromFtq_flushFromBpu_s2_bits_value(ifu_io_ftqInter_fromFtq_flushFromBpu_s2_bits_value),
    .io_ftqInter_fromFtq_flushFromBpu_s3_valid(ifu_io_ftqInter_fromFtq_flushFromBpu_s3_valid),
    .io_ftqInter_fromFtq_flushFromBpu_s3_bits_flag(ifu_io_ftqInter_fromFtq_flushFromBpu_s3_bits_flag),
    .io_ftqInter_fromFtq_flushFromBpu_s3_bits_value(ifu_io_ftqInter_fromFtq_flushFromBpu_s3_bits_value),
    .io_ftqInter_toFtq_pdWb_valid(ifu_io_ftqInter_toFtq_pdWb_valid),
    .io_ftqInter_toFtq_pdWb_bits_pc_0(ifu_io_ftqInter_toFtq_pdWb_bits_pc_0),
    .io_ftqInter_toFtq_pdWb_bits_pc_1(ifu_io_ftqInter_toFtq_pdWb_bits_pc_1),
    .io_ftqInter_toFtq_pdWb_bits_pc_2(ifu_io_ftqInter_toFtq_pdWb_bits_pc_2),
    .io_ftqInter_toFtq_pdWb_bits_pc_3(ifu_io_ftqInter_toFtq_pdWb_bits_pc_3),
    .io_ftqInter_toFtq_pdWb_bits_pc_4(ifu_io_ftqInter_toFtq_pdWb_bits_pc_4),
    .io_ftqInter_toFtq_pdWb_bits_pc_5(ifu_io_ftqInter_toFtq_pdWb_bits_pc_5),
    .io_ftqInter_toFtq_pdWb_bits_pc_6(ifu_io_ftqInter_toFtq_pdWb_bits_pc_6),
    .io_ftqInter_toFtq_pdWb_bits_pc_7(ifu_io_ftqInter_toFtq_pdWb_bits_pc_7),
    .io_ftqInter_toFtq_pdWb_bits_pd_0_valid(ifu_io_ftqInter_toFtq_pdWb_bits_pd_0_valid),
    .io_ftqInter_toFtq_pdWb_bits_pd_0_isRVC(ifu_io_ftqInter_toFtq_pdWb_bits_pd_0_isRVC),
    .io_ftqInter_toFtq_pdWb_bits_pd_0_brType(ifu_io_ftqInter_toFtq_pdWb_bits_pd_0_brType),
    .io_ftqInter_toFtq_pdWb_bits_pd_0_isCall(ifu_io_ftqInter_toFtq_pdWb_bits_pd_0_isCall),
    .io_ftqInter_toFtq_pdWb_bits_pd_0_isRet(ifu_io_ftqInter_toFtq_pdWb_bits_pd_0_isRet),
    .io_ftqInter_toFtq_pdWb_bits_pd_1_valid(ifu_io_ftqInter_toFtq_pdWb_bits_pd_1_valid),
    .io_ftqInter_toFtq_pdWb_bits_pd_1_isRVC(ifu_io_ftqInter_toFtq_pdWb_bits_pd_1_isRVC),
    .io_ftqInter_toFtq_pdWb_bits_pd_1_brType(ifu_io_ftqInter_toFtq_pdWb_bits_pd_1_brType),
    .io_ftqInter_toFtq_pdWb_bits_pd_1_isCall(ifu_io_ftqInter_toFtq_pdWb_bits_pd_1_isCall),
    .io_ftqInter_toFtq_pdWb_bits_pd_1_isRet(ifu_io_ftqInter_toFtq_pdWb_bits_pd_1_isRet),
    .io_ftqInter_toFtq_pdWb_bits_pd_2_valid(ifu_io_ftqInter_toFtq_pdWb_bits_pd_2_valid),
    .io_ftqInter_toFtq_pdWb_bits_pd_2_isRVC(ifu_io_ftqInter_toFtq_pdWb_bits_pd_2_isRVC),
    .io_ftqInter_toFtq_pdWb_bits_pd_2_brType(ifu_io_ftqInter_toFtq_pdWb_bits_pd_2_brType),
    .io_ftqInter_toFtq_pdWb_bits_pd_2_isCall(ifu_io_ftqInter_toFtq_pdWb_bits_pd_2_isCall),
    .io_ftqInter_toFtq_pdWb_bits_pd_2_isRet(ifu_io_ftqInter_toFtq_pdWb_bits_pd_2_isRet),
    .io_ftqInter_toFtq_pdWb_bits_pd_3_valid(ifu_io_ftqInter_toFtq_pdWb_bits_pd_3_valid),
    .io_ftqInter_toFtq_pdWb_bits_pd_3_isRVC(ifu_io_ftqInter_toFtq_pdWb_bits_pd_3_isRVC),
    .io_ftqInter_toFtq_pdWb_bits_pd_3_brType(ifu_io_ftqInter_toFtq_pdWb_bits_pd_3_brType),
    .io_ftqInter_toFtq_pdWb_bits_pd_3_isCall(ifu_io_ftqInter_toFtq_pdWb_bits_pd_3_isCall),
    .io_ftqInter_toFtq_pdWb_bits_pd_3_isRet(ifu_io_ftqInter_toFtq_pdWb_bits_pd_3_isRet),
    .io_ftqInter_toFtq_pdWb_bits_pd_4_valid(ifu_io_ftqInter_toFtq_pdWb_bits_pd_4_valid),
    .io_ftqInter_toFtq_pdWb_bits_pd_4_isRVC(ifu_io_ftqInter_toFtq_pdWb_bits_pd_4_isRVC),
    .io_ftqInter_toFtq_pdWb_bits_pd_4_brType(ifu_io_ftqInter_toFtq_pdWb_bits_pd_4_brType),
    .io_ftqInter_toFtq_pdWb_bits_pd_4_isCall(ifu_io_ftqInter_toFtq_pdWb_bits_pd_4_isCall),
    .io_ftqInter_toFtq_pdWb_bits_pd_4_isRet(ifu_io_ftqInter_toFtq_pdWb_bits_pd_4_isRet),
    .io_ftqInter_toFtq_pdWb_bits_pd_5_valid(ifu_io_ftqInter_toFtq_pdWb_bits_pd_5_valid),
    .io_ftqInter_toFtq_pdWb_bits_pd_5_isRVC(ifu_io_ftqInter_toFtq_pdWb_bits_pd_5_isRVC),
    .io_ftqInter_toFtq_pdWb_bits_pd_5_brType(ifu_io_ftqInter_toFtq_pdWb_bits_pd_5_brType),
    .io_ftqInter_toFtq_pdWb_bits_pd_5_isCall(ifu_io_ftqInter_toFtq_pdWb_bits_pd_5_isCall),
    .io_ftqInter_toFtq_pdWb_bits_pd_5_isRet(ifu_io_ftqInter_toFtq_pdWb_bits_pd_5_isRet),
    .io_ftqInter_toFtq_pdWb_bits_pd_6_valid(ifu_io_ftqInter_toFtq_pdWb_bits_pd_6_valid),
    .io_ftqInter_toFtq_pdWb_bits_pd_6_isRVC(ifu_io_ftqInter_toFtq_pdWb_bits_pd_6_isRVC),
    .io_ftqInter_toFtq_pdWb_bits_pd_6_brType(ifu_io_ftqInter_toFtq_pdWb_bits_pd_6_brType),
    .io_ftqInter_toFtq_pdWb_bits_pd_6_isCall(ifu_io_ftqInter_toFtq_pdWb_bits_pd_6_isCall),
    .io_ftqInter_toFtq_pdWb_bits_pd_6_isRet(ifu_io_ftqInter_toFtq_pdWb_bits_pd_6_isRet),
    .io_ftqInter_toFtq_pdWb_bits_pd_7_valid(ifu_io_ftqInter_toFtq_pdWb_bits_pd_7_valid),
    .io_ftqInter_toFtq_pdWb_bits_pd_7_isRVC(ifu_io_ftqInter_toFtq_pdWb_bits_pd_7_isRVC),
    .io_ftqInter_toFtq_pdWb_bits_pd_7_brType(ifu_io_ftqInter_toFtq_pdWb_bits_pd_7_brType),
    .io_ftqInter_toFtq_pdWb_bits_pd_7_isCall(ifu_io_ftqInter_toFtq_pdWb_bits_pd_7_isCall),
    .io_ftqInter_toFtq_pdWb_bits_pd_7_isRet(ifu_io_ftqInter_toFtq_pdWb_bits_pd_7_isRet),
    .io_ftqInter_toFtq_pdWb_bits_ftqIdx_flag(ifu_io_ftqInter_toFtq_pdWb_bits_ftqIdx_flag),
    .io_ftqInter_toFtq_pdWb_bits_ftqIdx_value(ifu_io_ftqInter_toFtq_pdWb_bits_ftqIdx_value),
    .io_ftqInter_toFtq_pdWb_bits_misOffset_valid(ifu_io_ftqInter_toFtq_pdWb_bits_misOffset_valid),
    .io_ftqInter_toFtq_pdWb_bits_misOffset_bits(ifu_io_ftqInter_toFtq_pdWb_bits_misOffset_bits),
    .io_ftqInter_toFtq_pdWb_bits_cfiOffset_valid(ifu_io_ftqInter_toFtq_pdWb_bits_cfiOffset_valid),
    .io_ftqInter_toFtq_pdWb_bits_target(ifu_io_ftqInter_toFtq_pdWb_bits_target),
    .io_ftqInter_toFtq_pdWb_bits_jalTarget(ifu_io_ftqInter_toFtq_pdWb_bits_jalTarget),
    .io_ftqInter_toFtq_pdWb_bits_instrRange_0(ifu_io_ftqInter_toFtq_pdWb_bits_instrRange_0),
    .io_ftqInter_toFtq_pdWb_bits_instrRange_1(ifu_io_ftqInter_toFtq_pdWb_bits_instrRange_1),
    .io_ftqInter_toFtq_pdWb_bits_instrRange_2(ifu_io_ftqInter_toFtq_pdWb_bits_instrRange_2),
    .io_ftqInter_toFtq_pdWb_bits_instrRange_3(ifu_io_ftqInter_toFtq_pdWb_bits_instrRange_3),
    .io_ftqInter_toFtq_pdWb_bits_instrRange_4(ifu_io_ftqInter_toFtq_pdWb_bits_instrRange_4),
    .io_ftqInter_toFtq_pdWb_bits_instrRange_5(ifu_io_ftqInter_toFtq_pdWb_bits_instrRange_5),
    .io_ftqInter_toFtq_pdWb_bits_instrRange_6(ifu_io_ftqInter_toFtq_pdWb_bits_instrRange_6),
    .io_ftqInter_toFtq_pdWb_bits_instrRange_7(ifu_io_ftqInter_toFtq_pdWb_bits_instrRange_7),
    .io_icacheInter_icacheReady(ifu_io_icacheInter_icacheReady),
    .io_icacheInter_resp_0_valid(ifu_io_icacheInter_resp_0_valid),
    .io_icacheInter_resp_0_bits_vaddr(ifu_io_icacheInter_resp_0_bits_vaddr),
    .io_icacheInter_resp_0_bits_registerData(ifu_io_icacheInter_resp_0_bits_registerData),
    .io_icacheInter_resp_0_bits_sramData(ifu_io_icacheInter_resp_0_bits_sramData),
    .io_icacheInter_resp_0_bits_select(ifu_io_icacheInter_resp_0_bits_select),
    .io_icacheInter_resp_0_bits_paddr(ifu_io_icacheInter_resp_0_bits_paddr),
    .io_icacheInter_resp_0_bits_tlbExcp_pageFault(ifu_io_icacheInter_resp_0_bits_tlbExcp_pageFault),
    .io_icacheInter_resp_0_bits_tlbExcp_accessFault(ifu_io_icacheInter_resp_0_bits_tlbExcp_accessFault),
    .io_icacheInter_resp_0_bits_tlbExcp_mmio(ifu_io_icacheInter_resp_0_bits_tlbExcp_mmio),
    .io_icacheInter_resp_1_valid(ifu_io_icacheInter_resp_1_valid),
    .io_icacheInter_resp_1_bits_vaddr(ifu_io_icacheInter_resp_1_bits_vaddr),
    .io_icacheInter_resp_1_bits_registerData(ifu_io_icacheInter_resp_1_bits_registerData),
    .io_icacheInter_resp_1_bits_sramData(ifu_io_icacheInter_resp_1_bits_sramData),
    .io_icacheInter_resp_1_bits_select(ifu_io_icacheInter_resp_1_bits_select),
    .io_icacheInter_resp_1_bits_tlbExcp_pageFault(ifu_io_icacheInter_resp_1_bits_tlbExcp_pageFault),
    .io_icacheInter_resp_1_bits_tlbExcp_accessFault(ifu_io_icacheInter_resp_1_bits_tlbExcp_accessFault),
    .io_icacheStop(ifu_io_icacheStop),
    .io_icachePerfInfo_only_0_hit(ifu_io_icachePerfInfo_only_0_hit),
    .io_icachePerfInfo_only_0_miss(ifu_io_icachePerfInfo_only_0_miss),
    .io_icachePerfInfo_hit_0_hit_1(ifu_io_icachePerfInfo_hit_0_hit_1),
    .io_icachePerfInfo_hit_0_miss_1(ifu_io_icachePerfInfo_hit_0_miss_1),
    .io_icachePerfInfo_miss_0_hit_1(ifu_io_icachePerfInfo_miss_0_hit_1),
    .io_icachePerfInfo_miss_0_miss_1(ifu_io_icachePerfInfo_miss_0_miss_1),
    .io_icachePerfInfo_hit_0_except_1(ifu_io_icachePerfInfo_hit_0_except_1),
    .io_icachePerfInfo_miss_0_except_1(ifu_io_icachePerfInfo_miss_0_except_1),
    .io_icachePerfInfo_except_0(ifu_io_icachePerfInfo_except_0),
    .io_icachePerfInfo_bank_hit_1(ifu_io_icachePerfInfo_bank_hit_1),
    .io_icachePerfInfo_hit(ifu_io_icachePerfInfo_hit),
    .io_toIbuffer_ready(ifu_io_toIbuffer_ready),
    .io_toIbuffer_valid(ifu_io_toIbuffer_valid),
    .io_toIbuffer_bits_instrs_0(ifu_io_toIbuffer_bits_instrs_0),
    .io_toIbuffer_bits_instrs_1(ifu_io_toIbuffer_bits_instrs_1),
    .io_toIbuffer_bits_instrs_2(ifu_io_toIbuffer_bits_instrs_2),
    .io_toIbuffer_bits_instrs_3(ifu_io_toIbuffer_bits_instrs_3),
    .io_toIbuffer_bits_instrs_4(ifu_io_toIbuffer_bits_instrs_4),
    .io_toIbuffer_bits_instrs_5(ifu_io_toIbuffer_bits_instrs_5),
    .io_toIbuffer_bits_instrs_6(ifu_io_toIbuffer_bits_instrs_6),
    .io_toIbuffer_bits_instrs_7(ifu_io_toIbuffer_bits_instrs_7),
    .io_toIbuffer_bits_valid(ifu_io_toIbuffer_bits_valid),
    .io_toIbuffer_bits_enqEnable(ifu_io_toIbuffer_bits_enqEnable),
    .io_toIbuffer_bits_pd_0_isRVC(ifu_io_toIbuffer_bits_pd_0_isRVC),
    .io_toIbuffer_bits_pd_0_brType(ifu_io_toIbuffer_bits_pd_0_brType),
    .io_toIbuffer_bits_pd_0_isCall(ifu_io_toIbuffer_bits_pd_0_isCall),
    .io_toIbuffer_bits_pd_0_isRet(ifu_io_toIbuffer_bits_pd_0_isRet),
    .io_toIbuffer_bits_pd_1_isRVC(ifu_io_toIbuffer_bits_pd_1_isRVC),
    .io_toIbuffer_bits_pd_1_brType(ifu_io_toIbuffer_bits_pd_1_brType),
    .io_toIbuffer_bits_pd_1_isCall(ifu_io_toIbuffer_bits_pd_1_isCall),
    .io_toIbuffer_bits_pd_1_isRet(ifu_io_toIbuffer_bits_pd_1_isRet),
    .io_toIbuffer_bits_pd_2_isRVC(ifu_io_toIbuffer_bits_pd_2_isRVC),
    .io_toIbuffer_bits_pd_2_brType(ifu_io_toIbuffer_bits_pd_2_brType),
    .io_toIbuffer_bits_pd_2_isCall(ifu_io_toIbuffer_bits_pd_2_isCall),
    .io_toIbuffer_bits_pd_2_isRet(ifu_io_toIbuffer_bits_pd_2_isRet),
    .io_toIbuffer_bits_pd_3_isRVC(ifu_io_toIbuffer_bits_pd_3_isRVC),
    .io_toIbuffer_bits_pd_3_brType(ifu_io_toIbuffer_bits_pd_3_brType),
    .io_toIbuffer_bits_pd_3_isCall(ifu_io_toIbuffer_bits_pd_3_isCall),
    .io_toIbuffer_bits_pd_3_isRet(ifu_io_toIbuffer_bits_pd_3_isRet),
    .io_toIbuffer_bits_pd_4_isRVC(ifu_io_toIbuffer_bits_pd_4_isRVC),
    .io_toIbuffer_bits_pd_4_brType(ifu_io_toIbuffer_bits_pd_4_brType),
    .io_toIbuffer_bits_pd_4_isCall(ifu_io_toIbuffer_bits_pd_4_isCall),
    .io_toIbuffer_bits_pd_4_isRet(ifu_io_toIbuffer_bits_pd_4_isRet),
    .io_toIbuffer_bits_pd_5_isRVC(ifu_io_toIbuffer_bits_pd_5_isRVC),
    .io_toIbuffer_bits_pd_5_brType(ifu_io_toIbuffer_bits_pd_5_brType),
    .io_toIbuffer_bits_pd_5_isCall(ifu_io_toIbuffer_bits_pd_5_isCall),
    .io_toIbuffer_bits_pd_5_isRet(ifu_io_toIbuffer_bits_pd_5_isRet),
    .io_toIbuffer_bits_pd_6_isRVC(ifu_io_toIbuffer_bits_pd_6_isRVC),
    .io_toIbuffer_bits_pd_6_brType(ifu_io_toIbuffer_bits_pd_6_brType),
    .io_toIbuffer_bits_pd_6_isCall(ifu_io_toIbuffer_bits_pd_6_isCall),
    .io_toIbuffer_bits_pd_6_isRet(ifu_io_toIbuffer_bits_pd_6_isRet),
    .io_toIbuffer_bits_pd_7_isRVC(ifu_io_toIbuffer_bits_pd_7_isRVC),
    .io_toIbuffer_bits_pd_7_brType(ifu_io_toIbuffer_bits_pd_7_brType),
    .io_toIbuffer_bits_pd_7_isCall(ifu_io_toIbuffer_bits_pd_7_isCall),
    .io_toIbuffer_bits_pd_7_isRet(ifu_io_toIbuffer_bits_pd_7_isRet),
    .io_toIbuffer_bits_foldpc_0(ifu_io_toIbuffer_bits_foldpc_0),
    .io_toIbuffer_bits_foldpc_1(ifu_io_toIbuffer_bits_foldpc_1),
    .io_toIbuffer_bits_foldpc_2(ifu_io_toIbuffer_bits_foldpc_2),
    .io_toIbuffer_bits_foldpc_3(ifu_io_toIbuffer_bits_foldpc_3),
    .io_toIbuffer_bits_foldpc_4(ifu_io_toIbuffer_bits_foldpc_4),
    .io_toIbuffer_bits_foldpc_5(ifu_io_toIbuffer_bits_foldpc_5),
    .io_toIbuffer_bits_foldpc_6(ifu_io_toIbuffer_bits_foldpc_6),
    .io_toIbuffer_bits_foldpc_7(ifu_io_toIbuffer_bits_foldpc_7),
    .io_toIbuffer_bits_ftqPtr_flag(ifu_io_toIbuffer_bits_ftqPtr_flag),
    .io_toIbuffer_bits_ftqPtr_value(ifu_io_toIbuffer_bits_ftqPtr_value),
    .io_toIbuffer_bits_ftqOffset_0_valid(ifu_io_toIbuffer_bits_ftqOffset_0_valid),
    .io_toIbuffer_bits_ftqOffset_1_valid(ifu_io_toIbuffer_bits_ftqOffset_1_valid),
    .io_toIbuffer_bits_ftqOffset_2_valid(ifu_io_toIbuffer_bits_ftqOffset_2_valid),
    .io_toIbuffer_bits_ftqOffset_3_valid(ifu_io_toIbuffer_bits_ftqOffset_3_valid),
    .io_toIbuffer_bits_ftqOffset_4_valid(ifu_io_toIbuffer_bits_ftqOffset_4_valid),
    .io_toIbuffer_bits_ftqOffset_5_valid(ifu_io_toIbuffer_bits_ftqOffset_5_valid),
    .io_toIbuffer_bits_ftqOffset_6_valid(ifu_io_toIbuffer_bits_ftqOffset_6_valid),
    .io_toIbuffer_bits_ftqOffset_7_valid(ifu_io_toIbuffer_bits_ftqOffset_7_valid),
    .io_toIbuffer_bits_ipf_0(ifu_io_toIbuffer_bits_ipf_0),
    .io_toIbuffer_bits_ipf_1(ifu_io_toIbuffer_bits_ipf_1),
    .io_toIbuffer_bits_ipf_2(ifu_io_toIbuffer_bits_ipf_2),
    .io_toIbuffer_bits_ipf_3(ifu_io_toIbuffer_bits_ipf_3),
    .io_toIbuffer_bits_ipf_4(ifu_io_toIbuffer_bits_ipf_4),
    .io_toIbuffer_bits_ipf_5(ifu_io_toIbuffer_bits_ipf_5),
    .io_toIbuffer_bits_ipf_6(ifu_io_toIbuffer_bits_ipf_6),
    .io_toIbuffer_bits_ipf_7(ifu_io_toIbuffer_bits_ipf_7),
    .io_toIbuffer_bits_acf_0(ifu_io_toIbuffer_bits_acf_0),
    .io_toIbuffer_bits_acf_1(ifu_io_toIbuffer_bits_acf_1),
    .io_toIbuffer_bits_acf_2(ifu_io_toIbuffer_bits_acf_2),
    .io_toIbuffer_bits_acf_3(ifu_io_toIbuffer_bits_acf_3),
    .io_toIbuffer_bits_acf_4(ifu_io_toIbuffer_bits_acf_4),
    .io_toIbuffer_bits_acf_5(ifu_io_toIbuffer_bits_acf_5),
    .io_toIbuffer_bits_acf_6(ifu_io_toIbuffer_bits_acf_6),
    .io_toIbuffer_bits_acf_7(ifu_io_toIbuffer_bits_acf_7),
    .io_toIbuffer_bits_crossPageIPFFix_0(ifu_io_toIbuffer_bits_crossPageIPFFix_0),
    .io_toIbuffer_bits_crossPageIPFFix_1(ifu_io_toIbuffer_bits_crossPageIPFFix_1),
    .io_toIbuffer_bits_crossPageIPFFix_2(ifu_io_toIbuffer_bits_crossPageIPFFix_2),
    .io_toIbuffer_bits_crossPageIPFFix_3(ifu_io_toIbuffer_bits_crossPageIPFFix_3),
    .io_toIbuffer_bits_crossPageIPFFix_4(ifu_io_toIbuffer_bits_crossPageIPFFix_4),
    .io_toIbuffer_bits_crossPageIPFFix_5(ifu_io_toIbuffer_bits_crossPageIPFFix_5),
    .io_toIbuffer_bits_crossPageIPFFix_6(ifu_io_toIbuffer_bits_crossPageIPFFix_6),
    .io_toIbuffer_bits_crossPageIPFFix_7(ifu_io_toIbuffer_bits_crossPageIPFFix_7),
    .io_toIbuffer_bits_triggered_0_frontendHit_0(ifu_io_toIbuffer_bits_triggered_0_frontendHit_0),
    .io_toIbuffer_bits_triggered_0_frontendHit_1(ifu_io_toIbuffer_bits_triggered_0_frontendHit_1),
    .io_toIbuffer_bits_triggered_0_frontendHit_2(ifu_io_toIbuffer_bits_triggered_0_frontendHit_2),
    .io_toIbuffer_bits_triggered_0_frontendHit_3(ifu_io_toIbuffer_bits_triggered_0_frontendHit_3),
    .io_toIbuffer_bits_triggered_0_backendEn_0(ifu_io_toIbuffer_bits_triggered_0_backendEn_0),
    .io_toIbuffer_bits_triggered_0_backendEn_1(ifu_io_toIbuffer_bits_triggered_0_backendEn_1),
    .io_toIbuffer_bits_triggered_1_frontendHit_0(ifu_io_toIbuffer_bits_triggered_1_frontendHit_0),
    .io_toIbuffer_bits_triggered_1_frontendHit_1(ifu_io_toIbuffer_bits_triggered_1_frontendHit_1),
    .io_toIbuffer_bits_triggered_1_frontendHit_2(ifu_io_toIbuffer_bits_triggered_1_frontendHit_2),
    .io_toIbuffer_bits_triggered_1_frontendHit_3(ifu_io_toIbuffer_bits_triggered_1_frontendHit_3),
    .io_toIbuffer_bits_triggered_1_backendEn_0(ifu_io_toIbuffer_bits_triggered_1_backendEn_0),
    .io_toIbuffer_bits_triggered_1_backendEn_1(ifu_io_toIbuffer_bits_triggered_1_backendEn_1),
    .io_toIbuffer_bits_triggered_2_frontendHit_0(ifu_io_toIbuffer_bits_triggered_2_frontendHit_0),
    .io_toIbuffer_bits_triggered_2_frontendHit_1(ifu_io_toIbuffer_bits_triggered_2_frontendHit_1),
    .io_toIbuffer_bits_triggered_2_frontendHit_2(ifu_io_toIbuffer_bits_triggered_2_frontendHit_2),
    .io_toIbuffer_bits_triggered_2_frontendHit_3(ifu_io_toIbuffer_bits_triggered_2_frontendHit_3),
    .io_toIbuffer_bits_triggered_2_backendEn_0(ifu_io_toIbuffer_bits_triggered_2_backendEn_0),
    .io_toIbuffer_bits_triggered_2_backendEn_1(ifu_io_toIbuffer_bits_triggered_2_backendEn_1),
    .io_toIbuffer_bits_triggered_3_frontendHit_0(ifu_io_toIbuffer_bits_triggered_3_frontendHit_0),
    .io_toIbuffer_bits_triggered_3_frontendHit_1(ifu_io_toIbuffer_bits_triggered_3_frontendHit_1),
    .io_toIbuffer_bits_triggered_3_frontendHit_2(ifu_io_toIbuffer_bits_triggered_3_frontendHit_2),
    .io_toIbuffer_bits_triggered_3_frontendHit_3(ifu_io_toIbuffer_bits_triggered_3_frontendHit_3),
    .io_toIbuffer_bits_triggered_3_backendEn_0(ifu_io_toIbuffer_bits_triggered_3_backendEn_0),
    .io_toIbuffer_bits_triggered_3_backendEn_1(ifu_io_toIbuffer_bits_triggered_3_backendEn_1),
    .io_toIbuffer_bits_triggered_4_frontendHit_0(ifu_io_toIbuffer_bits_triggered_4_frontendHit_0),
    .io_toIbuffer_bits_triggered_4_frontendHit_1(ifu_io_toIbuffer_bits_triggered_4_frontendHit_1),
    .io_toIbuffer_bits_triggered_4_frontendHit_2(ifu_io_toIbuffer_bits_triggered_4_frontendHit_2),
    .io_toIbuffer_bits_triggered_4_frontendHit_3(ifu_io_toIbuffer_bits_triggered_4_frontendHit_3),
    .io_toIbuffer_bits_triggered_4_backendEn_0(ifu_io_toIbuffer_bits_triggered_4_backendEn_0),
    .io_toIbuffer_bits_triggered_4_backendEn_1(ifu_io_toIbuffer_bits_triggered_4_backendEn_1),
    .io_toIbuffer_bits_triggered_5_frontendHit_0(ifu_io_toIbuffer_bits_triggered_5_frontendHit_0),
    .io_toIbuffer_bits_triggered_5_frontendHit_1(ifu_io_toIbuffer_bits_triggered_5_frontendHit_1),
    .io_toIbuffer_bits_triggered_5_frontendHit_2(ifu_io_toIbuffer_bits_triggered_5_frontendHit_2),
    .io_toIbuffer_bits_triggered_5_frontendHit_3(ifu_io_toIbuffer_bits_triggered_5_frontendHit_3),
    .io_toIbuffer_bits_triggered_5_backendEn_0(ifu_io_toIbuffer_bits_triggered_5_backendEn_0),
    .io_toIbuffer_bits_triggered_5_backendEn_1(ifu_io_toIbuffer_bits_triggered_5_backendEn_1),
    .io_toIbuffer_bits_triggered_6_frontendHit_0(ifu_io_toIbuffer_bits_triggered_6_frontendHit_0),
    .io_toIbuffer_bits_triggered_6_frontendHit_1(ifu_io_toIbuffer_bits_triggered_6_frontendHit_1),
    .io_toIbuffer_bits_triggered_6_frontendHit_2(ifu_io_toIbuffer_bits_triggered_6_frontendHit_2),
    .io_toIbuffer_bits_triggered_6_frontendHit_3(ifu_io_toIbuffer_bits_triggered_6_frontendHit_3),
    .io_toIbuffer_bits_triggered_6_backendEn_0(ifu_io_toIbuffer_bits_triggered_6_backendEn_0),
    .io_toIbuffer_bits_triggered_6_backendEn_1(ifu_io_toIbuffer_bits_triggered_6_backendEn_1),
    .io_toIbuffer_bits_triggered_7_frontendHit_0(ifu_io_toIbuffer_bits_triggered_7_frontendHit_0),
    .io_toIbuffer_bits_triggered_7_frontendHit_1(ifu_io_toIbuffer_bits_triggered_7_frontendHit_1),
    .io_toIbuffer_bits_triggered_7_frontendHit_2(ifu_io_toIbuffer_bits_triggered_7_frontendHit_2),
    .io_toIbuffer_bits_triggered_7_frontendHit_3(ifu_io_toIbuffer_bits_triggered_7_frontendHit_3),
    .io_toIbuffer_bits_triggered_7_backendEn_0(ifu_io_toIbuffer_bits_triggered_7_backendEn_0),
    .io_toIbuffer_bits_triggered_7_backendEn_1(ifu_io_toIbuffer_bits_triggered_7_backendEn_1),
    .io_uncacheInter_fromUncache_ready(ifu_io_uncacheInter_fromUncache_ready),
    .io_uncacheInter_fromUncache_valid(ifu_io_uncacheInter_fromUncache_valid),
    .io_uncacheInter_fromUncache_bits_data(ifu_io_uncacheInter_fromUncache_bits_data),
    .io_uncacheInter_toUncache_ready(ifu_io_uncacheInter_toUncache_ready),
    .io_uncacheInter_toUncache_valid(ifu_io_uncacheInter_toUncache_valid),
    .io_uncacheInter_toUncache_bits_addr(ifu_io_uncacheInter_toUncache_bits_addr),
    .io_frontendTrigger_t_valid(ifu_io_frontendTrigger_t_valid),
    .io_frontendTrigger_t_bits_addr(ifu_io_frontendTrigger_t_bits_addr),
    .io_frontendTrigger_t_bits_tdata_matchType(ifu_io_frontendTrigger_t_bits_tdata_matchType),
    .io_frontendTrigger_t_bits_tdata_select(ifu_io_frontendTrigger_t_bits_tdata_select),
    .io_frontendTrigger_t_bits_tdata_timing(ifu_io_frontendTrigger_t_bits_tdata_timing),
    .io_frontendTrigger_t_bits_tdata_chain(ifu_io_frontendTrigger_t_bits_tdata_chain),
    .io_frontendTrigger_t_bits_tdata_tdata2(ifu_io_frontendTrigger_t_bits_tdata_tdata2),
    .io_csrTriggerEnable_0(ifu_io_csrTriggerEnable_0),
    .io_csrTriggerEnable_1(ifu_io_csrTriggerEnable_1),
    .io_csrTriggerEnable_2(ifu_io_csrTriggerEnable_2),
    .io_csrTriggerEnable_3(ifu_io_csrTriggerEnable_3),
    .io_rob_commits_0_valid(ifu_io_rob_commits_0_valid),
    .io_rob_commits_0_bits_ftqIdx_flag(ifu_io_rob_commits_0_bits_ftqIdx_flag),
    .io_rob_commits_0_bits_ftqIdx_value(ifu_io_rob_commits_0_bits_ftqIdx_value),
    .io_rob_commits_0_bits_ftqOffset(ifu_io_rob_commits_0_bits_ftqOffset),
    .io_rob_commits_1_valid(ifu_io_rob_commits_1_valid),
    .io_rob_commits_1_bits_ftqIdx_flag(ifu_io_rob_commits_1_bits_ftqIdx_flag),
    .io_rob_commits_1_bits_ftqIdx_value(ifu_io_rob_commits_1_bits_ftqIdx_value),
    .io_rob_commits_1_bits_ftqOffset(ifu_io_rob_commits_1_bits_ftqOffset),
    .io_iTLBInter_req_valid(ifu_io_iTLBInter_req_valid),
    .io_iTLBInter_req_bits_vaddr(ifu_io_iTLBInter_req_bits_vaddr),
    .io_iTLBInter_resp_bits_paddr_0(ifu_io_iTLBInter_resp_bits_paddr_0),
    .io_iTLBInter_resp_bits_miss(ifu_io_iTLBInter_resp_bits_miss),
    .io_iTLBInter_resp_bits_excp_0_pf_instr(ifu_io_iTLBInter_resp_bits_excp_0_pf_instr),
    .io_iTLBInter_resp_bits_excp_0_af_instr(ifu_io_iTLBInter_resp_bits_excp_0_af_instr),
    .io_pmp_req_bits_addr(ifu_io_pmp_req_bits_addr),
    .io_pmp_resp_instr(ifu_io_pmp_resp_instr),
    .io_pmp_resp_mmio(ifu_io_pmp_resp_mmio),
    .io_mmioCommitRead_mmioFtqPtr_flag(ifu_io_mmioCommitRead_mmioFtqPtr_flag),
    .io_mmioCommitRead_mmioFtqPtr_value(ifu_io_mmioCommitRead_mmioFtqPtr_value),
    .io_mmioCommitRead_mmioLastCommit(ifu_io_mmioCommitRead_mmioLastCommit),
    .io_perf_0_value(ifu_io_perf_0_value),
    .io_perf_1_value(ifu_io_perf_1_value),
    .io_perf_2_value(ifu_io_perf_2_value),
    .io_perf_3_value(ifu_io_perf_3_value),
    .io_perf_4_value(ifu_io_perf_4_value),
    .io_perf_5_value(ifu_io_perf_5_value),
    .io_perf_6_value(ifu_io_perf_6_value),
    .io_perf_7_value(ifu_io_perf_7_value),
    .io_perf_8_value(ifu_io_perf_8_value),
    .io_perf_9_value(ifu_io_perf_9_value),
    .io_perf_10_value(ifu_io_perf_10_value),
    .io_perf_11_value(ifu_io_perf_11_value),
    .io_perf_12_value(ifu_io_perf_12_value)
  );
  Ibuffer ibuffer ( // @[Frontend.scala 68:24]
    .clock(ibuffer_clock),
    .reset(ibuffer_reset),
    .io_flush(ibuffer_io_flush),
    .io_in_ready(ibuffer_io_in_ready),
    .io_in_valid(ibuffer_io_in_valid),
    .io_in_bits_instrs_0(ibuffer_io_in_bits_instrs_0),
    .io_in_bits_instrs_1(ibuffer_io_in_bits_instrs_1),
    .io_in_bits_instrs_2(ibuffer_io_in_bits_instrs_2),
    .io_in_bits_instrs_3(ibuffer_io_in_bits_instrs_3),
    .io_in_bits_instrs_4(ibuffer_io_in_bits_instrs_4),
    .io_in_bits_instrs_5(ibuffer_io_in_bits_instrs_5),
    .io_in_bits_instrs_6(ibuffer_io_in_bits_instrs_6),
    .io_in_bits_instrs_7(ibuffer_io_in_bits_instrs_7),
    .io_in_bits_valid(ibuffer_io_in_bits_valid),
    .io_in_bits_enqEnable(ibuffer_io_in_bits_enqEnable),
    .io_in_bits_pd_0_isRVC(ibuffer_io_in_bits_pd_0_isRVC),
    .io_in_bits_pd_0_brType(ibuffer_io_in_bits_pd_0_brType),
    .io_in_bits_pd_0_isCall(ibuffer_io_in_bits_pd_0_isCall),
    .io_in_bits_pd_0_isRet(ibuffer_io_in_bits_pd_0_isRet),
    .io_in_bits_pd_1_isRVC(ibuffer_io_in_bits_pd_1_isRVC),
    .io_in_bits_pd_1_brType(ibuffer_io_in_bits_pd_1_brType),
    .io_in_bits_pd_1_isCall(ibuffer_io_in_bits_pd_1_isCall),
    .io_in_bits_pd_1_isRet(ibuffer_io_in_bits_pd_1_isRet),
    .io_in_bits_pd_2_isRVC(ibuffer_io_in_bits_pd_2_isRVC),
    .io_in_bits_pd_2_brType(ibuffer_io_in_bits_pd_2_brType),
    .io_in_bits_pd_2_isCall(ibuffer_io_in_bits_pd_2_isCall),
    .io_in_bits_pd_2_isRet(ibuffer_io_in_bits_pd_2_isRet),
    .io_in_bits_pd_3_isRVC(ibuffer_io_in_bits_pd_3_isRVC),
    .io_in_bits_pd_3_brType(ibuffer_io_in_bits_pd_3_brType),
    .io_in_bits_pd_3_isCall(ibuffer_io_in_bits_pd_3_isCall),
    .io_in_bits_pd_3_isRet(ibuffer_io_in_bits_pd_3_isRet),
    .io_in_bits_pd_4_isRVC(ibuffer_io_in_bits_pd_4_isRVC),
    .io_in_bits_pd_4_brType(ibuffer_io_in_bits_pd_4_brType),
    .io_in_bits_pd_4_isCall(ibuffer_io_in_bits_pd_4_isCall),
    .io_in_bits_pd_4_isRet(ibuffer_io_in_bits_pd_4_isRet),
    .io_in_bits_pd_5_isRVC(ibuffer_io_in_bits_pd_5_isRVC),
    .io_in_bits_pd_5_brType(ibuffer_io_in_bits_pd_5_brType),
    .io_in_bits_pd_5_isCall(ibuffer_io_in_bits_pd_5_isCall),
    .io_in_bits_pd_5_isRet(ibuffer_io_in_bits_pd_5_isRet),
    .io_in_bits_pd_6_isRVC(ibuffer_io_in_bits_pd_6_isRVC),
    .io_in_bits_pd_6_brType(ibuffer_io_in_bits_pd_6_brType),
    .io_in_bits_pd_6_isCall(ibuffer_io_in_bits_pd_6_isCall),
    .io_in_bits_pd_6_isRet(ibuffer_io_in_bits_pd_6_isRet),
    .io_in_bits_pd_7_isRVC(ibuffer_io_in_bits_pd_7_isRVC),
    .io_in_bits_pd_7_brType(ibuffer_io_in_bits_pd_7_brType),
    .io_in_bits_pd_7_isCall(ibuffer_io_in_bits_pd_7_isCall),
    .io_in_bits_pd_7_isRet(ibuffer_io_in_bits_pd_7_isRet),
    .io_in_bits_foldpc_0(ibuffer_io_in_bits_foldpc_0),
    .io_in_bits_foldpc_1(ibuffer_io_in_bits_foldpc_1),
    .io_in_bits_foldpc_2(ibuffer_io_in_bits_foldpc_2),
    .io_in_bits_foldpc_3(ibuffer_io_in_bits_foldpc_3),
    .io_in_bits_foldpc_4(ibuffer_io_in_bits_foldpc_4),
    .io_in_bits_foldpc_5(ibuffer_io_in_bits_foldpc_5),
    .io_in_bits_foldpc_6(ibuffer_io_in_bits_foldpc_6),
    .io_in_bits_foldpc_7(ibuffer_io_in_bits_foldpc_7),
    .io_in_bits_ftqPtr_flag(ibuffer_io_in_bits_ftqPtr_flag),
    .io_in_bits_ftqPtr_value(ibuffer_io_in_bits_ftqPtr_value),
    .io_in_bits_ftqOffset_0_valid(ibuffer_io_in_bits_ftqOffset_0_valid),
    .io_in_bits_ftqOffset_1_valid(ibuffer_io_in_bits_ftqOffset_1_valid),
    .io_in_bits_ftqOffset_2_valid(ibuffer_io_in_bits_ftqOffset_2_valid),
    .io_in_bits_ftqOffset_3_valid(ibuffer_io_in_bits_ftqOffset_3_valid),
    .io_in_bits_ftqOffset_4_valid(ibuffer_io_in_bits_ftqOffset_4_valid),
    .io_in_bits_ftqOffset_5_valid(ibuffer_io_in_bits_ftqOffset_5_valid),
    .io_in_bits_ftqOffset_6_valid(ibuffer_io_in_bits_ftqOffset_6_valid),
    .io_in_bits_ftqOffset_7_valid(ibuffer_io_in_bits_ftqOffset_7_valid),
    .io_in_bits_ipf_0(ibuffer_io_in_bits_ipf_0),
    .io_in_bits_ipf_1(ibuffer_io_in_bits_ipf_1),
    .io_in_bits_ipf_2(ibuffer_io_in_bits_ipf_2),
    .io_in_bits_ipf_3(ibuffer_io_in_bits_ipf_3),
    .io_in_bits_ipf_4(ibuffer_io_in_bits_ipf_4),
    .io_in_bits_ipf_5(ibuffer_io_in_bits_ipf_5),
    .io_in_bits_ipf_6(ibuffer_io_in_bits_ipf_6),
    .io_in_bits_ipf_7(ibuffer_io_in_bits_ipf_7),
    .io_in_bits_acf_0(ibuffer_io_in_bits_acf_0),
    .io_in_bits_acf_1(ibuffer_io_in_bits_acf_1),
    .io_in_bits_acf_2(ibuffer_io_in_bits_acf_2),
    .io_in_bits_acf_3(ibuffer_io_in_bits_acf_3),
    .io_in_bits_acf_4(ibuffer_io_in_bits_acf_4),
    .io_in_bits_acf_5(ibuffer_io_in_bits_acf_5),
    .io_in_bits_acf_6(ibuffer_io_in_bits_acf_6),
    .io_in_bits_acf_7(ibuffer_io_in_bits_acf_7),
    .io_in_bits_crossPageIPFFix_0(ibuffer_io_in_bits_crossPageIPFFix_0),
    .io_in_bits_crossPageIPFFix_1(ibuffer_io_in_bits_crossPageIPFFix_1),
    .io_in_bits_crossPageIPFFix_2(ibuffer_io_in_bits_crossPageIPFFix_2),
    .io_in_bits_crossPageIPFFix_3(ibuffer_io_in_bits_crossPageIPFFix_3),
    .io_in_bits_crossPageIPFFix_4(ibuffer_io_in_bits_crossPageIPFFix_4),
    .io_in_bits_crossPageIPFFix_5(ibuffer_io_in_bits_crossPageIPFFix_5),
    .io_in_bits_crossPageIPFFix_6(ibuffer_io_in_bits_crossPageIPFFix_6),
    .io_in_bits_crossPageIPFFix_7(ibuffer_io_in_bits_crossPageIPFFix_7),
    .io_in_bits_triggered_0_frontendHit_0(ibuffer_io_in_bits_triggered_0_frontendHit_0),
    .io_in_bits_triggered_0_frontendHit_1(ibuffer_io_in_bits_triggered_0_frontendHit_1),
    .io_in_bits_triggered_0_frontendHit_2(ibuffer_io_in_bits_triggered_0_frontendHit_2),
    .io_in_bits_triggered_0_frontendHit_3(ibuffer_io_in_bits_triggered_0_frontendHit_3),
    .io_in_bits_triggered_0_backendEn_0(ibuffer_io_in_bits_triggered_0_backendEn_0),
    .io_in_bits_triggered_0_backendEn_1(ibuffer_io_in_bits_triggered_0_backendEn_1),
    .io_in_bits_triggered_1_frontendHit_0(ibuffer_io_in_bits_triggered_1_frontendHit_0),
    .io_in_bits_triggered_1_frontendHit_1(ibuffer_io_in_bits_triggered_1_frontendHit_1),
    .io_in_bits_triggered_1_frontendHit_2(ibuffer_io_in_bits_triggered_1_frontendHit_2),
    .io_in_bits_triggered_1_frontendHit_3(ibuffer_io_in_bits_triggered_1_frontendHit_3),
    .io_in_bits_triggered_1_backendEn_0(ibuffer_io_in_bits_triggered_1_backendEn_0),
    .io_in_bits_triggered_1_backendEn_1(ibuffer_io_in_bits_triggered_1_backendEn_1),
    .io_in_bits_triggered_2_frontendHit_0(ibuffer_io_in_bits_triggered_2_frontendHit_0),
    .io_in_bits_triggered_2_frontendHit_1(ibuffer_io_in_bits_triggered_2_frontendHit_1),
    .io_in_bits_triggered_2_frontendHit_2(ibuffer_io_in_bits_triggered_2_frontendHit_2),
    .io_in_bits_triggered_2_frontendHit_3(ibuffer_io_in_bits_triggered_2_frontendHit_3),
    .io_in_bits_triggered_2_backendEn_0(ibuffer_io_in_bits_triggered_2_backendEn_0),
    .io_in_bits_triggered_2_backendEn_1(ibuffer_io_in_bits_triggered_2_backendEn_1),
    .io_in_bits_triggered_3_frontendHit_0(ibuffer_io_in_bits_triggered_3_frontendHit_0),
    .io_in_bits_triggered_3_frontendHit_1(ibuffer_io_in_bits_triggered_3_frontendHit_1),
    .io_in_bits_triggered_3_frontendHit_2(ibuffer_io_in_bits_triggered_3_frontendHit_2),
    .io_in_bits_triggered_3_frontendHit_3(ibuffer_io_in_bits_triggered_3_frontendHit_3),
    .io_in_bits_triggered_3_backendEn_0(ibuffer_io_in_bits_triggered_3_backendEn_0),
    .io_in_bits_triggered_3_backendEn_1(ibuffer_io_in_bits_triggered_3_backendEn_1),
    .io_in_bits_triggered_4_frontendHit_0(ibuffer_io_in_bits_triggered_4_frontendHit_0),
    .io_in_bits_triggered_4_frontendHit_1(ibuffer_io_in_bits_triggered_4_frontendHit_1),
    .io_in_bits_triggered_4_frontendHit_2(ibuffer_io_in_bits_triggered_4_frontendHit_2),
    .io_in_bits_triggered_4_frontendHit_3(ibuffer_io_in_bits_triggered_4_frontendHit_3),
    .io_in_bits_triggered_4_backendEn_0(ibuffer_io_in_bits_triggered_4_backendEn_0),
    .io_in_bits_triggered_4_backendEn_1(ibuffer_io_in_bits_triggered_4_backendEn_1),
    .io_in_bits_triggered_5_frontendHit_0(ibuffer_io_in_bits_triggered_5_frontendHit_0),
    .io_in_bits_triggered_5_frontendHit_1(ibuffer_io_in_bits_triggered_5_frontendHit_1),
    .io_in_bits_triggered_5_frontendHit_2(ibuffer_io_in_bits_triggered_5_frontendHit_2),
    .io_in_bits_triggered_5_frontendHit_3(ibuffer_io_in_bits_triggered_5_frontendHit_3),
    .io_in_bits_triggered_5_backendEn_0(ibuffer_io_in_bits_triggered_5_backendEn_0),
    .io_in_bits_triggered_5_backendEn_1(ibuffer_io_in_bits_triggered_5_backendEn_1),
    .io_in_bits_triggered_6_frontendHit_0(ibuffer_io_in_bits_triggered_6_frontendHit_0),
    .io_in_bits_triggered_6_frontendHit_1(ibuffer_io_in_bits_triggered_6_frontendHit_1),
    .io_in_bits_triggered_6_frontendHit_2(ibuffer_io_in_bits_triggered_6_frontendHit_2),
    .io_in_bits_triggered_6_frontendHit_3(ibuffer_io_in_bits_triggered_6_frontendHit_3),
    .io_in_bits_triggered_6_backendEn_0(ibuffer_io_in_bits_triggered_6_backendEn_0),
    .io_in_bits_triggered_6_backendEn_1(ibuffer_io_in_bits_triggered_6_backendEn_1),
    .io_in_bits_triggered_7_frontendHit_0(ibuffer_io_in_bits_triggered_7_frontendHit_0),
    .io_in_bits_triggered_7_frontendHit_1(ibuffer_io_in_bits_triggered_7_frontendHit_1),
    .io_in_bits_triggered_7_frontendHit_2(ibuffer_io_in_bits_triggered_7_frontendHit_2),
    .io_in_bits_triggered_7_frontendHit_3(ibuffer_io_in_bits_triggered_7_frontendHit_3),
    .io_in_bits_triggered_7_backendEn_0(ibuffer_io_in_bits_triggered_7_backendEn_0),
    .io_in_bits_triggered_7_backendEn_1(ibuffer_io_in_bits_triggered_7_backendEn_1),
    .io_out_0_ready(ibuffer_io_out_0_ready),
    .io_out_0_valid(ibuffer_io_out_0_valid),
    .io_out_0_bits_instr(ibuffer_io_out_0_bits_instr),
    .io_out_0_bits_foldpc(ibuffer_io_out_0_bits_foldpc),
    .io_out_0_bits_exceptionVec_1(ibuffer_io_out_0_bits_exceptionVec_1),
    .io_out_0_bits_exceptionVec_12(ibuffer_io_out_0_bits_exceptionVec_12),
    .io_out_0_bits_trigger_frontendHit_0(ibuffer_io_out_0_bits_trigger_frontendHit_0),
    .io_out_0_bits_trigger_frontendHit_1(ibuffer_io_out_0_bits_trigger_frontendHit_1),
    .io_out_0_bits_trigger_frontendHit_2(ibuffer_io_out_0_bits_trigger_frontendHit_2),
    .io_out_0_bits_trigger_frontendHit_3(ibuffer_io_out_0_bits_trigger_frontendHit_3),
    .io_out_0_bits_trigger_backendEn_0(ibuffer_io_out_0_bits_trigger_backendEn_0),
    .io_out_0_bits_trigger_backendEn_1(ibuffer_io_out_0_bits_trigger_backendEn_1),
    .io_out_0_bits_pd_isRVC(ibuffer_io_out_0_bits_pd_isRVC),
    .io_out_0_bits_pd_brType(ibuffer_io_out_0_bits_pd_brType),
    .io_out_0_bits_pd_isCall(ibuffer_io_out_0_bits_pd_isCall),
    .io_out_0_bits_pd_isRet(ibuffer_io_out_0_bits_pd_isRet),
    .io_out_0_bits_pred_taken(ibuffer_io_out_0_bits_pred_taken),
    .io_out_0_bits_crossPageIPFFix(ibuffer_io_out_0_bits_crossPageIPFFix),
    .io_out_0_bits_ftqPtr_flag(ibuffer_io_out_0_bits_ftqPtr_flag),
    .io_out_0_bits_ftqPtr_value(ibuffer_io_out_0_bits_ftqPtr_value),
    .io_out_0_bits_ftqOffset(ibuffer_io_out_0_bits_ftqOffset),
    .io_out_1_ready(ibuffer_io_out_1_ready),
    .io_out_1_valid(ibuffer_io_out_1_valid),
    .io_out_1_bits_instr(ibuffer_io_out_1_bits_instr),
    .io_out_1_bits_foldpc(ibuffer_io_out_1_bits_foldpc),
    .io_out_1_bits_exceptionVec_1(ibuffer_io_out_1_bits_exceptionVec_1),
    .io_out_1_bits_exceptionVec_12(ibuffer_io_out_1_bits_exceptionVec_12),
    .io_out_1_bits_trigger_frontendHit_0(ibuffer_io_out_1_bits_trigger_frontendHit_0),
    .io_out_1_bits_trigger_frontendHit_1(ibuffer_io_out_1_bits_trigger_frontendHit_1),
    .io_out_1_bits_trigger_frontendHit_2(ibuffer_io_out_1_bits_trigger_frontendHit_2),
    .io_out_1_bits_trigger_frontendHit_3(ibuffer_io_out_1_bits_trigger_frontendHit_3),
    .io_out_1_bits_trigger_backendEn_0(ibuffer_io_out_1_bits_trigger_backendEn_0),
    .io_out_1_bits_trigger_backendEn_1(ibuffer_io_out_1_bits_trigger_backendEn_1),
    .io_out_1_bits_pd_isRVC(ibuffer_io_out_1_bits_pd_isRVC),
    .io_out_1_bits_pd_brType(ibuffer_io_out_1_bits_pd_brType),
    .io_out_1_bits_pd_isCall(ibuffer_io_out_1_bits_pd_isCall),
    .io_out_1_bits_pd_isRet(ibuffer_io_out_1_bits_pd_isRet),
    .io_out_1_bits_pred_taken(ibuffer_io_out_1_bits_pred_taken),
    .io_out_1_bits_crossPageIPFFix(ibuffer_io_out_1_bits_crossPageIPFFix),
    .io_out_1_bits_ftqPtr_flag(ibuffer_io_out_1_bits_ftqPtr_flag),
    .io_out_1_bits_ftqPtr_value(ibuffer_io_out_1_bits_ftqPtr_value),
    .io_out_1_bits_ftqOffset(ibuffer_io_out_1_bits_ftqOffset),
    .io_perf_0_value(ibuffer_io_perf_0_value),
    .io_perf_1_value(ibuffer_io_perf_1_value),
    .io_perf_2_value(ibuffer_io_perf_2_value),
    .io_perf_3_value(ibuffer_io_perf_3_value),
    .io_perf_4_value(ibuffer_io_perf_4_value),
    .io_perf_5_value(ibuffer_io_perf_5_value),
    .io_perf_6_value(ibuffer_io_perf_6_value),
    .io_perf_7_value(ibuffer_io_perf_7_value)
  );
  Ftq ftq ( // @[Frontend.scala 69:19]
    .clock(ftq_clock),
    .reset(ftq_reset),
    .io_fromBpu_resp_ready(ftq_io_fromBpu_resp_ready),
    .io_fromBpu_resp_valid(ftq_io_fromBpu_resp_valid),
    .io_fromBpu_resp_bits_s1_pc(ftq_io_fromBpu_resp_bits_s1_pc),
    .io_fromBpu_resp_bits_s1_full_pred_br_taken_mask_0(ftq_io_fromBpu_resp_bits_s1_full_pred_br_taken_mask_0),
    .io_fromBpu_resp_bits_s1_full_pred_br_taken_mask_1(ftq_io_fromBpu_resp_bits_s1_full_pred_br_taken_mask_1),
    .io_fromBpu_resp_bits_s1_full_pred_slot_valids_0(ftq_io_fromBpu_resp_bits_s1_full_pred_slot_valids_0),
    .io_fromBpu_resp_bits_s1_full_pred_slot_valids_1(ftq_io_fromBpu_resp_bits_s1_full_pred_slot_valids_1),
    .io_fromBpu_resp_bits_s1_full_pred_targets_0(ftq_io_fromBpu_resp_bits_s1_full_pred_targets_0),
    .io_fromBpu_resp_bits_s1_full_pred_targets_1(ftq_io_fromBpu_resp_bits_s1_full_pred_targets_1),
    .io_fromBpu_resp_bits_s1_full_pred_offsets_0(ftq_io_fromBpu_resp_bits_s1_full_pred_offsets_0),
    .io_fromBpu_resp_bits_s1_full_pred_offsets_1(ftq_io_fromBpu_resp_bits_s1_full_pred_offsets_1),
    .io_fromBpu_resp_bits_s1_full_pred_fallThroughAddr(ftq_io_fromBpu_resp_bits_s1_full_pred_fallThroughAddr),
    .io_fromBpu_resp_bits_s1_full_pred_fallThroughErr(ftq_io_fromBpu_resp_bits_s1_full_pred_fallThroughErr),
    .io_fromBpu_resp_bits_s1_full_pred_is_br_sharing(ftq_io_fromBpu_resp_bits_s1_full_pred_is_br_sharing),
    .io_fromBpu_resp_bits_s1_full_pred_hit(ftq_io_fromBpu_resp_bits_s1_full_pred_hit),
    .io_fromBpu_resp_bits_s2_pc(ftq_io_fromBpu_resp_bits_s2_pc),
    .io_fromBpu_resp_bits_s2_valid(ftq_io_fromBpu_resp_bits_s2_valid),
    .io_fromBpu_resp_bits_s2_hasRedirect(ftq_io_fromBpu_resp_bits_s2_hasRedirect),
    .io_fromBpu_resp_bits_s2_ftq_idx_flag(ftq_io_fromBpu_resp_bits_s2_ftq_idx_flag),
    .io_fromBpu_resp_bits_s2_ftq_idx_value(ftq_io_fromBpu_resp_bits_s2_ftq_idx_value),
    .io_fromBpu_resp_bits_s2_full_pred_br_taken_mask_0(ftq_io_fromBpu_resp_bits_s2_full_pred_br_taken_mask_0),
    .io_fromBpu_resp_bits_s2_full_pred_br_taken_mask_1(ftq_io_fromBpu_resp_bits_s2_full_pred_br_taken_mask_1),
    .io_fromBpu_resp_bits_s2_full_pred_slot_valids_0(ftq_io_fromBpu_resp_bits_s2_full_pred_slot_valids_0),
    .io_fromBpu_resp_bits_s2_full_pred_slot_valids_1(ftq_io_fromBpu_resp_bits_s2_full_pred_slot_valids_1),
    .io_fromBpu_resp_bits_s2_full_pred_targets_0(ftq_io_fromBpu_resp_bits_s2_full_pred_targets_0),
    .io_fromBpu_resp_bits_s2_full_pred_targets_1(ftq_io_fromBpu_resp_bits_s2_full_pred_targets_1),
    .io_fromBpu_resp_bits_s2_full_pred_offsets_0(ftq_io_fromBpu_resp_bits_s2_full_pred_offsets_0),
    .io_fromBpu_resp_bits_s2_full_pred_offsets_1(ftq_io_fromBpu_resp_bits_s2_full_pred_offsets_1),
    .io_fromBpu_resp_bits_s2_full_pred_fallThroughAddr(ftq_io_fromBpu_resp_bits_s2_full_pred_fallThroughAddr),
    .io_fromBpu_resp_bits_s2_full_pred_fallThroughErr(ftq_io_fromBpu_resp_bits_s2_full_pred_fallThroughErr),
    .io_fromBpu_resp_bits_s2_full_pred_is_br_sharing(ftq_io_fromBpu_resp_bits_s2_full_pred_is_br_sharing),
    .io_fromBpu_resp_bits_s2_full_pred_hit(ftq_io_fromBpu_resp_bits_s2_full_pred_hit),
    .io_fromBpu_resp_bits_s3_pc(ftq_io_fromBpu_resp_bits_s3_pc),
    .io_fromBpu_resp_bits_s3_valid(ftq_io_fromBpu_resp_bits_s3_valid),
    .io_fromBpu_resp_bits_s3_hasRedirect(ftq_io_fromBpu_resp_bits_s3_hasRedirect),
    .io_fromBpu_resp_bits_s3_ftq_idx_flag(ftq_io_fromBpu_resp_bits_s3_ftq_idx_flag),
    .io_fromBpu_resp_bits_s3_ftq_idx_value(ftq_io_fromBpu_resp_bits_s3_ftq_idx_value),
    .io_fromBpu_resp_bits_s3_full_pred_br_taken_mask_0(ftq_io_fromBpu_resp_bits_s3_full_pred_br_taken_mask_0),
    .io_fromBpu_resp_bits_s3_full_pred_br_taken_mask_1(ftq_io_fromBpu_resp_bits_s3_full_pred_br_taken_mask_1),
    .io_fromBpu_resp_bits_s3_full_pred_slot_valids_0(ftq_io_fromBpu_resp_bits_s3_full_pred_slot_valids_0),
    .io_fromBpu_resp_bits_s3_full_pred_slot_valids_1(ftq_io_fromBpu_resp_bits_s3_full_pred_slot_valids_1),
    .io_fromBpu_resp_bits_s3_full_pred_targets_0(ftq_io_fromBpu_resp_bits_s3_full_pred_targets_0),
    .io_fromBpu_resp_bits_s3_full_pred_targets_1(ftq_io_fromBpu_resp_bits_s3_full_pred_targets_1),
    .io_fromBpu_resp_bits_s3_full_pred_offsets_0(ftq_io_fromBpu_resp_bits_s3_full_pred_offsets_0),
    .io_fromBpu_resp_bits_s3_full_pred_offsets_1(ftq_io_fromBpu_resp_bits_s3_full_pred_offsets_1),
    .io_fromBpu_resp_bits_s3_full_pred_fallThroughAddr(ftq_io_fromBpu_resp_bits_s3_full_pred_fallThroughAddr),
    .io_fromBpu_resp_bits_s3_full_pred_fallThroughErr(ftq_io_fromBpu_resp_bits_s3_full_pred_fallThroughErr),
    .io_fromBpu_resp_bits_s3_full_pred_is_br_sharing(ftq_io_fromBpu_resp_bits_s3_full_pred_is_br_sharing),
    .io_fromBpu_resp_bits_s3_full_pred_hit(ftq_io_fromBpu_resp_bits_s3_full_pred_hit),
    .io_fromBpu_resp_bits_last_stage_meta(ftq_io_fromBpu_resp_bits_last_stage_meta),
    .io_fromBpu_resp_bits_last_stage_spec_info_folded_hist_hist_17_folded_hist(
      ftq_io_fromBpu_resp_bits_last_stage_spec_info_folded_hist_hist_17_folded_hist),
    .io_fromBpu_resp_bits_last_stage_spec_info_folded_hist_hist_16_folded_hist(
      ftq_io_fromBpu_resp_bits_last_stage_spec_info_folded_hist_hist_16_folded_hist),
    .io_fromBpu_resp_bits_last_stage_spec_info_folded_hist_hist_15_folded_hist(
      ftq_io_fromBpu_resp_bits_last_stage_spec_info_folded_hist_hist_15_folded_hist),
    .io_fromBpu_resp_bits_last_stage_spec_info_folded_hist_hist_14_folded_hist(
      ftq_io_fromBpu_resp_bits_last_stage_spec_info_folded_hist_hist_14_folded_hist),
    .io_fromBpu_resp_bits_last_stage_spec_info_folded_hist_hist_13_folded_hist(
      ftq_io_fromBpu_resp_bits_last_stage_spec_info_folded_hist_hist_13_folded_hist),
    .io_fromBpu_resp_bits_last_stage_spec_info_folded_hist_hist_12_folded_hist(
      ftq_io_fromBpu_resp_bits_last_stage_spec_info_folded_hist_hist_12_folded_hist),
    .io_fromBpu_resp_bits_last_stage_spec_info_folded_hist_hist_11_folded_hist(
      ftq_io_fromBpu_resp_bits_last_stage_spec_info_folded_hist_hist_11_folded_hist),
    .io_fromBpu_resp_bits_last_stage_spec_info_folded_hist_hist_10_folded_hist(
      ftq_io_fromBpu_resp_bits_last_stage_spec_info_folded_hist_hist_10_folded_hist),
    .io_fromBpu_resp_bits_last_stage_spec_info_folded_hist_hist_9_folded_hist(
      ftq_io_fromBpu_resp_bits_last_stage_spec_info_folded_hist_hist_9_folded_hist),
    .io_fromBpu_resp_bits_last_stage_spec_info_folded_hist_hist_8_folded_hist(
      ftq_io_fromBpu_resp_bits_last_stage_spec_info_folded_hist_hist_8_folded_hist),
    .io_fromBpu_resp_bits_last_stage_spec_info_folded_hist_hist_7_folded_hist(
      ftq_io_fromBpu_resp_bits_last_stage_spec_info_folded_hist_hist_7_folded_hist),
    .io_fromBpu_resp_bits_last_stage_spec_info_folded_hist_hist_6_folded_hist(
      ftq_io_fromBpu_resp_bits_last_stage_spec_info_folded_hist_hist_6_folded_hist),
    .io_fromBpu_resp_bits_last_stage_spec_info_folded_hist_hist_5_folded_hist(
      ftq_io_fromBpu_resp_bits_last_stage_spec_info_folded_hist_hist_5_folded_hist),
    .io_fromBpu_resp_bits_last_stage_spec_info_folded_hist_hist_4_folded_hist(
      ftq_io_fromBpu_resp_bits_last_stage_spec_info_folded_hist_hist_4_folded_hist),
    .io_fromBpu_resp_bits_last_stage_spec_info_folded_hist_hist_3_folded_hist(
      ftq_io_fromBpu_resp_bits_last_stage_spec_info_folded_hist_hist_3_folded_hist),
    .io_fromBpu_resp_bits_last_stage_spec_info_folded_hist_hist_2_folded_hist(
      ftq_io_fromBpu_resp_bits_last_stage_spec_info_folded_hist_hist_2_folded_hist),
    .io_fromBpu_resp_bits_last_stage_spec_info_folded_hist_hist_1_folded_hist(
      ftq_io_fromBpu_resp_bits_last_stage_spec_info_folded_hist_hist_1_folded_hist),
    .io_fromBpu_resp_bits_last_stage_spec_info_folded_hist_hist_0_folded_hist(
      ftq_io_fromBpu_resp_bits_last_stage_spec_info_folded_hist_hist_0_folded_hist),
    .io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_5_bits_0(
      ftq_io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_5_bits_0),
    .io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_5_bits_1(
      ftq_io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_5_bits_1),
    .io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_5_bits_2(
      ftq_io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_5_bits_2),
    .io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_5_bits_3(
      ftq_io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_5_bits_3),
    .io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_4_bits_0(
      ftq_io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_4_bits_0),
    .io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_4_bits_1(
      ftq_io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_4_bits_1),
    .io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_4_bits_2(
      ftq_io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_4_bits_2),
    .io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_4_bits_3(
      ftq_io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_4_bits_3),
    .io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_3_bits_0(
      ftq_io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_3_bits_0),
    .io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_3_bits_1(
      ftq_io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_3_bits_1),
    .io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_3_bits_2(
      ftq_io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_3_bits_2),
    .io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_3_bits_3(
      ftq_io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_3_bits_3),
    .io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_2_bits_0(
      ftq_io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_2_bits_0),
    .io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_2_bits_1(
      ftq_io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_2_bits_1),
    .io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_2_bits_2(
      ftq_io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_2_bits_2),
    .io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_2_bits_3(
      ftq_io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_2_bits_3),
    .io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_1_bits_0(
      ftq_io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_1_bits_0),
    .io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_1_bits_1(
      ftq_io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_1_bits_1),
    .io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_1_bits_2(
      ftq_io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_1_bits_2),
    .io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_1_bits_3(
      ftq_io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_1_bits_3),
    .io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_0_bits_0(
      ftq_io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_0_bits_0),
    .io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_0_bits_1(
      ftq_io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_0_bits_1),
    .io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_0_bits_2(
      ftq_io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_0_bits_2),
    .io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_0_bits_3(
      ftq_io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_0_bits_3),
    .io_fromBpu_resp_bits_last_stage_spec_info_lastBrNumOH(ftq_io_fromBpu_resp_bits_last_stage_spec_info_lastBrNumOH),
    .io_fromBpu_resp_bits_last_stage_spec_info_histPtr_flag(ftq_io_fromBpu_resp_bits_last_stage_spec_info_histPtr_flag),
    .io_fromBpu_resp_bits_last_stage_spec_info_histPtr_value(ftq_io_fromBpu_resp_bits_last_stage_spec_info_histPtr_value
      ),
    .io_fromBpu_resp_bits_last_stage_spec_info_rasSp(ftq_io_fromBpu_resp_bits_last_stage_spec_info_rasSp),
    .io_fromBpu_resp_bits_last_stage_spec_info_rasTop_retAddr(
      ftq_io_fromBpu_resp_bits_last_stage_spec_info_rasTop_retAddr),
    .io_fromBpu_resp_bits_last_stage_spec_info_rasTop_ctr(ftq_io_fromBpu_resp_bits_last_stage_spec_info_rasTop_ctr),
    .io_fromBpu_resp_bits_last_stage_ftb_entry_valid(ftq_io_fromBpu_resp_bits_last_stage_ftb_entry_valid),
    .io_fromBpu_resp_bits_last_stage_ftb_entry_brSlots_0_offset(
      ftq_io_fromBpu_resp_bits_last_stage_ftb_entry_brSlots_0_offset),
    .io_fromBpu_resp_bits_last_stage_ftb_entry_brSlots_0_lower(
      ftq_io_fromBpu_resp_bits_last_stage_ftb_entry_brSlots_0_lower),
    .io_fromBpu_resp_bits_last_stage_ftb_entry_brSlots_0_tarStat(
      ftq_io_fromBpu_resp_bits_last_stage_ftb_entry_brSlots_0_tarStat),
    .io_fromBpu_resp_bits_last_stage_ftb_entry_brSlots_0_sharing(
      ftq_io_fromBpu_resp_bits_last_stage_ftb_entry_brSlots_0_sharing),
    .io_fromBpu_resp_bits_last_stage_ftb_entry_brSlots_0_valid(
      ftq_io_fromBpu_resp_bits_last_stage_ftb_entry_brSlots_0_valid),
    .io_fromBpu_resp_bits_last_stage_ftb_entry_tailSlot_offset(
      ftq_io_fromBpu_resp_bits_last_stage_ftb_entry_tailSlot_offset),
    .io_fromBpu_resp_bits_last_stage_ftb_entry_tailSlot_lower(
      ftq_io_fromBpu_resp_bits_last_stage_ftb_entry_tailSlot_lower),
    .io_fromBpu_resp_bits_last_stage_ftb_entry_tailSlot_tarStat(
      ftq_io_fromBpu_resp_bits_last_stage_ftb_entry_tailSlot_tarStat),
    .io_fromBpu_resp_bits_last_stage_ftb_entry_tailSlot_sharing(
      ftq_io_fromBpu_resp_bits_last_stage_ftb_entry_tailSlot_sharing),
    .io_fromBpu_resp_bits_last_stage_ftb_entry_tailSlot_valid(
      ftq_io_fromBpu_resp_bits_last_stage_ftb_entry_tailSlot_valid),
    .io_fromBpu_resp_bits_last_stage_ftb_entry_pftAddr(ftq_io_fromBpu_resp_bits_last_stage_ftb_entry_pftAddr),
    .io_fromBpu_resp_bits_last_stage_ftb_entry_carry(ftq_io_fromBpu_resp_bits_last_stage_ftb_entry_carry),
    .io_fromBpu_resp_bits_last_stage_ftb_entry_isCall(ftq_io_fromBpu_resp_bits_last_stage_ftb_entry_isCall),
    .io_fromBpu_resp_bits_last_stage_ftb_entry_isRet(ftq_io_fromBpu_resp_bits_last_stage_ftb_entry_isRet),
    .io_fromBpu_resp_bits_last_stage_ftb_entry_isJalr(ftq_io_fromBpu_resp_bits_last_stage_ftb_entry_isJalr),
    .io_fromBpu_resp_bits_last_stage_ftb_entry_last_may_be_rvi_call(
      ftq_io_fromBpu_resp_bits_last_stage_ftb_entry_last_may_be_rvi_call),
    .io_fromBpu_resp_bits_last_stage_ftb_entry_always_taken_0(
      ftq_io_fromBpu_resp_bits_last_stage_ftb_entry_always_taken_0),
    .io_fromBpu_resp_bits_last_stage_ftb_entry_always_taken_1(
      ftq_io_fromBpu_resp_bits_last_stage_ftb_entry_always_taken_1),
    .io_fromIfu_pdWb_valid(ftq_io_fromIfu_pdWb_valid),
    .io_fromIfu_pdWb_bits_pc_0(ftq_io_fromIfu_pdWb_bits_pc_0),
    .io_fromIfu_pdWb_bits_pc_1(ftq_io_fromIfu_pdWb_bits_pc_1),
    .io_fromIfu_pdWb_bits_pc_2(ftq_io_fromIfu_pdWb_bits_pc_2),
    .io_fromIfu_pdWb_bits_pc_3(ftq_io_fromIfu_pdWb_bits_pc_3),
    .io_fromIfu_pdWb_bits_pc_4(ftq_io_fromIfu_pdWb_bits_pc_4),
    .io_fromIfu_pdWb_bits_pc_5(ftq_io_fromIfu_pdWb_bits_pc_5),
    .io_fromIfu_pdWb_bits_pc_6(ftq_io_fromIfu_pdWb_bits_pc_6),
    .io_fromIfu_pdWb_bits_pc_7(ftq_io_fromIfu_pdWb_bits_pc_7),
    .io_fromIfu_pdWb_bits_pd_0_valid(ftq_io_fromIfu_pdWb_bits_pd_0_valid),
    .io_fromIfu_pdWb_bits_pd_0_isRVC(ftq_io_fromIfu_pdWb_bits_pd_0_isRVC),
    .io_fromIfu_pdWb_bits_pd_0_brType(ftq_io_fromIfu_pdWb_bits_pd_0_brType),
    .io_fromIfu_pdWb_bits_pd_0_isCall(ftq_io_fromIfu_pdWb_bits_pd_0_isCall),
    .io_fromIfu_pdWb_bits_pd_0_isRet(ftq_io_fromIfu_pdWb_bits_pd_0_isRet),
    .io_fromIfu_pdWb_bits_pd_1_valid(ftq_io_fromIfu_pdWb_bits_pd_1_valid),
    .io_fromIfu_pdWb_bits_pd_1_isRVC(ftq_io_fromIfu_pdWb_bits_pd_1_isRVC),
    .io_fromIfu_pdWb_bits_pd_1_brType(ftq_io_fromIfu_pdWb_bits_pd_1_brType),
    .io_fromIfu_pdWb_bits_pd_1_isCall(ftq_io_fromIfu_pdWb_bits_pd_1_isCall),
    .io_fromIfu_pdWb_bits_pd_1_isRet(ftq_io_fromIfu_pdWb_bits_pd_1_isRet),
    .io_fromIfu_pdWb_bits_pd_2_valid(ftq_io_fromIfu_pdWb_bits_pd_2_valid),
    .io_fromIfu_pdWb_bits_pd_2_isRVC(ftq_io_fromIfu_pdWb_bits_pd_2_isRVC),
    .io_fromIfu_pdWb_bits_pd_2_brType(ftq_io_fromIfu_pdWb_bits_pd_2_brType),
    .io_fromIfu_pdWb_bits_pd_2_isCall(ftq_io_fromIfu_pdWb_bits_pd_2_isCall),
    .io_fromIfu_pdWb_bits_pd_2_isRet(ftq_io_fromIfu_pdWb_bits_pd_2_isRet),
    .io_fromIfu_pdWb_bits_pd_3_valid(ftq_io_fromIfu_pdWb_bits_pd_3_valid),
    .io_fromIfu_pdWb_bits_pd_3_isRVC(ftq_io_fromIfu_pdWb_bits_pd_3_isRVC),
    .io_fromIfu_pdWb_bits_pd_3_brType(ftq_io_fromIfu_pdWb_bits_pd_3_brType),
    .io_fromIfu_pdWb_bits_pd_3_isCall(ftq_io_fromIfu_pdWb_bits_pd_3_isCall),
    .io_fromIfu_pdWb_bits_pd_3_isRet(ftq_io_fromIfu_pdWb_bits_pd_3_isRet),
    .io_fromIfu_pdWb_bits_pd_4_valid(ftq_io_fromIfu_pdWb_bits_pd_4_valid),
    .io_fromIfu_pdWb_bits_pd_4_isRVC(ftq_io_fromIfu_pdWb_bits_pd_4_isRVC),
    .io_fromIfu_pdWb_bits_pd_4_brType(ftq_io_fromIfu_pdWb_bits_pd_4_brType),
    .io_fromIfu_pdWb_bits_pd_4_isCall(ftq_io_fromIfu_pdWb_bits_pd_4_isCall),
    .io_fromIfu_pdWb_bits_pd_4_isRet(ftq_io_fromIfu_pdWb_bits_pd_4_isRet),
    .io_fromIfu_pdWb_bits_pd_5_valid(ftq_io_fromIfu_pdWb_bits_pd_5_valid),
    .io_fromIfu_pdWb_bits_pd_5_isRVC(ftq_io_fromIfu_pdWb_bits_pd_5_isRVC),
    .io_fromIfu_pdWb_bits_pd_5_brType(ftq_io_fromIfu_pdWb_bits_pd_5_brType),
    .io_fromIfu_pdWb_bits_pd_5_isCall(ftq_io_fromIfu_pdWb_bits_pd_5_isCall),
    .io_fromIfu_pdWb_bits_pd_5_isRet(ftq_io_fromIfu_pdWb_bits_pd_5_isRet),
    .io_fromIfu_pdWb_bits_pd_6_valid(ftq_io_fromIfu_pdWb_bits_pd_6_valid),
    .io_fromIfu_pdWb_bits_pd_6_isRVC(ftq_io_fromIfu_pdWb_bits_pd_6_isRVC),
    .io_fromIfu_pdWb_bits_pd_6_brType(ftq_io_fromIfu_pdWb_bits_pd_6_brType),
    .io_fromIfu_pdWb_bits_pd_6_isCall(ftq_io_fromIfu_pdWb_bits_pd_6_isCall),
    .io_fromIfu_pdWb_bits_pd_6_isRet(ftq_io_fromIfu_pdWb_bits_pd_6_isRet),
    .io_fromIfu_pdWb_bits_pd_7_valid(ftq_io_fromIfu_pdWb_bits_pd_7_valid),
    .io_fromIfu_pdWb_bits_pd_7_isRVC(ftq_io_fromIfu_pdWb_bits_pd_7_isRVC),
    .io_fromIfu_pdWb_bits_pd_7_brType(ftq_io_fromIfu_pdWb_bits_pd_7_brType),
    .io_fromIfu_pdWb_bits_pd_7_isCall(ftq_io_fromIfu_pdWb_bits_pd_7_isCall),
    .io_fromIfu_pdWb_bits_pd_7_isRet(ftq_io_fromIfu_pdWb_bits_pd_7_isRet),
    .io_fromIfu_pdWb_bits_ftqIdx_flag(ftq_io_fromIfu_pdWb_bits_ftqIdx_flag),
    .io_fromIfu_pdWb_bits_ftqIdx_value(ftq_io_fromIfu_pdWb_bits_ftqIdx_value),
    .io_fromIfu_pdWb_bits_misOffset_valid(ftq_io_fromIfu_pdWb_bits_misOffset_valid),
    .io_fromIfu_pdWb_bits_misOffset_bits(ftq_io_fromIfu_pdWb_bits_misOffset_bits),
    .io_fromIfu_pdWb_bits_cfiOffset_valid(ftq_io_fromIfu_pdWb_bits_cfiOffset_valid),
    .io_fromIfu_pdWb_bits_target(ftq_io_fromIfu_pdWb_bits_target),
    .io_fromIfu_pdWb_bits_jalTarget(ftq_io_fromIfu_pdWb_bits_jalTarget),
    .io_fromIfu_pdWb_bits_instrRange_0(ftq_io_fromIfu_pdWb_bits_instrRange_0),
    .io_fromIfu_pdWb_bits_instrRange_1(ftq_io_fromIfu_pdWb_bits_instrRange_1),
    .io_fromIfu_pdWb_bits_instrRange_2(ftq_io_fromIfu_pdWb_bits_instrRange_2),
    .io_fromIfu_pdWb_bits_instrRange_3(ftq_io_fromIfu_pdWb_bits_instrRange_3),
    .io_fromIfu_pdWb_bits_instrRange_4(ftq_io_fromIfu_pdWb_bits_instrRange_4),
    .io_fromIfu_pdWb_bits_instrRange_5(ftq_io_fromIfu_pdWb_bits_instrRange_5),
    .io_fromIfu_pdWb_bits_instrRange_6(ftq_io_fromIfu_pdWb_bits_instrRange_6),
    .io_fromIfu_pdWb_bits_instrRange_7(ftq_io_fromIfu_pdWb_bits_instrRange_7),
    .io_fromBackend_rob_commits_0_valid(ftq_io_fromBackend_rob_commits_0_valid),
    .io_fromBackend_rob_commits_0_bits_commitType(ftq_io_fromBackend_rob_commits_0_bits_commitType),
    .io_fromBackend_rob_commits_0_bits_ftqIdx_flag(ftq_io_fromBackend_rob_commits_0_bits_ftqIdx_flag),
    .io_fromBackend_rob_commits_0_bits_ftqIdx_value(ftq_io_fromBackend_rob_commits_0_bits_ftqIdx_value),
    .io_fromBackend_rob_commits_0_bits_ftqOffset(ftq_io_fromBackend_rob_commits_0_bits_ftqOffset),
    .io_fromBackend_rob_commits_1_valid(ftq_io_fromBackend_rob_commits_1_valid),
    .io_fromBackend_rob_commits_1_bits_commitType(ftq_io_fromBackend_rob_commits_1_bits_commitType),
    .io_fromBackend_rob_commits_1_bits_ftqIdx_flag(ftq_io_fromBackend_rob_commits_1_bits_ftqIdx_flag),
    .io_fromBackend_rob_commits_1_bits_ftqIdx_value(ftq_io_fromBackend_rob_commits_1_bits_ftqIdx_value),
    .io_fromBackend_rob_commits_1_bits_ftqOffset(ftq_io_fromBackend_rob_commits_1_bits_ftqOffset),
    .io_fromBackend_redirect_valid(ftq_io_fromBackend_redirect_valid),
    .io_fromBackend_redirect_bits_ftqIdx_flag(ftq_io_fromBackend_redirect_bits_ftqIdx_flag),
    .io_fromBackend_redirect_bits_ftqIdx_value(ftq_io_fromBackend_redirect_bits_ftqIdx_value),
    .io_fromBackend_redirect_bits_ftqOffset(ftq_io_fromBackend_redirect_bits_ftqOffset),
    .io_fromBackend_redirect_bits_level(ftq_io_fromBackend_redirect_bits_level),
    .io_fromBackend_redirect_bits_cfiUpdate_pc(ftq_io_fromBackend_redirect_bits_cfiUpdate_pc),
    .io_fromBackend_redirect_bits_cfiUpdate_pd_isRVC(ftq_io_fromBackend_redirect_bits_cfiUpdate_pd_isRVC),
    .io_fromBackend_redirect_bits_cfiUpdate_pd_brType(ftq_io_fromBackend_redirect_bits_cfiUpdate_pd_brType),
    .io_fromBackend_redirect_bits_cfiUpdate_pd_isCall(ftq_io_fromBackend_redirect_bits_cfiUpdate_pd_isCall),
    .io_fromBackend_redirect_bits_cfiUpdate_pd_isRet(ftq_io_fromBackend_redirect_bits_cfiUpdate_pd_isRet),
    .io_fromBackend_redirect_bits_cfiUpdate_target(ftq_io_fromBackend_redirect_bits_cfiUpdate_target),
    .io_fromBackend_redirect_bits_cfiUpdate_taken(ftq_io_fromBackend_redirect_bits_cfiUpdate_taken),
    .io_fromBackend_redirect_bits_cfiUpdate_isMisPred(ftq_io_fromBackend_redirect_bits_cfiUpdate_isMisPred),
    .io_toBpu_redirect_valid(ftq_io_toBpu_redirect_valid),
    .io_toBpu_redirect_bits_level(ftq_io_toBpu_redirect_bits_level),
    .io_toBpu_redirect_bits_cfiUpdate_pc(ftq_io_toBpu_redirect_bits_cfiUpdate_pc),
    .io_toBpu_redirect_bits_cfiUpdate_pd_isRVC(ftq_io_toBpu_redirect_bits_cfiUpdate_pd_isRVC),
    .io_toBpu_redirect_bits_cfiUpdate_pd_isCall(ftq_io_toBpu_redirect_bits_cfiUpdate_pd_isCall),
    .io_toBpu_redirect_bits_cfiUpdate_pd_isRet(ftq_io_toBpu_redirect_bits_cfiUpdate_pd_isRet),
    .io_toBpu_redirect_bits_cfiUpdate_rasSp(ftq_io_toBpu_redirect_bits_cfiUpdate_rasSp),
    .io_toBpu_redirect_bits_cfiUpdate_rasEntry_retAddr(ftq_io_toBpu_redirect_bits_cfiUpdate_rasEntry_retAddr),
    .io_toBpu_redirect_bits_cfiUpdate_rasEntry_ctr(ftq_io_toBpu_redirect_bits_cfiUpdate_rasEntry_ctr),
    .io_toBpu_redirect_bits_cfiUpdate_folded_hist_hist_17_folded_hist(
      ftq_io_toBpu_redirect_bits_cfiUpdate_folded_hist_hist_17_folded_hist),
    .io_toBpu_redirect_bits_cfiUpdate_folded_hist_hist_16_folded_hist(
      ftq_io_toBpu_redirect_bits_cfiUpdate_folded_hist_hist_16_folded_hist),
    .io_toBpu_redirect_bits_cfiUpdate_folded_hist_hist_15_folded_hist(
      ftq_io_toBpu_redirect_bits_cfiUpdate_folded_hist_hist_15_folded_hist),
    .io_toBpu_redirect_bits_cfiUpdate_folded_hist_hist_14_folded_hist(
      ftq_io_toBpu_redirect_bits_cfiUpdate_folded_hist_hist_14_folded_hist),
    .io_toBpu_redirect_bits_cfiUpdate_folded_hist_hist_13_folded_hist(
      ftq_io_toBpu_redirect_bits_cfiUpdate_folded_hist_hist_13_folded_hist),
    .io_toBpu_redirect_bits_cfiUpdate_folded_hist_hist_12_folded_hist(
      ftq_io_toBpu_redirect_bits_cfiUpdate_folded_hist_hist_12_folded_hist),
    .io_toBpu_redirect_bits_cfiUpdate_folded_hist_hist_11_folded_hist(
      ftq_io_toBpu_redirect_bits_cfiUpdate_folded_hist_hist_11_folded_hist),
    .io_toBpu_redirect_bits_cfiUpdate_folded_hist_hist_10_folded_hist(
      ftq_io_toBpu_redirect_bits_cfiUpdate_folded_hist_hist_10_folded_hist),
    .io_toBpu_redirect_bits_cfiUpdate_folded_hist_hist_9_folded_hist(
      ftq_io_toBpu_redirect_bits_cfiUpdate_folded_hist_hist_9_folded_hist),
    .io_toBpu_redirect_bits_cfiUpdate_folded_hist_hist_8_folded_hist(
      ftq_io_toBpu_redirect_bits_cfiUpdate_folded_hist_hist_8_folded_hist),
    .io_toBpu_redirect_bits_cfiUpdate_folded_hist_hist_7_folded_hist(
      ftq_io_toBpu_redirect_bits_cfiUpdate_folded_hist_hist_7_folded_hist),
    .io_toBpu_redirect_bits_cfiUpdate_folded_hist_hist_6_folded_hist(
      ftq_io_toBpu_redirect_bits_cfiUpdate_folded_hist_hist_6_folded_hist),
    .io_toBpu_redirect_bits_cfiUpdate_folded_hist_hist_5_folded_hist(
      ftq_io_toBpu_redirect_bits_cfiUpdate_folded_hist_hist_5_folded_hist),
    .io_toBpu_redirect_bits_cfiUpdate_folded_hist_hist_4_folded_hist(
      ftq_io_toBpu_redirect_bits_cfiUpdate_folded_hist_hist_4_folded_hist),
    .io_toBpu_redirect_bits_cfiUpdate_folded_hist_hist_3_folded_hist(
      ftq_io_toBpu_redirect_bits_cfiUpdate_folded_hist_hist_3_folded_hist),
    .io_toBpu_redirect_bits_cfiUpdate_folded_hist_hist_2_folded_hist(
      ftq_io_toBpu_redirect_bits_cfiUpdate_folded_hist_hist_2_folded_hist),
    .io_toBpu_redirect_bits_cfiUpdate_folded_hist_hist_1_folded_hist(
      ftq_io_toBpu_redirect_bits_cfiUpdate_folded_hist_hist_1_folded_hist),
    .io_toBpu_redirect_bits_cfiUpdate_folded_hist_hist_0_folded_hist(
      ftq_io_toBpu_redirect_bits_cfiUpdate_folded_hist_hist_0_folded_hist),
    .io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_5_bits_0(ftq_io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_5_bits_0),
    .io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_5_bits_1(ftq_io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_5_bits_1),
    .io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_5_bits_2(ftq_io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_5_bits_2),
    .io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_5_bits_3(ftq_io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_5_bits_3),
    .io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_4_bits_0(ftq_io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_4_bits_0),
    .io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_4_bits_1(ftq_io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_4_bits_1),
    .io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_4_bits_2(ftq_io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_4_bits_2),
    .io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_3_bits_0(ftq_io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_3_bits_0),
    .io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_3_bits_1(ftq_io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_3_bits_1),
    .io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_3_bits_2(ftq_io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_3_bits_2),
    .io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_3_bits_3(ftq_io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_3_bits_3),
    .io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_2_bits_0(ftq_io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_2_bits_0),
    .io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_2_bits_1(ftq_io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_2_bits_1),
    .io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_2_bits_2(ftq_io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_2_bits_2),
    .io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_2_bits_3(ftq_io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_2_bits_3),
    .io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_1_bits_0(ftq_io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_1_bits_0),
    .io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_1_bits_1(ftq_io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_1_bits_1),
    .io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_1_bits_2(ftq_io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_1_bits_2),
    .io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_1_bits_3(ftq_io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_1_bits_3),
    .io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_0_bits_0(ftq_io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_0_bits_0),
    .io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_0_bits_1(ftq_io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_0_bits_1),
    .io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_0_bits_2(ftq_io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_0_bits_2),
    .io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_0_bits_3(ftq_io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_0_bits_3),
    .io_toBpu_redirect_bits_cfiUpdate_lastBrNumOH(ftq_io_toBpu_redirect_bits_cfiUpdate_lastBrNumOH),
    .io_toBpu_redirect_bits_cfiUpdate_histPtr_flag(ftq_io_toBpu_redirect_bits_cfiUpdate_histPtr_flag),
    .io_toBpu_redirect_bits_cfiUpdate_histPtr_value(ftq_io_toBpu_redirect_bits_cfiUpdate_histPtr_value),
    .io_toBpu_redirect_bits_cfiUpdate_target(ftq_io_toBpu_redirect_bits_cfiUpdate_target),
    .io_toBpu_redirect_bits_cfiUpdate_taken(ftq_io_toBpu_redirect_bits_cfiUpdate_taken),
    .io_toBpu_redirect_bits_cfiUpdate_shift(ftq_io_toBpu_redirect_bits_cfiUpdate_shift),
    .io_toBpu_redirect_bits_cfiUpdate_addIntoHist(ftq_io_toBpu_redirect_bits_cfiUpdate_addIntoHist),
    .io_toBpu_update_valid(ftq_io_toBpu_update_valid),
    .io_toBpu_update_bits_pc(ftq_io_toBpu_update_bits_pc),
    .io_toBpu_update_bits_spec_info_folded_hist_hist_17_folded_hist(
      ftq_io_toBpu_update_bits_spec_info_folded_hist_hist_17_folded_hist),
    .io_toBpu_update_bits_spec_info_folded_hist_hist_16_folded_hist(
      ftq_io_toBpu_update_bits_spec_info_folded_hist_hist_16_folded_hist),
    .io_toBpu_update_bits_spec_info_folded_hist_hist_15_folded_hist(
      ftq_io_toBpu_update_bits_spec_info_folded_hist_hist_15_folded_hist),
    .io_toBpu_update_bits_spec_info_folded_hist_hist_14_folded_hist(
      ftq_io_toBpu_update_bits_spec_info_folded_hist_hist_14_folded_hist),
    .io_toBpu_update_bits_spec_info_folded_hist_hist_13_folded_hist(
      ftq_io_toBpu_update_bits_spec_info_folded_hist_hist_13_folded_hist),
    .io_toBpu_update_bits_spec_info_folded_hist_hist_12_folded_hist(
      ftq_io_toBpu_update_bits_spec_info_folded_hist_hist_12_folded_hist),
    .io_toBpu_update_bits_spec_info_folded_hist_hist_10_folded_hist(
      ftq_io_toBpu_update_bits_spec_info_folded_hist_hist_10_folded_hist),
    .io_toBpu_update_bits_spec_info_folded_hist_hist_9_folded_hist(
      ftq_io_toBpu_update_bits_spec_info_folded_hist_hist_9_folded_hist),
    .io_toBpu_update_bits_spec_info_folded_hist_hist_8_folded_hist(
      ftq_io_toBpu_update_bits_spec_info_folded_hist_hist_8_folded_hist),
    .io_toBpu_update_bits_spec_info_folded_hist_hist_7_folded_hist(
      ftq_io_toBpu_update_bits_spec_info_folded_hist_hist_7_folded_hist),
    .io_toBpu_update_bits_spec_info_folded_hist_hist_6_folded_hist(
      ftq_io_toBpu_update_bits_spec_info_folded_hist_hist_6_folded_hist),
    .io_toBpu_update_bits_spec_info_folded_hist_hist_5_folded_hist(
      ftq_io_toBpu_update_bits_spec_info_folded_hist_hist_5_folded_hist),
    .io_toBpu_update_bits_spec_info_folded_hist_hist_4_folded_hist(
      ftq_io_toBpu_update_bits_spec_info_folded_hist_hist_4_folded_hist),
    .io_toBpu_update_bits_spec_info_folded_hist_hist_3_folded_hist(
      ftq_io_toBpu_update_bits_spec_info_folded_hist_hist_3_folded_hist),
    .io_toBpu_update_bits_spec_info_folded_hist_hist_2_folded_hist(
      ftq_io_toBpu_update_bits_spec_info_folded_hist_hist_2_folded_hist),
    .io_toBpu_update_bits_spec_info_folded_hist_hist_1_folded_hist(
      ftq_io_toBpu_update_bits_spec_info_folded_hist_hist_1_folded_hist),
    .io_toBpu_update_bits_spec_info_folded_hist_hist_0_folded_hist(
      ftq_io_toBpu_update_bits_spec_info_folded_hist_hist_0_folded_hist),
    .io_toBpu_update_bits_ftb_entry_valid(ftq_io_toBpu_update_bits_ftb_entry_valid),
    .io_toBpu_update_bits_ftb_entry_brSlots_0_offset(ftq_io_toBpu_update_bits_ftb_entry_brSlots_0_offset),
    .io_toBpu_update_bits_ftb_entry_brSlots_0_lower(ftq_io_toBpu_update_bits_ftb_entry_brSlots_0_lower),
    .io_toBpu_update_bits_ftb_entry_brSlots_0_tarStat(ftq_io_toBpu_update_bits_ftb_entry_brSlots_0_tarStat),
    .io_toBpu_update_bits_ftb_entry_brSlots_0_sharing(ftq_io_toBpu_update_bits_ftb_entry_brSlots_0_sharing),
    .io_toBpu_update_bits_ftb_entry_brSlots_0_valid(ftq_io_toBpu_update_bits_ftb_entry_brSlots_0_valid),
    .io_toBpu_update_bits_ftb_entry_tailSlot_offset(ftq_io_toBpu_update_bits_ftb_entry_tailSlot_offset),
    .io_toBpu_update_bits_ftb_entry_tailSlot_lower(ftq_io_toBpu_update_bits_ftb_entry_tailSlot_lower),
    .io_toBpu_update_bits_ftb_entry_tailSlot_tarStat(ftq_io_toBpu_update_bits_ftb_entry_tailSlot_tarStat),
    .io_toBpu_update_bits_ftb_entry_tailSlot_sharing(ftq_io_toBpu_update_bits_ftb_entry_tailSlot_sharing),
    .io_toBpu_update_bits_ftb_entry_tailSlot_valid(ftq_io_toBpu_update_bits_ftb_entry_tailSlot_valid),
    .io_toBpu_update_bits_ftb_entry_pftAddr(ftq_io_toBpu_update_bits_ftb_entry_pftAddr),
    .io_toBpu_update_bits_ftb_entry_carry(ftq_io_toBpu_update_bits_ftb_entry_carry),
    .io_toBpu_update_bits_ftb_entry_isCall(ftq_io_toBpu_update_bits_ftb_entry_isCall),
    .io_toBpu_update_bits_ftb_entry_isRet(ftq_io_toBpu_update_bits_ftb_entry_isRet),
    .io_toBpu_update_bits_ftb_entry_isJalr(ftq_io_toBpu_update_bits_ftb_entry_isJalr),
    .io_toBpu_update_bits_ftb_entry_last_may_be_rvi_call(ftq_io_toBpu_update_bits_ftb_entry_last_may_be_rvi_call),
    .io_toBpu_update_bits_ftb_entry_always_taken_0(ftq_io_toBpu_update_bits_ftb_entry_always_taken_0),
    .io_toBpu_update_bits_ftb_entry_always_taken_1(ftq_io_toBpu_update_bits_ftb_entry_always_taken_1),
    .io_toBpu_update_bits_br_taken_mask_0(ftq_io_toBpu_update_bits_br_taken_mask_0),
    .io_toBpu_update_bits_br_taken_mask_1(ftq_io_toBpu_update_bits_br_taken_mask_1),
    .io_toBpu_update_bits_jmp_taken(ftq_io_toBpu_update_bits_jmp_taken),
    .io_toBpu_update_bits_mispred_mask_0(ftq_io_toBpu_update_bits_mispred_mask_0),
    .io_toBpu_update_bits_mispred_mask_1(ftq_io_toBpu_update_bits_mispred_mask_1),
    .io_toBpu_update_bits_mispred_mask_2(ftq_io_toBpu_update_bits_mispred_mask_2),
    .io_toBpu_update_bits_false_hit(ftq_io_toBpu_update_bits_false_hit),
    .io_toBpu_update_bits_old_entry(ftq_io_toBpu_update_bits_old_entry),
    .io_toBpu_update_bits_meta(ftq_io_toBpu_update_bits_meta),
    .io_toBpu_update_bits_full_target(ftq_io_toBpu_update_bits_full_target),
    .io_toBpu_enq_ptr_flag(ftq_io_toBpu_enq_ptr_flag),
    .io_toBpu_enq_ptr_value(ftq_io_toBpu_enq_ptr_value),
    .io_toIfu_req_ready(ftq_io_toIfu_req_ready),
    .io_toIfu_req_valid(ftq_io_toIfu_req_valid),
    .io_toIfu_req_bits_startAddr(ftq_io_toIfu_req_bits_startAddr),
    .io_toIfu_req_bits_nextlineStart(ftq_io_toIfu_req_bits_nextlineStart),
    .io_toIfu_req_bits_nextStartAddr(ftq_io_toIfu_req_bits_nextStartAddr),
    .io_toIfu_req_bits_ftqIdx_flag(ftq_io_toIfu_req_bits_ftqIdx_flag),
    .io_toIfu_req_bits_ftqIdx_value(ftq_io_toIfu_req_bits_ftqIdx_value),
    .io_toIfu_req_bits_ftqOffset_valid(ftq_io_toIfu_req_bits_ftqOffset_valid),
    .io_toIfu_req_bits_ftqOffset_bits(ftq_io_toIfu_req_bits_ftqOffset_bits),
    .io_toIfu_redirect_valid(ftq_io_toIfu_redirect_valid),
    .io_toIfu_redirect_bits_ftqIdx_flag(ftq_io_toIfu_redirect_bits_ftqIdx_flag),
    .io_toIfu_redirect_bits_ftqIdx_value(ftq_io_toIfu_redirect_bits_ftqIdx_value),
    .io_toIfu_redirect_bits_ftqOffset(ftq_io_toIfu_redirect_bits_ftqOffset),
    .io_toIfu_redirect_bits_level(ftq_io_toIfu_redirect_bits_level),
    .io_toIfu_flushFromBpu_s2_valid(ftq_io_toIfu_flushFromBpu_s2_valid),
    .io_toIfu_flushFromBpu_s2_bits_flag(ftq_io_toIfu_flushFromBpu_s2_bits_flag),
    .io_toIfu_flushFromBpu_s2_bits_value(ftq_io_toIfu_flushFromBpu_s2_bits_value),
    .io_toIfu_flushFromBpu_s3_valid(ftq_io_toIfu_flushFromBpu_s3_valid),
    .io_toIfu_flushFromBpu_s3_bits_flag(ftq_io_toIfu_flushFromBpu_s3_bits_flag),
    .io_toIfu_flushFromBpu_s3_bits_value(ftq_io_toIfu_flushFromBpu_s3_bits_value),
    .io_toICache_req_valid(ftq_io_toICache_req_valid),
    .io_toICache_req_bits_pcMemRead_0_startAddr(ftq_io_toICache_req_bits_pcMemRead_0_startAddr),
    .io_toICache_req_bits_pcMemRead_0_nextlineStart(ftq_io_toICache_req_bits_pcMemRead_0_nextlineStart),
    .io_toICache_req_bits_pcMemRead_1_startAddr(ftq_io_toICache_req_bits_pcMemRead_1_startAddr),
    .io_toICache_req_bits_pcMemRead_1_nextlineStart(ftq_io_toICache_req_bits_pcMemRead_1_nextlineStart),
    .io_toICache_req_bits_pcMemRead_2_startAddr(ftq_io_toICache_req_bits_pcMemRead_2_startAddr),
    .io_toICache_req_bits_pcMemRead_2_nextlineStart(ftq_io_toICache_req_bits_pcMemRead_2_nextlineStart),
    .io_toICache_req_bits_pcMemRead_3_startAddr(ftq_io_toICache_req_bits_pcMemRead_3_startAddr),
    .io_toICache_req_bits_pcMemRead_3_nextlineStart(ftq_io_toICache_req_bits_pcMemRead_3_nextlineStart),
    .io_toICache_req_bits_pcMemRead_4_startAddr(ftq_io_toICache_req_bits_pcMemRead_4_startAddr),
    .io_toICache_req_bits_pcMemRead_4_nextlineStart(ftq_io_toICache_req_bits_pcMemRead_4_nextlineStart),
    .io_toICache_req_bits_readValid_0(ftq_io_toICache_req_bits_readValid_0),
    .io_toICache_req_bits_readValid_1(ftq_io_toICache_req_bits_readValid_1),
    .io_toICache_req_bits_readValid_2(ftq_io_toICache_req_bits_readValid_2),
    .io_toICache_req_bits_readValid_3(ftq_io_toICache_req_bits_readValid_3),
    .io_toICache_req_bits_readValid_4(ftq_io_toICache_req_bits_readValid_4),
    .io_toBackend_pc_mem_wen(ftq_io_toBackend_pc_mem_wen),
    .io_toBackend_pc_mem_waddr(ftq_io_toBackend_pc_mem_waddr),
    .io_toBackend_pc_mem_wdata_startAddr(ftq_io_toBackend_pc_mem_wdata_startAddr),
    .io_toBackend_pc_mem_wdata_nextLineAddr(ftq_io_toBackend_pc_mem_wdata_nextLineAddr),
    .io_toBackend_pc_mem_wdata_isNextMask_0(ftq_io_toBackend_pc_mem_wdata_isNextMask_0),
    .io_toBackend_pc_mem_wdata_isNextMask_1(ftq_io_toBackend_pc_mem_wdata_isNextMask_1),
    .io_toBackend_pc_mem_wdata_isNextMask_2(ftq_io_toBackend_pc_mem_wdata_isNextMask_2),
    .io_toBackend_pc_mem_wdata_isNextMask_3(ftq_io_toBackend_pc_mem_wdata_isNextMask_3),
    .io_toBackend_pc_mem_wdata_isNextMask_4(ftq_io_toBackend_pc_mem_wdata_isNextMask_4),
    .io_toBackend_pc_mem_wdata_isNextMask_5(ftq_io_toBackend_pc_mem_wdata_isNextMask_5),
    .io_toBackend_pc_mem_wdata_isNextMask_6(ftq_io_toBackend_pc_mem_wdata_isNextMask_6),
    .io_toBackend_pc_mem_wdata_isNextMask_7(ftq_io_toBackend_pc_mem_wdata_isNextMask_7),
    .io_toBackend_newest_entry_target(ftq_io_toBackend_newest_entry_target),
    .io_toBackend_newest_entry_ptr_flag(ftq_io_toBackend_newest_entry_ptr_flag),
    .io_toBackend_newest_entry_ptr_value(ftq_io_toBackend_newest_entry_ptr_value),
    .io_mmioCommitRead_mmioFtqPtr_flag(ftq_io_mmioCommitRead_mmioFtqPtr_flag),
    .io_mmioCommitRead_mmioFtqPtr_value(ftq_io_mmioCommitRead_mmioFtqPtr_value),
    .io_mmioCommitRead_mmioLastCommit(ftq_io_mmioCommitRead_mmioLastCommit),
    .io_perf_0_value(ftq_io_perf_0_value),
    .io_perf_1_value(ftq_io_perf_1_value),
    .io_perf_2_value(ftq_io_perf_2_value),
    .io_perf_3_value(ftq_io_perf_3_value),
    .io_perf_4_value(ftq_io_perf_4_value),
    .io_perf_5_value(ftq_io_perf_5_value),
    .io_perf_6_value(ftq_io_perf_6_value),
    .io_perf_7_value(ftq_io_perf_7_value),
    .io_perf_8_value(ftq_io_perf_8_value),
    .io_perf_9_value(ftq_io_perf_9_value),
    .io_perf_10_value(ftq_io_perf_10_value),
    .io_perf_11_value(ftq_io_perf_11_value),
    .io_perf_12_value(ftq_io_perf_12_value),
    .io_perf_13_value(ftq_io_perf_13_value),
    .io_perf_14_value(ftq_io_perf_14_value),
    .io_perf_15_value(ftq_io_perf_15_value),
    .io_perf_16_value(ftq_io_perf_16_value),
    .io_perf_17_value(ftq_io_perf_17_value),
    .io_perf_18_value(ftq_io_perf_18_value),
    .io_perf_19_value(ftq_io_perf_19_value),
    .io_perf_20_value(ftq_io_perf_20_value),
    .io_perf_21_value(ftq_io_perf_21_value),
    .io_perf_22_value(ftq_io_perf_22_value),
    .io_perf_23_value(ftq_io_perf_23_value)
  );
  DelayN_17 tlbCsr_delay ( // @[Hold.scala 97:23]
    .clock(tlbCsr_delay_clock),
    .io_in_satp_mode(tlbCsr_delay_io_in_satp_mode),
    .io_in_satp_asid(tlbCsr_delay_io_in_satp_asid),
    .io_in_satp_ppn(tlbCsr_delay_io_in_satp_ppn),
    .io_in_satp_changed(tlbCsr_delay_io_in_satp_changed),
    .io_in_priv_mxr(tlbCsr_delay_io_in_priv_mxr),
    .io_in_priv_sum(tlbCsr_delay_io_in_priv_sum),
    .io_in_priv_imode(tlbCsr_delay_io_in_priv_imode),
    .io_in_priv_dmode(tlbCsr_delay_io_in_priv_dmode),
    .io_out_satp_mode(tlbCsr_delay_io_out_satp_mode),
    .io_out_satp_asid(tlbCsr_delay_io_out_satp_asid),
    .io_out_satp_ppn(tlbCsr_delay_io_out_satp_ppn),
    .io_out_satp_changed(tlbCsr_delay_io_out_satp_changed),
    .io_out_priv_mxr(tlbCsr_delay_io_out_priv_mxr),
    .io_out_priv_sum(tlbCsr_delay_io_out_priv_sum),
    .io_out_priv_imode(tlbCsr_delay_io_out_priv_imode),
    .io_out_priv_dmode(tlbCsr_delay_io_out_priv_dmode)
  );
  DelayN_18 csrCtrl_delay ( // @[Hold.scala 97:23]
    .clock(csrCtrl_delay_clock),
    .io_in_icache_parity_enable(csrCtrl_delay_io_in_icache_parity_enable),
    .io_in_lvpred_disable(csrCtrl_delay_io_in_lvpred_disable),
    .io_in_no_spec_load(csrCtrl_delay_io_in_no_spec_load),
    .io_in_storeset_wait_store(csrCtrl_delay_io_in_storeset_wait_store),
    .io_in_lvpred_timeout(csrCtrl_delay_io_in_lvpred_timeout),
    .io_in_bp_ctrl_ubtb_enable(csrCtrl_delay_io_in_bp_ctrl_ubtb_enable),
    .io_in_bp_ctrl_btb_enable(csrCtrl_delay_io_in_bp_ctrl_btb_enable),
    .io_in_bp_ctrl_tage_enable(csrCtrl_delay_io_in_bp_ctrl_tage_enable),
    .io_in_bp_ctrl_sc_enable(csrCtrl_delay_io_in_bp_ctrl_sc_enable),
    .io_in_bp_ctrl_ras_enable(csrCtrl_delay_io_in_bp_ctrl_ras_enable),
    .io_in_sbuffer_threshold(csrCtrl_delay_io_in_sbuffer_threshold),
    .io_in_ldld_vio_check_enable(csrCtrl_delay_io_in_ldld_vio_check_enable),
    .io_in_cache_error_enable(csrCtrl_delay_io_in_cache_error_enable),
    .io_in_uncache_write_outstanding_enable(csrCtrl_delay_io_in_uncache_write_outstanding_enable),
    .io_in_fusion_enable(csrCtrl_delay_io_in_fusion_enable),
    .io_in_wfi_enable(csrCtrl_delay_io_in_wfi_enable),
    .io_in_svinval_enable(csrCtrl_delay_io_in_svinval_enable),
    .io_in_distribute_csr_wvalid(csrCtrl_delay_io_in_distribute_csr_wvalid),
    .io_in_distribute_csr_waddr(csrCtrl_delay_io_in_distribute_csr_waddr),
    .io_in_distribute_csr_wdata(csrCtrl_delay_io_in_distribute_csr_wdata),
    .io_in_singlestep(csrCtrl_delay_io_in_singlestep),
    .io_in_frontend_trigger_t_valid(csrCtrl_delay_io_in_frontend_trigger_t_valid),
    .io_in_frontend_trigger_t_bits_addr(csrCtrl_delay_io_in_frontend_trigger_t_bits_addr),
    .io_in_frontend_trigger_t_bits_tdata_matchType(csrCtrl_delay_io_in_frontend_trigger_t_bits_tdata_matchType),
    .io_in_frontend_trigger_t_bits_tdata_select(csrCtrl_delay_io_in_frontend_trigger_t_bits_tdata_select),
    .io_in_frontend_trigger_t_bits_tdata_timing(csrCtrl_delay_io_in_frontend_trigger_t_bits_tdata_timing),
    .io_in_frontend_trigger_t_bits_tdata_chain(csrCtrl_delay_io_in_frontend_trigger_t_bits_tdata_chain),
    .io_in_frontend_trigger_t_bits_tdata_tdata2(csrCtrl_delay_io_in_frontend_trigger_t_bits_tdata_tdata2),
    .io_in_mem_trigger_t_valid(csrCtrl_delay_io_in_mem_trigger_t_valid),
    .io_in_mem_trigger_t_bits_addr(csrCtrl_delay_io_in_mem_trigger_t_bits_addr),
    .io_in_mem_trigger_t_bits_tdata_matchType(csrCtrl_delay_io_in_mem_trigger_t_bits_tdata_matchType),
    .io_in_mem_trigger_t_bits_tdata_select(csrCtrl_delay_io_in_mem_trigger_t_bits_tdata_select),
    .io_in_mem_trigger_t_bits_tdata_chain(csrCtrl_delay_io_in_mem_trigger_t_bits_tdata_chain),
    .io_in_mem_trigger_t_bits_tdata_tdata2(csrCtrl_delay_io_in_mem_trigger_t_bits_tdata_tdata2),
    .io_in_trigger_enable_0(csrCtrl_delay_io_in_trigger_enable_0),
    .io_in_trigger_enable_1(csrCtrl_delay_io_in_trigger_enable_1),
    .io_in_trigger_enable_2(csrCtrl_delay_io_in_trigger_enable_2),
    .io_in_trigger_enable_3(csrCtrl_delay_io_in_trigger_enable_3),
    .io_in_trigger_enable_4(csrCtrl_delay_io_in_trigger_enable_4),
    .io_in_trigger_enable_5(csrCtrl_delay_io_in_trigger_enable_5),
    .io_in_trigger_enable_6(csrCtrl_delay_io_in_trigger_enable_6),
    .io_in_trigger_enable_7(csrCtrl_delay_io_in_trigger_enable_7),
    .io_in_trigger_enable_8(csrCtrl_delay_io_in_trigger_enable_8),
    .io_in_trigger_enable_9(csrCtrl_delay_io_in_trigger_enable_9),
    .io_out_icache_parity_enable(csrCtrl_delay_io_out_icache_parity_enable),
    .io_out_lvpred_disable(csrCtrl_delay_io_out_lvpred_disable),
    .io_out_no_spec_load(csrCtrl_delay_io_out_no_spec_load),
    .io_out_storeset_wait_store(csrCtrl_delay_io_out_storeset_wait_store),
    .io_out_lvpred_timeout(csrCtrl_delay_io_out_lvpred_timeout),
    .io_out_bp_ctrl_ubtb_enable(csrCtrl_delay_io_out_bp_ctrl_ubtb_enable),
    .io_out_bp_ctrl_btb_enable(csrCtrl_delay_io_out_bp_ctrl_btb_enable),
    .io_out_bp_ctrl_tage_enable(csrCtrl_delay_io_out_bp_ctrl_tage_enable),
    .io_out_bp_ctrl_sc_enable(csrCtrl_delay_io_out_bp_ctrl_sc_enable),
    .io_out_bp_ctrl_ras_enable(csrCtrl_delay_io_out_bp_ctrl_ras_enable),
    .io_out_sbuffer_threshold(csrCtrl_delay_io_out_sbuffer_threshold),
    .io_out_ldld_vio_check_enable(csrCtrl_delay_io_out_ldld_vio_check_enable),
    .io_out_cache_error_enable(csrCtrl_delay_io_out_cache_error_enable),
    .io_out_uncache_write_outstanding_enable(csrCtrl_delay_io_out_uncache_write_outstanding_enable),
    .io_out_fusion_enable(csrCtrl_delay_io_out_fusion_enable),
    .io_out_wfi_enable(csrCtrl_delay_io_out_wfi_enable),
    .io_out_svinval_enable(csrCtrl_delay_io_out_svinval_enable),
    .io_out_distribute_csr_wvalid(csrCtrl_delay_io_out_distribute_csr_wvalid),
    .io_out_distribute_csr_waddr(csrCtrl_delay_io_out_distribute_csr_waddr),
    .io_out_distribute_csr_wdata(csrCtrl_delay_io_out_distribute_csr_wdata),
    .io_out_singlestep(csrCtrl_delay_io_out_singlestep),
    .io_out_frontend_trigger_t_valid(csrCtrl_delay_io_out_frontend_trigger_t_valid),
    .io_out_frontend_trigger_t_bits_addr(csrCtrl_delay_io_out_frontend_trigger_t_bits_addr),
    .io_out_frontend_trigger_t_bits_tdata_matchType(csrCtrl_delay_io_out_frontend_trigger_t_bits_tdata_matchType),
    .io_out_frontend_trigger_t_bits_tdata_select(csrCtrl_delay_io_out_frontend_trigger_t_bits_tdata_select),
    .io_out_frontend_trigger_t_bits_tdata_timing(csrCtrl_delay_io_out_frontend_trigger_t_bits_tdata_timing),
    .io_out_frontend_trigger_t_bits_tdata_chain(csrCtrl_delay_io_out_frontend_trigger_t_bits_tdata_chain),
    .io_out_frontend_trigger_t_bits_tdata_tdata2(csrCtrl_delay_io_out_frontend_trigger_t_bits_tdata_tdata2),
    .io_out_mem_trigger_t_valid(csrCtrl_delay_io_out_mem_trigger_t_valid),
    .io_out_mem_trigger_t_bits_addr(csrCtrl_delay_io_out_mem_trigger_t_bits_addr),
    .io_out_mem_trigger_t_bits_tdata_matchType(csrCtrl_delay_io_out_mem_trigger_t_bits_tdata_matchType),
    .io_out_mem_trigger_t_bits_tdata_select(csrCtrl_delay_io_out_mem_trigger_t_bits_tdata_select),
    .io_out_mem_trigger_t_bits_tdata_chain(csrCtrl_delay_io_out_mem_trigger_t_bits_tdata_chain),
    .io_out_mem_trigger_t_bits_tdata_tdata2(csrCtrl_delay_io_out_mem_trigger_t_bits_tdata_tdata2),
    .io_out_trigger_enable_0(csrCtrl_delay_io_out_trigger_enable_0),
    .io_out_trigger_enable_1(csrCtrl_delay_io_out_trigger_enable_1),
    .io_out_trigger_enable_2(csrCtrl_delay_io_out_trigger_enable_2),
    .io_out_trigger_enable_3(csrCtrl_delay_io_out_trigger_enable_3),
    .io_out_trigger_enable_4(csrCtrl_delay_io_out_trigger_enable_4),
    .io_out_trigger_enable_5(csrCtrl_delay_io_out_trigger_enable_5),
    .io_out_trigger_enable_6(csrCtrl_delay_io_out_trigger_enable_6),
    .io_out_trigger_enable_7(csrCtrl_delay_io_out_trigger_enable_7),
    .io_out_trigger_enable_8(csrCtrl_delay_io_out_trigger_enable_8),
    .io_out_trigger_enable_9(csrCtrl_delay_io_out_trigger_enable_9)
  );
  PMP pmp ( // @[Frontend.scala 87:19]
    .clock(pmp_clock),
    .reset(pmp_reset),
    .io_distribute_csr_wvalid(pmp_io_distribute_csr_wvalid),
    .io_distribute_csr_waddr(pmp_io_distribute_csr_waddr),
    .io_distribute_csr_wdata(pmp_io_distribute_csr_wdata),
    .io_pmp_0_cfg_l(pmp_io_pmp_0_cfg_l),
    .io_pmp_0_cfg_a(pmp_io_pmp_0_cfg_a),
    .io_pmp_0_cfg_x(pmp_io_pmp_0_cfg_x),
    .io_pmp_0_cfg_w(pmp_io_pmp_0_cfg_w),
    .io_pmp_0_cfg_r(pmp_io_pmp_0_cfg_r),
    .io_pmp_0_addr(pmp_io_pmp_0_addr),
    .io_pmp_0_mask(pmp_io_pmp_0_mask),
    .io_pmp_1_cfg_l(pmp_io_pmp_1_cfg_l),
    .io_pmp_1_cfg_a(pmp_io_pmp_1_cfg_a),
    .io_pmp_1_cfg_x(pmp_io_pmp_1_cfg_x),
    .io_pmp_1_cfg_w(pmp_io_pmp_1_cfg_w),
    .io_pmp_1_cfg_r(pmp_io_pmp_1_cfg_r),
    .io_pmp_1_addr(pmp_io_pmp_1_addr),
    .io_pmp_1_mask(pmp_io_pmp_1_mask),
    .io_pmp_2_cfg_l(pmp_io_pmp_2_cfg_l),
    .io_pmp_2_cfg_a(pmp_io_pmp_2_cfg_a),
    .io_pmp_2_cfg_x(pmp_io_pmp_2_cfg_x),
    .io_pmp_2_cfg_w(pmp_io_pmp_2_cfg_w),
    .io_pmp_2_cfg_r(pmp_io_pmp_2_cfg_r),
    .io_pmp_2_addr(pmp_io_pmp_2_addr),
    .io_pmp_2_mask(pmp_io_pmp_2_mask),
    .io_pmp_3_cfg_l(pmp_io_pmp_3_cfg_l),
    .io_pmp_3_cfg_a(pmp_io_pmp_3_cfg_a),
    .io_pmp_3_cfg_x(pmp_io_pmp_3_cfg_x),
    .io_pmp_3_cfg_w(pmp_io_pmp_3_cfg_w),
    .io_pmp_3_cfg_r(pmp_io_pmp_3_cfg_r),
    .io_pmp_3_addr(pmp_io_pmp_3_addr),
    .io_pmp_3_mask(pmp_io_pmp_3_mask),
    .io_pmp_4_cfg_l(pmp_io_pmp_4_cfg_l),
    .io_pmp_4_cfg_a(pmp_io_pmp_4_cfg_a),
    .io_pmp_4_cfg_x(pmp_io_pmp_4_cfg_x),
    .io_pmp_4_cfg_w(pmp_io_pmp_4_cfg_w),
    .io_pmp_4_cfg_r(pmp_io_pmp_4_cfg_r),
    .io_pmp_4_addr(pmp_io_pmp_4_addr),
    .io_pmp_4_mask(pmp_io_pmp_4_mask),
    .io_pmp_5_cfg_l(pmp_io_pmp_5_cfg_l),
    .io_pmp_5_cfg_a(pmp_io_pmp_5_cfg_a),
    .io_pmp_5_cfg_x(pmp_io_pmp_5_cfg_x),
    .io_pmp_5_cfg_w(pmp_io_pmp_5_cfg_w),
    .io_pmp_5_cfg_r(pmp_io_pmp_5_cfg_r),
    .io_pmp_5_addr(pmp_io_pmp_5_addr),
    .io_pmp_5_mask(pmp_io_pmp_5_mask),
    .io_pmp_6_cfg_l(pmp_io_pmp_6_cfg_l),
    .io_pmp_6_cfg_a(pmp_io_pmp_6_cfg_a),
    .io_pmp_6_cfg_x(pmp_io_pmp_6_cfg_x),
    .io_pmp_6_cfg_w(pmp_io_pmp_6_cfg_w),
    .io_pmp_6_cfg_r(pmp_io_pmp_6_cfg_r),
    .io_pmp_6_addr(pmp_io_pmp_6_addr),
    .io_pmp_6_mask(pmp_io_pmp_6_mask),
    .io_pmp_7_cfg_l(pmp_io_pmp_7_cfg_l),
    .io_pmp_7_cfg_a(pmp_io_pmp_7_cfg_a),
    .io_pmp_7_cfg_x(pmp_io_pmp_7_cfg_x),
    .io_pmp_7_cfg_w(pmp_io_pmp_7_cfg_w),
    .io_pmp_7_cfg_r(pmp_io_pmp_7_cfg_r),
    .io_pmp_7_addr(pmp_io_pmp_7_addr),
    .io_pmp_7_mask(pmp_io_pmp_7_mask),
    .io_pmp_8_cfg_l(pmp_io_pmp_8_cfg_l),
    .io_pmp_8_cfg_a(pmp_io_pmp_8_cfg_a),
    .io_pmp_8_cfg_x(pmp_io_pmp_8_cfg_x),
    .io_pmp_8_cfg_w(pmp_io_pmp_8_cfg_w),
    .io_pmp_8_cfg_r(pmp_io_pmp_8_cfg_r),
    .io_pmp_8_addr(pmp_io_pmp_8_addr),
    .io_pmp_8_mask(pmp_io_pmp_8_mask),
    .io_pmp_9_cfg_l(pmp_io_pmp_9_cfg_l),
    .io_pmp_9_cfg_a(pmp_io_pmp_9_cfg_a),
    .io_pmp_9_cfg_x(pmp_io_pmp_9_cfg_x),
    .io_pmp_9_cfg_w(pmp_io_pmp_9_cfg_w),
    .io_pmp_9_cfg_r(pmp_io_pmp_9_cfg_r),
    .io_pmp_9_addr(pmp_io_pmp_9_addr),
    .io_pmp_9_mask(pmp_io_pmp_9_mask),
    .io_pmp_10_cfg_l(pmp_io_pmp_10_cfg_l),
    .io_pmp_10_cfg_a(pmp_io_pmp_10_cfg_a),
    .io_pmp_10_cfg_x(pmp_io_pmp_10_cfg_x),
    .io_pmp_10_cfg_w(pmp_io_pmp_10_cfg_w),
    .io_pmp_10_cfg_r(pmp_io_pmp_10_cfg_r),
    .io_pmp_10_addr(pmp_io_pmp_10_addr),
    .io_pmp_10_mask(pmp_io_pmp_10_mask),
    .io_pmp_11_cfg_l(pmp_io_pmp_11_cfg_l),
    .io_pmp_11_cfg_a(pmp_io_pmp_11_cfg_a),
    .io_pmp_11_cfg_x(pmp_io_pmp_11_cfg_x),
    .io_pmp_11_cfg_w(pmp_io_pmp_11_cfg_w),
    .io_pmp_11_cfg_r(pmp_io_pmp_11_cfg_r),
    .io_pmp_11_addr(pmp_io_pmp_11_addr),
    .io_pmp_11_mask(pmp_io_pmp_11_mask),
    .io_pmp_12_cfg_l(pmp_io_pmp_12_cfg_l),
    .io_pmp_12_cfg_a(pmp_io_pmp_12_cfg_a),
    .io_pmp_12_cfg_x(pmp_io_pmp_12_cfg_x),
    .io_pmp_12_cfg_w(pmp_io_pmp_12_cfg_w),
    .io_pmp_12_cfg_r(pmp_io_pmp_12_cfg_r),
    .io_pmp_12_addr(pmp_io_pmp_12_addr),
    .io_pmp_12_mask(pmp_io_pmp_12_mask),
    .io_pmp_13_cfg_l(pmp_io_pmp_13_cfg_l),
    .io_pmp_13_cfg_a(pmp_io_pmp_13_cfg_a),
    .io_pmp_13_cfg_x(pmp_io_pmp_13_cfg_x),
    .io_pmp_13_cfg_w(pmp_io_pmp_13_cfg_w),
    .io_pmp_13_cfg_r(pmp_io_pmp_13_cfg_r),
    .io_pmp_13_addr(pmp_io_pmp_13_addr),
    .io_pmp_13_mask(pmp_io_pmp_13_mask),
    .io_pmp_14_cfg_l(pmp_io_pmp_14_cfg_l),
    .io_pmp_14_cfg_a(pmp_io_pmp_14_cfg_a),
    .io_pmp_14_cfg_x(pmp_io_pmp_14_cfg_x),
    .io_pmp_14_cfg_w(pmp_io_pmp_14_cfg_w),
    .io_pmp_14_cfg_r(pmp_io_pmp_14_cfg_r),
    .io_pmp_14_addr(pmp_io_pmp_14_addr),
    .io_pmp_14_mask(pmp_io_pmp_14_mask),
    .io_pmp_15_cfg_l(pmp_io_pmp_15_cfg_l),
    .io_pmp_15_cfg_a(pmp_io_pmp_15_cfg_a),
    .io_pmp_15_cfg_x(pmp_io_pmp_15_cfg_x),
    .io_pmp_15_cfg_w(pmp_io_pmp_15_cfg_w),
    .io_pmp_15_cfg_r(pmp_io_pmp_15_cfg_r),
    .io_pmp_15_addr(pmp_io_pmp_15_addr),
    .io_pmp_15_mask(pmp_io_pmp_15_mask),
    .io_pma_0_cfg_c(pmp_io_pma_0_cfg_c),
    .io_pma_0_cfg_atomic(pmp_io_pma_0_cfg_atomic),
    .io_pma_0_cfg_a(pmp_io_pma_0_cfg_a),
    .io_pma_0_cfg_x(pmp_io_pma_0_cfg_x),
    .io_pma_0_cfg_w(pmp_io_pma_0_cfg_w),
    .io_pma_0_cfg_r(pmp_io_pma_0_cfg_r),
    .io_pma_0_addr(pmp_io_pma_0_addr),
    .io_pma_0_mask(pmp_io_pma_0_mask),
    .io_pma_1_cfg_c(pmp_io_pma_1_cfg_c),
    .io_pma_1_cfg_atomic(pmp_io_pma_1_cfg_atomic),
    .io_pma_1_cfg_a(pmp_io_pma_1_cfg_a),
    .io_pma_1_cfg_x(pmp_io_pma_1_cfg_x),
    .io_pma_1_cfg_w(pmp_io_pma_1_cfg_w),
    .io_pma_1_cfg_r(pmp_io_pma_1_cfg_r),
    .io_pma_1_addr(pmp_io_pma_1_addr),
    .io_pma_1_mask(pmp_io_pma_1_mask),
    .io_pma_2_cfg_c(pmp_io_pma_2_cfg_c),
    .io_pma_2_cfg_atomic(pmp_io_pma_2_cfg_atomic),
    .io_pma_2_cfg_a(pmp_io_pma_2_cfg_a),
    .io_pma_2_cfg_x(pmp_io_pma_2_cfg_x),
    .io_pma_2_cfg_w(pmp_io_pma_2_cfg_w),
    .io_pma_2_cfg_r(pmp_io_pma_2_cfg_r),
    .io_pma_2_addr(pmp_io_pma_2_addr),
    .io_pma_2_mask(pmp_io_pma_2_mask),
    .io_pma_3_cfg_c(pmp_io_pma_3_cfg_c),
    .io_pma_3_cfg_atomic(pmp_io_pma_3_cfg_atomic),
    .io_pma_3_cfg_a(pmp_io_pma_3_cfg_a),
    .io_pma_3_cfg_x(pmp_io_pma_3_cfg_x),
    .io_pma_3_cfg_w(pmp_io_pma_3_cfg_w),
    .io_pma_3_cfg_r(pmp_io_pma_3_cfg_r),
    .io_pma_3_addr(pmp_io_pma_3_addr),
    .io_pma_3_mask(pmp_io_pma_3_mask),
    .io_pma_4_cfg_c(pmp_io_pma_4_cfg_c),
    .io_pma_4_cfg_atomic(pmp_io_pma_4_cfg_atomic),
    .io_pma_4_cfg_a(pmp_io_pma_4_cfg_a),
    .io_pma_4_cfg_x(pmp_io_pma_4_cfg_x),
    .io_pma_4_cfg_w(pmp_io_pma_4_cfg_w),
    .io_pma_4_cfg_r(pmp_io_pma_4_cfg_r),
    .io_pma_4_addr(pmp_io_pma_4_addr),
    .io_pma_4_mask(pmp_io_pma_4_mask),
    .io_pma_5_cfg_c(pmp_io_pma_5_cfg_c),
    .io_pma_5_cfg_atomic(pmp_io_pma_5_cfg_atomic),
    .io_pma_5_cfg_a(pmp_io_pma_5_cfg_a),
    .io_pma_5_cfg_x(pmp_io_pma_5_cfg_x),
    .io_pma_5_cfg_w(pmp_io_pma_5_cfg_w),
    .io_pma_5_cfg_r(pmp_io_pma_5_cfg_r),
    .io_pma_5_addr(pmp_io_pma_5_addr),
    .io_pma_5_mask(pmp_io_pma_5_mask),
    .io_pma_6_cfg_c(pmp_io_pma_6_cfg_c),
    .io_pma_6_cfg_atomic(pmp_io_pma_6_cfg_atomic),
    .io_pma_6_cfg_a(pmp_io_pma_6_cfg_a),
    .io_pma_6_cfg_x(pmp_io_pma_6_cfg_x),
    .io_pma_6_cfg_w(pmp_io_pma_6_cfg_w),
    .io_pma_6_cfg_r(pmp_io_pma_6_cfg_r),
    .io_pma_6_addr(pmp_io_pma_6_addr),
    .io_pma_6_mask(pmp_io_pma_6_mask),
    .io_pma_7_cfg_c(pmp_io_pma_7_cfg_c),
    .io_pma_7_cfg_atomic(pmp_io_pma_7_cfg_atomic),
    .io_pma_7_cfg_a(pmp_io_pma_7_cfg_a),
    .io_pma_7_cfg_x(pmp_io_pma_7_cfg_x),
    .io_pma_7_cfg_w(pmp_io_pma_7_cfg_w),
    .io_pma_7_cfg_r(pmp_io_pma_7_cfg_r),
    .io_pma_7_addr(pmp_io_pma_7_addr),
    .io_pma_7_mask(pmp_io_pma_7_mask),
    .io_pma_8_cfg_c(pmp_io_pma_8_cfg_c),
    .io_pma_8_cfg_atomic(pmp_io_pma_8_cfg_atomic),
    .io_pma_8_cfg_a(pmp_io_pma_8_cfg_a),
    .io_pma_8_cfg_x(pmp_io_pma_8_cfg_x),
    .io_pma_8_cfg_w(pmp_io_pma_8_cfg_w),
    .io_pma_8_cfg_r(pmp_io_pma_8_cfg_r),
    .io_pma_8_addr(pmp_io_pma_8_addr),
    .io_pma_8_mask(pmp_io_pma_8_mask),
    .io_pma_9_cfg_c(pmp_io_pma_9_cfg_c),
    .io_pma_9_cfg_atomic(pmp_io_pma_9_cfg_atomic),
    .io_pma_9_cfg_a(pmp_io_pma_9_cfg_a),
    .io_pma_9_cfg_x(pmp_io_pma_9_cfg_x),
    .io_pma_9_cfg_w(pmp_io_pma_9_cfg_w),
    .io_pma_9_cfg_r(pmp_io_pma_9_cfg_r),
    .io_pma_9_addr(pmp_io_pma_9_addr),
    .io_pma_9_mask(pmp_io_pma_9_mask),
    .io_pma_10_cfg_c(pmp_io_pma_10_cfg_c),
    .io_pma_10_cfg_atomic(pmp_io_pma_10_cfg_atomic),
    .io_pma_10_cfg_a(pmp_io_pma_10_cfg_a),
    .io_pma_10_cfg_x(pmp_io_pma_10_cfg_x),
    .io_pma_10_cfg_w(pmp_io_pma_10_cfg_w),
    .io_pma_10_cfg_r(pmp_io_pma_10_cfg_r),
    .io_pma_10_addr(pmp_io_pma_10_addr),
    .io_pma_10_mask(pmp_io_pma_10_mask),
    .io_pma_11_cfg_c(pmp_io_pma_11_cfg_c),
    .io_pma_11_cfg_atomic(pmp_io_pma_11_cfg_atomic),
    .io_pma_11_cfg_a(pmp_io_pma_11_cfg_a),
    .io_pma_11_cfg_x(pmp_io_pma_11_cfg_x),
    .io_pma_11_cfg_w(pmp_io_pma_11_cfg_w),
    .io_pma_11_cfg_r(pmp_io_pma_11_cfg_r),
    .io_pma_11_addr(pmp_io_pma_11_addr),
    .io_pma_11_mask(pmp_io_pma_11_mask),
    .io_pma_12_cfg_c(pmp_io_pma_12_cfg_c),
    .io_pma_12_cfg_atomic(pmp_io_pma_12_cfg_atomic),
    .io_pma_12_cfg_a(pmp_io_pma_12_cfg_a),
    .io_pma_12_cfg_x(pmp_io_pma_12_cfg_x),
    .io_pma_12_cfg_w(pmp_io_pma_12_cfg_w),
    .io_pma_12_cfg_r(pmp_io_pma_12_cfg_r),
    .io_pma_12_addr(pmp_io_pma_12_addr),
    .io_pma_12_mask(pmp_io_pma_12_mask),
    .io_pma_13_cfg_c(pmp_io_pma_13_cfg_c),
    .io_pma_13_cfg_atomic(pmp_io_pma_13_cfg_atomic),
    .io_pma_13_cfg_a(pmp_io_pma_13_cfg_a),
    .io_pma_13_cfg_x(pmp_io_pma_13_cfg_x),
    .io_pma_13_cfg_w(pmp_io_pma_13_cfg_w),
    .io_pma_13_cfg_r(pmp_io_pma_13_cfg_r),
    .io_pma_13_addr(pmp_io_pma_13_addr),
    .io_pma_13_mask(pmp_io_pma_13_mask),
    .io_pma_14_cfg_c(pmp_io_pma_14_cfg_c),
    .io_pma_14_cfg_atomic(pmp_io_pma_14_cfg_atomic),
    .io_pma_14_cfg_a(pmp_io_pma_14_cfg_a),
    .io_pma_14_cfg_x(pmp_io_pma_14_cfg_x),
    .io_pma_14_cfg_w(pmp_io_pma_14_cfg_w),
    .io_pma_14_cfg_r(pmp_io_pma_14_cfg_r),
    .io_pma_14_addr(pmp_io_pma_14_addr),
    .io_pma_14_mask(pmp_io_pma_14_mask),
    .io_pma_15_cfg_c(pmp_io_pma_15_cfg_c),
    .io_pma_15_cfg_atomic(pmp_io_pma_15_cfg_atomic),
    .io_pma_15_cfg_a(pmp_io_pma_15_cfg_a),
    .io_pma_15_cfg_x(pmp_io_pma_15_cfg_x),
    .io_pma_15_cfg_w(pmp_io_pma_15_cfg_w),
    .io_pma_15_cfg_r(pmp_io_pma_15_cfg_r),
    .io_pma_15_addr(pmp_io_pma_15_addr),
    .io_pma_15_mask(pmp_io_pma_15_mask)
  );
  PMPChecker PMPChecker ( // @[Frontend.scala 88:45]
    .io_check_env_mode(PMPChecker_io_check_env_mode),
    .io_check_env_pmp_0_cfg_l(PMPChecker_io_check_env_pmp_0_cfg_l),
    .io_check_env_pmp_0_cfg_a(PMPChecker_io_check_env_pmp_0_cfg_a),
    .io_check_env_pmp_0_cfg_x(PMPChecker_io_check_env_pmp_0_cfg_x),
    .io_check_env_pmp_0_cfg_w(PMPChecker_io_check_env_pmp_0_cfg_w),
    .io_check_env_pmp_0_cfg_r(PMPChecker_io_check_env_pmp_0_cfg_r),
    .io_check_env_pmp_0_addr(PMPChecker_io_check_env_pmp_0_addr),
    .io_check_env_pmp_0_mask(PMPChecker_io_check_env_pmp_0_mask),
    .io_check_env_pmp_1_cfg_l(PMPChecker_io_check_env_pmp_1_cfg_l),
    .io_check_env_pmp_1_cfg_a(PMPChecker_io_check_env_pmp_1_cfg_a),
    .io_check_env_pmp_1_cfg_x(PMPChecker_io_check_env_pmp_1_cfg_x),
    .io_check_env_pmp_1_cfg_w(PMPChecker_io_check_env_pmp_1_cfg_w),
    .io_check_env_pmp_1_cfg_r(PMPChecker_io_check_env_pmp_1_cfg_r),
    .io_check_env_pmp_1_addr(PMPChecker_io_check_env_pmp_1_addr),
    .io_check_env_pmp_1_mask(PMPChecker_io_check_env_pmp_1_mask),
    .io_check_env_pmp_2_cfg_l(PMPChecker_io_check_env_pmp_2_cfg_l),
    .io_check_env_pmp_2_cfg_a(PMPChecker_io_check_env_pmp_2_cfg_a),
    .io_check_env_pmp_2_cfg_x(PMPChecker_io_check_env_pmp_2_cfg_x),
    .io_check_env_pmp_2_cfg_w(PMPChecker_io_check_env_pmp_2_cfg_w),
    .io_check_env_pmp_2_cfg_r(PMPChecker_io_check_env_pmp_2_cfg_r),
    .io_check_env_pmp_2_addr(PMPChecker_io_check_env_pmp_2_addr),
    .io_check_env_pmp_2_mask(PMPChecker_io_check_env_pmp_2_mask),
    .io_check_env_pmp_3_cfg_l(PMPChecker_io_check_env_pmp_3_cfg_l),
    .io_check_env_pmp_3_cfg_a(PMPChecker_io_check_env_pmp_3_cfg_a),
    .io_check_env_pmp_3_cfg_x(PMPChecker_io_check_env_pmp_3_cfg_x),
    .io_check_env_pmp_3_cfg_w(PMPChecker_io_check_env_pmp_3_cfg_w),
    .io_check_env_pmp_3_cfg_r(PMPChecker_io_check_env_pmp_3_cfg_r),
    .io_check_env_pmp_3_addr(PMPChecker_io_check_env_pmp_3_addr),
    .io_check_env_pmp_3_mask(PMPChecker_io_check_env_pmp_3_mask),
    .io_check_env_pmp_4_cfg_l(PMPChecker_io_check_env_pmp_4_cfg_l),
    .io_check_env_pmp_4_cfg_a(PMPChecker_io_check_env_pmp_4_cfg_a),
    .io_check_env_pmp_4_cfg_x(PMPChecker_io_check_env_pmp_4_cfg_x),
    .io_check_env_pmp_4_cfg_w(PMPChecker_io_check_env_pmp_4_cfg_w),
    .io_check_env_pmp_4_cfg_r(PMPChecker_io_check_env_pmp_4_cfg_r),
    .io_check_env_pmp_4_addr(PMPChecker_io_check_env_pmp_4_addr),
    .io_check_env_pmp_4_mask(PMPChecker_io_check_env_pmp_4_mask),
    .io_check_env_pmp_5_cfg_l(PMPChecker_io_check_env_pmp_5_cfg_l),
    .io_check_env_pmp_5_cfg_a(PMPChecker_io_check_env_pmp_5_cfg_a),
    .io_check_env_pmp_5_cfg_x(PMPChecker_io_check_env_pmp_5_cfg_x),
    .io_check_env_pmp_5_cfg_w(PMPChecker_io_check_env_pmp_5_cfg_w),
    .io_check_env_pmp_5_cfg_r(PMPChecker_io_check_env_pmp_5_cfg_r),
    .io_check_env_pmp_5_addr(PMPChecker_io_check_env_pmp_5_addr),
    .io_check_env_pmp_5_mask(PMPChecker_io_check_env_pmp_5_mask),
    .io_check_env_pmp_6_cfg_l(PMPChecker_io_check_env_pmp_6_cfg_l),
    .io_check_env_pmp_6_cfg_a(PMPChecker_io_check_env_pmp_6_cfg_a),
    .io_check_env_pmp_6_cfg_x(PMPChecker_io_check_env_pmp_6_cfg_x),
    .io_check_env_pmp_6_cfg_w(PMPChecker_io_check_env_pmp_6_cfg_w),
    .io_check_env_pmp_6_cfg_r(PMPChecker_io_check_env_pmp_6_cfg_r),
    .io_check_env_pmp_6_addr(PMPChecker_io_check_env_pmp_6_addr),
    .io_check_env_pmp_6_mask(PMPChecker_io_check_env_pmp_6_mask),
    .io_check_env_pmp_7_cfg_l(PMPChecker_io_check_env_pmp_7_cfg_l),
    .io_check_env_pmp_7_cfg_a(PMPChecker_io_check_env_pmp_7_cfg_a),
    .io_check_env_pmp_7_cfg_x(PMPChecker_io_check_env_pmp_7_cfg_x),
    .io_check_env_pmp_7_cfg_w(PMPChecker_io_check_env_pmp_7_cfg_w),
    .io_check_env_pmp_7_cfg_r(PMPChecker_io_check_env_pmp_7_cfg_r),
    .io_check_env_pmp_7_addr(PMPChecker_io_check_env_pmp_7_addr),
    .io_check_env_pmp_7_mask(PMPChecker_io_check_env_pmp_7_mask),
    .io_check_env_pmp_8_cfg_l(PMPChecker_io_check_env_pmp_8_cfg_l),
    .io_check_env_pmp_8_cfg_a(PMPChecker_io_check_env_pmp_8_cfg_a),
    .io_check_env_pmp_8_cfg_x(PMPChecker_io_check_env_pmp_8_cfg_x),
    .io_check_env_pmp_8_cfg_w(PMPChecker_io_check_env_pmp_8_cfg_w),
    .io_check_env_pmp_8_cfg_r(PMPChecker_io_check_env_pmp_8_cfg_r),
    .io_check_env_pmp_8_addr(PMPChecker_io_check_env_pmp_8_addr),
    .io_check_env_pmp_8_mask(PMPChecker_io_check_env_pmp_8_mask),
    .io_check_env_pmp_9_cfg_l(PMPChecker_io_check_env_pmp_9_cfg_l),
    .io_check_env_pmp_9_cfg_a(PMPChecker_io_check_env_pmp_9_cfg_a),
    .io_check_env_pmp_9_cfg_x(PMPChecker_io_check_env_pmp_9_cfg_x),
    .io_check_env_pmp_9_cfg_w(PMPChecker_io_check_env_pmp_9_cfg_w),
    .io_check_env_pmp_9_cfg_r(PMPChecker_io_check_env_pmp_9_cfg_r),
    .io_check_env_pmp_9_addr(PMPChecker_io_check_env_pmp_9_addr),
    .io_check_env_pmp_9_mask(PMPChecker_io_check_env_pmp_9_mask),
    .io_check_env_pmp_10_cfg_l(PMPChecker_io_check_env_pmp_10_cfg_l),
    .io_check_env_pmp_10_cfg_a(PMPChecker_io_check_env_pmp_10_cfg_a),
    .io_check_env_pmp_10_cfg_x(PMPChecker_io_check_env_pmp_10_cfg_x),
    .io_check_env_pmp_10_cfg_w(PMPChecker_io_check_env_pmp_10_cfg_w),
    .io_check_env_pmp_10_cfg_r(PMPChecker_io_check_env_pmp_10_cfg_r),
    .io_check_env_pmp_10_addr(PMPChecker_io_check_env_pmp_10_addr),
    .io_check_env_pmp_10_mask(PMPChecker_io_check_env_pmp_10_mask),
    .io_check_env_pmp_11_cfg_l(PMPChecker_io_check_env_pmp_11_cfg_l),
    .io_check_env_pmp_11_cfg_a(PMPChecker_io_check_env_pmp_11_cfg_a),
    .io_check_env_pmp_11_cfg_x(PMPChecker_io_check_env_pmp_11_cfg_x),
    .io_check_env_pmp_11_cfg_w(PMPChecker_io_check_env_pmp_11_cfg_w),
    .io_check_env_pmp_11_cfg_r(PMPChecker_io_check_env_pmp_11_cfg_r),
    .io_check_env_pmp_11_addr(PMPChecker_io_check_env_pmp_11_addr),
    .io_check_env_pmp_11_mask(PMPChecker_io_check_env_pmp_11_mask),
    .io_check_env_pmp_12_cfg_l(PMPChecker_io_check_env_pmp_12_cfg_l),
    .io_check_env_pmp_12_cfg_a(PMPChecker_io_check_env_pmp_12_cfg_a),
    .io_check_env_pmp_12_cfg_x(PMPChecker_io_check_env_pmp_12_cfg_x),
    .io_check_env_pmp_12_cfg_w(PMPChecker_io_check_env_pmp_12_cfg_w),
    .io_check_env_pmp_12_cfg_r(PMPChecker_io_check_env_pmp_12_cfg_r),
    .io_check_env_pmp_12_addr(PMPChecker_io_check_env_pmp_12_addr),
    .io_check_env_pmp_12_mask(PMPChecker_io_check_env_pmp_12_mask),
    .io_check_env_pmp_13_cfg_l(PMPChecker_io_check_env_pmp_13_cfg_l),
    .io_check_env_pmp_13_cfg_a(PMPChecker_io_check_env_pmp_13_cfg_a),
    .io_check_env_pmp_13_cfg_x(PMPChecker_io_check_env_pmp_13_cfg_x),
    .io_check_env_pmp_13_cfg_w(PMPChecker_io_check_env_pmp_13_cfg_w),
    .io_check_env_pmp_13_cfg_r(PMPChecker_io_check_env_pmp_13_cfg_r),
    .io_check_env_pmp_13_addr(PMPChecker_io_check_env_pmp_13_addr),
    .io_check_env_pmp_13_mask(PMPChecker_io_check_env_pmp_13_mask),
    .io_check_env_pmp_14_cfg_l(PMPChecker_io_check_env_pmp_14_cfg_l),
    .io_check_env_pmp_14_cfg_a(PMPChecker_io_check_env_pmp_14_cfg_a),
    .io_check_env_pmp_14_cfg_x(PMPChecker_io_check_env_pmp_14_cfg_x),
    .io_check_env_pmp_14_cfg_w(PMPChecker_io_check_env_pmp_14_cfg_w),
    .io_check_env_pmp_14_cfg_r(PMPChecker_io_check_env_pmp_14_cfg_r),
    .io_check_env_pmp_14_addr(PMPChecker_io_check_env_pmp_14_addr),
    .io_check_env_pmp_14_mask(PMPChecker_io_check_env_pmp_14_mask),
    .io_check_env_pmp_15_cfg_l(PMPChecker_io_check_env_pmp_15_cfg_l),
    .io_check_env_pmp_15_cfg_a(PMPChecker_io_check_env_pmp_15_cfg_a),
    .io_check_env_pmp_15_cfg_x(PMPChecker_io_check_env_pmp_15_cfg_x),
    .io_check_env_pmp_15_cfg_w(PMPChecker_io_check_env_pmp_15_cfg_w),
    .io_check_env_pmp_15_cfg_r(PMPChecker_io_check_env_pmp_15_cfg_r),
    .io_check_env_pmp_15_addr(PMPChecker_io_check_env_pmp_15_addr),
    .io_check_env_pmp_15_mask(PMPChecker_io_check_env_pmp_15_mask),
    .io_check_env_pma_0_cfg_c(PMPChecker_io_check_env_pma_0_cfg_c),
    .io_check_env_pma_0_cfg_atomic(PMPChecker_io_check_env_pma_0_cfg_atomic),
    .io_check_env_pma_0_cfg_a(PMPChecker_io_check_env_pma_0_cfg_a),
    .io_check_env_pma_0_cfg_x(PMPChecker_io_check_env_pma_0_cfg_x),
    .io_check_env_pma_0_cfg_w(PMPChecker_io_check_env_pma_0_cfg_w),
    .io_check_env_pma_0_cfg_r(PMPChecker_io_check_env_pma_0_cfg_r),
    .io_check_env_pma_0_addr(PMPChecker_io_check_env_pma_0_addr),
    .io_check_env_pma_0_mask(PMPChecker_io_check_env_pma_0_mask),
    .io_check_env_pma_1_cfg_c(PMPChecker_io_check_env_pma_1_cfg_c),
    .io_check_env_pma_1_cfg_atomic(PMPChecker_io_check_env_pma_1_cfg_atomic),
    .io_check_env_pma_1_cfg_a(PMPChecker_io_check_env_pma_1_cfg_a),
    .io_check_env_pma_1_cfg_x(PMPChecker_io_check_env_pma_1_cfg_x),
    .io_check_env_pma_1_cfg_w(PMPChecker_io_check_env_pma_1_cfg_w),
    .io_check_env_pma_1_cfg_r(PMPChecker_io_check_env_pma_1_cfg_r),
    .io_check_env_pma_1_addr(PMPChecker_io_check_env_pma_1_addr),
    .io_check_env_pma_1_mask(PMPChecker_io_check_env_pma_1_mask),
    .io_check_env_pma_2_cfg_c(PMPChecker_io_check_env_pma_2_cfg_c),
    .io_check_env_pma_2_cfg_atomic(PMPChecker_io_check_env_pma_2_cfg_atomic),
    .io_check_env_pma_2_cfg_a(PMPChecker_io_check_env_pma_2_cfg_a),
    .io_check_env_pma_2_cfg_x(PMPChecker_io_check_env_pma_2_cfg_x),
    .io_check_env_pma_2_cfg_w(PMPChecker_io_check_env_pma_2_cfg_w),
    .io_check_env_pma_2_cfg_r(PMPChecker_io_check_env_pma_2_cfg_r),
    .io_check_env_pma_2_addr(PMPChecker_io_check_env_pma_2_addr),
    .io_check_env_pma_2_mask(PMPChecker_io_check_env_pma_2_mask),
    .io_check_env_pma_3_cfg_c(PMPChecker_io_check_env_pma_3_cfg_c),
    .io_check_env_pma_3_cfg_atomic(PMPChecker_io_check_env_pma_3_cfg_atomic),
    .io_check_env_pma_3_cfg_a(PMPChecker_io_check_env_pma_3_cfg_a),
    .io_check_env_pma_3_cfg_x(PMPChecker_io_check_env_pma_3_cfg_x),
    .io_check_env_pma_3_cfg_w(PMPChecker_io_check_env_pma_3_cfg_w),
    .io_check_env_pma_3_cfg_r(PMPChecker_io_check_env_pma_3_cfg_r),
    .io_check_env_pma_3_addr(PMPChecker_io_check_env_pma_3_addr),
    .io_check_env_pma_3_mask(PMPChecker_io_check_env_pma_3_mask),
    .io_check_env_pma_4_cfg_c(PMPChecker_io_check_env_pma_4_cfg_c),
    .io_check_env_pma_4_cfg_atomic(PMPChecker_io_check_env_pma_4_cfg_atomic),
    .io_check_env_pma_4_cfg_a(PMPChecker_io_check_env_pma_4_cfg_a),
    .io_check_env_pma_4_cfg_x(PMPChecker_io_check_env_pma_4_cfg_x),
    .io_check_env_pma_4_cfg_w(PMPChecker_io_check_env_pma_4_cfg_w),
    .io_check_env_pma_4_cfg_r(PMPChecker_io_check_env_pma_4_cfg_r),
    .io_check_env_pma_4_addr(PMPChecker_io_check_env_pma_4_addr),
    .io_check_env_pma_4_mask(PMPChecker_io_check_env_pma_4_mask),
    .io_check_env_pma_5_cfg_c(PMPChecker_io_check_env_pma_5_cfg_c),
    .io_check_env_pma_5_cfg_atomic(PMPChecker_io_check_env_pma_5_cfg_atomic),
    .io_check_env_pma_5_cfg_a(PMPChecker_io_check_env_pma_5_cfg_a),
    .io_check_env_pma_5_cfg_x(PMPChecker_io_check_env_pma_5_cfg_x),
    .io_check_env_pma_5_cfg_w(PMPChecker_io_check_env_pma_5_cfg_w),
    .io_check_env_pma_5_cfg_r(PMPChecker_io_check_env_pma_5_cfg_r),
    .io_check_env_pma_5_addr(PMPChecker_io_check_env_pma_5_addr),
    .io_check_env_pma_5_mask(PMPChecker_io_check_env_pma_5_mask),
    .io_check_env_pma_6_cfg_c(PMPChecker_io_check_env_pma_6_cfg_c),
    .io_check_env_pma_6_cfg_atomic(PMPChecker_io_check_env_pma_6_cfg_atomic),
    .io_check_env_pma_6_cfg_a(PMPChecker_io_check_env_pma_6_cfg_a),
    .io_check_env_pma_6_cfg_x(PMPChecker_io_check_env_pma_6_cfg_x),
    .io_check_env_pma_6_cfg_w(PMPChecker_io_check_env_pma_6_cfg_w),
    .io_check_env_pma_6_cfg_r(PMPChecker_io_check_env_pma_6_cfg_r),
    .io_check_env_pma_6_addr(PMPChecker_io_check_env_pma_6_addr),
    .io_check_env_pma_6_mask(PMPChecker_io_check_env_pma_6_mask),
    .io_check_env_pma_7_cfg_c(PMPChecker_io_check_env_pma_7_cfg_c),
    .io_check_env_pma_7_cfg_atomic(PMPChecker_io_check_env_pma_7_cfg_atomic),
    .io_check_env_pma_7_cfg_a(PMPChecker_io_check_env_pma_7_cfg_a),
    .io_check_env_pma_7_cfg_x(PMPChecker_io_check_env_pma_7_cfg_x),
    .io_check_env_pma_7_cfg_w(PMPChecker_io_check_env_pma_7_cfg_w),
    .io_check_env_pma_7_cfg_r(PMPChecker_io_check_env_pma_7_cfg_r),
    .io_check_env_pma_7_addr(PMPChecker_io_check_env_pma_7_addr),
    .io_check_env_pma_7_mask(PMPChecker_io_check_env_pma_7_mask),
    .io_check_env_pma_8_cfg_c(PMPChecker_io_check_env_pma_8_cfg_c),
    .io_check_env_pma_8_cfg_atomic(PMPChecker_io_check_env_pma_8_cfg_atomic),
    .io_check_env_pma_8_cfg_a(PMPChecker_io_check_env_pma_8_cfg_a),
    .io_check_env_pma_8_cfg_x(PMPChecker_io_check_env_pma_8_cfg_x),
    .io_check_env_pma_8_cfg_w(PMPChecker_io_check_env_pma_8_cfg_w),
    .io_check_env_pma_8_cfg_r(PMPChecker_io_check_env_pma_8_cfg_r),
    .io_check_env_pma_8_addr(PMPChecker_io_check_env_pma_8_addr),
    .io_check_env_pma_8_mask(PMPChecker_io_check_env_pma_8_mask),
    .io_check_env_pma_9_cfg_c(PMPChecker_io_check_env_pma_9_cfg_c),
    .io_check_env_pma_9_cfg_atomic(PMPChecker_io_check_env_pma_9_cfg_atomic),
    .io_check_env_pma_9_cfg_a(PMPChecker_io_check_env_pma_9_cfg_a),
    .io_check_env_pma_9_cfg_x(PMPChecker_io_check_env_pma_9_cfg_x),
    .io_check_env_pma_9_cfg_w(PMPChecker_io_check_env_pma_9_cfg_w),
    .io_check_env_pma_9_cfg_r(PMPChecker_io_check_env_pma_9_cfg_r),
    .io_check_env_pma_9_addr(PMPChecker_io_check_env_pma_9_addr),
    .io_check_env_pma_9_mask(PMPChecker_io_check_env_pma_9_mask),
    .io_check_env_pma_10_cfg_c(PMPChecker_io_check_env_pma_10_cfg_c),
    .io_check_env_pma_10_cfg_atomic(PMPChecker_io_check_env_pma_10_cfg_atomic),
    .io_check_env_pma_10_cfg_a(PMPChecker_io_check_env_pma_10_cfg_a),
    .io_check_env_pma_10_cfg_x(PMPChecker_io_check_env_pma_10_cfg_x),
    .io_check_env_pma_10_cfg_w(PMPChecker_io_check_env_pma_10_cfg_w),
    .io_check_env_pma_10_cfg_r(PMPChecker_io_check_env_pma_10_cfg_r),
    .io_check_env_pma_10_addr(PMPChecker_io_check_env_pma_10_addr),
    .io_check_env_pma_10_mask(PMPChecker_io_check_env_pma_10_mask),
    .io_check_env_pma_11_cfg_c(PMPChecker_io_check_env_pma_11_cfg_c),
    .io_check_env_pma_11_cfg_atomic(PMPChecker_io_check_env_pma_11_cfg_atomic),
    .io_check_env_pma_11_cfg_a(PMPChecker_io_check_env_pma_11_cfg_a),
    .io_check_env_pma_11_cfg_x(PMPChecker_io_check_env_pma_11_cfg_x),
    .io_check_env_pma_11_cfg_w(PMPChecker_io_check_env_pma_11_cfg_w),
    .io_check_env_pma_11_cfg_r(PMPChecker_io_check_env_pma_11_cfg_r),
    .io_check_env_pma_11_addr(PMPChecker_io_check_env_pma_11_addr),
    .io_check_env_pma_11_mask(PMPChecker_io_check_env_pma_11_mask),
    .io_check_env_pma_12_cfg_c(PMPChecker_io_check_env_pma_12_cfg_c),
    .io_check_env_pma_12_cfg_atomic(PMPChecker_io_check_env_pma_12_cfg_atomic),
    .io_check_env_pma_12_cfg_a(PMPChecker_io_check_env_pma_12_cfg_a),
    .io_check_env_pma_12_cfg_x(PMPChecker_io_check_env_pma_12_cfg_x),
    .io_check_env_pma_12_cfg_w(PMPChecker_io_check_env_pma_12_cfg_w),
    .io_check_env_pma_12_cfg_r(PMPChecker_io_check_env_pma_12_cfg_r),
    .io_check_env_pma_12_addr(PMPChecker_io_check_env_pma_12_addr),
    .io_check_env_pma_12_mask(PMPChecker_io_check_env_pma_12_mask),
    .io_check_env_pma_13_cfg_c(PMPChecker_io_check_env_pma_13_cfg_c),
    .io_check_env_pma_13_cfg_atomic(PMPChecker_io_check_env_pma_13_cfg_atomic),
    .io_check_env_pma_13_cfg_a(PMPChecker_io_check_env_pma_13_cfg_a),
    .io_check_env_pma_13_cfg_x(PMPChecker_io_check_env_pma_13_cfg_x),
    .io_check_env_pma_13_cfg_w(PMPChecker_io_check_env_pma_13_cfg_w),
    .io_check_env_pma_13_cfg_r(PMPChecker_io_check_env_pma_13_cfg_r),
    .io_check_env_pma_13_addr(PMPChecker_io_check_env_pma_13_addr),
    .io_check_env_pma_13_mask(PMPChecker_io_check_env_pma_13_mask),
    .io_check_env_pma_14_cfg_c(PMPChecker_io_check_env_pma_14_cfg_c),
    .io_check_env_pma_14_cfg_atomic(PMPChecker_io_check_env_pma_14_cfg_atomic),
    .io_check_env_pma_14_cfg_a(PMPChecker_io_check_env_pma_14_cfg_a),
    .io_check_env_pma_14_cfg_x(PMPChecker_io_check_env_pma_14_cfg_x),
    .io_check_env_pma_14_cfg_w(PMPChecker_io_check_env_pma_14_cfg_w),
    .io_check_env_pma_14_cfg_r(PMPChecker_io_check_env_pma_14_cfg_r),
    .io_check_env_pma_14_addr(PMPChecker_io_check_env_pma_14_addr),
    .io_check_env_pma_14_mask(PMPChecker_io_check_env_pma_14_mask),
    .io_check_env_pma_15_cfg_c(PMPChecker_io_check_env_pma_15_cfg_c),
    .io_check_env_pma_15_cfg_atomic(PMPChecker_io_check_env_pma_15_cfg_atomic),
    .io_check_env_pma_15_cfg_a(PMPChecker_io_check_env_pma_15_cfg_a),
    .io_check_env_pma_15_cfg_x(PMPChecker_io_check_env_pma_15_cfg_x),
    .io_check_env_pma_15_cfg_w(PMPChecker_io_check_env_pma_15_cfg_w),
    .io_check_env_pma_15_cfg_r(PMPChecker_io_check_env_pma_15_cfg_r),
    .io_check_env_pma_15_addr(PMPChecker_io_check_env_pma_15_addr),
    .io_check_env_pma_15_mask(PMPChecker_io_check_env_pma_15_mask),
    .io_req_bits_addr(PMPChecker_io_req_bits_addr),
    .io_req_bits_cmd(PMPChecker_io_req_bits_cmd),
    .io_resp_ld(PMPChecker_io_resp_ld),
    .io_resp_st(PMPChecker_io_resp_st),
    .io_resp_instr(PMPChecker_io_resp_instr),
    .io_resp_mmio(PMPChecker_io_resp_mmio),
    .io_resp_atomic(PMPChecker_io_resp_atomic)
  );
  PMPChecker PMPChecker_1 ( // @[Frontend.scala 88:45]
    .io_check_env_mode(PMPChecker_1_io_check_env_mode),
    .io_check_env_pmp_0_cfg_l(PMPChecker_1_io_check_env_pmp_0_cfg_l),
    .io_check_env_pmp_0_cfg_a(PMPChecker_1_io_check_env_pmp_0_cfg_a),
    .io_check_env_pmp_0_cfg_x(PMPChecker_1_io_check_env_pmp_0_cfg_x),
    .io_check_env_pmp_0_cfg_w(PMPChecker_1_io_check_env_pmp_0_cfg_w),
    .io_check_env_pmp_0_cfg_r(PMPChecker_1_io_check_env_pmp_0_cfg_r),
    .io_check_env_pmp_0_addr(PMPChecker_1_io_check_env_pmp_0_addr),
    .io_check_env_pmp_0_mask(PMPChecker_1_io_check_env_pmp_0_mask),
    .io_check_env_pmp_1_cfg_l(PMPChecker_1_io_check_env_pmp_1_cfg_l),
    .io_check_env_pmp_1_cfg_a(PMPChecker_1_io_check_env_pmp_1_cfg_a),
    .io_check_env_pmp_1_cfg_x(PMPChecker_1_io_check_env_pmp_1_cfg_x),
    .io_check_env_pmp_1_cfg_w(PMPChecker_1_io_check_env_pmp_1_cfg_w),
    .io_check_env_pmp_1_cfg_r(PMPChecker_1_io_check_env_pmp_1_cfg_r),
    .io_check_env_pmp_1_addr(PMPChecker_1_io_check_env_pmp_1_addr),
    .io_check_env_pmp_1_mask(PMPChecker_1_io_check_env_pmp_1_mask),
    .io_check_env_pmp_2_cfg_l(PMPChecker_1_io_check_env_pmp_2_cfg_l),
    .io_check_env_pmp_2_cfg_a(PMPChecker_1_io_check_env_pmp_2_cfg_a),
    .io_check_env_pmp_2_cfg_x(PMPChecker_1_io_check_env_pmp_2_cfg_x),
    .io_check_env_pmp_2_cfg_w(PMPChecker_1_io_check_env_pmp_2_cfg_w),
    .io_check_env_pmp_2_cfg_r(PMPChecker_1_io_check_env_pmp_2_cfg_r),
    .io_check_env_pmp_2_addr(PMPChecker_1_io_check_env_pmp_2_addr),
    .io_check_env_pmp_2_mask(PMPChecker_1_io_check_env_pmp_2_mask),
    .io_check_env_pmp_3_cfg_l(PMPChecker_1_io_check_env_pmp_3_cfg_l),
    .io_check_env_pmp_3_cfg_a(PMPChecker_1_io_check_env_pmp_3_cfg_a),
    .io_check_env_pmp_3_cfg_x(PMPChecker_1_io_check_env_pmp_3_cfg_x),
    .io_check_env_pmp_3_cfg_w(PMPChecker_1_io_check_env_pmp_3_cfg_w),
    .io_check_env_pmp_3_cfg_r(PMPChecker_1_io_check_env_pmp_3_cfg_r),
    .io_check_env_pmp_3_addr(PMPChecker_1_io_check_env_pmp_3_addr),
    .io_check_env_pmp_3_mask(PMPChecker_1_io_check_env_pmp_3_mask),
    .io_check_env_pmp_4_cfg_l(PMPChecker_1_io_check_env_pmp_4_cfg_l),
    .io_check_env_pmp_4_cfg_a(PMPChecker_1_io_check_env_pmp_4_cfg_a),
    .io_check_env_pmp_4_cfg_x(PMPChecker_1_io_check_env_pmp_4_cfg_x),
    .io_check_env_pmp_4_cfg_w(PMPChecker_1_io_check_env_pmp_4_cfg_w),
    .io_check_env_pmp_4_cfg_r(PMPChecker_1_io_check_env_pmp_4_cfg_r),
    .io_check_env_pmp_4_addr(PMPChecker_1_io_check_env_pmp_4_addr),
    .io_check_env_pmp_4_mask(PMPChecker_1_io_check_env_pmp_4_mask),
    .io_check_env_pmp_5_cfg_l(PMPChecker_1_io_check_env_pmp_5_cfg_l),
    .io_check_env_pmp_5_cfg_a(PMPChecker_1_io_check_env_pmp_5_cfg_a),
    .io_check_env_pmp_5_cfg_x(PMPChecker_1_io_check_env_pmp_5_cfg_x),
    .io_check_env_pmp_5_cfg_w(PMPChecker_1_io_check_env_pmp_5_cfg_w),
    .io_check_env_pmp_5_cfg_r(PMPChecker_1_io_check_env_pmp_5_cfg_r),
    .io_check_env_pmp_5_addr(PMPChecker_1_io_check_env_pmp_5_addr),
    .io_check_env_pmp_5_mask(PMPChecker_1_io_check_env_pmp_5_mask),
    .io_check_env_pmp_6_cfg_l(PMPChecker_1_io_check_env_pmp_6_cfg_l),
    .io_check_env_pmp_6_cfg_a(PMPChecker_1_io_check_env_pmp_6_cfg_a),
    .io_check_env_pmp_6_cfg_x(PMPChecker_1_io_check_env_pmp_6_cfg_x),
    .io_check_env_pmp_6_cfg_w(PMPChecker_1_io_check_env_pmp_6_cfg_w),
    .io_check_env_pmp_6_cfg_r(PMPChecker_1_io_check_env_pmp_6_cfg_r),
    .io_check_env_pmp_6_addr(PMPChecker_1_io_check_env_pmp_6_addr),
    .io_check_env_pmp_6_mask(PMPChecker_1_io_check_env_pmp_6_mask),
    .io_check_env_pmp_7_cfg_l(PMPChecker_1_io_check_env_pmp_7_cfg_l),
    .io_check_env_pmp_7_cfg_a(PMPChecker_1_io_check_env_pmp_7_cfg_a),
    .io_check_env_pmp_7_cfg_x(PMPChecker_1_io_check_env_pmp_7_cfg_x),
    .io_check_env_pmp_7_cfg_w(PMPChecker_1_io_check_env_pmp_7_cfg_w),
    .io_check_env_pmp_7_cfg_r(PMPChecker_1_io_check_env_pmp_7_cfg_r),
    .io_check_env_pmp_7_addr(PMPChecker_1_io_check_env_pmp_7_addr),
    .io_check_env_pmp_7_mask(PMPChecker_1_io_check_env_pmp_7_mask),
    .io_check_env_pmp_8_cfg_l(PMPChecker_1_io_check_env_pmp_8_cfg_l),
    .io_check_env_pmp_8_cfg_a(PMPChecker_1_io_check_env_pmp_8_cfg_a),
    .io_check_env_pmp_8_cfg_x(PMPChecker_1_io_check_env_pmp_8_cfg_x),
    .io_check_env_pmp_8_cfg_w(PMPChecker_1_io_check_env_pmp_8_cfg_w),
    .io_check_env_pmp_8_cfg_r(PMPChecker_1_io_check_env_pmp_8_cfg_r),
    .io_check_env_pmp_8_addr(PMPChecker_1_io_check_env_pmp_8_addr),
    .io_check_env_pmp_8_mask(PMPChecker_1_io_check_env_pmp_8_mask),
    .io_check_env_pmp_9_cfg_l(PMPChecker_1_io_check_env_pmp_9_cfg_l),
    .io_check_env_pmp_9_cfg_a(PMPChecker_1_io_check_env_pmp_9_cfg_a),
    .io_check_env_pmp_9_cfg_x(PMPChecker_1_io_check_env_pmp_9_cfg_x),
    .io_check_env_pmp_9_cfg_w(PMPChecker_1_io_check_env_pmp_9_cfg_w),
    .io_check_env_pmp_9_cfg_r(PMPChecker_1_io_check_env_pmp_9_cfg_r),
    .io_check_env_pmp_9_addr(PMPChecker_1_io_check_env_pmp_9_addr),
    .io_check_env_pmp_9_mask(PMPChecker_1_io_check_env_pmp_9_mask),
    .io_check_env_pmp_10_cfg_l(PMPChecker_1_io_check_env_pmp_10_cfg_l),
    .io_check_env_pmp_10_cfg_a(PMPChecker_1_io_check_env_pmp_10_cfg_a),
    .io_check_env_pmp_10_cfg_x(PMPChecker_1_io_check_env_pmp_10_cfg_x),
    .io_check_env_pmp_10_cfg_w(PMPChecker_1_io_check_env_pmp_10_cfg_w),
    .io_check_env_pmp_10_cfg_r(PMPChecker_1_io_check_env_pmp_10_cfg_r),
    .io_check_env_pmp_10_addr(PMPChecker_1_io_check_env_pmp_10_addr),
    .io_check_env_pmp_10_mask(PMPChecker_1_io_check_env_pmp_10_mask),
    .io_check_env_pmp_11_cfg_l(PMPChecker_1_io_check_env_pmp_11_cfg_l),
    .io_check_env_pmp_11_cfg_a(PMPChecker_1_io_check_env_pmp_11_cfg_a),
    .io_check_env_pmp_11_cfg_x(PMPChecker_1_io_check_env_pmp_11_cfg_x),
    .io_check_env_pmp_11_cfg_w(PMPChecker_1_io_check_env_pmp_11_cfg_w),
    .io_check_env_pmp_11_cfg_r(PMPChecker_1_io_check_env_pmp_11_cfg_r),
    .io_check_env_pmp_11_addr(PMPChecker_1_io_check_env_pmp_11_addr),
    .io_check_env_pmp_11_mask(PMPChecker_1_io_check_env_pmp_11_mask),
    .io_check_env_pmp_12_cfg_l(PMPChecker_1_io_check_env_pmp_12_cfg_l),
    .io_check_env_pmp_12_cfg_a(PMPChecker_1_io_check_env_pmp_12_cfg_a),
    .io_check_env_pmp_12_cfg_x(PMPChecker_1_io_check_env_pmp_12_cfg_x),
    .io_check_env_pmp_12_cfg_w(PMPChecker_1_io_check_env_pmp_12_cfg_w),
    .io_check_env_pmp_12_cfg_r(PMPChecker_1_io_check_env_pmp_12_cfg_r),
    .io_check_env_pmp_12_addr(PMPChecker_1_io_check_env_pmp_12_addr),
    .io_check_env_pmp_12_mask(PMPChecker_1_io_check_env_pmp_12_mask),
    .io_check_env_pmp_13_cfg_l(PMPChecker_1_io_check_env_pmp_13_cfg_l),
    .io_check_env_pmp_13_cfg_a(PMPChecker_1_io_check_env_pmp_13_cfg_a),
    .io_check_env_pmp_13_cfg_x(PMPChecker_1_io_check_env_pmp_13_cfg_x),
    .io_check_env_pmp_13_cfg_w(PMPChecker_1_io_check_env_pmp_13_cfg_w),
    .io_check_env_pmp_13_cfg_r(PMPChecker_1_io_check_env_pmp_13_cfg_r),
    .io_check_env_pmp_13_addr(PMPChecker_1_io_check_env_pmp_13_addr),
    .io_check_env_pmp_13_mask(PMPChecker_1_io_check_env_pmp_13_mask),
    .io_check_env_pmp_14_cfg_l(PMPChecker_1_io_check_env_pmp_14_cfg_l),
    .io_check_env_pmp_14_cfg_a(PMPChecker_1_io_check_env_pmp_14_cfg_a),
    .io_check_env_pmp_14_cfg_x(PMPChecker_1_io_check_env_pmp_14_cfg_x),
    .io_check_env_pmp_14_cfg_w(PMPChecker_1_io_check_env_pmp_14_cfg_w),
    .io_check_env_pmp_14_cfg_r(PMPChecker_1_io_check_env_pmp_14_cfg_r),
    .io_check_env_pmp_14_addr(PMPChecker_1_io_check_env_pmp_14_addr),
    .io_check_env_pmp_14_mask(PMPChecker_1_io_check_env_pmp_14_mask),
    .io_check_env_pmp_15_cfg_l(PMPChecker_1_io_check_env_pmp_15_cfg_l),
    .io_check_env_pmp_15_cfg_a(PMPChecker_1_io_check_env_pmp_15_cfg_a),
    .io_check_env_pmp_15_cfg_x(PMPChecker_1_io_check_env_pmp_15_cfg_x),
    .io_check_env_pmp_15_cfg_w(PMPChecker_1_io_check_env_pmp_15_cfg_w),
    .io_check_env_pmp_15_cfg_r(PMPChecker_1_io_check_env_pmp_15_cfg_r),
    .io_check_env_pmp_15_addr(PMPChecker_1_io_check_env_pmp_15_addr),
    .io_check_env_pmp_15_mask(PMPChecker_1_io_check_env_pmp_15_mask),
    .io_check_env_pma_0_cfg_c(PMPChecker_1_io_check_env_pma_0_cfg_c),
    .io_check_env_pma_0_cfg_atomic(PMPChecker_1_io_check_env_pma_0_cfg_atomic),
    .io_check_env_pma_0_cfg_a(PMPChecker_1_io_check_env_pma_0_cfg_a),
    .io_check_env_pma_0_cfg_x(PMPChecker_1_io_check_env_pma_0_cfg_x),
    .io_check_env_pma_0_cfg_w(PMPChecker_1_io_check_env_pma_0_cfg_w),
    .io_check_env_pma_0_cfg_r(PMPChecker_1_io_check_env_pma_0_cfg_r),
    .io_check_env_pma_0_addr(PMPChecker_1_io_check_env_pma_0_addr),
    .io_check_env_pma_0_mask(PMPChecker_1_io_check_env_pma_0_mask),
    .io_check_env_pma_1_cfg_c(PMPChecker_1_io_check_env_pma_1_cfg_c),
    .io_check_env_pma_1_cfg_atomic(PMPChecker_1_io_check_env_pma_1_cfg_atomic),
    .io_check_env_pma_1_cfg_a(PMPChecker_1_io_check_env_pma_1_cfg_a),
    .io_check_env_pma_1_cfg_x(PMPChecker_1_io_check_env_pma_1_cfg_x),
    .io_check_env_pma_1_cfg_w(PMPChecker_1_io_check_env_pma_1_cfg_w),
    .io_check_env_pma_1_cfg_r(PMPChecker_1_io_check_env_pma_1_cfg_r),
    .io_check_env_pma_1_addr(PMPChecker_1_io_check_env_pma_1_addr),
    .io_check_env_pma_1_mask(PMPChecker_1_io_check_env_pma_1_mask),
    .io_check_env_pma_2_cfg_c(PMPChecker_1_io_check_env_pma_2_cfg_c),
    .io_check_env_pma_2_cfg_atomic(PMPChecker_1_io_check_env_pma_2_cfg_atomic),
    .io_check_env_pma_2_cfg_a(PMPChecker_1_io_check_env_pma_2_cfg_a),
    .io_check_env_pma_2_cfg_x(PMPChecker_1_io_check_env_pma_2_cfg_x),
    .io_check_env_pma_2_cfg_w(PMPChecker_1_io_check_env_pma_2_cfg_w),
    .io_check_env_pma_2_cfg_r(PMPChecker_1_io_check_env_pma_2_cfg_r),
    .io_check_env_pma_2_addr(PMPChecker_1_io_check_env_pma_2_addr),
    .io_check_env_pma_2_mask(PMPChecker_1_io_check_env_pma_2_mask),
    .io_check_env_pma_3_cfg_c(PMPChecker_1_io_check_env_pma_3_cfg_c),
    .io_check_env_pma_3_cfg_atomic(PMPChecker_1_io_check_env_pma_3_cfg_atomic),
    .io_check_env_pma_3_cfg_a(PMPChecker_1_io_check_env_pma_3_cfg_a),
    .io_check_env_pma_3_cfg_x(PMPChecker_1_io_check_env_pma_3_cfg_x),
    .io_check_env_pma_3_cfg_w(PMPChecker_1_io_check_env_pma_3_cfg_w),
    .io_check_env_pma_3_cfg_r(PMPChecker_1_io_check_env_pma_3_cfg_r),
    .io_check_env_pma_3_addr(PMPChecker_1_io_check_env_pma_3_addr),
    .io_check_env_pma_3_mask(PMPChecker_1_io_check_env_pma_3_mask),
    .io_check_env_pma_4_cfg_c(PMPChecker_1_io_check_env_pma_4_cfg_c),
    .io_check_env_pma_4_cfg_atomic(PMPChecker_1_io_check_env_pma_4_cfg_atomic),
    .io_check_env_pma_4_cfg_a(PMPChecker_1_io_check_env_pma_4_cfg_a),
    .io_check_env_pma_4_cfg_x(PMPChecker_1_io_check_env_pma_4_cfg_x),
    .io_check_env_pma_4_cfg_w(PMPChecker_1_io_check_env_pma_4_cfg_w),
    .io_check_env_pma_4_cfg_r(PMPChecker_1_io_check_env_pma_4_cfg_r),
    .io_check_env_pma_4_addr(PMPChecker_1_io_check_env_pma_4_addr),
    .io_check_env_pma_4_mask(PMPChecker_1_io_check_env_pma_4_mask),
    .io_check_env_pma_5_cfg_c(PMPChecker_1_io_check_env_pma_5_cfg_c),
    .io_check_env_pma_5_cfg_atomic(PMPChecker_1_io_check_env_pma_5_cfg_atomic),
    .io_check_env_pma_5_cfg_a(PMPChecker_1_io_check_env_pma_5_cfg_a),
    .io_check_env_pma_5_cfg_x(PMPChecker_1_io_check_env_pma_5_cfg_x),
    .io_check_env_pma_5_cfg_w(PMPChecker_1_io_check_env_pma_5_cfg_w),
    .io_check_env_pma_5_cfg_r(PMPChecker_1_io_check_env_pma_5_cfg_r),
    .io_check_env_pma_5_addr(PMPChecker_1_io_check_env_pma_5_addr),
    .io_check_env_pma_5_mask(PMPChecker_1_io_check_env_pma_5_mask),
    .io_check_env_pma_6_cfg_c(PMPChecker_1_io_check_env_pma_6_cfg_c),
    .io_check_env_pma_6_cfg_atomic(PMPChecker_1_io_check_env_pma_6_cfg_atomic),
    .io_check_env_pma_6_cfg_a(PMPChecker_1_io_check_env_pma_6_cfg_a),
    .io_check_env_pma_6_cfg_x(PMPChecker_1_io_check_env_pma_6_cfg_x),
    .io_check_env_pma_6_cfg_w(PMPChecker_1_io_check_env_pma_6_cfg_w),
    .io_check_env_pma_6_cfg_r(PMPChecker_1_io_check_env_pma_6_cfg_r),
    .io_check_env_pma_6_addr(PMPChecker_1_io_check_env_pma_6_addr),
    .io_check_env_pma_6_mask(PMPChecker_1_io_check_env_pma_6_mask),
    .io_check_env_pma_7_cfg_c(PMPChecker_1_io_check_env_pma_7_cfg_c),
    .io_check_env_pma_7_cfg_atomic(PMPChecker_1_io_check_env_pma_7_cfg_atomic),
    .io_check_env_pma_7_cfg_a(PMPChecker_1_io_check_env_pma_7_cfg_a),
    .io_check_env_pma_7_cfg_x(PMPChecker_1_io_check_env_pma_7_cfg_x),
    .io_check_env_pma_7_cfg_w(PMPChecker_1_io_check_env_pma_7_cfg_w),
    .io_check_env_pma_7_cfg_r(PMPChecker_1_io_check_env_pma_7_cfg_r),
    .io_check_env_pma_7_addr(PMPChecker_1_io_check_env_pma_7_addr),
    .io_check_env_pma_7_mask(PMPChecker_1_io_check_env_pma_7_mask),
    .io_check_env_pma_8_cfg_c(PMPChecker_1_io_check_env_pma_8_cfg_c),
    .io_check_env_pma_8_cfg_atomic(PMPChecker_1_io_check_env_pma_8_cfg_atomic),
    .io_check_env_pma_8_cfg_a(PMPChecker_1_io_check_env_pma_8_cfg_a),
    .io_check_env_pma_8_cfg_x(PMPChecker_1_io_check_env_pma_8_cfg_x),
    .io_check_env_pma_8_cfg_w(PMPChecker_1_io_check_env_pma_8_cfg_w),
    .io_check_env_pma_8_cfg_r(PMPChecker_1_io_check_env_pma_8_cfg_r),
    .io_check_env_pma_8_addr(PMPChecker_1_io_check_env_pma_8_addr),
    .io_check_env_pma_8_mask(PMPChecker_1_io_check_env_pma_8_mask),
    .io_check_env_pma_9_cfg_c(PMPChecker_1_io_check_env_pma_9_cfg_c),
    .io_check_env_pma_9_cfg_atomic(PMPChecker_1_io_check_env_pma_9_cfg_atomic),
    .io_check_env_pma_9_cfg_a(PMPChecker_1_io_check_env_pma_9_cfg_a),
    .io_check_env_pma_9_cfg_x(PMPChecker_1_io_check_env_pma_9_cfg_x),
    .io_check_env_pma_9_cfg_w(PMPChecker_1_io_check_env_pma_9_cfg_w),
    .io_check_env_pma_9_cfg_r(PMPChecker_1_io_check_env_pma_9_cfg_r),
    .io_check_env_pma_9_addr(PMPChecker_1_io_check_env_pma_9_addr),
    .io_check_env_pma_9_mask(PMPChecker_1_io_check_env_pma_9_mask),
    .io_check_env_pma_10_cfg_c(PMPChecker_1_io_check_env_pma_10_cfg_c),
    .io_check_env_pma_10_cfg_atomic(PMPChecker_1_io_check_env_pma_10_cfg_atomic),
    .io_check_env_pma_10_cfg_a(PMPChecker_1_io_check_env_pma_10_cfg_a),
    .io_check_env_pma_10_cfg_x(PMPChecker_1_io_check_env_pma_10_cfg_x),
    .io_check_env_pma_10_cfg_w(PMPChecker_1_io_check_env_pma_10_cfg_w),
    .io_check_env_pma_10_cfg_r(PMPChecker_1_io_check_env_pma_10_cfg_r),
    .io_check_env_pma_10_addr(PMPChecker_1_io_check_env_pma_10_addr),
    .io_check_env_pma_10_mask(PMPChecker_1_io_check_env_pma_10_mask),
    .io_check_env_pma_11_cfg_c(PMPChecker_1_io_check_env_pma_11_cfg_c),
    .io_check_env_pma_11_cfg_atomic(PMPChecker_1_io_check_env_pma_11_cfg_atomic),
    .io_check_env_pma_11_cfg_a(PMPChecker_1_io_check_env_pma_11_cfg_a),
    .io_check_env_pma_11_cfg_x(PMPChecker_1_io_check_env_pma_11_cfg_x),
    .io_check_env_pma_11_cfg_w(PMPChecker_1_io_check_env_pma_11_cfg_w),
    .io_check_env_pma_11_cfg_r(PMPChecker_1_io_check_env_pma_11_cfg_r),
    .io_check_env_pma_11_addr(PMPChecker_1_io_check_env_pma_11_addr),
    .io_check_env_pma_11_mask(PMPChecker_1_io_check_env_pma_11_mask),
    .io_check_env_pma_12_cfg_c(PMPChecker_1_io_check_env_pma_12_cfg_c),
    .io_check_env_pma_12_cfg_atomic(PMPChecker_1_io_check_env_pma_12_cfg_atomic),
    .io_check_env_pma_12_cfg_a(PMPChecker_1_io_check_env_pma_12_cfg_a),
    .io_check_env_pma_12_cfg_x(PMPChecker_1_io_check_env_pma_12_cfg_x),
    .io_check_env_pma_12_cfg_w(PMPChecker_1_io_check_env_pma_12_cfg_w),
    .io_check_env_pma_12_cfg_r(PMPChecker_1_io_check_env_pma_12_cfg_r),
    .io_check_env_pma_12_addr(PMPChecker_1_io_check_env_pma_12_addr),
    .io_check_env_pma_12_mask(PMPChecker_1_io_check_env_pma_12_mask),
    .io_check_env_pma_13_cfg_c(PMPChecker_1_io_check_env_pma_13_cfg_c),
    .io_check_env_pma_13_cfg_atomic(PMPChecker_1_io_check_env_pma_13_cfg_atomic),
    .io_check_env_pma_13_cfg_a(PMPChecker_1_io_check_env_pma_13_cfg_a),
    .io_check_env_pma_13_cfg_x(PMPChecker_1_io_check_env_pma_13_cfg_x),
    .io_check_env_pma_13_cfg_w(PMPChecker_1_io_check_env_pma_13_cfg_w),
    .io_check_env_pma_13_cfg_r(PMPChecker_1_io_check_env_pma_13_cfg_r),
    .io_check_env_pma_13_addr(PMPChecker_1_io_check_env_pma_13_addr),
    .io_check_env_pma_13_mask(PMPChecker_1_io_check_env_pma_13_mask),
    .io_check_env_pma_14_cfg_c(PMPChecker_1_io_check_env_pma_14_cfg_c),
    .io_check_env_pma_14_cfg_atomic(PMPChecker_1_io_check_env_pma_14_cfg_atomic),
    .io_check_env_pma_14_cfg_a(PMPChecker_1_io_check_env_pma_14_cfg_a),
    .io_check_env_pma_14_cfg_x(PMPChecker_1_io_check_env_pma_14_cfg_x),
    .io_check_env_pma_14_cfg_w(PMPChecker_1_io_check_env_pma_14_cfg_w),
    .io_check_env_pma_14_cfg_r(PMPChecker_1_io_check_env_pma_14_cfg_r),
    .io_check_env_pma_14_addr(PMPChecker_1_io_check_env_pma_14_addr),
    .io_check_env_pma_14_mask(PMPChecker_1_io_check_env_pma_14_mask),
    .io_check_env_pma_15_cfg_c(PMPChecker_1_io_check_env_pma_15_cfg_c),
    .io_check_env_pma_15_cfg_atomic(PMPChecker_1_io_check_env_pma_15_cfg_atomic),
    .io_check_env_pma_15_cfg_a(PMPChecker_1_io_check_env_pma_15_cfg_a),
    .io_check_env_pma_15_cfg_x(PMPChecker_1_io_check_env_pma_15_cfg_x),
    .io_check_env_pma_15_cfg_w(PMPChecker_1_io_check_env_pma_15_cfg_w),
    .io_check_env_pma_15_cfg_r(PMPChecker_1_io_check_env_pma_15_cfg_r),
    .io_check_env_pma_15_addr(PMPChecker_1_io_check_env_pma_15_addr),
    .io_check_env_pma_15_mask(PMPChecker_1_io_check_env_pma_15_mask),
    .io_req_bits_addr(PMPChecker_1_io_req_bits_addr),
    .io_req_bits_cmd(PMPChecker_1_io_req_bits_cmd),
    .io_resp_ld(PMPChecker_1_io_resp_ld),
    .io_resp_st(PMPChecker_1_io_resp_st),
    .io_resp_instr(PMPChecker_1_io_resp_instr),
    .io_resp_mmio(PMPChecker_1_io_resp_mmio),
    .io_resp_atomic(PMPChecker_1_io_resp_atomic)
  );
  PMPChecker PMPChecker_2 ( // @[Frontend.scala 88:45]
    .io_check_env_mode(PMPChecker_2_io_check_env_mode),
    .io_check_env_pmp_0_cfg_l(PMPChecker_2_io_check_env_pmp_0_cfg_l),
    .io_check_env_pmp_0_cfg_a(PMPChecker_2_io_check_env_pmp_0_cfg_a),
    .io_check_env_pmp_0_cfg_x(PMPChecker_2_io_check_env_pmp_0_cfg_x),
    .io_check_env_pmp_0_cfg_w(PMPChecker_2_io_check_env_pmp_0_cfg_w),
    .io_check_env_pmp_0_cfg_r(PMPChecker_2_io_check_env_pmp_0_cfg_r),
    .io_check_env_pmp_0_addr(PMPChecker_2_io_check_env_pmp_0_addr),
    .io_check_env_pmp_0_mask(PMPChecker_2_io_check_env_pmp_0_mask),
    .io_check_env_pmp_1_cfg_l(PMPChecker_2_io_check_env_pmp_1_cfg_l),
    .io_check_env_pmp_1_cfg_a(PMPChecker_2_io_check_env_pmp_1_cfg_a),
    .io_check_env_pmp_1_cfg_x(PMPChecker_2_io_check_env_pmp_1_cfg_x),
    .io_check_env_pmp_1_cfg_w(PMPChecker_2_io_check_env_pmp_1_cfg_w),
    .io_check_env_pmp_1_cfg_r(PMPChecker_2_io_check_env_pmp_1_cfg_r),
    .io_check_env_pmp_1_addr(PMPChecker_2_io_check_env_pmp_1_addr),
    .io_check_env_pmp_1_mask(PMPChecker_2_io_check_env_pmp_1_mask),
    .io_check_env_pmp_2_cfg_l(PMPChecker_2_io_check_env_pmp_2_cfg_l),
    .io_check_env_pmp_2_cfg_a(PMPChecker_2_io_check_env_pmp_2_cfg_a),
    .io_check_env_pmp_2_cfg_x(PMPChecker_2_io_check_env_pmp_2_cfg_x),
    .io_check_env_pmp_2_cfg_w(PMPChecker_2_io_check_env_pmp_2_cfg_w),
    .io_check_env_pmp_2_cfg_r(PMPChecker_2_io_check_env_pmp_2_cfg_r),
    .io_check_env_pmp_2_addr(PMPChecker_2_io_check_env_pmp_2_addr),
    .io_check_env_pmp_2_mask(PMPChecker_2_io_check_env_pmp_2_mask),
    .io_check_env_pmp_3_cfg_l(PMPChecker_2_io_check_env_pmp_3_cfg_l),
    .io_check_env_pmp_3_cfg_a(PMPChecker_2_io_check_env_pmp_3_cfg_a),
    .io_check_env_pmp_3_cfg_x(PMPChecker_2_io_check_env_pmp_3_cfg_x),
    .io_check_env_pmp_3_cfg_w(PMPChecker_2_io_check_env_pmp_3_cfg_w),
    .io_check_env_pmp_3_cfg_r(PMPChecker_2_io_check_env_pmp_3_cfg_r),
    .io_check_env_pmp_3_addr(PMPChecker_2_io_check_env_pmp_3_addr),
    .io_check_env_pmp_3_mask(PMPChecker_2_io_check_env_pmp_3_mask),
    .io_check_env_pmp_4_cfg_l(PMPChecker_2_io_check_env_pmp_4_cfg_l),
    .io_check_env_pmp_4_cfg_a(PMPChecker_2_io_check_env_pmp_4_cfg_a),
    .io_check_env_pmp_4_cfg_x(PMPChecker_2_io_check_env_pmp_4_cfg_x),
    .io_check_env_pmp_4_cfg_w(PMPChecker_2_io_check_env_pmp_4_cfg_w),
    .io_check_env_pmp_4_cfg_r(PMPChecker_2_io_check_env_pmp_4_cfg_r),
    .io_check_env_pmp_4_addr(PMPChecker_2_io_check_env_pmp_4_addr),
    .io_check_env_pmp_4_mask(PMPChecker_2_io_check_env_pmp_4_mask),
    .io_check_env_pmp_5_cfg_l(PMPChecker_2_io_check_env_pmp_5_cfg_l),
    .io_check_env_pmp_5_cfg_a(PMPChecker_2_io_check_env_pmp_5_cfg_a),
    .io_check_env_pmp_5_cfg_x(PMPChecker_2_io_check_env_pmp_5_cfg_x),
    .io_check_env_pmp_5_cfg_w(PMPChecker_2_io_check_env_pmp_5_cfg_w),
    .io_check_env_pmp_5_cfg_r(PMPChecker_2_io_check_env_pmp_5_cfg_r),
    .io_check_env_pmp_5_addr(PMPChecker_2_io_check_env_pmp_5_addr),
    .io_check_env_pmp_5_mask(PMPChecker_2_io_check_env_pmp_5_mask),
    .io_check_env_pmp_6_cfg_l(PMPChecker_2_io_check_env_pmp_6_cfg_l),
    .io_check_env_pmp_6_cfg_a(PMPChecker_2_io_check_env_pmp_6_cfg_a),
    .io_check_env_pmp_6_cfg_x(PMPChecker_2_io_check_env_pmp_6_cfg_x),
    .io_check_env_pmp_6_cfg_w(PMPChecker_2_io_check_env_pmp_6_cfg_w),
    .io_check_env_pmp_6_cfg_r(PMPChecker_2_io_check_env_pmp_6_cfg_r),
    .io_check_env_pmp_6_addr(PMPChecker_2_io_check_env_pmp_6_addr),
    .io_check_env_pmp_6_mask(PMPChecker_2_io_check_env_pmp_6_mask),
    .io_check_env_pmp_7_cfg_l(PMPChecker_2_io_check_env_pmp_7_cfg_l),
    .io_check_env_pmp_7_cfg_a(PMPChecker_2_io_check_env_pmp_7_cfg_a),
    .io_check_env_pmp_7_cfg_x(PMPChecker_2_io_check_env_pmp_7_cfg_x),
    .io_check_env_pmp_7_cfg_w(PMPChecker_2_io_check_env_pmp_7_cfg_w),
    .io_check_env_pmp_7_cfg_r(PMPChecker_2_io_check_env_pmp_7_cfg_r),
    .io_check_env_pmp_7_addr(PMPChecker_2_io_check_env_pmp_7_addr),
    .io_check_env_pmp_7_mask(PMPChecker_2_io_check_env_pmp_7_mask),
    .io_check_env_pmp_8_cfg_l(PMPChecker_2_io_check_env_pmp_8_cfg_l),
    .io_check_env_pmp_8_cfg_a(PMPChecker_2_io_check_env_pmp_8_cfg_a),
    .io_check_env_pmp_8_cfg_x(PMPChecker_2_io_check_env_pmp_8_cfg_x),
    .io_check_env_pmp_8_cfg_w(PMPChecker_2_io_check_env_pmp_8_cfg_w),
    .io_check_env_pmp_8_cfg_r(PMPChecker_2_io_check_env_pmp_8_cfg_r),
    .io_check_env_pmp_8_addr(PMPChecker_2_io_check_env_pmp_8_addr),
    .io_check_env_pmp_8_mask(PMPChecker_2_io_check_env_pmp_8_mask),
    .io_check_env_pmp_9_cfg_l(PMPChecker_2_io_check_env_pmp_9_cfg_l),
    .io_check_env_pmp_9_cfg_a(PMPChecker_2_io_check_env_pmp_9_cfg_a),
    .io_check_env_pmp_9_cfg_x(PMPChecker_2_io_check_env_pmp_9_cfg_x),
    .io_check_env_pmp_9_cfg_w(PMPChecker_2_io_check_env_pmp_9_cfg_w),
    .io_check_env_pmp_9_cfg_r(PMPChecker_2_io_check_env_pmp_9_cfg_r),
    .io_check_env_pmp_9_addr(PMPChecker_2_io_check_env_pmp_9_addr),
    .io_check_env_pmp_9_mask(PMPChecker_2_io_check_env_pmp_9_mask),
    .io_check_env_pmp_10_cfg_l(PMPChecker_2_io_check_env_pmp_10_cfg_l),
    .io_check_env_pmp_10_cfg_a(PMPChecker_2_io_check_env_pmp_10_cfg_a),
    .io_check_env_pmp_10_cfg_x(PMPChecker_2_io_check_env_pmp_10_cfg_x),
    .io_check_env_pmp_10_cfg_w(PMPChecker_2_io_check_env_pmp_10_cfg_w),
    .io_check_env_pmp_10_cfg_r(PMPChecker_2_io_check_env_pmp_10_cfg_r),
    .io_check_env_pmp_10_addr(PMPChecker_2_io_check_env_pmp_10_addr),
    .io_check_env_pmp_10_mask(PMPChecker_2_io_check_env_pmp_10_mask),
    .io_check_env_pmp_11_cfg_l(PMPChecker_2_io_check_env_pmp_11_cfg_l),
    .io_check_env_pmp_11_cfg_a(PMPChecker_2_io_check_env_pmp_11_cfg_a),
    .io_check_env_pmp_11_cfg_x(PMPChecker_2_io_check_env_pmp_11_cfg_x),
    .io_check_env_pmp_11_cfg_w(PMPChecker_2_io_check_env_pmp_11_cfg_w),
    .io_check_env_pmp_11_cfg_r(PMPChecker_2_io_check_env_pmp_11_cfg_r),
    .io_check_env_pmp_11_addr(PMPChecker_2_io_check_env_pmp_11_addr),
    .io_check_env_pmp_11_mask(PMPChecker_2_io_check_env_pmp_11_mask),
    .io_check_env_pmp_12_cfg_l(PMPChecker_2_io_check_env_pmp_12_cfg_l),
    .io_check_env_pmp_12_cfg_a(PMPChecker_2_io_check_env_pmp_12_cfg_a),
    .io_check_env_pmp_12_cfg_x(PMPChecker_2_io_check_env_pmp_12_cfg_x),
    .io_check_env_pmp_12_cfg_w(PMPChecker_2_io_check_env_pmp_12_cfg_w),
    .io_check_env_pmp_12_cfg_r(PMPChecker_2_io_check_env_pmp_12_cfg_r),
    .io_check_env_pmp_12_addr(PMPChecker_2_io_check_env_pmp_12_addr),
    .io_check_env_pmp_12_mask(PMPChecker_2_io_check_env_pmp_12_mask),
    .io_check_env_pmp_13_cfg_l(PMPChecker_2_io_check_env_pmp_13_cfg_l),
    .io_check_env_pmp_13_cfg_a(PMPChecker_2_io_check_env_pmp_13_cfg_a),
    .io_check_env_pmp_13_cfg_x(PMPChecker_2_io_check_env_pmp_13_cfg_x),
    .io_check_env_pmp_13_cfg_w(PMPChecker_2_io_check_env_pmp_13_cfg_w),
    .io_check_env_pmp_13_cfg_r(PMPChecker_2_io_check_env_pmp_13_cfg_r),
    .io_check_env_pmp_13_addr(PMPChecker_2_io_check_env_pmp_13_addr),
    .io_check_env_pmp_13_mask(PMPChecker_2_io_check_env_pmp_13_mask),
    .io_check_env_pmp_14_cfg_l(PMPChecker_2_io_check_env_pmp_14_cfg_l),
    .io_check_env_pmp_14_cfg_a(PMPChecker_2_io_check_env_pmp_14_cfg_a),
    .io_check_env_pmp_14_cfg_x(PMPChecker_2_io_check_env_pmp_14_cfg_x),
    .io_check_env_pmp_14_cfg_w(PMPChecker_2_io_check_env_pmp_14_cfg_w),
    .io_check_env_pmp_14_cfg_r(PMPChecker_2_io_check_env_pmp_14_cfg_r),
    .io_check_env_pmp_14_addr(PMPChecker_2_io_check_env_pmp_14_addr),
    .io_check_env_pmp_14_mask(PMPChecker_2_io_check_env_pmp_14_mask),
    .io_check_env_pmp_15_cfg_l(PMPChecker_2_io_check_env_pmp_15_cfg_l),
    .io_check_env_pmp_15_cfg_a(PMPChecker_2_io_check_env_pmp_15_cfg_a),
    .io_check_env_pmp_15_cfg_x(PMPChecker_2_io_check_env_pmp_15_cfg_x),
    .io_check_env_pmp_15_cfg_w(PMPChecker_2_io_check_env_pmp_15_cfg_w),
    .io_check_env_pmp_15_cfg_r(PMPChecker_2_io_check_env_pmp_15_cfg_r),
    .io_check_env_pmp_15_addr(PMPChecker_2_io_check_env_pmp_15_addr),
    .io_check_env_pmp_15_mask(PMPChecker_2_io_check_env_pmp_15_mask),
    .io_check_env_pma_0_cfg_c(PMPChecker_2_io_check_env_pma_0_cfg_c),
    .io_check_env_pma_0_cfg_atomic(PMPChecker_2_io_check_env_pma_0_cfg_atomic),
    .io_check_env_pma_0_cfg_a(PMPChecker_2_io_check_env_pma_0_cfg_a),
    .io_check_env_pma_0_cfg_x(PMPChecker_2_io_check_env_pma_0_cfg_x),
    .io_check_env_pma_0_cfg_w(PMPChecker_2_io_check_env_pma_0_cfg_w),
    .io_check_env_pma_0_cfg_r(PMPChecker_2_io_check_env_pma_0_cfg_r),
    .io_check_env_pma_0_addr(PMPChecker_2_io_check_env_pma_0_addr),
    .io_check_env_pma_0_mask(PMPChecker_2_io_check_env_pma_0_mask),
    .io_check_env_pma_1_cfg_c(PMPChecker_2_io_check_env_pma_1_cfg_c),
    .io_check_env_pma_1_cfg_atomic(PMPChecker_2_io_check_env_pma_1_cfg_atomic),
    .io_check_env_pma_1_cfg_a(PMPChecker_2_io_check_env_pma_1_cfg_a),
    .io_check_env_pma_1_cfg_x(PMPChecker_2_io_check_env_pma_1_cfg_x),
    .io_check_env_pma_1_cfg_w(PMPChecker_2_io_check_env_pma_1_cfg_w),
    .io_check_env_pma_1_cfg_r(PMPChecker_2_io_check_env_pma_1_cfg_r),
    .io_check_env_pma_1_addr(PMPChecker_2_io_check_env_pma_1_addr),
    .io_check_env_pma_1_mask(PMPChecker_2_io_check_env_pma_1_mask),
    .io_check_env_pma_2_cfg_c(PMPChecker_2_io_check_env_pma_2_cfg_c),
    .io_check_env_pma_2_cfg_atomic(PMPChecker_2_io_check_env_pma_2_cfg_atomic),
    .io_check_env_pma_2_cfg_a(PMPChecker_2_io_check_env_pma_2_cfg_a),
    .io_check_env_pma_2_cfg_x(PMPChecker_2_io_check_env_pma_2_cfg_x),
    .io_check_env_pma_2_cfg_w(PMPChecker_2_io_check_env_pma_2_cfg_w),
    .io_check_env_pma_2_cfg_r(PMPChecker_2_io_check_env_pma_2_cfg_r),
    .io_check_env_pma_2_addr(PMPChecker_2_io_check_env_pma_2_addr),
    .io_check_env_pma_2_mask(PMPChecker_2_io_check_env_pma_2_mask),
    .io_check_env_pma_3_cfg_c(PMPChecker_2_io_check_env_pma_3_cfg_c),
    .io_check_env_pma_3_cfg_atomic(PMPChecker_2_io_check_env_pma_3_cfg_atomic),
    .io_check_env_pma_3_cfg_a(PMPChecker_2_io_check_env_pma_3_cfg_a),
    .io_check_env_pma_3_cfg_x(PMPChecker_2_io_check_env_pma_3_cfg_x),
    .io_check_env_pma_3_cfg_w(PMPChecker_2_io_check_env_pma_3_cfg_w),
    .io_check_env_pma_3_cfg_r(PMPChecker_2_io_check_env_pma_3_cfg_r),
    .io_check_env_pma_3_addr(PMPChecker_2_io_check_env_pma_3_addr),
    .io_check_env_pma_3_mask(PMPChecker_2_io_check_env_pma_3_mask),
    .io_check_env_pma_4_cfg_c(PMPChecker_2_io_check_env_pma_4_cfg_c),
    .io_check_env_pma_4_cfg_atomic(PMPChecker_2_io_check_env_pma_4_cfg_atomic),
    .io_check_env_pma_4_cfg_a(PMPChecker_2_io_check_env_pma_4_cfg_a),
    .io_check_env_pma_4_cfg_x(PMPChecker_2_io_check_env_pma_4_cfg_x),
    .io_check_env_pma_4_cfg_w(PMPChecker_2_io_check_env_pma_4_cfg_w),
    .io_check_env_pma_4_cfg_r(PMPChecker_2_io_check_env_pma_4_cfg_r),
    .io_check_env_pma_4_addr(PMPChecker_2_io_check_env_pma_4_addr),
    .io_check_env_pma_4_mask(PMPChecker_2_io_check_env_pma_4_mask),
    .io_check_env_pma_5_cfg_c(PMPChecker_2_io_check_env_pma_5_cfg_c),
    .io_check_env_pma_5_cfg_atomic(PMPChecker_2_io_check_env_pma_5_cfg_atomic),
    .io_check_env_pma_5_cfg_a(PMPChecker_2_io_check_env_pma_5_cfg_a),
    .io_check_env_pma_5_cfg_x(PMPChecker_2_io_check_env_pma_5_cfg_x),
    .io_check_env_pma_5_cfg_w(PMPChecker_2_io_check_env_pma_5_cfg_w),
    .io_check_env_pma_5_cfg_r(PMPChecker_2_io_check_env_pma_5_cfg_r),
    .io_check_env_pma_5_addr(PMPChecker_2_io_check_env_pma_5_addr),
    .io_check_env_pma_5_mask(PMPChecker_2_io_check_env_pma_5_mask),
    .io_check_env_pma_6_cfg_c(PMPChecker_2_io_check_env_pma_6_cfg_c),
    .io_check_env_pma_6_cfg_atomic(PMPChecker_2_io_check_env_pma_6_cfg_atomic),
    .io_check_env_pma_6_cfg_a(PMPChecker_2_io_check_env_pma_6_cfg_a),
    .io_check_env_pma_6_cfg_x(PMPChecker_2_io_check_env_pma_6_cfg_x),
    .io_check_env_pma_6_cfg_w(PMPChecker_2_io_check_env_pma_6_cfg_w),
    .io_check_env_pma_6_cfg_r(PMPChecker_2_io_check_env_pma_6_cfg_r),
    .io_check_env_pma_6_addr(PMPChecker_2_io_check_env_pma_6_addr),
    .io_check_env_pma_6_mask(PMPChecker_2_io_check_env_pma_6_mask),
    .io_check_env_pma_7_cfg_c(PMPChecker_2_io_check_env_pma_7_cfg_c),
    .io_check_env_pma_7_cfg_atomic(PMPChecker_2_io_check_env_pma_7_cfg_atomic),
    .io_check_env_pma_7_cfg_a(PMPChecker_2_io_check_env_pma_7_cfg_a),
    .io_check_env_pma_7_cfg_x(PMPChecker_2_io_check_env_pma_7_cfg_x),
    .io_check_env_pma_7_cfg_w(PMPChecker_2_io_check_env_pma_7_cfg_w),
    .io_check_env_pma_7_cfg_r(PMPChecker_2_io_check_env_pma_7_cfg_r),
    .io_check_env_pma_7_addr(PMPChecker_2_io_check_env_pma_7_addr),
    .io_check_env_pma_7_mask(PMPChecker_2_io_check_env_pma_7_mask),
    .io_check_env_pma_8_cfg_c(PMPChecker_2_io_check_env_pma_8_cfg_c),
    .io_check_env_pma_8_cfg_atomic(PMPChecker_2_io_check_env_pma_8_cfg_atomic),
    .io_check_env_pma_8_cfg_a(PMPChecker_2_io_check_env_pma_8_cfg_a),
    .io_check_env_pma_8_cfg_x(PMPChecker_2_io_check_env_pma_8_cfg_x),
    .io_check_env_pma_8_cfg_w(PMPChecker_2_io_check_env_pma_8_cfg_w),
    .io_check_env_pma_8_cfg_r(PMPChecker_2_io_check_env_pma_8_cfg_r),
    .io_check_env_pma_8_addr(PMPChecker_2_io_check_env_pma_8_addr),
    .io_check_env_pma_8_mask(PMPChecker_2_io_check_env_pma_8_mask),
    .io_check_env_pma_9_cfg_c(PMPChecker_2_io_check_env_pma_9_cfg_c),
    .io_check_env_pma_9_cfg_atomic(PMPChecker_2_io_check_env_pma_9_cfg_atomic),
    .io_check_env_pma_9_cfg_a(PMPChecker_2_io_check_env_pma_9_cfg_a),
    .io_check_env_pma_9_cfg_x(PMPChecker_2_io_check_env_pma_9_cfg_x),
    .io_check_env_pma_9_cfg_w(PMPChecker_2_io_check_env_pma_9_cfg_w),
    .io_check_env_pma_9_cfg_r(PMPChecker_2_io_check_env_pma_9_cfg_r),
    .io_check_env_pma_9_addr(PMPChecker_2_io_check_env_pma_9_addr),
    .io_check_env_pma_9_mask(PMPChecker_2_io_check_env_pma_9_mask),
    .io_check_env_pma_10_cfg_c(PMPChecker_2_io_check_env_pma_10_cfg_c),
    .io_check_env_pma_10_cfg_atomic(PMPChecker_2_io_check_env_pma_10_cfg_atomic),
    .io_check_env_pma_10_cfg_a(PMPChecker_2_io_check_env_pma_10_cfg_a),
    .io_check_env_pma_10_cfg_x(PMPChecker_2_io_check_env_pma_10_cfg_x),
    .io_check_env_pma_10_cfg_w(PMPChecker_2_io_check_env_pma_10_cfg_w),
    .io_check_env_pma_10_cfg_r(PMPChecker_2_io_check_env_pma_10_cfg_r),
    .io_check_env_pma_10_addr(PMPChecker_2_io_check_env_pma_10_addr),
    .io_check_env_pma_10_mask(PMPChecker_2_io_check_env_pma_10_mask),
    .io_check_env_pma_11_cfg_c(PMPChecker_2_io_check_env_pma_11_cfg_c),
    .io_check_env_pma_11_cfg_atomic(PMPChecker_2_io_check_env_pma_11_cfg_atomic),
    .io_check_env_pma_11_cfg_a(PMPChecker_2_io_check_env_pma_11_cfg_a),
    .io_check_env_pma_11_cfg_x(PMPChecker_2_io_check_env_pma_11_cfg_x),
    .io_check_env_pma_11_cfg_w(PMPChecker_2_io_check_env_pma_11_cfg_w),
    .io_check_env_pma_11_cfg_r(PMPChecker_2_io_check_env_pma_11_cfg_r),
    .io_check_env_pma_11_addr(PMPChecker_2_io_check_env_pma_11_addr),
    .io_check_env_pma_11_mask(PMPChecker_2_io_check_env_pma_11_mask),
    .io_check_env_pma_12_cfg_c(PMPChecker_2_io_check_env_pma_12_cfg_c),
    .io_check_env_pma_12_cfg_atomic(PMPChecker_2_io_check_env_pma_12_cfg_atomic),
    .io_check_env_pma_12_cfg_a(PMPChecker_2_io_check_env_pma_12_cfg_a),
    .io_check_env_pma_12_cfg_x(PMPChecker_2_io_check_env_pma_12_cfg_x),
    .io_check_env_pma_12_cfg_w(PMPChecker_2_io_check_env_pma_12_cfg_w),
    .io_check_env_pma_12_cfg_r(PMPChecker_2_io_check_env_pma_12_cfg_r),
    .io_check_env_pma_12_addr(PMPChecker_2_io_check_env_pma_12_addr),
    .io_check_env_pma_12_mask(PMPChecker_2_io_check_env_pma_12_mask),
    .io_check_env_pma_13_cfg_c(PMPChecker_2_io_check_env_pma_13_cfg_c),
    .io_check_env_pma_13_cfg_atomic(PMPChecker_2_io_check_env_pma_13_cfg_atomic),
    .io_check_env_pma_13_cfg_a(PMPChecker_2_io_check_env_pma_13_cfg_a),
    .io_check_env_pma_13_cfg_x(PMPChecker_2_io_check_env_pma_13_cfg_x),
    .io_check_env_pma_13_cfg_w(PMPChecker_2_io_check_env_pma_13_cfg_w),
    .io_check_env_pma_13_cfg_r(PMPChecker_2_io_check_env_pma_13_cfg_r),
    .io_check_env_pma_13_addr(PMPChecker_2_io_check_env_pma_13_addr),
    .io_check_env_pma_13_mask(PMPChecker_2_io_check_env_pma_13_mask),
    .io_check_env_pma_14_cfg_c(PMPChecker_2_io_check_env_pma_14_cfg_c),
    .io_check_env_pma_14_cfg_atomic(PMPChecker_2_io_check_env_pma_14_cfg_atomic),
    .io_check_env_pma_14_cfg_a(PMPChecker_2_io_check_env_pma_14_cfg_a),
    .io_check_env_pma_14_cfg_x(PMPChecker_2_io_check_env_pma_14_cfg_x),
    .io_check_env_pma_14_cfg_w(PMPChecker_2_io_check_env_pma_14_cfg_w),
    .io_check_env_pma_14_cfg_r(PMPChecker_2_io_check_env_pma_14_cfg_r),
    .io_check_env_pma_14_addr(PMPChecker_2_io_check_env_pma_14_addr),
    .io_check_env_pma_14_mask(PMPChecker_2_io_check_env_pma_14_mask),
    .io_check_env_pma_15_cfg_c(PMPChecker_2_io_check_env_pma_15_cfg_c),
    .io_check_env_pma_15_cfg_atomic(PMPChecker_2_io_check_env_pma_15_cfg_atomic),
    .io_check_env_pma_15_cfg_a(PMPChecker_2_io_check_env_pma_15_cfg_a),
    .io_check_env_pma_15_cfg_x(PMPChecker_2_io_check_env_pma_15_cfg_x),
    .io_check_env_pma_15_cfg_w(PMPChecker_2_io_check_env_pma_15_cfg_w),
    .io_check_env_pma_15_cfg_r(PMPChecker_2_io_check_env_pma_15_cfg_r),
    .io_check_env_pma_15_addr(PMPChecker_2_io_check_env_pma_15_addr),
    .io_check_env_pma_15_mask(PMPChecker_2_io_check_env_pma_15_mask),
    .io_req_bits_addr(PMPChecker_2_io_req_bits_addr),
    .io_req_bits_cmd(PMPChecker_2_io_req_bits_cmd),
    .io_resp_ld(PMPChecker_2_io_resp_ld),
    .io_resp_st(PMPChecker_2_io_resp_st),
    .io_resp_instr(PMPChecker_2_io_resp_instr),
    .io_resp_mmio(PMPChecker_2_io_resp_mmio),
    .io_resp_atomic(PMPChecker_2_io_resp_atomic)
  );
  PMPChecker PMPChecker_3 ( // @[Frontend.scala 88:45]
    .io_check_env_mode(PMPChecker_3_io_check_env_mode),
    .io_check_env_pmp_0_cfg_l(PMPChecker_3_io_check_env_pmp_0_cfg_l),
    .io_check_env_pmp_0_cfg_a(PMPChecker_3_io_check_env_pmp_0_cfg_a),
    .io_check_env_pmp_0_cfg_x(PMPChecker_3_io_check_env_pmp_0_cfg_x),
    .io_check_env_pmp_0_cfg_w(PMPChecker_3_io_check_env_pmp_0_cfg_w),
    .io_check_env_pmp_0_cfg_r(PMPChecker_3_io_check_env_pmp_0_cfg_r),
    .io_check_env_pmp_0_addr(PMPChecker_3_io_check_env_pmp_0_addr),
    .io_check_env_pmp_0_mask(PMPChecker_3_io_check_env_pmp_0_mask),
    .io_check_env_pmp_1_cfg_l(PMPChecker_3_io_check_env_pmp_1_cfg_l),
    .io_check_env_pmp_1_cfg_a(PMPChecker_3_io_check_env_pmp_1_cfg_a),
    .io_check_env_pmp_1_cfg_x(PMPChecker_3_io_check_env_pmp_1_cfg_x),
    .io_check_env_pmp_1_cfg_w(PMPChecker_3_io_check_env_pmp_1_cfg_w),
    .io_check_env_pmp_1_cfg_r(PMPChecker_3_io_check_env_pmp_1_cfg_r),
    .io_check_env_pmp_1_addr(PMPChecker_3_io_check_env_pmp_1_addr),
    .io_check_env_pmp_1_mask(PMPChecker_3_io_check_env_pmp_1_mask),
    .io_check_env_pmp_2_cfg_l(PMPChecker_3_io_check_env_pmp_2_cfg_l),
    .io_check_env_pmp_2_cfg_a(PMPChecker_3_io_check_env_pmp_2_cfg_a),
    .io_check_env_pmp_2_cfg_x(PMPChecker_3_io_check_env_pmp_2_cfg_x),
    .io_check_env_pmp_2_cfg_w(PMPChecker_3_io_check_env_pmp_2_cfg_w),
    .io_check_env_pmp_2_cfg_r(PMPChecker_3_io_check_env_pmp_2_cfg_r),
    .io_check_env_pmp_2_addr(PMPChecker_3_io_check_env_pmp_2_addr),
    .io_check_env_pmp_2_mask(PMPChecker_3_io_check_env_pmp_2_mask),
    .io_check_env_pmp_3_cfg_l(PMPChecker_3_io_check_env_pmp_3_cfg_l),
    .io_check_env_pmp_3_cfg_a(PMPChecker_3_io_check_env_pmp_3_cfg_a),
    .io_check_env_pmp_3_cfg_x(PMPChecker_3_io_check_env_pmp_3_cfg_x),
    .io_check_env_pmp_3_cfg_w(PMPChecker_3_io_check_env_pmp_3_cfg_w),
    .io_check_env_pmp_3_cfg_r(PMPChecker_3_io_check_env_pmp_3_cfg_r),
    .io_check_env_pmp_3_addr(PMPChecker_3_io_check_env_pmp_3_addr),
    .io_check_env_pmp_3_mask(PMPChecker_3_io_check_env_pmp_3_mask),
    .io_check_env_pmp_4_cfg_l(PMPChecker_3_io_check_env_pmp_4_cfg_l),
    .io_check_env_pmp_4_cfg_a(PMPChecker_3_io_check_env_pmp_4_cfg_a),
    .io_check_env_pmp_4_cfg_x(PMPChecker_3_io_check_env_pmp_4_cfg_x),
    .io_check_env_pmp_4_cfg_w(PMPChecker_3_io_check_env_pmp_4_cfg_w),
    .io_check_env_pmp_4_cfg_r(PMPChecker_3_io_check_env_pmp_4_cfg_r),
    .io_check_env_pmp_4_addr(PMPChecker_3_io_check_env_pmp_4_addr),
    .io_check_env_pmp_4_mask(PMPChecker_3_io_check_env_pmp_4_mask),
    .io_check_env_pmp_5_cfg_l(PMPChecker_3_io_check_env_pmp_5_cfg_l),
    .io_check_env_pmp_5_cfg_a(PMPChecker_3_io_check_env_pmp_5_cfg_a),
    .io_check_env_pmp_5_cfg_x(PMPChecker_3_io_check_env_pmp_5_cfg_x),
    .io_check_env_pmp_5_cfg_w(PMPChecker_3_io_check_env_pmp_5_cfg_w),
    .io_check_env_pmp_5_cfg_r(PMPChecker_3_io_check_env_pmp_5_cfg_r),
    .io_check_env_pmp_5_addr(PMPChecker_3_io_check_env_pmp_5_addr),
    .io_check_env_pmp_5_mask(PMPChecker_3_io_check_env_pmp_5_mask),
    .io_check_env_pmp_6_cfg_l(PMPChecker_3_io_check_env_pmp_6_cfg_l),
    .io_check_env_pmp_6_cfg_a(PMPChecker_3_io_check_env_pmp_6_cfg_a),
    .io_check_env_pmp_6_cfg_x(PMPChecker_3_io_check_env_pmp_6_cfg_x),
    .io_check_env_pmp_6_cfg_w(PMPChecker_3_io_check_env_pmp_6_cfg_w),
    .io_check_env_pmp_6_cfg_r(PMPChecker_3_io_check_env_pmp_6_cfg_r),
    .io_check_env_pmp_6_addr(PMPChecker_3_io_check_env_pmp_6_addr),
    .io_check_env_pmp_6_mask(PMPChecker_3_io_check_env_pmp_6_mask),
    .io_check_env_pmp_7_cfg_l(PMPChecker_3_io_check_env_pmp_7_cfg_l),
    .io_check_env_pmp_7_cfg_a(PMPChecker_3_io_check_env_pmp_7_cfg_a),
    .io_check_env_pmp_7_cfg_x(PMPChecker_3_io_check_env_pmp_7_cfg_x),
    .io_check_env_pmp_7_cfg_w(PMPChecker_3_io_check_env_pmp_7_cfg_w),
    .io_check_env_pmp_7_cfg_r(PMPChecker_3_io_check_env_pmp_7_cfg_r),
    .io_check_env_pmp_7_addr(PMPChecker_3_io_check_env_pmp_7_addr),
    .io_check_env_pmp_7_mask(PMPChecker_3_io_check_env_pmp_7_mask),
    .io_check_env_pmp_8_cfg_l(PMPChecker_3_io_check_env_pmp_8_cfg_l),
    .io_check_env_pmp_8_cfg_a(PMPChecker_3_io_check_env_pmp_8_cfg_a),
    .io_check_env_pmp_8_cfg_x(PMPChecker_3_io_check_env_pmp_8_cfg_x),
    .io_check_env_pmp_8_cfg_w(PMPChecker_3_io_check_env_pmp_8_cfg_w),
    .io_check_env_pmp_8_cfg_r(PMPChecker_3_io_check_env_pmp_8_cfg_r),
    .io_check_env_pmp_8_addr(PMPChecker_3_io_check_env_pmp_8_addr),
    .io_check_env_pmp_8_mask(PMPChecker_3_io_check_env_pmp_8_mask),
    .io_check_env_pmp_9_cfg_l(PMPChecker_3_io_check_env_pmp_9_cfg_l),
    .io_check_env_pmp_9_cfg_a(PMPChecker_3_io_check_env_pmp_9_cfg_a),
    .io_check_env_pmp_9_cfg_x(PMPChecker_3_io_check_env_pmp_9_cfg_x),
    .io_check_env_pmp_9_cfg_w(PMPChecker_3_io_check_env_pmp_9_cfg_w),
    .io_check_env_pmp_9_cfg_r(PMPChecker_3_io_check_env_pmp_9_cfg_r),
    .io_check_env_pmp_9_addr(PMPChecker_3_io_check_env_pmp_9_addr),
    .io_check_env_pmp_9_mask(PMPChecker_3_io_check_env_pmp_9_mask),
    .io_check_env_pmp_10_cfg_l(PMPChecker_3_io_check_env_pmp_10_cfg_l),
    .io_check_env_pmp_10_cfg_a(PMPChecker_3_io_check_env_pmp_10_cfg_a),
    .io_check_env_pmp_10_cfg_x(PMPChecker_3_io_check_env_pmp_10_cfg_x),
    .io_check_env_pmp_10_cfg_w(PMPChecker_3_io_check_env_pmp_10_cfg_w),
    .io_check_env_pmp_10_cfg_r(PMPChecker_3_io_check_env_pmp_10_cfg_r),
    .io_check_env_pmp_10_addr(PMPChecker_3_io_check_env_pmp_10_addr),
    .io_check_env_pmp_10_mask(PMPChecker_3_io_check_env_pmp_10_mask),
    .io_check_env_pmp_11_cfg_l(PMPChecker_3_io_check_env_pmp_11_cfg_l),
    .io_check_env_pmp_11_cfg_a(PMPChecker_3_io_check_env_pmp_11_cfg_a),
    .io_check_env_pmp_11_cfg_x(PMPChecker_3_io_check_env_pmp_11_cfg_x),
    .io_check_env_pmp_11_cfg_w(PMPChecker_3_io_check_env_pmp_11_cfg_w),
    .io_check_env_pmp_11_cfg_r(PMPChecker_3_io_check_env_pmp_11_cfg_r),
    .io_check_env_pmp_11_addr(PMPChecker_3_io_check_env_pmp_11_addr),
    .io_check_env_pmp_11_mask(PMPChecker_3_io_check_env_pmp_11_mask),
    .io_check_env_pmp_12_cfg_l(PMPChecker_3_io_check_env_pmp_12_cfg_l),
    .io_check_env_pmp_12_cfg_a(PMPChecker_3_io_check_env_pmp_12_cfg_a),
    .io_check_env_pmp_12_cfg_x(PMPChecker_3_io_check_env_pmp_12_cfg_x),
    .io_check_env_pmp_12_cfg_w(PMPChecker_3_io_check_env_pmp_12_cfg_w),
    .io_check_env_pmp_12_cfg_r(PMPChecker_3_io_check_env_pmp_12_cfg_r),
    .io_check_env_pmp_12_addr(PMPChecker_3_io_check_env_pmp_12_addr),
    .io_check_env_pmp_12_mask(PMPChecker_3_io_check_env_pmp_12_mask),
    .io_check_env_pmp_13_cfg_l(PMPChecker_3_io_check_env_pmp_13_cfg_l),
    .io_check_env_pmp_13_cfg_a(PMPChecker_3_io_check_env_pmp_13_cfg_a),
    .io_check_env_pmp_13_cfg_x(PMPChecker_3_io_check_env_pmp_13_cfg_x),
    .io_check_env_pmp_13_cfg_w(PMPChecker_3_io_check_env_pmp_13_cfg_w),
    .io_check_env_pmp_13_cfg_r(PMPChecker_3_io_check_env_pmp_13_cfg_r),
    .io_check_env_pmp_13_addr(PMPChecker_3_io_check_env_pmp_13_addr),
    .io_check_env_pmp_13_mask(PMPChecker_3_io_check_env_pmp_13_mask),
    .io_check_env_pmp_14_cfg_l(PMPChecker_3_io_check_env_pmp_14_cfg_l),
    .io_check_env_pmp_14_cfg_a(PMPChecker_3_io_check_env_pmp_14_cfg_a),
    .io_check_env_pmp_14_cfg_x(PMPChecker_3_io_check_env_pmp_14_cfg_x),
    .io_check_env_pmp_14_cfg_w(PMPChecker_3_io_check_env_pmp_14_cfg_w),
    .io_check_env_pmp_14_cfg_r(PMPChecker_3_io_check_env_pmp_14_cfg_r),
    .io_check_env_pmp_14_addr(PMPChecker_3_io_check_env_pmp_14_addr),
    .io_check_env_pmp_14_mask(PMPChecker_3_io_check_env_pmp_14_mask),
    .io_check_env_pmp_15_cfg_l(PMPChecker_3_io_check_env_pmp_15_cfg_l),
    .io_check_env_pmp_15_cfg_a(PMPChecker_3_io_check_env_pmp_15_cfg_a),
    .io_check_env_pmp_15_cfg_x(PMPChecker_3_io_check_env_pmp_15_cfg_x),
    .io_check_env_pmp_15_cfg_w(PMPChecker_3_io_check_env_pmp_15_cfg_w),
    .io_check_env_pmp_15_cfg_r(PMPChecker_3_io_check_env_pmp_15_cfg_r),
    .io_check_env_pmp_15_addr(PMPChecker_3_io_check_env_pmp_15_addr),
    .io_check_env_pmp_15_mask(PMPChecker_3_io_check_env_pmp_15_mask),
    .io_check_env_pma_0_cfg_c(PMPChecker_3_io_check_env_pma_0_cfg_c),
    .io_check_env_pma_0_cfg_atomic(PMPChecker_3_io_check_env_pma_0_cfg_atomic),
    .io_check_env_pma_0_cfg_a(PMPChecker_3_io_check_env_pma_0_cfg_a),
    .io_check_env_pma_0_cfg_x(PMPChecker_3_io_check_env_pma_0_cfg_x),
    .io_check_env_pma_0_cfg_w(PMPChecker_3_io_check_env_pma_0_cfg_w),
    .io_check_env_pma_0_cfg_r(PMPChecker_3_io_check_env_pma_0_cfg_r),
    .io_check_env_pma_0_addr(PMPChecker_3_io_check_env_pma_0_addr),
    .io_check_env_pma_0_mask(PMPChecker_3_io_check_env_pma_0_mask),
    .io_check_env_pma_1_cfg_c(PMPChecker_3_io_check_env_pma_1_cfg_c),
    .io_check_env_pma_1_cfg_atomic(PMPChecker_3_io_check_env_pma_1_cfg_atomic),
    .io_check_env_pma_1_cfg_a(PMPChecker_3_io_check_env_pma_1_cfg_a),
    .io_check_env_pma_1_cfg_x(PMPChecker_3_io_check_env_pma_1_cfg_x),
    .io_check_env_pma_1_cfg_w(PMPChecker_3_io_check_env_pma_1_cfg_w),
    .io_check_env_pma_1_cfg_r(PMPChecker_3_io_check_env_pma_1_cfg_r),
    .io_check_env_pma_1_addr(PMPChecker_3_io_check_env_pma_1_addr),
    .io_check_env_pma_1_mask(PMPChecker_3_io_check_env_pma_1_mask),
    .io_check_env_pma_2_cfg_c(PMPChecker_3_io_check_env_pma_2_cfg_c),
    .io_check_env_pma_2_cfg_atomic(PMPChecker_3_io_check_env_pma_2_cfg_atomic),
    .io_check_env_pma_2_cfg_a(PMPChecker_3_io_check_env_pma_2_cfg_a),
    .io_check_env_pma_2_cfg_x(PMPChecker_3_io_check_env_pma_2_cfg_x),
    .io_check_env_pma_2_cfg_w(PMPChecker_3_io_check_env_pma_2_cfg_w),
    .io_check_env_pma_2_cfg_r(PMPChecker_3_io_check_env_pma_2_cfg_r),
    .io_check_env_pma_2_addr(PMPChecker_3_io_check_env_pma_2_addr),
    .io_check_env_pma_2_mask(PMPChecker_3_io_check_env_pma_2_mask),
    .io_check_env_pma_3_cfg_c(PMPChecker_3_io_check_env_pma_3_cfg_c),
    .io_check_env_pma_3_cfg_atomic(PMPChecker_3_io_check_env_pma_3_cfg_atomic),
    .io_check_env_pma_3_cfg_a(PMPChecker_3_io_check_env_pma_3_cfg_a),
    .io_check_env_pma_3_cfg_x(PMPChecker_3_io_check_env_pma_3_cfg_x),
    .io_check_env_pma_3_cfg_w(PMPChecker_3_io_check_env_pma_3_cfg_w),
    .io_check_env_pma_3_cfg_r(PMPChecker_3_io_check_env_pma_3_cfg_r),
    .io_check_env_pma_3_addr(PMPChecker_3_io_check_env_pma_3_addr),
    .io_check_env_pma_3_mask(PMPChecker_3_io_check_env_pma_3_mask),
    .io_check_env_pma_4_cfg_c(PMPChecker_3_io_check_env_pma_4_cfg_c),
    .io_check_env_pma_4_cfg_atomic(PMPChecker_3_io_check_env_pma_4_cfg_atomic),
    .io_check_env_pma_4_cfg_a(PMPChecker_3_io_check_env_pma_4_cfg_a),
    .io_check_env_pma_4_cfg_x(PMPChecker_3_io_check_env_pma_4_cfg_x),
    .io_check_env_pma_4_cfg_w(PMPChecker_3_io_check_env_pma_4_cfg_w),
    .io_check_env_pma_4_cfg_r(PMPChecker_3_io_check_env_pma_4_cfg_r),
    .io_check_env_pma_4_addr(PMPChecker_3_io_check_env_pma_4_addr),
    .io_check_env_pma_4_mask(PMPChecker_3_io_check_env_pma_4_mask),
    .io_check_env_pma_5_cfg_c(PMPChecker_3_io_check_env_pma_5_cfg_c),
    .io_check_env_pma_5_cfg_atomic(PMPChecker_3_io_check_env_pma_5_cfg_atomic),
    .io_check_env_pma_5_cfg_a(PMPChecker_3_io_check_env_pma_5_cfg_a),
    .io_check_env_pma_5_cfg_x(PMPChecker_3_io_check_env_pma_5_cfg_x),
    .io_check_env_pma_5_cfg_w(PMPChecker_3_io_check_env_pma_5_cfg_w),
    .io_check_env_pma_5_cfg_r(PMPChecker_3_io_check_env_pma_5_cfg_r),
    .io_check_env_pma_5_addr(PMPChecker_3_io_check_env_pma_5_addr),
    .io_check_env_pma_5_mask(PMPChecker_3_io_check_env_pma_5_mask),
    .io_check_env_pma_6_cfg_c(PMPChecker_3_io_check_env_pma_6_cfg_c),
    .io_check_env_pma_6_cfg_atomic(PMPChecker_3_io_check_env_pma_6_cfg_atomic),
    .io_check_env_pma_6_cfg_a(PMPChecker_3_io_check_env_pma_6_cfg_a),
    .io_check_env_pma_6_cfg_x(PMPChecker_3_io_check_env_pma_6_cfg_x),
    .io_check_env_pma_6_cfg_w(PMPChecker_3_io_check_env_pma_6_cfg_w),
    .io_check_env_pma_6_cfg_r(PMPChecker_3_io_check_env_pma_6_cfg_r),
    .io_check_env_pma_6_addr(PMPChecker_3_io_check_env_pma_6_addr),
    .io_check_env_pma_6_mask(PMPChecker_3_io_check_env_pma_6_mask),
    .io_check_env_pma_7_cfg_c(PMPChecker_3_io_check_env_pma_7_cfg_c),
    .io_check_env_pma_7_cfg_atomic(PMPChecker_3_io_check_env_pma_7_cfg_atomic),
    .io_check_env_pma_7_cfg_a(PMPChecker_3_io_check_env_pma_7_cfg_a),
    .io_check_env_pma_7_cfg_x(PMPChecker_3_io_check_env_pma_7_cfg_x),
    .io_check_env_pma_7_cfg_w(PMPChecker_3_io_check_env_pma_7_cfg_w),
    .io_check_env_pma_7_cfg_r(PMPChecker_3_io_check_env_pma_7_cfg_r),
    .io_check_env_pma_7_addr(PMPChecker_3_io_check_env_pma_7_addr),
    .io_check_env_pma_7_mask(PMPChecker_3_io_check_env_pma_7_mask),
    .io_check_env_pma_8_cfg_c(PMPChecker_3_io_check_env_pma_8_cfg_c),
    .io_check_env_pma_8_cfg_atomic(PMPChecker_3_io_check_env_pma_8_cfg_atomic),
    .io_check_env_pma_8_cfg_a(PMPChecker_3_io_check_env_pma_8_cfg_a),
    .io_check_env_pma_8_cfg_x(PMPChecker_3_io_check_env_pma_8_cfg_x),
    .io_check_env_pma_8_cfg_w(PMPChecker_3_io_check_env_pma_8_cfg_w),
    .io_check_env_pma_8_cfg_r(PMPChecker_3_io_check_env_pma_8_cfg_r),
    .io_check_env_pma_8_addr(PMPChecker_3_io_check_env_pma_8_addr),
    .io_check_env_pma_8_mask(PMPChecker_3_io_check_env_pma_8_mask),
    .io_check_env_pma_9_cfg_c(PMPChecker_3_io_check_env_pma_9_cfg_c),
    .io_check_env_pma_9_cfg_atomic(PMPChecker_3_io_check_env_pma_9_cfg_atomic),
    .io_check_env_pma_9_cfg_a(PMPChecker_3_io_check_env_pma_9_cfg_a),
    .io_check_env_pma_9_cfg_x(PMPChecker_3_io_check_env_pma_9_cfg_x),
    .io_check_env_pma_9_cfg_w(PMPChecker_3_io_check_env_pma_9_cfg_w),
    .io_check_env_pma_9_cfg_r(PMPChecker_3_io_check_env_pma_9_cfg_r),
    .io_check_env_pma_9_addr(PMPChecker_3_io_check_env_pma_9_addr),
    .io_check_env_pma_9_mask(PMPChecker_3_io_check_env_pma_9_mask),
    .io_check_env_pma_10_cfg_c(PMPChecker_3_io_check_env_pma_10_cfg_c),
    .io_check_env_pma_10_cfg_atomic(PMPChecker_3_io_check_env_pma_10_cfg_atomic),
    .io_check_env_pma_10_cfg_a(PMPChecker_3_io_check_env_pma_10_cfg_a),
    .io_check_env_pma_10_cfg_x(PMPChecker_3_io_check_env_pma_10_cfg_x),
    .io_check_env_pma_10_cfg_w(PMPChecker_3_io_check_env_pma_10_cfg_w),
    .io_check_env_pma_10_cfg_r(PMPChecker_3_io_check_env_pma_10_cfg_r),
    .io_check_env_pma_10_addr(PMPChecker_3_io_check_env_pma_10_addr),
    .io_check_env_pma_10_mask(PMPChecker_3_io_check_env_pma_10_mask),
    .io_check_env_pma_11_cfg_c(PMPChecker_3_io_check_env_pma_11_cfg_c),
    .io_check_env_pma_11_cfg_atomic(PMPChecker_3_io_check_env_pma_11_cfg_atomic),
    .io_check_env_pma_11_cfg_a(PMPChecker_3_io_check_env_pma_11_cfg_a),
    .io_check_env_pma_11_cfg_x(PMPChecker_3_io_check_env_pma_11_cfg_x),
    .io_check_env_pma_11_cfg_w(PMPChecker_3_io_check_env_pma_11_cfg_w),
    .io_check_env_pma_11_cfg_r(PMPChecker_3_io_check_env_pma_11_cfg_r),
    .io_check_env_pma_11_addr(PMPChecker_3_io_check_env_pma_11_addr),
    .io_check_env_pma_11_mask(PMPChecker_3_io_check_env_pma_11_mask),
    .io_check_env_pma_12_cfg_c(PMPChecker_3_io_check_env_pma_12_cfg_c),
    .io_check_env_pma_12_cfg_atomic(PMPChecker_3_io_check_env_pma_12_cfg_atomic),
    .io_check_env_pma_12_cfg_a(PMPChecker_3_io_check_env_pma_12_cfg_a),
    .io_check_env_pma_12_cfg_x(PMPChecker_3_io_check_env_pma_12_cfg_x),
    .io_check_env_pma_12_cfg_w(PMPChecker_3_io_check_env_pma_12_cfg_w),
    .io_check_env_pma_12_cfg_r(PMPChecker_3_io_check_env_pma_12_cfg_r),
    .io_check_env_pma_12_addr(PMPChecker_3_io_check_env_pma_12_addr),
    .io_check_env_pma_12_mask(PMPChecker_3_io_check_env_pma_12_mask),
    .io_check_env_pma_13_cfg_c(PMPChecker_3_io_check_env_pma_13_cfg_c),
    .io_check_env_pma_13_cfg_atomic(PMPChecker_3_io_check_env_pma_13_cfg_atomic),
    .io_check_env_pma_13_cfg_a(PMPChecker_3_io_check_env_pma_13_cfg_a),
    .io_check_env_pma_13_cfg_x(PMPChecker_3_io_check_env_pma_13_cfg_x),
    .io_check_env_pma_13_cfg_w(PMPChecker_3_io_check_env_pma_13_cfg_w),
    .io_check_env_pma_13_cfg_r(PMPChecker_3_io_check_env_pma_13_cfg_r),
    .io_check_env_pma_13_addr(PMPChecker_3_io_check_env_pma_13_addr),
    .io_check_env_pma_13_mask(PMPChecker_3_io_check_env_pma_13_mask),
    .io_check_env_pma_14_cfg_c(PMPChecker_3_io_check_env_pma_14_cfg_c),
    .io_check_env_pma_14_cfg_atomic(PMPChecker_3_io_check_env_pma_14_cfg_atomic),
    .io_check_env_pma_14_cfg_a(PMPChecker_3_io_check_env_pma_14_cfg_a),
    .io_check_env_pma_14_cfg_x(PMPChecker_3_io_check_env_pma_14_cfg_x),
    .io_check_env_pma_14_cfg_w(PMPChecker_3_io_check_env_pma_14_cfg_w),
    .io_check_env_pma_14_cfg_r(PMPChecker_3_io_check_env_pma_14_cfg_r),
    .io_check_env_pma_14_addr(PMPChecker_3_io_check_env_pma_14_addr),
    .io_check_env_pma_14_mask(PMPChecker_3_io_check_env_pma_14_mask),
    .io_check_env_pma_15_cfg_c(PMPChecker_3_io_check_env_pma_15_cfg_c),
    .io_check_env_pma_15_cfg_atomic(PMPChecker_3_io_check_env_pma_15_cfg_atomic),
    .io_check_env_pma_15_cfg_a(PMPChecker_3_io_check_env_pma_15_cfg_a),
    .io_check_env_pma_15_cfg_x(PMPChecker_3_io_check_env_pma_15_cfg_x),
    .io_check_env_pma_15_cfg_w(PMPChecker_3_io_check_env_pma_15_cfg_w),
    .io_check_env_pma_15_cfg_r(PMPChecker_3_io_check_env_pma_15_cfg_r),
    .io_check_env_pma_15_addr(PMPChecker_3_io_check_env_pma_15_addr),
    .io_check_env_pma_15_mask(PMPChecker_3_io_check_env_pma_15_mask),
    .io_req_bits_addr(PMPChecker_3_io_req_bits_addr),
    .io_req_bits_cmd(PMPChecker_3_io_req_bits_cmd),
    .io_resp_ld(PMPChecker_3_io_resp_ld),
    .io_resp_st(PMPChecker_3_io_resp_st),
    .io_resp_instr(PMPChecker_3_io_resp_instr),
    .io_resp_mmio(PMPChecker_3_io_resp_mmio),
    .io_resp_atomic(PMPChecker_3_io_resp_atomic)
  );
  TLB itlb ( // @[Frontend.scala 104:20]
    .clock(itlb_clock),
    .reset(itlb_reset),
    .io_sfence_valid(itlb_io_sfence_valid),
    .io_sfence_bits_rs1(itlb_io_sfence_bits_rs1),
    .io_sfence_bits_rs2(itlb_io_sfence_bits_rs2),
    .io_sfence_bits_addr(itlb_io_sfence_bits_addr),
    .io_sfence_bits_asid(itlb_io_sfence_bits_asid),
    .io_csr_satp_mode(itlb_io_csr_satp_mode),
    .io_csr_satp_asid(itlb_io_csr_satp_asid),
    .io_csr_satp_changed(itlb_io_csr_satp_changed),
    .io_csr_priv_imode(itlb_io_csr_priv_imode),
    .io_requestor_0_req_ready(itlb_io_requestor_0_req_ready),
    .io_requestor_0_req_valid(itlb_io_requestor_0_req_valid),
    .io_requestor_0_req_bits_vaddr(itlb_io_requestor_0_req_bits_vaddr),
    .io_requestor_0_req_bits_kill(itlb_io_requestor_0_req_bits_kill),
    .io_requestor_0_resp_ready(itlb_io_requestor_0_resp_ready),
    .io_requestor_0_resp_valid(itlb_io_requestor_0_resp_valid),
    .io_requestor_0_resp_bits_paddr_0(itlb_io_requestor_0_resp_bits_paddr_0),
    .io_requestor_0_resp_bits_excp_0_pf_instr(itlb_io_requestor_0_resp_bits_excp_0_pf_instr),
    .io_requestor_0_resp_bits_excp_0_af_instr(itlb_io_requestor_0_resp_bits_excp_0_af_instr),
    .io_requestor_1_req_ready(itlb_io_requestor_1_req_ready),
    .io_requestor_1_req_valid(itlb_io_requestor_1_req_valid),
    .io_requestor_1_req_bits_vaddr(itlb_io_requestor_1_req_bits_vaddr),
    .io_requestor_1_req_bits_kill(itlb_io_requestor_1_req_bits_kill),
    .io_requestor_1_resp_ready(itlb_io_requestor_1_resp_ready),
    .io_requestor_1_resp_valid(itlb_io_requestor_1_resp_valid),
    .io_requestor_1_resp_bits_paddr_0(itlb_io_requestor_1_resp_bits_paddr_0),
    .io_requestor_1_resp_bits_excp_0_pf_instr(itlb_io_requestor_1_resp_bits_excp_0_pf_instr),
    .io_requestor_1_resp_bits_excp_0_af_instr(itlb_io_requestor_1_resp_bits_excp_0_af_instr),
    .io_requestor_3_req_ready(itlb_io_requestor_3_req_ready),
    .io_requestor_3_req_valid(itlb_io_requestor_3_req_valid),
    .io_requestor_3_req_bits_vaddr(itlb_io_requestor_3_req_bits_vaddr),
    .io_requestor_3_resp_valid(itlb_io_requestor_3_resp_valid),
    .io_requestor_3_resp_bits_paddr_0(itlb_io_requestor_3_resp_bits_paddr_0),
    .io_requestor_3_resp_bits_miss(itlb_io_requestor_3_resp_bits_miss),
    .io_requestor_3_resp_bits_excp_0_pf_instr(itlb_io_requestor_3_resp_bits_excp_0_pf_instr),
    .io_requestor_3_resp_bits_excp_0_af_instr(itlb_io_requestor_3_resp_bits_excp_0_af_instr),
    .io_flushPipe_0(itlb_io_flushPipe_0),
    .io_flushPipe_1(itlb_io_flushPipe_1),
    .io_flushPipe_3(itlb_io_flushPipe_3),
    .io_ptw_req_0_ready(itlb_io_ptw_req_0_ready),
    .io_ptw_req_0_valid(itlb_io_ptw_req_0_valid),
    .io_ptw_req_0_bits_vpn(itlb_io_ptw_req_0_bits_vpn),
    .io_ptw_req_1_ready(itlb_io_ptw_req_1_ready),
    .io_ptw_req_1_valid(itlb_io_ptw_req_1_valid),
    .io_ptw_req_1_bits_vpn(itlb_io_ptw_req_1_bits_vpn),
    .io_ptw_req_3_ready(itlb_io_ptw_req_3_ready),
    .io_ptw_req_3_valid(itlb_io_ptw_req_3_valid),
    .io_ptw_req_3_bits_vpn(itlb_io_ptw_req_3_bits_vpn),
    .io_ptw_resp_ready(itlb_io_ptw_resp_ready),
    .io_ptw_resp_valid(itlb_io_ptw_resp_valid),
    .io_ptw_resp_bits_entry_tag(itlb_io_ptw_resp_bits_entry_tag),
    .io_ptw_resp_bits_entry_asid(itlb_io_ptw_resp_bits_entry_asid),
    .io_ptw_resp_bits_entry_ppn(itlb_io_ptw_resp_bits_entry_ppn),
    .io_ptw_resp_bits_entry_perm_d(itlb_io_ptw_resp_bits_entry_perm_d),
    .io_ptw_resp_bits_entry_perm_a(itlb_io_ptw_resp_bits_entry_perm_a),
    .io_ptw_resp_bits_entry_perm_g(itlb_io_ptw_resp_bits_entry_perm_g),
    .io_ptw_resp_bits_entry_perm_u(itlb_io_ptw_resp_bits_entry_perm_u),
    .io_ptw_resp_bits_entry_perm_x(itlb_io_ptw_resp_bits_entry_perm_x),
    .io_ptw_resp_bits_entry_perm_w(itlb_io_ptw_resp_bits_entry_perm_w),
    .io_ptw_resp_bits_entry_perm_r(itlb_io_ptw_resp_bits_entry_perm_r),
    .io_ptw_resp_bits_entry_level(itlb_io_ptw_resp_bits_entry_level),
    .io_ptw_resp_bits_pf(itlb_io_ptw_resp_bits_pf),
    .io_ptw_resp_bits_af(itlb_io_ptw_resp_bits_af)
  );
  PFEvent pfevent ( // @[Frontend.scala 165:23]
    .clock(pfevent_clock),
    .reset(pfevent_reset),
    .io_distribute_csr_wvalid(pfevent_io_distribute_csr_wvalid),
    .io_distribute_csr_waddr(pfevent_io_distribute_csr_waddr),
    .io_distribute_csr_wdata(pfevent_io_distribute_csr_wdata),
    .io_hpmevent_0(pfevent_io_hpmevent_0),
    .io_hpmevent_1(pfevent_io_hpmevent_1),
    .io_hpmevent_2(pfevent_io_hpmevent_2),
    .io_hpmevent_3(pfevent_io_hpmevent_3),
    .io_hpmevent_4(pfevent_io_hpmevent_4),
    .io_hpmevent_5(pfevent_io_hpmevent_5),
    .io_hpmevent_6(pfevent_io_hpmevent_6),
    .io_hpmevent_7(pfevent_io_hpmevent_7),
    .io_hpmevent_8(pfevent_io_hpmevent_8),
    .io_hpmevent_9(pfevent_io_hpmevent_9),
    .io_hpmevent_10(pfevent_io_hpmevent_10),
    .io_hpmevent_11(pfevent_io_hpmevent_11),
    .io_hpmevent_12(pfevent_io_hpmevent_12),
    .io_hpmevent_13(pfevent_io_hpmevent_13),
    .io_hpmevent_14(pfevent_io_hpmevent_14),
    .io_hpmevent_15(pfevent_io_hpmevent_15),
    .io_hpmevent_16(pfevent_io_hpmevent_16),
    .io_hpmevent_17(pfevent_io_hpmevent_17),
    .io_hpmevent_18(pfevent_io_hpmevent_18),
    .io_hpmevent_19(pfevent_io_hpmevent_19),
    .io_hpmevent_20(pfevent_io_hpmevent_20),
    .io_hpmevent_21(pfevent_io_hpmevent_21),
    .io_hpmevent_22(pfevent_io_hpmevent_22),
    .io_hpmevent_23(pfevent_io_hpmevent_23)
  );
  HPerfMonitor hpm ( // @[PerfCounterUtils.scala 255:21]
    .clock(hpm_clock),
    .io_hpm_event_0(hpm_io_hpm_event_0),
    .io_hpm_event_1(hpm_io_hpm_event_1),
    .io_hpm_event_2(hpm_io_hpm_event_2),
    .io_hpm_event_3(hpm_io_hpm_event_3),
    .io_hpm_event_4(hpm_io_hpm_event_4),
    .io_hpm_event_5(hpm_io_hpm_event_5),
    .io_hpm_event_6(hpm_io_hpm_event_6),
    .io_hpm_event_7(hpm_io_hpm_event_7),
    .io_events_sets_0_value(hpm_io_events_sets_0_value),
    .io_events_sets_1_value(hpm_io_events_sets_1_value),
    .io_events_sets_2_value(hpm_io_events_sets_2_value),
    .io_events_sets_3_value(hpm_io_events_sets_3_value),
    .io_events_sets_4_value(hpm_io_events_sets_4_value),
    .io_events_sets_5_value(hpm_io_events_sets_5_value),
    .io_events_sets_6_value(hpm_io_events_sets_6_value),
    .io_events_sets_7_value(hpm_io_events_sets_7_value),
    .io_events_sets_8_value(hpm_io_events_sets_8_value),
    .io_events_sets_9_value(hpm_io_events_sets_9_value),
    .io_events_sets_10_value(hpm_io_events_sets_10_value),
    .io_events_sets_11_value(hpm_io_events_sets_11_value),
    .io_events_sets_12_value(hpm_io_events_sets_12_value),
    .io_events_sets_13_value(hpm_io_events_sets_13_value),
    .io_events_sets_14_value(hpm_io_events_sets_14_value),
    .io_events_sets_15_value(hpm_io_events_sets_15_value),
    .io_events_sets_16_value(hpm_io_events_sets_16_value),
    .io_events_sets_17_value(hpm_io_events_sets_17_value),
    .io_events_sets_18_value(hpm_io_events_sets_18_value),
    .io_events_sets_19_value(hpm_io_events_sets_19_value),
    .io_events_sets_20_value(hpm_io_events_sets_20_value),
    .io_events_sets_23_value(hpm_io_events_sets_23_value),
    .io_events_sets_24_value(hpm_io_events_sets_24_value),
    .io_events_sets_25_value(hpm_io_events_sets_25_value),
    .io_events_sets_26_value(hpm_io_events_sets_26_value),
    .io_events_sets_27_value(hpm_io_events_sets_27_value),
    .io_events_sets_28_value(hpm_io_events_sets_28_value),
    .io_events_sets_29_value(hpm_io_events_sets_29_value),
    .io_events_sets_30_value(hpm_io_events_sets_30_value),
    .io_events_sets_31_value(hpm_io_events_sets_31_value),
    .io_events_sets_32_value(hpm_io_events_sets_32_value),
    .io_events_sets_33_value(hpm_io_events_sets_33_value),
    .io_events_sets_34_value(hpm_io_events_sets_34_value),
    .io_events_sets_35_value(hpm_io_events_sets_35_value),
    .io_events_sets_36_value(hpm_io_events_sets_36_value),
    .io_events_sets_37_value(hpm_io_events_sets_37_value),
    .io_events_sets_38_value(hpm_io_events_sets_38_value),
    .io_events_sets_39_value(hpm_io_events_sets_39_value),
    .io_events_sets_40_value(hpm_io_events_sets_40_value),
    .io_events_sets_41_value(hpm_io_events_sets_41_value),
    .io_events_sets_42_value(hpm_io_events_sets_42_value),
    .io_events_sets_43_value(hpm_io_events_sets_43_value),
    .io_events_sets_44_value(hpm_io_events_sets_44_value),
    .io_events_sets_45_value(hpm_io_events_sets_45_value),
    .io_events_sets_46_value(hpm_io_events_sets_46_value),
    .io_events_sets_47_value(hpm_io_events_sets_47_value),
    .io_events_sets_48_value(hpm_io_events_sets_48_value),
    .io_events_sets_49_value(hpm_io_events_sets_49_value),
    .io_events_sets_50_value(hpm_io_events_sets_50_value),
    .io_events_sets_51_value(hpm_io_events_sets_51_value),
    .io_events_sets_52_value(hpm_io_events_sets_52_value),
    .io_events_sets_53_value(hpm_io_events_sets_53_value),
    .io_perf_0_value(hpm_io_perf_0_value),
    .io_perf_1_value(hpm_io_perf_1_value),
    .io_perf_2_value(hpm_io_perf_2_value),
    .io_perf_3_value(hpm_io_perf_3_value),
    .io_perf_4_value(hpm_io_perf_4_value),
    .io_perf_5_value(hpm_io_perf_5_value),
    .io_perf_6_value(hpm_io_perf_6_value),
    .io_perf_7_value(hpm_io_perf_7_value)
  );
  assign auto_icache_client_out_a_valid = icache_auto_client_out_a_valid; // @[LazyModule.scala 311:12]
  assign auto_icache_client_out_a_bits_opcode = icache_auto_client_out_a_bits_opcode; // @[LazyModule.scala 311:12]
  assign auto_icache_client_out_a_bits_size = icache_auto_client_out_a_bits_size; // @[LazyModule.scala 311:12]
  assign auto_icache_client_out_a_bits_source = icache_auto_client_out_a_bits_source; // @[LazyModule.scala 311:12]
  assign auto_icache_client_out_a_bits_address = icache_auto_client_out_a_bits_address; // @[LazyModule.scala 311:12]
  assign auto_icache_client_out_a_bits_mask = icache_auto_client_out_a_bits_mask; // @[LazyModule.scala 311:12]
  assign auto_icache_client_out_bready = icache_auto_client_out_bready; // @[LazyModule.scala 311:12]
  assign auto_icache_client_out_c_valid = icache_auto_client_out_c_valid; // @[LazyModule.scala 311:12]
  assign auto_icache_client_out_c_bits_opcode = icache_auto_client_out_c_bits_opcode; // @[LazyModule.scala 311:12]
  assign auto_icache_client_out_c_bits_param = icache_auto_client_out_c_bits_param; // @[LazyModule.scala 311:12]
  assign auto_icache_client_out_c_bits_address = icache_auto_client_out_c_bits_address; // @[LazyModule.scala 311:12]
  assign auto_icache_client_out_c_bits_echo_blockisdirty = icache_auto_client_out_c_bits_echo_blockisdirty; // @[LazyModule.scala 311:12]
  assign auto_icache_client_out_c_bits_data = icache_auto_client_out_c_bits_data; // @[LazyModule.scala 311:12]
  assign auto_icache_client_out_d_ready = icache_auto_client_out_d_ready; // @[LazyModule.scala 311:12]
  assign auto_icache_client_out_e_valid = icache_auto_client_out_e_valid; // @[LazyModule.scala 311:12]
  assign auto_icache_client_out_e_bits_sink = icache_auto_client_out_e_bits_sink; // @[LazyModule.scala 311:12]
  assign auto_instrUncache_client_out_a_valid = instrUncache_auto_client_out_a_valid; // @[LazyModule.scala 311:12]
  assign auto_instrUncache_client_out_a_bits_address = instrUncache_auto_client_out_a_bits_address; // @[LazyModule.scala 311:12]
  assign auto_instrUncache_client_out_d_ready = instrUncache_auto_client_out_d_ready; // @[LazyModule.scala 311:12]
  assign io_ptw_req_0_valid = itlb_io_ptw_req_0_valid; // @[MMUBundle.scala 487:9]
  assign io_ptw_req_0_bits_vpn = itlb_io_ptw_req_0_bits_vpn; // @[MMUBundle.scala 487:9]
  assign io_ptw_req_1_valid = itlb_io_ptw_req_1_valid; // @[MMUBundle.scala 487:9]
  assign io_ptw_req_1_bits_vpn = itlb_io_ptw_req_1_bits_vpn; // @[MMUBundle.scala 487:9]
  assign io_ptw_req_3_valid = itlb_io_ptw_req_3_valid; // @[MMUBundle.scala 487:9]
  assign io_ptw_req_3_bits_vpn = itlb_io_ptw_req_3_bits_vpn; // @[MMUBundle.scala 487:9]
  assign io_backend_cfVec_0_valid = ibuffer_io_out_0_valid; // @[Frontend.scala 151:20]
  assign io_backend_cfVec_0_bits_instr = ibuffer_io_out_0_bits_instr; // @[Frontend.scala 151:20]
  assign io_backend_cfVec_0_bits_foldpc = ibuffer_io_out_0_bits_foldpc; // @[Frontend.scala 151:20]
  assign io_backend_cfVec_0_bits_exceptionVec_1 = ibuffer_io_out_0_bits_exceptionVec_1; // @[Frontend.scala 151:20]
  assign io_backend_cfVec_0_bits_exceptionVec_12 = ibuffer_io_out_0_bits_exceptionVec_12; // @[Frontend.scala 151:20]
  assign io_backend_cfVec_0_bits_trigger_frontendHit_0 = ibuffer_io_out_0_bits_trigger_frontendHit_0; // @[Frontend.scala 151:20]
  assign io_backend_cfVec_0_bits_trigger_frontendHit_1 = ibuffer_io_out_0_bits_trigger_frontendHit_1; // @[Frontend.scala 151:20]
  assign io_backend_cfVec_0_bits_trigger_frontendHit_2 = ibuffer_io_out_0_bits_trigger_frontendHit_2; // @[Frontend.scala 151:20]
  assign io_backend_cfVec_0_bits_trigger_frontendHit_3 = ibuffer_io_out_0_bits_trigger_frontendHit_3; // @[Frontend.scala 151:20]
  assign io_backend_cfVec_0_bits_trigger_backendEn_0 = ibuffer_io_out_0_bits_trigger_backendEn_0; // @[Frontend.scala 151:20]
  assign io_backend_cfVec_0_bits_trigger_backendEn_1 = ibuffer_io_out_0_bits_trigger_backendEn_1; // @[Frontend.scala 151:20]
  assign io_backend_cfVec_0_bits_pd_isRVC = ibuffer_io_out_0_bits_pd_isRVC; // @[Frontend.scala 151:20]
  assign io_backend_cfVec_0_bits_pd_brType = ibuffer_io_out_0_bits_pd_brType; // @[Frontend.scala 151:20]
  assign io_backend_cfVec_0_bits_pd_isCall = ibuffer_io_out_0_bits_pd_isCall; // @[Frontend.scala 151:20]
  assign io_backend_cfVec_0_bits_pd_isRet = ibuffer_io_out_0_bits_pd_isRet; // @[Frontend.scala 151:20]
  assign io_backend_cfVec_0_bits_pred_taken = ibuffer_io_out_0_bits_pred_taken; // @[Frontend.scala 151:20]
  assign io_backend_cfVec_0_bits_crossPageIPFFix = ibuffer_io_out_0_bits_crossPageIPFFix; // @[Frontend.scala 151:20]
  assign io_backend_cfVec_0_bits_ftqPtr_flag = ibuffer_io_out_0_bits_ftqPtr_flag; // @[Frontend.scala 151:20]
  assign io_backend_cfVec_0_bits_ftqPtr_value = ibuffer_io_out_0_bits_ftqPtr_value; // @[Frontend.scala 151:20]
  assign io_backend_cfVec_0_bits_ftqOffset = ibuffer_io_out_0_bits_ftqOffset; // @[Frontend.scala 151:20]
  assign io_backend_cfVec_1_valid = ibuffer_io_out_1_valid; // @[Frontend.scala 151:20]
  assign io_backend_cfVec_1_bits_instr = ibuffer_io_out_1_bits_instr; // @[Frontend.scala 151:20]
  assign io_backend_cfVec_1_bits_foldpc = ibuffer_io_out_1_bits_foldpc; // @[Frontend.scala 151:20]
  assign io_backend_cfVec_1_bits_exceptionVec_1 = ibuffer_io_out_1_bits_exceptionVec_1; // @[Frontend.scala 151:20]
  assign io_backend_cfVec_1_bits_exceptionVec_12 = ibuffer_io_out_1_bits_exceptionVec_12; // @[Frontend.scala 151:20]
  assign io_backend_cfVec_1_bits_trigger_frontendHit_0 = ibuffer_io_out_1_bits_trigger_frontendHit_0; // @[Frontend.scala 151:20]
  assign io_backend_cfVec_1_bits_trigger_frontendHit_1 = ibuffer_io_out_1_bits_trigger_frontendHit_1; // @[Frontend.scala 151:20]
  assign io_backend_cfVec_1_bits_trigger_frontendHit_2 = ibuffer_io_out_1_bits_trigger_frontendHit_2; // @[Frontend.scala 151:20]
  assign io_backend_cfVec_1_bits_trigger_frontendHit_3 = ibuffer_io_out_1_bits_trigger_frontendHit_3; // @[Frontend.scala 151:20]
  assign io_backend_cfVec_1_bits_trigger_backendEn_0 = ibuffer_io_out_1_bits_trigger_backendEn_0; // @[Frontend.scala 151:20]
  assign io_backend_cfVec_1_bits_trigger_backendEn_1 = ibuffer_io_out_1_bits_trigger_backendEn_1; // @[Frontend.scala 151:20]
  assign io_backend_cfVec_1_bits_pd_isRVC = ibuffer_io_out_1_bits_pd_isRVC; // @[Frontend.scala 151:20]
  assign io_backend_cfVec_1_bits_pd_brType = ibuffer_io_out_1_bits_pd_brType; // @[Frontend.scala 151:20]
  assign io_backend_cfVec_1_bits_pd_isCall = ibuffer_io_out_1_bits_pd_isCall; // @[Frontend.scala 151:20]
  assign io_backend_cfVec_1_bits_pd_isRet = ibuffer_io_out_1_bits_pd_isRet; // @[Frontend.scala 151:20]
  assign io_backend_cfVec_1_bits_pred_taken = ibuffer_io_out_1_bits_pred_taken; // @[Frontend.scala 151:20]
  assign io_backend_cfVec_1_bits_crossPageIPFFix = ibuffer_io_out_1_bits_crossPageIPFFix; // @[Frontend.scala 151:20]
  assign io_backend_cfVec_1_bits_ftqPtr_flag = ibuffer_io_out_1_bits_ftqPtr_flag; // @[Frontend.scala 151:20]
  assign io_backend_cfVec_1_bits_ftqPtr_value = ibuffer_io_out_1_bits_ftqPtr_value; // @[Frontend.scala 151:20]
  assign io_backend_cfVec_1_bits_ftqOffset = ibuffer_io_out_1_bits_ftqOffset; // @[Frontend.scala 151:20]
  assign io_backend_fromFtq_pc_mem_wen = ftq_io_toBackend_pc_mem_wen; // @[Frontend.scala 145:22]
  assign io_backend_fromFtq_pc_mem_waddr = ftq_io_toBackend_pc_mem_waddr; // @[Frontend.scala 145:22]
  assign io_backend_fromFtq_pc_mem_wdata_startAddr = ftq_io_toBackend_pc_mem_wdata_startAddr; // @[Frontend.scala 145:22]
  assign io_backend_fromFtq_pc_mem_wdata_nextLineAddr = ftq_io_toBackend_pc_mem_wdata_nextLineAddr; // @[Frontend.scala 145:22]
  assign io_backend_fromFtq_pc_mem_wdata_isNextMask_0 = ftq_io_toBackend_pc_mem_wdata_isNextMask_0; // @[Frontend.scala 145:22]
  assign io_backend_fromFtq_pc_mem_wdata_isNextMask_1 = ftq_io_toBackend_pc_mem_wdata_isNextMask_1; // @[Frontend.scala 145:22]
  assign io_backend_fromFtq_pc_mem_wdata_isNextMask_2 = ftq_io_toBackend_pc_mem_wdata_isNextMask_2; // @[Frontend.scala 145:22]
  assign io_backend_fromFtq_pc_mem_wdata_isNextMask_3 = ftq_io_toBackend_pc_mem_wdata_isNextMask_3; // @[Frontend.scala 145:22]
  assign io_backend_fromFtq_pc_mem_wdata_isNextMask_4 = ftq_io_toBackend_pc_mem_wdata_isNextMask_4; // @[Frontend.scala 145:22]
  assign io_backend_fromFtq_pc_mem_wdata_isNextMask_5 = ftq_io_toBackend_pc_mem_wdata_isNextMask_5; // @[Frontend.scala 145:22]
  assign io_backend_fromFtq_pc_mem_wdata_isNextMask_6 = ftq_io_toBackend_pc_mem_wdata_isNextMask_6; // @[Frontend.scala 145:22]
  assign io_backend_fromFtq_pc_mem_wdata_isNextMask_7 = ftq_io_toBackend_pc_mem_wdata_isNextMask_7; // @[Frontend.scala 145:22]
  assign io_backend_fromFtq_newest_entry_target = ftq_io_toBackend_newest_entry_target; // @[Frontend.scala 145:22]
  assign io_backend_fromFtq_newest_entry_ptr_flag = ftq_io_toBackend_newest_entry_ptr_flag; // @[Frontend.scala 145:22]
  assign io_backend_fromFtq_newest_entry_ptr_value = ftq_io_toBackend_newest_entry_ptr_value; // @[Frontend.scala 145:22]
  assign io_csrUpdate_wvalid = io_csrUpdate_REG_wvalid; // @[Frontend.scala 136:16]
  assign io_csrUpdate_waddr = io_csrUpdate_REG_waddr; // @[Frontend.scala 136:16]
  assign io_csrUpdate_wdata = io_csrUpdate_REG_wdata; // @[Frontend.scala 136:16]
  assign io_error_paddr = io_error_REG_1_paddr; // @[Frontend.scala 156:12]
  assign io_error_report_to_beu = io_error_REG_1_report_to_beu; // @[Frontend.scala 156:12]
  assign io_perf_0_value = io_perf_0_value_REG_1; // @[PerfCounterUtils.scala 188:17]
  assign io_perf_1_value = io_perf_1_value_REG_1; // @[PerfCounterUtils.scala 188:17]
  assign io_perf_2_value = io_perf_2_value_REG_1; // @[PerfCounterUtils.scala 188:17]
  assign io_perf_3_value = io_perf_3_value_REG_1; // @[PerfCounterUtils.scala 188:17]
  assign io_perf_4_value = io_perf_4_value_REG_1; // @[PerfCounterUtils.scala 188:17]
  assign io_perf_5_value = io_perf_5_value_REG_1; // @[PerfCounterUtils.scala 188:17]
  assign io_perf_6_value = io_perf_6_value_REG_1; // @[PerfCounterUtils.scala 188:17]
  assign io_perf_7_value = io_perf_7_value_REG_1; // @[PerfCounterUtils.scala 188:17]
  assign instrUncache_clock = clock;
  assign instrUncache_reset = reset;
  assign instrUncache_auto_client_out_a_ready = auto_instrUncache_client_out_a_ready; // @[LazyModule.scala 311:12]
  assign instrUncache_auto_client_out_d_valid = auto_instrUncache_client_out_d_valid; // @[LazyModule.scala 311:12]
  assign instrUncache_auto_client_out_d_bits_source = auto_instrUncache_client_out_d_bits_source; // @[LazyModule.scala 311:12]
  assign instrUncache_auto_client_out_d_bits_data = auto_instrUncache_client_out_d_bits_data; // @[LazyModule.scala 311:12]
  assign instrUncache_io_req_valid = ifu_io_uncacheInter_toUncache_valid; // @[Frontend.scala 153:25]
  assign instrUncache_io_req_bits_addr = ifu_io_uncacheInter_toUncache_bits_addr; // @[Frontend.scala 153:25]
  assign icache_clock = clock;
  assign icache_reset = reset;
  assign icache_auto_client_out_a_ready = auto_icache_client_out_a_ready; // @[LazyModule.scala 311:12]
  assign icache_auto_client_out_bvalid = auto_icache_client_out_bvalid; // @[LazyModule.scala 311:12]
  assign icache_auto_client_out_bparam = auto_icache_client_out_bparam; // @[LazyModule.scala 311:12]
  assign icache_auto_client_out_baddress = auto_icache_client_out_baddress; // @[LazyModule.scala 311:12]
  assign icache_auto_client_out_bdata = auto_icache_client_out_bdata; // @[LazyModule.scala 311:12]
  assign icache_auto_client_out_c_ready = auto_icache_client_out_c_ready; // @[LazyModule.scala 311:12]
  assign icache_auto_client_out_d_valid = auto_icache_client_out_d_valid; // @[LazyModule.scala 311:12]
  assign icache_auto_client_out_d_bits_opcode = auto_icache_client_out_d_bits_opcode; // @[LazyModule.scala 311:12]
  assign icache_auto_client_out_d_bits_param = auto_icache_client_out_d_bits_param; // @[LazyModule.scala 311:12]
  assign icache_auto_client_out_d_bits_source = auto_icache_client_out_d_bits_source; // @[LazyModule.scala 311:12]
  assign icache_auto_client_out_d_bits_sink = auto_icache_client_out_d_bits_sink; // @[LazyModule.scala 311:12]
  assign icache_auto_client_out_d_bits_echo_blockisdirty = auto_icache_client_out_d_bits_echo_blockisdirty; // @[LazyModule.scala 311:12]
  assign icache_auto_client_out_d_bits_data = auto_icache_client_out_d_bits_data; // @[LazyModule.scala 311:12]
  assign icache_auto_client_out_d_bits_corrupt = auto_icache_client_out_d_bits_corrupt; // @[LazyModule.scala 311:12]
  assign icache_auto_client_out_e_ready = auto_icache_client_out_e_ready; // @[LazyModule.scala 311:12]
  assign icache_io_stop = ifu_io_icacheStop; // @[Frontend.scala 131:18]
  assign icache_io_fetch_req_valid = ftq_io_toICache_req_valid; // @[Frontend.scala 126:23]
  assign icache_io_fetch_req_bits_pcMemRead_0_startAddr = ftq_io_toICache_req_bits_pcMemRead_0_startAddr; // @[Frontend.scala 126:23]
  assign icache_io_fetch_req_bits_pcMemRead_0_nextlineStart = ftq_io_toICache_req_bits_pcMemRead_0_nextlineStart; // @[Frontend.scala 126:23]
  assign icache_io_fetch_req_bits_pcMemRead_1_startAddr = ftq_io_toICache_req_bits_pcMemRead_1_startAddr; // @[Frontend.scala 126:23]
  assign icache_io_fetch_req_bits_pcMemRead_1_nextlineStart = ftq_io_toICache_req_bits_pcMemRead_1_nextlineStart; // @[Frontend.scala 126:23]
  assign icache_io_fetch_req_bits_pcMemRead_2_startAddr = ftq_io_toICache_req_bits_pcMemRead_2_startAddr; // @[Frontend.scala 126:23]
  assign icache_io_fetch_req_bits_pcMemRead_2_nextlineStart = ftq_io_toICache_req_bits_pcMemRead_2_nextlineStart; // @[Frontend.scala 126:23]
  assign icache_io_fetch_req_bits_pcMemRead_3_startAddr = ftq_io_toICache_req_bits_pcMemRead_3_startAddr; // @[Frontend.scala 126:23]
  assign icache_io_fetch_req_bits_pcMemRead_3_nextlineStart = ftq_io_toICache_req_bits_pcMemRead_3_nextlineStart; // @[Frontend.scala 126:23]
  assign icache_io_fetch_req_bits_pcMemRead_4_startAddr = ftq_io_toICache_req_bits_pcMemRead_4_startAddr; // @[Frontend.scala 126:23]
  assign icache_io_fetch_req_bits_pcMemRead_4_nextlineStart = ftq_io_toICache_req_bits_pcMemRead_4_nextlineStart; // @[Frontend.scala 126:23]
  assign icache_io_fetch_req_bits_readValid_0 = ftq_io_toICache_req_bits_readValid_0; // @[Frontend.scala 126:23]
  assign icache_io_fetch_req_bits_readValid_1 = ftq_io_toICache_req_bits_readValid_1; // @[Frontend.scala 126:23]
  assign icache_io_fetch_req_bits_readValid_2 = ftq_io_toICache_req_bits_readValid_2; // @[Frontend.scala 126:23]
  assign icache_io_fetch_req_bits_readValid_3 = ftq_io_toICache_req_bits_readValid_3; // @[Frontend.scala 126:23]
  assign icache_io_fetch_req_bits_readValid_4 = ftq_io_toICache_req_bits_readValid_4; // @[Frontend.scala 126:23]
  assign icache_io_pmp_0_resp_instr = PMPChecker_io_resp_instr; // @[Frontend.scala 88:{26,26}]
  assign icache_io_pmp_0_resp_mmio = PMPChecker_io_resp_mmio; // @[Frontend.scala 88:{26,26}]
  assign icache_io_pmp_1_resp_instr = PMPChecker_1_io_resp_instr; // @[Frontend.scala 88:{26,26}]
  assign icache_io_itlb_0_req_ready = itlb_io_requestor_0_req_ready; // @[Frontend.scala 105:73]
  assign icache_io_itlb_0_resp_valid = itlb_io_requestor_0_resp_valid; // @[Frontend.scala 105:73]
  assign icache_io_itlb_0_resp_bits_paddr_0 = itlb_io_requestor_0_resp_bits_paddr_0; // @[Frontend.scala 105:73]
  assign icache_io_itlb_0_resp_bits_excp_0_pf_instr = itlb_io_requestor_0_resp_bits_excp_0_pf_instr; // @[Frontend.scala 105:73]
  assign icache_io_itlb_0_resp_bits_excp_0_af_instr = itlb_io_requestor_0_resp_bits_excp_0_af_instr; // @[Frontend.scala 105:73]
  assign icache_io_itlb_1_req_ready = itlb_io_requestor_1_req_ready; // @[Frontend.scala 105:73]
  assign icache_io_itlb_1_resp_valid = itlb_io_requestor_1_resp_valid; // @[Frontend.scala 105:73]
  assign icache_io_itlb_1_resp_bits_paddr_0 = itlb_io_requestor_1_resp_bits_paddr_0; // @[Frontend.scala 105:73]
  assign icache_io_itlb_1_resp_bits_excp_0_pf_instr = itlb_io_requestor_1_resp_bits_excp_0_pf_instr; // @[Frontend.scala 105:73]
  assign icache_io_itlb_1_resp_bits_excp_0_af_instr = itlb_io_requestor_1_resp_bits_excp_0_af_instr; // @[Frontend.scala 105:73]
  assign icache_io_csr_distribute_csr_wvalid = csrCtrl_delay_io_out_distribute_csr_wvalid; // @[Frontend.scala 135:32]
  assign icache_io_csr_distribute_csr_waddr = csrCtrl_delay_io_out_distribute_csr_waddr; // @[Frontend.scala 135:32]
  assign icache_io_csr_distribute_csr_wdata = csrCtrl_delay_io_out_distribute_csr_wdata; // @[Frontend.scala 135:32]
  assign icache_io_csr_parity_enable = icache_io_csr_parity_enable_REG; // @[Frontend.scala 139:31]
  assign bpu_clock = clock;
  assign bpu_reset = reset;
  assign bpu_io_bpu_to_ftq_resp_ready = ftq_io_fromBpu_resp_ready; // @[Frontend.scala 121:27]
  assign bpu_io_ftq_to_bpu_redirect_valid = ftq_io_toBpu_redirect_valid; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_redirect_bits_level = ftq_io_toBpu_redirect_bits_level; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_pc = ftq_io_toBpu_redirect_bits_cfiUpdate_pc; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_pd_isRVC = ftq_io_toBpu_redirect_bits_cfiUpdate_pd_isRVC; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_pd_isCall = ftq_io_toBpu_redirect_bits_cfiUpdate_pd_isCall; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_pd_isRet = ftq_io_toBpu_redirect_bits_cfiUpdate_pd_isRet; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_rasSp = ftq_io_toBpu_redirect_bits_cfiUpdate_rasSp; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_rasEntry_retAddr =
    ftq_io_toBpu_redirect_bits_cfiUpdate_rasEntry_retAddr; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_rasEntry_ctr = ftq_io_toBpu_redirect_bits_cfiUpdate_rasEntry_ctr; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_17_folded_hist =
    ftq_io_toBpu_redirect_bits_cfiUpdate_folded_hist_hist_17_folded_hist; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_16_folded_hist =
    ftq_io_toBpu_redirect_bits_cfiUpdate_folded_hist_hist_16_folded_hist; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_15_folded_hist =
    ftq_io_toBpu_redirect_bits_cfiUpdate_folded_hist_hist_15_folded_hist; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_14_folded_hist =
    ftq_io_toBpu_redirect_bits_cfiUpdate_folded_hist_hist_14_folded_hist; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_13_folded_hist =
    ftq_io_toBpu_redirect_bits_cfiUpdate_folded_hist_hist_13_folded_hist; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_12_folded_hist =
    ftq_io_toBpu_redirect_bits_cfiUpdate_folded_hist_hist_12_folded_hist; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_11_folded_hist =
    ftq_io_toBpu_redirect_bits_cfiUpdate_folded_hist_hist_11_folded_hist; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_10_folded_hist =
    ftq_io_toBpu_redirect_bits_cfiUpdate_folded_hist_hist_10_folded_hist; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_9_folded_hist =
    ftq_io_toBpu_redirect_bits_cfiUpdate_folded_hist_hist_9_folded_hist; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_8_folded_hist =
    ftq_io_toBpu_redirect_bits_cfiUpdate_folded_hist_hist_8_folded_hist; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_7_folded_hist =
    ftq_io_toBpu_redirect_bits_cfiUpdate_folded_hist_hist_7_folded_hist; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_6_folded_hist =
    ftq_io_toBpu_redirect_bits_cfiUpdate_folded_hist_hist_6_folded_hist; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_5_folded_hist =
    ftq_io_toBpu_redirect_bits_cfiUpdate_folded_hist_hist_5_folded_hist; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_4_folded_hist =
    ftq_io_toBpu_redirect_bits_cfiUpdate_folded_hist_hist_4_folded_hist; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_3_folded_hist =
    ftq_io_toBpu_redirect_bits_cfiUpdate_folded_hist_hist_3_folded_hist; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_2_folded_hist =
    ftq_io_toBpu_redirect_bits_cfiUpdate_folded_hist_hist_2_folded_hist; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_1_folded_hist =
    ftq_io_toBpu_redirect_bits_cfiUpdate_folded_hist_hist_1_folded_hist; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_folded_hist_hist_0_folded_hist =
    ftq_io_toBpu_redirect_bits_cfiUpdate_folded_hist_hist_0_folded_hist; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_5_bits_0 =
    ftq_io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_5_bits_0; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_5_bits_1 =
    ftq_io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_5_bits_1; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_5_bits_2 =
    ftq_io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_5_bits_2; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_5_bits_3 =
    ftq_io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_5_bits_3; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_4_bits_0 =
    ftq_io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_4_bits_0; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_4_bits_1 =
    ftq_io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_4_bits_1; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_4_bits_2 =
    ftq_io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_4_bits_2; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_3_bits_0 =
    ftq_io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_3_bits_0; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_3_bits_1 =
    ftq_io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_3_bits_1; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_3_bits_2 =
    ftq_io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_3_bits_2; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_3_bits_3 =
    ftq_io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_3_bits_3; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_2_bits_0 =
    ftq_io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_2_bits_0; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_2_bits_1 =
    ftq_io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_2_bits_1; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_2_bits_2 =
    ftq_io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_2_bits_2; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_2_bits_3 =
    ftq_io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_2_bits_3; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_1_bits_0 =
    ftq_io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_1_bits_0; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_1_bits_1 =
    ftq_io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_1_bits_1; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_1_bits_2 =
    ftq_io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_1_bits_2; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_1_bits_3 =
    ftq_io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_1_bits_3; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_0_bits_0 =
    ftq_io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_0_bits_0; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_0_bits_1 =
    ftq_io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_0_bits_1; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_0_bits_2 =
    ftq_io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_0_bits_2; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_afhob_afhob_0_bits_3 =
    ftq_io_toBpu_redirect_bits_cfiUpdate_afhob_afhob_0_bits_3; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_lastBrNumOH = ftq_io_toBpu_redirect_bits_cfiUpdate_lastBrNumOH; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_histPtr_flag = ftq_io_toBpu_redirect_bits_cfiUpdate_histPtr_flag; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_histPtr_value = ftq_io_toBpu_redirect_bits_cfiUpdate_histPtr_value; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_target = ftq_io_toBpu_redirect_bits_cfiUpdate_target; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_taken = ftq_io_toBpu_redirect_bits_cfiUpdate_taken; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_shift = ftq_io_toBpu_redirect_bits_cfiUpdate_shift; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_redirect_bits_cfiUpdate_addIntoHist = ftq_io_toBpu_redirect_bits_cfiUpdate_addIntoHist; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_update_valid = ftq_io_toBpu_update_valid; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_update_bits_pc = ftq_io_toBpu_update_bits_pc; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_17_folded_hist =
    ftq_io_toBpu_update_bits_spec_info_folded_hist_hist_17_folded_hist; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_16_folded_hist =
    ftq_io_toBpu_update_bits_spec_info_folded_hist_hist_16_folded_hist; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_15_folded_hist =
    ftq_io_toBpu_update_bits_spec_info_folded_hist_hist_15_folded_hist; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_14_folded_hist =
    ftq_io_toBpu_update_bits_spec_info_folded_hist_hist_14_folded_hist; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_13_folded_hist =
    ftq_io_toBpu_update_bits_spec_info_folded_hist_hist_13_folded_hist; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_12_folded_hist =
    ftq_io_toBpu_update_bits_spec_info_folded_hist_hist_12_folded_hist; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_10_folded_hist =
    ftq_io_toBpu_update_bits_spec_info_folded_hist_hist_10_folded_hist; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_9_folded_hist =
    ftq_io_toBpu_update_bits_spec_info_folded_hist_hist_9_folded_hist; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_8_folded_hist =
    ftq_io_toBpu_update_bits_spec_info_folded_hist_hist_8_folded_hist; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_7_folded_hist =
    ftq_io_toBpu_update_bits_spec_info_folded_hist_hist_7_folded_hist; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_6_folded_hist =
    ftq_io_toBpu_update_bits_spec_info_folded_hist_hist_6_folded_hist; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_5_folded_hist =
    ftq_io_toBpu_update_bits_spec_info_folded_hist_hist_5_folded_hist; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_4_folded_hist =
    ftq_io_toBpu_update_bits_spec_info_folded_hist_hist_4_folded_hist; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_3_folded_hist =
    ftq_io_toBpu_update_bits_spec_info_folded_hist_hist_3_folded_hist; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_2_folded_hist =
    ftq_io_toBpu_update_bits_spec_info_folded_hist_hist_2_folded_hist; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_1_folded_hist =
    ftq_io_toBpu_update_bits_spec_info_folded_hist_hist_1_folded_hist; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_update_bits_spec_info_folded_hist_hist_0_folded_hist =
    ftq_io_toBpu_update_bits_spec_info_folded_hist_hist_0_folded_hist; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_update_bits_ftb_entry_valid = ftq_io_toBpu_update_bits_ftb_entry_valid; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_update_bits_ftb_entry_brSlots_0_offset = ftq_io_toBpu_update_bits_ftb_entry_brSlots_0_offset; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_update_bits_ftb_entry_brSlots_0_lower = ftq_io_toBpu_update_bits_ftb_entry_brSlots_0_lower; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_update_bits_ftb_entry_brSlots_0_tarStat =
    ftq_io_toBpu_update_bits_ftb_entry_brSlots_0_tarStat; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_update_bits_ftb_entry_brSlots_0_sharing =
    ftq_io_toBpu_update_bits_ftb_entry_brSlots_0_sharing; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_update_bits_ftb_entry_brSlots_0_valid = ftq_io_toBpu_update_bits_ftb_entry_brSlots_0_valid; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_update_bits_ftb_entry_tailSlot_offset = ftq_io_toBpu_update_bits_ftb_entry_tailSlot_offset; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_update_bits_ftb_entry_tailSlot_lower = ftq_io_toBpu_update_bits_ftb_entry_tailSlot_lower; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_update_bits_ftb_entry_tailSlot_tarStat = ftq_io_toBpu_update_bits_ftb_entry_tailSlot_tarStat; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_update_bits_ftb_entry_tailSlot_sharing = ftq_io_toBpu_update_bits_ftb_entry_tailSlot_sharing; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_update_bits_ftb_entry_tailSlot_valid = ftq_io_toBpu_update_bits_ftb_entry_tailSlot_valid; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_update_bits_ftb_entry_pftAddr = ftq_io_toBpu_update_bits_ftb_entry_pftAddr; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_update_bits_ftb_entry_carry = ftq_io_toBpu_update_bits_ftb_entry_carry; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_update_bits_ftb_entry_isCall = ftq_io_toBpu_update_bits_ftb_entry_isCall; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_update_bits_ftb_entry_isRet = ftq_io_toBpu_update_bits_ftb_entry_isRet; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_update_bits_ftb_entry_isJalr = ftq_io_toBpu_update_bits_ftb_entry_isJalr; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_update_bits_ftb_entry_last_may_be_rvi_call =
    ftq_io_toBpu_update_bits_ftb_entry_last_may_be_rvi_call; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_update_bits_ftb_entry_always_taken_0 = ftq_io_toBpu_update_bits_ftb_entry_always_taken_0; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_update_bits_ftb_entry_always_taken_1 = ftq_io_toBpu_update_bits_ftb_entry_always_taken_1; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_update_bits_br_taken_mask_0 = ftq_io_toBpu_update_bits_br_taken_mask_0; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_update_bits_br_taken_mask_1 = ftq_io_toBpu_update_bits_br_taken_mask_1; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_update_bits_jmp_taken = ftq_io_toBpu_update_bits_jmp_taken; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_update_bits_mispred_mask_0 = ftq_io_toBpu_update_bits_mispred_mask_0; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_update_bits_mispred_mask_1 = ftq_io_toBpu_update_bits_mispred_mask_1; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_update_bits_mispred_mask_2 = ftq_io_toBpu_update_bits_mispred_mask_2; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_update_bits_old_entry = ftq_io_toBpu_update_bits_old_entry; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_update_bits_meta = ftq_io_toBpu_update_bits_meta; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_update_bits_full_target = ftq_io_toBpu_update_bits_full_target; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_enq_ptr_flag = ftq_io_toBpu_enq_ptr_flag; // @[Frontend.scala 120:27]
  assign bpu_io_ftq_to_bpu_enq_ptr_value = ftq_io_toBpu_enq_ptr_value; // @[Frontend.scala 120:27]
  assign bpu_io_ctrl_ubtb_enable = csrCtrl_delay_io_out_bp_ctrl_ubtb_enable; // @[Frontend.scala 83:15]
  assign bpu_io_ctrl_btb_enable = csrCtrl_delay_io_out_bp_ctrl_btb_enable; // @[Frontend.scala 83:15]
  assign bpu_io_ctrl_tage_enable = csrCtrl_delay_io_out_bp_ctrl_tage_enable; // @[Frontend.scala 83:15]
  assign bpu_io_ctrl_sc_enable = csrCtrl_delay_io_out_bp_ctrl_sc_enable; // @[Frontend.scala 83:15]
  assign bpu_io_ctrl_ras_enable = csrCtrl_delay_io_out_bp_ctrl_ras_enable; // @[Frontend.scala 83:15]
  assign bpu_io_reset_vector = io_reset_vector; // @[Frontend.scala 84:23]
  assign ifu_clock = clock;
  assign ifu_reset = reset;
  assign ifu_io_ftqInter_fromFtq_req_valid = ftq_io_toIfu_req_valid; // @[Frontend.scala 116:27]
  assign ifu_io_ftqInter_fromFtq_req_bits_startAddr = ftq_io_toIfu_req_bits_startAddr; // @[Frontend.scala 116:27]
  assign ifu_io_ftqInter_fromFtq_req_bits_nextlineStart = ftq_io_toIfu_req_bits_nextlineStart; // @[Frontend.scala 116:27]
  assign ifu_io_ftqInter_fromFtq_req_bits_nextStartAddr = ftq_io_toIfu_req_bits_nextStartAddr; // @[Frontend.scala 116:27]
  assign ifu_io_ftqInter_fromFtq_req_bits_ftqIdx_flag = ftq_io_toIfu_req_bits_ftqIdx_flag; // @[Frontend.scala 116:27]
  assign ifu_io_ftqInter_fromFtq_req_bits_ftqIdx_value = ftq_io_toIfu_req_bits_ftqIdx_value; // @[Frontend.scala 116:27]
  assign ifu_io_ftqInter_fromFtq_req_bits_ftqOffset_valid = ftq_io_toIfu_req_bits_ftqOffset_valid; // @[Frontend.scala 116:27]
  assign ifu_io_ftqInter_fromFtq_req_bits_ftqOffset_bits = ftq_io_toIfu_req_bits_ftqOffset_bits; // @[Frontend.scala 116:27]
  assign ifu_io_ftqInter_fromFtq_redirect_valid = ftq_io_toIfu_redirect_valid; // @[Frontend.scala 116:27]
  assign ifu_io_ftqInter_fromFtq_redirect_bits_ftqIdx_flag = ftq_io_toIfu_redirect_bits_ftqIdx_flag; // @[Frontend.scala 116:27]
  assign ifu_io_ftqInter_fromFtq_redirect_bits_ftqIdx_value = ftq_io_toIfu_redirect_bits_ftqIdx_value; // @[Frontend.scala 116:27]
  assign ifu_io_ftqInter_fromFtq_redirect_bits_ftqOffset = ftq_io_toIfu_redirect_bits_ftqOffset; // @[Frontend.scala 116:27]
  assign ifu_io_ftqInter_fromFtq_redirect_bits_level = ftq_io_toIfu_redirect_bits_level; // @[Frontend.scala 116:27]
  assign ifu_io_ftqInter_fromFtq_flushFromBpu_s2_valid = ftq_io_toIfu_flushFromBpu_s2_valid; // @[Frontend.scala 116:27]
  assign ifu_io_ftqInter_fromFtq_flushFromBpu_s2_bits_flag = ftq_io_toIfu_flushFromBpu_s2_bits_flag; // @[Frontend.scala 116:27]
  assign ifu_io_ftqInter_fromFtq_flushFromBpu_s2_bits_value = ftq_io_toIfu_flushFromBpu_s2_bits_value; // @[Frontend.scala 116:27]
  assign ifu_io_ftqInter_fromFtq_flushFromBpu_s3_valid = ftq_io_toIfu_flushFromBpu_s3_valid; // @[Frontend.scala 116:27]
  assign ifu_io_ftqInter_fromFtq_flushFromBpu_s3_bits_flag = ftq_io_toIfu_flushFromBpu_s3_bits_flag; // @[Frontend.scala 116:27]
  assign ifu_io_ftqInter_fromFtq_flushFromBpu_s3_bits_value = ftq_io_toIfu_flushFromBpu_s3_bits_value; // @[Frontend.scala 116:27]
  assign ifu_io_icacheInter_icacheReady = icache_io_toIFU; // @[Frontend.scala 130:34]
  assign ifu_io_icacheInter_resp_0_valid = icache_io_fetch_resp_0_valid; // @[Frontend.scala 129:27]
  assign ifu_io_icacheInter_resp_0_bits_vaddr = icache_io_fetch_resp_0_bits_vaddr; // @[Frontend.scala 129:27]
  assign ifu_io_icacheInter_resp_0_bits_registerData = icache_io_fetch_resp_0_bits_registerData; // @[Frontend.scala 129:27]
  assign ifu_io_icacheInter_resp_0_bits_sramData = icache_io_fetch_resp_0_bits_sramData; // @[Frontend.scala 129:27]
  assign ifu_io_icacheInter_resp_0_bits_select = icache_io_fetch_resp_0_bits_select; // @[Frontend.scala 129:27]
  assign ifu_io_icacheInter_resp_0_bits_paddr = icache_io_fetch_resp_0_bits_paddr; // @[Frontend.scala 129:27]
  assign ifu_io_icacheInter_resp_0_bits_tlbExcp_pageFault = icache_io_fetch_resp_0_bits_tlbExcp_pageFault; // @[Frontend.scala 129:27]
  assign ifu_io_icacheInter_resp_0_bits_tlbExcp_accessFault = icache_io_fetch_resp_0_bits_tlbExcp_accessFault; // @[Frontend.scala 129:27]
  assign ifu_io_icacheInter_resp_0_bits_tlbExcp_mmio = icache_io_fetch_resp_0_bits_tlbExcp_mmio; // @[Frontend.scala 129:27]
  assign ifu_io_icacheInter_resp_1_valid = icache_io_fetch_resp_1_valid; // @[Frontend.scala 129:27]
  assign ifu_io_icacheInter_resp_1_bits_vaddr = icache_io_fetch_resp_1_bits_vaddr; // @[Frontend.scala 129:27]
  assign ifu_io_icacheInter_resp_1_bits_registerData = icache_io_fetch_resp_1_bits_registerData; // @[Frontend.scala 129:27]
  assign ifu_io_icacheInter_resp_1_bits_sramData = icache_io_fetch_resp_1_bits_sramData; // @[Frontend.scala 129:27]
  assign ifu_io_icacheInter_resp_1_bits_select = icache_io_fetch_resp_1_bits_select; // @[Frontend.scala 129:27]
  assign ifu_io_icacheInter_resp_1_bits_tlbExcp_pageFault = icache_io_fetch_resp_1_bits_tlbExcp_pageFault; // @[Frontend.scala 129:27]
  assign ifu_io_icacheInter_resp_1_bits_tlbExcp_accessFault = icache_io_fetch_resp_1_bits_tlbExcp_accessFault; // @[Frontend.scala 129:27]
  assign ifu_io_icachePerfInfo_only_0_hit = icache_io_perfInfo_only_0_hit; // @[Frontend.scala 133:25]
  assign ifu_io_icachePerfInfo_only_0_miss = icache_io_perfInfo_only_0_miss; // @[Frontend.scala 133:25]
  assign ifu_io_icachePerfInfo_hit_0_hit_1 = icache_io_perfInfo_hit_0_hit_1; // @[Frontend.scala 133:25]
  assign ifu_io_icachePerfInfo_hit_0_miss_1 = icache_io_perfInfo_hit_0_miss_1; // @[Frontend.scala 133:25]
  assign ifu_io_icachePerfInfo_miss_0_hit_1 = icache_io_perfInfo_miss_0_hit_1; // @[Frontend.scala 133:25]
  assign ifu_io_icachePerfInfo_miss_0_miss_1 = icache_io_perfInfo_miss_0_miss_1; // @[Frontend.scala 133:25]
  assign ifu_io_icachePerfInfo_hit_0_except_1 = icache_io_perfInfo_hit_0_except_1; // @[Frontend.scala 133:25]
  assign ifu_io_icachePerfInfo_miss_0_except_1 = icache_io_perfInfo_miss_0_except_1; // @[Frontend.scala 133:25]
  assign ifu_io_icachePerfInfo_except_0 = icache_io_perfInfo_except_0; // @[Frontend.scala 133:25]
  assign ifu_io_icachePerfInfo_bank_hit_1 = icache_io_perfInfo_bank_hit_1; // @[Frontend.scala 133:25]
  assign ifu_io_icachePerfInfo_hit = icache_io_perfInfo_hit; // @[Frontend.scala 133:25]
  assign ifu_io_toIbuffer_ready = ibuffer_io_in_ready; // @[Frontend.scala 142:23]
  assign ifu_io_uncacheInter_fromUncache_valid = instrUncache_io_resp_valid; // @[Frontend.scala 154:35]
  assign ifu_io_uncacheInter_fromUncache_bits_data = instrUncache_io_resp_bits_data; // @[Frontend.scala 154:35]
  assign ifu_io_uncacheInter_toUncache_ready = instrUncache_io_req_ready; // @[Frontend.scala 153:25]
  assign ifu_io_frontendTrigger_t_valid = csrCtrl_delay_io_out_frontend_trigger_t_valid; // @[Frontend.scala 78:26]
  assign ifu_io_frontendTrigger_t_bits_addr = csrCtrl_delay_io_out_frontend_trigger_t_bits_addr; // @[Frontend.scala 78:26]
  assign ifu_io_frontendTrigger_t_bits_tdata_matchType = csrCtrl_delay_io_out_frontend_trigger_t_bits_tdata_matchType; // @[Frontend.scala 78:26]
  assign ifu_io_frontendTrigger_t_bits_tdata_select = csrCtrl_delay_io_out_frontend_trigger_t_bits_tdata_select; // @[Frontend.scala 78:26]
  assign ifu_io_frontendTrigger_t_bits_tdata_timing = csrCtrl_delay_io_out_frontend_trigger_t_bits_tdata_timing; // @[Frontend.scala 78:26]
  assign ifu_io_frontendTrigger_t_bits_tdata_chain = csrCtrl_delay_io_out_frontend_trigger_t_bits_tdata_chain; // @[Frontend.scala 78:26]
  assign ifu_io_frontendTrigger_t_bits_tdata_tdata2 = csrCtrl_delay_io_out_frontend_trigger_t_bits_tdata_tdata2; // @[Frontend.scala 78:26]
  assign ifu_io_csrTriggerEnable_0 = csrCtrl_delay_io_out_trigger_enable_0; // @[Frontend.scala 80:{37,37}]
  assign ifu_io_csrTriggerEnable_1 = csrCtrl_delay_io_out_trigger_enable_1; // @[Frontend.scala 80:{37,37}]
  assign ifu_io_csrTriggerEnable_2 = csrCtrl_delay_io_out_trigger_enable_6; // @[Frontend.scala 80:{37,37}]
  assign ifu_io_csrTriggerEnable_3 = csrCtrl_delay_io_out_trigger_enable_8; // @[Frontend.scala 80:{37,37}]
  assign ifu_io_rob_commits_0_valid = io_backend_toFtq_rob_commits_0_valid; // @[Frontend.scala 148:22]
  assign ifu_io_rob_commits_0_bits_ftqIdx_flag = io_backend_toFtq_rob_commits_0_bits_ftqIdx_flag; // @[Frontend.scala 148:22]
  assign ifu_io_rob_commits_0_bits_ftqIdx_value = io_backend_toFtq_rob_commits_0_bits_ftqIdx_value; // @[Frontend.scala 148:22]
  assign ifu_io_rob_commits_0_bits_ftqOffset = io_backend_toFtq_rob_commits_0_bits_ftqOffset; // @[Frontend.scala 148:22]
  assign ifu_io_rob_commits_1_valid = io_backend_toFtq_rob_commits_1_valid; // @[Frontend.scala 148:22]
  assign ifu_io_rob_commits_1_bits_ftqIdx_flag = io_backend_toFtq_rob_commits_1_bits_ftqIdx_flag; // @[Frontend.scala 148:22]
  assign ifu_io_rob_commits_1_bits_ftqIdx_value = io_backend_toFtq_rob_commits_1_bits_ftqIdx_value; // @[Frontend.scala 148:22]
  assign ifu_io_rob_commits_1_bits_ftqOffset = io_backend_toFtq_rob_commits_1_bits_ftqOffset; // @[Frontend.scala 148:22]
  assign ifu_io_iTLBInter_resp_bits_paddr_0 = itlb_io_requestor_3_resp_bits_paddr_0; // @[Frontend.scala 106:24]
  assign ifu_io_iTLBInter_resp_bits_miss = itlb_io_requestor_3_resp_bits_miss; // @[Frontend.scala 106:24]
  assign ifu_io_iTLBInter_resp_bits_excp_0_pf_instr = itlb_io_requestor_3_resp_bits_excp_0_pf_instr; // @[Frontend.scala 106:24]
  assign ifu_io_iTLBInter_resp_bits_excp_0_af_instr = itlb_io_requestor_3_resp_bits_excp_0_af_instr; // @[Frontend.scala 106:24]
  assign ifu_io_pmp_resp_instr = PMPChecker_3_io_resp_instr; // @[Frontend.scala 88:{26,26}]
  assign ifu_io_pmp_resp_mmio = PMPChecker_3_io_resp_mmio; // @[Frontend.scala 88:{26,26}]
  assign ifu_io_mmioCommitRead_mmioLastCommit = ftq_io_mmioCommitRead_mmioLastCommit; // @[Frontend.scala 123:27]
  assign ibuffer_clock = clock;
  assign ibuffer_reset = reset;
  assign ibuffer_io_flush = needFlush; // @[Frontend.scala 150:20]
  assign ibuffer_io_in_valid = ifu_io_toIbuffer_valid; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_instrs_0 = ifu_io_toIbuffer_bits_instrs_0; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_instrs_1 = ifu_io_toIbuffer_bits_instrs_1; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_instrs_2 = ifu_io_toIbuffer_bits_instrs_2; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_instrs_3 = ifu_io_toIbuffer_bits_instrs_3; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_instrs_4 = ifu_io_toIbuffer_bits_instrs_4; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_instrs_5 = ifu_io_toIbuffer_bits_instrs_5; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_instrs_6 = ifu_io_toIbuffer_bits_instrs_6; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_instrs_7 = ifu_io_toIbuffer_bits_instrs_7; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_valid = ifu_io_toIbuffer_bits_valid; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_enqEnable = ifu_io_toIbuffer_bits_enqEnable; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_pd_0_isRVC = ifu_io_toIbuffer_bits_pd_0_isRVC; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_pd_0_brType = ifu_io_toIbuffer_bits_pd_0_brType; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_pd_0_isCall = ifu_io_toIbuffer_bits_pd_0_isCall; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_pd_0_isRet = ifu_io_toIbuffer_bits_pd_0_isRet; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_pd_1_isRVC = ifu_io_toIbuffer_bits_pd_1_isRVC; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_pd_1_brType = ifu_io_toIbuffer_bits_pd_1_brType; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_pd_1_isCall = ifu_io_toIbuffer_bits_pd_1_isCall; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_pd_1_isRet = ifu_io_toIbuffer_bits_pd_1_isRet; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_pd_2_isRVC = ifu_io_toIbuffer_bits_pd_2_isRVC; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_pd_2_brType = ifu_io_toIbuffer_bits_pd_2_brType; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_pd_2_isCall = ifu_io_toIbuffer_bits_pd_2_isCall; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_pd_2_isRet = ifu_io_toIbuffer_bits_pd_2_isRet; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_pd_3_isRVC = ifu_io_toIbuffer_bits_pd_3_isRVC; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_pd_3_brType = ifu_io_toIbuffer_bits_pd_3_brType; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_pd_3_isCall = ifu_io_toIbuffer_bits_pd_3_isCall; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_pd_3_isRet = ifu_io_toIbuffer_bits_pd_3_isRet; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_pd_4_isRVC = ifu_io_toIbuffer_bits_pd_4_isRVC; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_pd_4_brType = ifu_io_toIbuffer_bits_pd_4_brType; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_pd_4_isCall = ifu_io_toIbuffer_bits_pd_4_isCall; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_pd_4_isRet = ifu_io_toIbuffer_bits_pd_4_isRet; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_pd_5_isRVC = ifu_io_toIbuffer_bits_pd_5_isRVC; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_pd_5_brType = ifu_io_toIbuffer_bits_pd_5_brType; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_pd_5_isCall = ifu_io_toIbuffer_bits_pd_5_isCall; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_pd_5_isRet = ifu_io_toIbuffer_bits_pd_5_isRet; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_pd_6_isRVC = ifu_io_toIbuffer_bits_pd_6_isRVC; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_pd_6_brType = ifu_io_toIbuffer_bits_pd_6_brType; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_pd_6_isCall = ifu_io_toIbuffer_bits_pd_6_isCall; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_pd_6_isRet = ifu_io_toIbuffer_bits_pd_6_isRet; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_pd_7_isRVC = ifu_io_toIbuffer_bits_pd_7_isRVC; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_pd_7_brType = ifu_io_toIbuffer_bits_pd_7_brType; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_pd_7_isCall = ifu_io_toIbuffer_bits_pd_7_isCall; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_pd_7_isRet = ifu_io_toIbuffer_bits_pd_7_isRet; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_foldpc_0 = ifu_io_toIbuffer_bits_foldpc_0; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_foldpc_1 = ifu_io_toIbuffer_bits_foldpc_1; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_foldpc_2 = ifu_io_toIbuffer_bits_foldpc_2; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_foldpc_3 = ifu_io_toIbuffer_bits_foldpc_3; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_foldpc_4 = ifu_io_toIbuffer_bits_foldpc_4; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_foldpc_5 = ifu_io_toIbuffer_bits_foldpc_5; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_foldpc_6 = ifu_io_toIbuffer_bits_foldpc_6; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_foldpc_7 = ifu_io_toIbuffer_bits_foldpc_7; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_ftqPtr_flag = ifu_io_toIbuffer_bits_ftqPtr_flag; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_ftqPtr_value = ifu_io_toIbuffer_bits_ftqPtr_value; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_ftqOffset_0_valid = ifu_io_toIbuffer_bits_ftqOffset_0_valid; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_ftqOffset_1_valid = ifu_io_toIbuffer_bits_ftqOffset_1_valid; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_ftqOffset_2_valid = ifu_io_toIbuffer_bits_ftqOffset_2_valid; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_ftqOffset_3_valid = ifu_io_toIbuffer_bits_ftqOffset_3_valid; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_ftqOffset_4_valid = ifu_io_toIbuffer_bits_ftqOffset_4_valid; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_ftqOffset_5_valid = ifu_io_toIbuffer_bits_ftqOffset_5_valid; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_ftqOffset_6_valid = ifu_io_toIbuffer_bits_ftqOffset_6_valid; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_ftqOffset_7_valid = ifu_io_toIbuffer_bits_ftqOffset_7_valid; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_ipf_0 = ifu_io_toIbuffer_bits_ipf_0; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_ipf_1 = ifu_io_toIbuffer_bits_ipf_1; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_ipf_2 = ifu_io_toIbuffer_bits_ipf_2; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_ipf_3 = ifu_io_toIbuffer_bits_ipf_3; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_ipf_4 = ifu_io_toIbuffer_bits_ipf_4; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_ipf_5 = ifu_io_toIbuffer_bits_ipf_5; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_ipf_6 = ifu_io_toIbuffer_bits_ipf_6; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_ipf_7 = ifu_io_toIbuffer_bits_ipf_7; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_acf_0 = ifu_io_toIbuffer_bits_acf_0; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_acf_1 = ifu_io_toIbuffer_bits_acf_1; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_acf_2 = ifu_io_toIbuffer_bits_acf_2; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_acf_3 = ifu_io_toIbuffer_bits_acf_3; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_acf_4 = ifu_io_toIbuffer_bits_acf_4; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_acf_5 = ifu_io_toIbuffer_bits_acf_5; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_acf_6 = ifu_io_toIbuffer_bits_acf_6; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_acf_7 = ifu_io_toIbuffer_bits_acf_7; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_crossPageIPFFix_0 = ifu_io_toIbuffer_bits_crossPageIPFFix_0; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_crossPageIPFFix_1 = ifu_io_toIbuffer_bits_crossPageIPFFix_1; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_crossPageIPFFix_2 = ifu_io_toIbuffer_bits_crossPageIPFFix_2; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_crossPageIPFFix_3 = ifu_io_toIbuffer_bits_crossPageIPFFix_3; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_crossPageIPFFix_4 = ifu_io_toIbuffer_bits_crossPageIPFFix_4; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_crossPageIPFFix_5 = ifu_io_toIbuffer_bits_crossPageIPFFix_5; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_crossPageIPFFix_6 = ifu_io_toIbuffer_bits_crossPageIPFFix_6; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_crossPageIPFFix_7 = ifu_io_toIbuffer_bits_crossPageIPFFix_7; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_triggered_0_frontendHit_0 = ifu_io_toIbuffer_bits_triggered_0_frontendHit_0; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_triggered_0_frontendHit_1 = ifu_io_toIbuffer_bits_triggered_0_frontendHit_1; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_triggered_0_frontendHit_2 = ifu_io_toIbuffer_bits_triggered_0_frontendHit_2; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_triggered_0_frontendHit_3 = ifu_io_toIbuffer_bits_triggered_0_frontendHit_3; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_triggered_0_backendEn_0 = ifu_io_toIbuffer_bits_triggered_0_backendEn_0; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_triggered_0_backendEn_1 = ifu_io_toIbuffer_bits_triggered_0_backendEn_1; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_triggered_1_frontendHit_0 = ifu_io_toIbuffer_bits_triggered_1_frontendHit_0; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_triggered_1_frontendHit_1 = ifu_io_toIbuffer_bits_triggered_1_frontendHit_1; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_triggered_1_frontendHit_2 = ifu_io_toIbuffer_bits_triggered_1_frontendHit_2; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_triggered_1_frontendHit_3 = ifu_io_toIbuffer_bits_triggered_1_frontendHit_3; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_triggered_1_backendEn_0 = ifu_io_toIbuffer_bits_triggered_1_backendEn_0; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_triggered_1_backendEn_1 = ifu_io_toIbuffer_bits_triggered_1_backendEn_1; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_triggered_2_frontendHit_0 = ifu_io_toIbuffer_bits_triggered_2_frontendHit_0; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_triggered_2_frontendHit_1 = ifu_io_toIbuffer_bits_triggered_2_frontendHit_1; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_triggered_2_frontendHit_2 = ifu_io_toIbuffer_bits_triggered_2_frontendHit_2; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_triggered_2_frontendHit_3 = ifu_io_toIbuffer_bits_triggered_2_frontendHit_3; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_triggered_2_backendEn_0 = ifu_io_toIbuffer_bits_triggered_2_backendEn_0; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_triggered_2_backendEn_1 = ifu_io_toIbuffer_bits_triggered_2_backendEn_1; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_triggered_3_frontendHit_0 = ifu_io_toIbuffer_bits_triggered_3_frontendHit_0; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_triggered_3_frontendHit_1 = ifu_io_toIbuffer_bits_triggered_3_frontendHit_1; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_triggered_3_frontendHit_2 = ifu_io_toIbuffer_bits_triggered_3_frontendHit_2; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_triggered_3_frontendHit_3 = ifu_io_toIbuffer_bits_triggered_3_frontendHit_3; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_triggered_3_backendEn_0 = ifu_io_toIbuffer_bits_triggered_3_backendEn_0; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_triggered_3_backendEn_1 = ifu_io_toIbuffer_bits_triggered_3_backendEn_1; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_triggered_4_frontendHit_0 = ifu_io_toIbuffer_bits_triggered_4_frontendHit_0; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_triggered_4_frontendHit_1 = ifu_io_toIbuffer_bits_triggered_4_frontendHit_1; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_triggered_4_frontendHit_2 = ifu_io_toIbuffer_bits_triggered_4_frontendHit_2; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_triggered_4_frontendHit_3 = ifu_io_toIbuffer_bits_triggered_4_frontendHit_3; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_triggered_4_backendEn_0 = ifu_io_toIbuffer_bits_triggered_4_backendEn_0; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_triggered_4_backendEn_1 = ifu_io_toIbuffer_bits_triggered_4_backendEn_1; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_triggered_5_frontendHit_0 = ifu_io_toIbuffer_bits_triggered_5_frontendHit_0; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_triggered_5_frontendHit_1 = ifu_io_toIbuffer_bits_triggered_5_frontendHit_1; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_triggered_5_frontendHit_2 = ifu_io_toIbuffer_bits_triggered_5_frontendHit_2; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_triggered_5_frontendHit_3 = ifu_io_toIbuffer_bits_triggered_5_frontendHit_3; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_triggered_5_backendEn_0 = ifu_io_toIbuffer_bits_triggered_5_backendEn_0; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_triggered_5_backendEn_1 = ifu_io_toIbuffer_bits_triggered_5_backendEn_1; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_triggered_6_frontendHit_0 = ifu_io_toIbuffer_bits_triggered_6_frontendHit_0; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_triggered_6_frontendHit_1 = ifu_io_toIbuffer_bits_triggered_6_frontendHit_1; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_triggered_6_frontendHit_2 = ifu_io_toIbuffer_bits_triggered_6_frontendHit_2; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_triggered_6_frontendHit_3 = ifu_io_toIbuffer_bits_triggered_6_frontendHit_3; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_triggered_6_backendEn_0 = ifu_io_toIbuffer_bits_triggered_6_backendEn_0; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_triggered_6_backendEn_1 = ifu_io_toIbuffer_bits_triggered_6_backendEn_1; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_triggered_7_frontendHit_0 = ifu_io_toIbuffer_bits_triggered_7_frontendHit_0; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_triggered_7_frontendHit_1 = ifu_io_toIbuffer_bits_triggered_7_frontendHit_1; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_triggered_7_frontendHit_2 = ifu_io_toIbuffer_bits_triggered_7_frontendHit_2; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_triggered_7_frontendHit_3 = ifu_io_toIbuffer_bits_triggered_7_frontendHit_3; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_triggered_7_backendEn_0 = ifu_io_toIbuffer_bits_triggered_7_backendEn_0; // @[Frontend.scala 142:23]
  assign ibuffer_io_in_bits_triggered_7_backendEn_1 = ifu_io_toIbuffer_bits_triggered_7_backendEn_1; // @[Frontend.scala 142:23]
  assign ibuffer_io_out_0_ready = io_backend_cfVec_0_ready; // @[Frontend.scala 151:20]
  assign ibuffer_io_out_1_ready = io_backend_cfVec_1_ready; // @[Frontend.scala 151:20]
  assign ftq_clock = clock;
  assign ftq_reset = reset;
  assign ftq_io_fromBpu_resp_valid = bpu_io_bpu_to_ftq_resp_valid; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_s1_pc = bpu_io_bpu_to_ftq_resp_bits_s1_pc; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_s1_full_pred_br_taken_mask_0 =
    bpu_io_bpu_to_ftq_resp_bits_s1_full_pred_br_taken_mask_0; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_s1_full_pred_br_taken_mask_1 =
    bpu_io_bpu_to_ftq_resp_bits_s1_full_pred_br_taken_mask_1; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_s1_full_pred_slot_valids_0 = bpu_io_bpu_to_ftq_resp_bits_s1_full_pred_slot_valids_0; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_s1_full_pred_slot_valids_1 = bpu_io_bpu_to_ftq_resp_bits_s1_full_pred_slot_valids_1; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_s1_full_pred_targets_0 = bpu_io_bpu_to_ftq_resp_bits_s1_full_pred_targets_0; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_s1_full_pred_targets_1 = bpu_io_bpu_to_ftq_resp_bits_s1_full_pred_targets_1; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_s1_full_pred_offsets_0 = bpu_io_bpu_to_ftq_resp_bits_s1_full_pred_offsets_0; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_s1_full_pred_offsets_1 = bpu_io_bpu_to_ftq_resp_bits_s1_full_pred_offsets_1; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_s1_full_pred_fallThroughAddr =
    bpu_io_bpu_to_ftq_resp_bits_s1_full_pred_fallThroughAddr; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_s1_full_pred_fallThroughErr = bpu_io_bpu_to_ftq_resp_bits_s1_full_pred_fallThroughErr; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_s1_full_pred_is_br_sharing = bpu_io_bpu_to_ftq_resp_bits_s1_full_pred_is_br_sharing; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_s1_full_pred_hit = bpu_io_bpu_to_ftq_resp_bits_s1_full_pred_hit; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_s2_pc = bpu_io_bpu_to_ftq_resp_bits_s2_pc; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_s2_valid = bpu_io_bpu_to_ftq_resp_bits_s2_valid; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_s2_hasRedirect = bpu_io_bpu_to_ftq_resp_bits_s2_hasRedirect; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_s2_ftq_idx_flag = bpu_io_bpu_to_ftq_resp_bits_s2_ftq_idx_flag; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_s2_ftq_idx_value = bpu_io_bpu_to_ftq_resp_bits_s2_ftq_idx_value; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_s2_full_pred_br_taken_mask_0 =
    bpu_io_bpu_to_ftq_resp_bits_s2_full_pred_br_taken_mask_0; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_s2_full_pred_br_taken_mask_1 =
    bpu_io_bpu_to_ftq_resp_bits_s2_full_pred_br_taken_mask_1; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_s2_full_pred_slot_valids_0 = bpu_io_bpu_to_ftq_resp_bits_s2_full_pred_slot_valids_0; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_s2_full_pred_slot_valids_1 = bpu_io_bpu_to_ftq_resp_bits_s2_full_pred_slot_valids_1; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_s2_full_pred_targets_0 = bpu_io_bpu_to_ftq_resp_bits_s2_full_pred_targets_0; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_s2_full_pred_targets_1 = bpu_io_bpu_to_ftq_resp_bits_s2_full_pred_targets_1; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_s2_full_pred_offsets_0 = bpu_io_bpu_to_ftq_resp_bits_s2_full_pred_offsets_0; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_s2_full_pred_offsets_1 = bpu_io_bpu_to_ftq_resp_bits_s2_full_pred_offsets_1; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_s2_full_pred_fallThroughAddr =
    bpu_io_bpu_to_ftq_resp_bits_s2_full_pred_fallThroughAddr; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_s2_full_pred_fallThroughErr = bpu_io_bpu_to_ftq_resp_bits_s2_full_pred_fallThroughErr; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_s2_full_pred_is_br_sharing = bpu_io_bpu_to_ftq_resp_bits_s2_full_pred_is_br_sharing; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_s2_full_pred_hit = bpu_io_bpu_to_ftq_resp_bits_s2_full_pred_hit; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_s3_pc = bpu_io_bpu_to_ftq_resp_bits_s3_pc; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_s3_valid = bpu_io_bpu_to_ftq_resp_bits_s3_valid; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_s3_hasRedirect = bpu_io_bpu_to_ftq_resp_bits_s3_hasRedirect; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_s3_ftq_idx_flag = bpu_io_bpu_to_ftq_resp_bits_s3_ftq_idx_flag; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_s3_ftq_idx_value = bpu_io_bpu_to_ftq_resp_bits_s3_ftq_idx_value; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_s3_full_pred_br_taken_mask_0 =
    bpu_io_bpu_to_ftq_resp_bits_s3_full_pred_br_taken_mask_0; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_s3_full_pred_br_taken_mask_1 =
    bpu_io_bpu_to_ftq_resp_bits_s3_full_pred_br_taken_mask_1; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_s3_full_pred_slot_valids_0 = bpu_io_bpu_to_ftq_resp_bits_s3_full_pred_slot_valids_0; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_s3_full_pred_slot_valids_1 = bpu_io_bpu_to_ftq_resp_bits_s3_full_pred_slot_valids_1; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_s3_full_pred_targets_0 = bpu_io_bpu_to_ftq_resp_bits_s3_full_pred_targets_0; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_s3_full_pred_targets_1 = bpu_io_bpu_to_ftq_resp_bits_s3_full_pred_targets_1; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_s3_full_pred_offsets_0 = bpu_io_bpu_to_ftq_resp_bits_s3_full_pred_offsets_0; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_s3_full_pred_offsets_1 = bpu_io_bpu_to_ftq_resp_bits_s3_full_pred_offsets_1; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_s3_full_pred_fallThroughAddr =
    bpu_io_bpu_to_ftq_resp_bits_s3_full_pred_fallThroughAddr; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_s3_full_pred_fallThroughErr = bpu_io_bpu_to_ftq_resp_bits_s3_full_pred_fallThroughErr; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_s3_full_pred_is_br_sharing = bpu_io_bpu_to_ftq_resp_bits_s3_full_pred_is_br_sharing; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_s3_full_pred_hit = bpu_io_bpu_to_ftq_resp_bits_s3_full_pred_hit; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_last_stage_meta = bpu_io_bpu_to_ftq_resp_bits_last_stage_meta; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_last_stage_spec_info_folded_hist_hist_17_folded_hist =
    bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_17_folded_hist; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_last_stage_spec_info_folded_hist_hist_16_folded_hist =
    bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_16_folded_hist; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_last_stage_spec_info_folded_hist_hist_15_folded_hist =
    bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_15_folded_hist; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_last_stage_spec_info_folded_hist_hist_14_folded_hist =
    bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_14_folded_hist; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_last_stage_spec_info_folded_hist_hist_13_folded_hist =
    bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_13_folded_hist; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_last_stage_spec_info_folded_hist_hist_12_folded_hist =
    bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_12_folded_hist; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_last_stage_spec_info_folded_hist_hist_11_folded_hist =
    bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_11_folded_hist; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_last_stage_spec_info_folded_hist_hist_10_folded_hist =
    bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_10_folded_hist; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_last_stage_spec_info_folded_hist_hist_9_folded_hist =
    bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_9_folded_hist; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_last_stage_spec_info_folded_hist_hist_8_folded_hist =
    bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_8_folded_hist; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_last_stage_spec_info_folded_hist_hist_7_folded_hist =
    bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_7_folded_hist; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_last_stage_spec_info_folded_hist_hist_6_folded_hist =
    bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_6_folded_hist; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_last_stage_spec_info_folded_hist_hist_5_folded_hist =
    bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_5_folded_hist; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_last_stage_spec_info_folded_hist_hist_4_folded_hist =
    bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_4_folded_hist; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_last_stage_spec_info_folded_hist_hist_3_folded_hist =
    bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_3_folded_hist; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_last_stage_spec_info_folded_hist_hist_2_folded_hist =
    bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_2_folded_hist; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_last_stage_spec_info_folded_hist_hist_1_folded_hist =
    bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_1_folded_hist; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_last_stage_spec_info_folded_hist_hist_0_folded_hist =
    bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_folded_hist_hist_0_folded_hist; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_5_bits_0 =
    bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_5_bits_0; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_5_bits_1 =
    bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_5_bits_1; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_5_bits_2 =
    bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_5_bits_2; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_5_bits_3 =
    bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_5_bits_3; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_4_bits_0 =
    bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_4_bits_0; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_4_bits_1 =
    bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_4_bits_1; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_4_bits_2 =
    bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_4_bits_2; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_4_bits_3 =
    bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_4_bits_3; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_3_bits_0 =
    bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_3_bits_0; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_3_bits_1 =
    bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_3_bits_1; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_3_bits_2 =
    bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_3_bits_2; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_3_bits_3 =
    bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_3_bits_3; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_2_bits_0 =
    bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_2_bits_0; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_2_bits_1 =
    bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_2_bits_1; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_2_bits_2 =
    bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_2_bits_2; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_2_bits_3 =
    bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_2_bits_3; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_1_bits_0 =
    bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_1_bits_0; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_1_bits_1 =
    bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_1_bits_1; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_1_bits_2 =
    bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_1_bits_2; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_1_bits_3 =
    bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_1_bits_3; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_0_bits_0 =
    bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_0_bits_0; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_0_bits_1 =
    bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_0_bits_1; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_0_bits_2 =
    bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_0_bits_2; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_last_stage_spec_info_afhob_afhob_0_bits_3 =
    bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_afhob_afhob_0_bits_3; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_last_stage_spec_info_lastBrNumOH =
    bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_lastBrNumOH; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_last_stage_spec_info_histPtr_flag =
    bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_histPtr_flag; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_last_stage_spec_info_histPtr_value =
    bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_histPtr_value; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_last_stage_spec_info_rasSp = bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_rasSp; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_last_stage_spec_info_rasTop_retAddr =
    bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_rasTop_retAddr; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_last_stage_spec_info_rasTop_ctr =
    bpu_io_bpu_to_ftq_resp_bits_last_stage_spec_info_rasTop_ctr; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_last_stage_ftb_entry_valid = bpu_io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_valid; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_last_stage_ftb_entry_brSlots_0_offset =
    bpu_io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_brSlots_0_offset; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_last_stage_ftb_entry_brSlots_0_lower =
    bpu_io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_brSlots_0_lower; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_last_stage_ftb_entry_brSlots_0_tarStat =
    bpu_io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_brSlots_0_tarStat; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_last_stage_ftb_entry_brSlots_0_sharing =
    bpu_io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_brSlots_0_sharing; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_last_stage_ftb_entry_brSlots_0_valid =
    bpu_io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_brSlots_0_valid; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_last_stage_ftb_entry_tailSlot_offset =
    bpu_io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_tailSlot_offset; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_last_stage_ftb_entry_tailSlot_lower =
    bpu_io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_tailSlot_lower; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_last_stage_ftb_entry_tailSlot_tarStat =
    bpu_io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_tailSlot_tarStat; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_last_stage_ftb_entry_tailSlot_sharing =
    bpu_io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_tailSlot_sharing; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_last_stage_ftb_entry_tailSlot_valid =
    bpu_io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_tailSlot_valid; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_last_stage_ftb_entry_pftAddr =
    bpu_io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_pftAddr; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_last_stage_ftb_entry_carry = bpu_io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_carry; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_last_stage_ftb_entry_isCall = bpu_io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_isCall; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_last_stage_ftb_entry_isRet = bpu_io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_isRet; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_last_stage_ftb_entry_isJalr = bpu_io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_isJalr; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_last_stage_ftb_entry_last_may_be_rvi_call =
    bpu_io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_last_may_be_rvi_call; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_last_stage_ftb_entry_always_taken_0 =
    bpu_io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_always_taken_0; // @[Frontend.scala 121:27]
  assign ftq_io_fromBpu_resp_bits_last_stage_ftb_entry_always_taken_1 =
    bpu_io_bpu_to_ftq_resp_bits_last_stage_ftb_entry_always_taken_1; // @[Frontend.scala 121:27]
  assign ftq_io_fromIfu_pdWb_valid = ifu_io_ftqInter_toFtq_pdWb_valid; // @[Frontend.scala 119:27]
  assign ftq_io_fromIfu_pdWb_bits_pc_0 = ifu_io_ftqInter_toFtq_pdWb_bits_pc_0; // @[Frontend.scala 119:27]
  assign ftq_io_fromIfu_pdWb_bits_pc_1 = ifu_io_ftqInter_toFtq_pdWb_bits_pc_1; // @[Frontend.scala 119:27]
  assign ftq_io_fromIfu_pdWb_bits_pc_2 = ifu_io_ftqInter_toFtq_pdWb_bits_pc_2; // @[Frontend.scala 119:27]
  assign ftq_io_fromIfu_pdWb_bits_pc_3 = ifu_io_ftqInter_toFtq_pdWb_bits_pc_3; // @[Frontend.scala 119:27]
  assign ftq_io_fromIfu_pdWb_bits_pc_4 = ifu_io_ftqInter_toFtq_pdWb_bits_pc_4; // @[Frontend.scala 119:27]
  assign ftq_io_fromIfu_pdWb_bits_pc_5 = ifu_io_ftqInter_toFtq_pdWb_bits_pc_5; // @[Frontend.scala 119:27]
  assign ftq_io_fromIfu_pdWb_bits_pc_6 = ifu_io_ftqInter_toFtq_pdWb_bits_pc_6; // @[Frontend.scala 119:27]
  assign ftq_io_fromIfu_pdWb_bits_pc_7 = ifu_io_ftqInter_toFtq_pdWb_bits_pc_7; // @[Frontend.scala 119:27]
  assign ftq_io_fromIfu_pdWb_bits_pd_0_valid = ifu_io_ftqInter_toFtq_pdWb_bits_pd_0_valid; // @[Frontend.scala 119:27]
  assign ftq_io_fromIfu_pdWb_bits_pd_0_isRVC = ifu_io_ftqInter_toFtq_pdWb_bits_pd_0_isRVC; // @[Frontend.scala 119:27]
  assign ftq_io_fromIfu_pdWb_bits_pd_0_brType = ifu_io_ftqInter_toFtq_pdWb_bits_pd_0_brType; // @[Frontend.scala 119:27]
  assign ftq_io_fromIfu_pdWb_bits_pd_0_isCall = ifu_io_ftqInter_toFtq_pdWb_bits_pd_0_isCall; // @[Frontend.scala 119:27]
  assign ftq_io_fromIfu_pdWb_bits_pd_0_isRet = ifu_io_ftqInter_toFtq_pdWb_bits_pd_0_isRet; // @[Frontend.scala 119:27]
  assign ftq_io_fromIfu_pdWb_bits_pd_1_valid = ifu_io_ftqInter_toFtq_pdWb_bits_pd_1_valid; // @[Frontend.scala 119:27]
  assign ftq_io_fromIfu_pdWb_bits_pd_1_isRVC = ifu_io_ftqInter_toFtq_pdWb_bits_pd_1_isRVC; // @[Frontend.scala 119:27]
  assign ftq_io_fromIfu_pdWb_bits_pd_1_brType = ifu_io_ftqInter_toFtq_pdWb_bits_pd_1_brType; // @[Frontend.scala 119:27]
  assign ftq_io_fromIfu_pdWb_bits_pd_1_isCall = ifu_io_ftqInter_toFtq_pdWb_bits_pd_1_isCall; // @[Frontend.scala 119:27]
  assign ftq_io_fromIfu_pdWb_bits_pd_1_isRet = ifu_io_ftqInter_toFtq_pdWb_bits_pd_1_isRet; // @[Frontend.scala 119:27]
  assign ftq_io_fromIfu_pdWb_bits_pd_2_valid = ifu_io_ftqInter_toFtq_pdWb_bits_pd_2_valid; // @[Frontend.scala 119:27]
  assign ftq_io_fromIfu_pdWb_bits_pd_2_isRVC = ifu_io_ftqInter_toFtq_pdWb_bits_pd_2_isRVC; // @[Frontend.scala 119:27]
  assign ftq_io_fromIfu_pdWb_bits_pd_2_brType = ifu_io_ftqInter_toFtq_pdWb_bits_pd_2_brType; // @[Frontend.scala 119:27]
  assign ftq_io_fromIfu_pdWb_bits_pd_2_isCall = ifu_io_ftqInter_toFtq_pdWb_bits_pd_2_isCall; // @[Frontend.scala 119:27]
  assign ftq_io_fromIfu_pdWb_bits_pd_2_isRet = ifu_io_ftqInter_toFtq_pdWb_bits_pd_2_isRet; // @[Frontend.scala 119:27]
  assign ftq_io_fromIfu_pdWb_bits_pd_3_valid = ifu_io_ftqInter_toFtq_pdWb_bits_pd_3_valid; // @[Frontend.scala 119:27]
  assign ftq_io_fromIfu_pdWb_bits_pd_3_isRVC = ifu_io_ftqInter_toFtq_pdWb_bits_pd_3_isRVC; // @[Frontend.scala 119:27]
  assign ftq_io_fromIfu_pdWb_bits_pd_3_brType = ifu_io_ftqInter_toFtq_pdWb_bits_pd_3_brType; // @[Frontend.scala 119:27]
  assign ftq_io_fromIfu_pdWb_bits_pd_3_isCall = ifu_io_ftqInter_toFtq_pdWb_bits_pd_3_isCall; // @[Frontend.scala 119:27]
  assign ftq_io_fromIfu_pdWb_bits_pd_3_isRet = ifu_io_ftqInter_toFtq_pdWb_bits_pd_3_isRet; // @[Frontend.scala 119:27]
  assign ftq_io_fromIfu_pdWb_bits_pd_4_valid = ifu_io_ftqInter_toFtq_pdWb_bits_pd_4_valid; // @[Frontend.scala 119:27]
  assign ftq_io_fromIfu_pdWb_bits_pd_4_isRVC = ifu_io_ftqInter_toFtq_pdWb_bits_pd_4_isRVC; // @[Frontend.scala 119:27]
  assign ftq_io_fromIfu_pdWb_bits_pd_4_brType = ifu_io_ftqInter_toFtq_pdWb_bits_pd_4_brType; // @[Frontend.scala 119:27]
  assign ftq_io_fromIfu_pdWb_bits_pd_4_isCall = ifu_io_ftqInter_toFtq_pdWb_bits_pd_4_isCall; // @[Frontend.scala 119:27]
  assign ftq_io_fromIfu_pdWb_bits_pd_4_isRet = ifu_io_ftqInter_toFtq_pdWb_bits_pd_4_isRet; // @[Frontend.scala 119:27]
  assign ftq_io_fromIfu_pdWb_bits_pd_5_valid = ifu_io_ftqInter_toFtq_pdWb_bits_pd_5_valid; // @[Frontend.scala 119:27]
  assign ftq_io_fromIfu_pdWb_bits_pd_5_isRVC = ifu_io_ftqInter_toFtq_pdWb_bits_pd_5_isRVC; // @[Frontend.scala 119:27]
  assign ftq_io_fromIfu_pdWb_bits_pd_5_brType = ifu_io_ftqInter_toFtq_pdWb_bits_pd_5_brType; // @[Frontend.scala 119:27]
  assign ftq_io_fromIfu_pdWb_bits_pd_5_isCall = ifu_io_ftqInter_toFtq_pdWb_bits_pd_5_isCall; // @[Frontend.scala 119:27]
  assign ftq_io_fromIfu_pdWb_bits_pd_5_isRet = ifu_io_ftqInter_toFtq_pdWb_bits_pd_5_isRet; // @[Frontend.scala 119:27]
  assign ftq_io_fromIfu_pdWb_bits_pd_6_valid = ifu_io_ftqInter_toFtq_pdWb_bits_pd_6_valid; // @[Frontend.scala 119:27]
  assign ftq_io_fromIfu_pdWb_bits_pd_6_isRVC = ifu_io_ftqInter_toFtq_pdWb_bits_pd_6_isRVC; // @[Frontend.scala 119:27]
  assign ftq_io_fromIfu_pdWb_bits_pd_6_brType = ifu_io_ftqInter_toFtq_pdWb_bits_pd_6_brType; // @[Frontend.scala 119:27]
  assign ftq_io_fromIfu_pdWb_bits_pd_6_isCall = ifu_io_ftqInter_toFtq_pdWb_bits_pd_6_isCall; // @[Frontend.scala 119:27]
  assign ftq_io_fromIfu_pdWb_bits_pd_6_isRet = ifu_io_ftqInter_toFtq_pdWb_bits_pd_6_isRet; // @[Frontend.scala 119:27]
  assign ftq_io_fromIfu_pdWb_bits_pd_7_valid = ifu_io_ftqInter_toFtq_pdWb_bits_pd_7_valid; // @[Frontend.scala 119:27]
  assign ftq_io_fromIfu_pdWb_bits_pd_7_isRVC = ifu_io_ftqInter_toFtq_pdWb_bits_pd_7_isRVC; // @[Frontend.scala 119:27]
  assign ftq_io_fromIfu_pdWb_bits_pd_7_brType = ifu_io_ftqInter_toFtq_pdWb_bits_pd_7_brType; // @[Frontend.scala 119:27]
  assign ftq_io_fromIfu_pdWb_bits_pd_7_isCall = ifu_io_ftqInter_toFtq_pdWb_bits_pd_7_isCall; // @[Frontend.scala 119:27]
  assign ftq_io_fromIfu_pdWb_bits_pd_7_isRet = ifu_io_ftqInter_toFtq_pdWb_bits_pd_7_isRet; // @[Frontend.scala 119:27]
  assign ftq_io_fromIfu_pdWb_bits_ftqIdx_flag = ifu_io_ftqInter_toFtq_pdWb_bits_ftqIdx_flag; // @[Frontend.scala 119:27]
  assign ftq_io_fromIfu_pdWb_bits_ftqIdx_value = ifu_io_ftqInter_toFtq_pdWb_bits_ftqIdx_value; // @[Frontend.scala 119:27]
  assign ftq_io_fromIfu_pdWb_bits_misOffset_valid = ifu_io_ftqInter_toFtq_pdWb_bits_misOffset_valid; // @[Frontend.scala 119:27]
  assign ftq_io_fromIfu_pdWb_bits_misOffset_bits = ifu_io_ftqInter_toFtq_pdWb_bits_misOffset_bits; // @[Frontend.scala 119:27]
  assign ftq_io_fromIfu_pdWb_bits_cfiOffset_valid = ifu_io_ftqInter_toFtq_pdWb_bits_cfiOffset_valid; // @[Frontend.scala 119:27]
  assign ftq_io_fromIfu_pdWb_bits_target = ifu_io_ftqInter_toFtq_pdWb_bits_target; // @[Frontend.scala 119:27]
  assign ftq_io_fromIfu_pdWb_bits_jalTarget = ifu_io_ftqInter_toFtq_pdWb_bits_jalTarget; // @[Frontend.scala 119:27]
  assign ftq_io_fromIfu_pdWb_bits_instrRange_0 = ifu_io_ftqInter_toFtq_pdWb_bits_instrRange_0; // @[Frontend.scala 119:27]
  assign ftq_io_fromIfu_pdWb_bits_instrRange_1 = ifu_io_ftqInter_toFtq_pdWb_bits_instrRange_1; // @[Frontend.scala 119:27]
  assign ftq_io_fromIfu_pdWb_bits_instrRange_2 = ifu_io_ftqInter_toFtq_pdWb_bits_instrRange_2; // @[Frontend.scala 119:27]
  assign ftq_io_fromIfu_pdWb_bits_instrRange_3 = ifu_io_ftqInter_toFtq_pdWb_bits_instrRange_3; // @[Frontend.scala 119:27]
  assign ftq_io_fromIfu_pdWb_bits_instrRange_4 = ifu_io_ftqInter_toFtq_pdWb_bits_instrRange_4; // @[Frontend.scala 119:27]
  assign ftq_io_fromIfu_pdWb_bits_instrRange_5 = ifu_io_ftqInter_toFtq_pdWb_bits_instrRange_5; // @[Frontend.scala 119:27]
  assign ftq_io_fromIfu_pdWb_bits_instrRange_6 = ifu_io_ftqInter_toFtq_pdWb_bits_instrRange_6; // @[Frontend.scala 119:27]
  assign ftq_io_fromIfu_pdWb_bits_instrRange_7 = ifu_io_ftqInter_toFtq_pdWb_bits_instrRange_7; // @[Frontend.scala 119:27]
  assign ftq_io_fromBackend_rob_commits_0_valid = io_backend_toFtq_rob_commits_0_valid; // @[Frontend.scala 144:22]
  assign ftq_io_fromBackend_rob_commits_0_bits_commitType = io_backend_toFtq_rob_commits_0_bits_commitType; // @[Frontend.scala 144:22]
  assign ftq_io_fromBackend_rob_commits_0_bits_ftqIdx_flag = io_backend_toFtq_rob_commits_0_bits_ftqIdx_flag; // @[Frontend.scala 144:22]
  assign ftq_io_fromBackend_rob_commits_0_bits_ftqIdx_value = io_backend_toFtq_rob_commits_0_bits_ftqIdx_value; // @[Frontend.scala 144:22]
  assign ftq_io_fromBackend_rob_commits_0_bits_ftqOffset = io_backend_toFtq_rob_commits_0_bits_ftqOffset; // @[Frontend.scala 144:22]
  assign ftq_io_fromBackend_rob_commits_1_valid = io_backend_toFtq_rob_commits_1_valid; // @[Frontend.scala 144:22]
  assign ftq_io_fromBackend_rob_commits_1_bits_commitType = io_backend_toFtq_rob_commits_1_bits_commitType; // @[Frontend.scala 144:22]
  assign ftq_io_fromBackend_rob_commits_1_bits_ftqIdx_flag = io_backend_toFtq_rob_commits_1_bits_ftqIdx_flag; // @[Frontend.scala 144:22]
  assign ftq_io_fromBackend_rob_commits_1_bits_ftqIdx_value = io_backend_toFtq_rob_commits_1_bits_ftqIdx_value; // @[Frontend.scala 144:22]
  assign ftq_io_fromBackend_rob_commits_1_bits_ftqOffset = io_backend_toFtq_rob_commits_1_bits_ftqOffset; // @[Frontend.scala 144:22]
  assign ftq_io_fromBackend_redirect_valid = io_backend_toFtq_redirect_valid; // @[Frontend.scala 144:22]
  assign ftq_io_fromBackend_redirect_bits_ftqIdx_flag = io_backend_toFtq_redirect_bits_ftqIdx_flag; // @[Frontend.scala 144:22]
  assign ftq_io_fromBackend_redirect_bits_ftqIdx_value = io_backend_toFtq_redirect_bits_ftqIdx_value; // @[Frontend.scala 144:22]
  assign ftq_io_fromBackend_redirect_bits_ftqOffset = io_backend_toFtq_redirect_bits_ftqOffset; // @[Frontend.scala 144:22]
  assign ftq_io_fromBackend_redirect_bits_level = io_backend_toFtq_redirect_bits_level; // @[Frontend.scala 144:22]
  assign ftq_io_fromBackend_redirect_bits_cfiUpdate_pc = io_backend_toFtq_redirect_bits_cfiUpdate_pc; // @[Frontend.scala 144:22]
  assign ftq_io_fromBackend_redirect_bits_cfiUpdate_pd_isRVC = io_backend_toFtq_redirect_bits_cfiUpdate_pd_isRVC; // @[Frontend.scala 144:22]
  assign ftq_io_fromBackend_redirect_bits_cfiUpdate_pd_brType = io_backend_toFtq_redirect_bits_cfiUpdate_pd_brType; // @[Frontend.scala 144:22]
  assign ftq_io_fromBackend_redirect_bits_cfiUpdate_pd_isCall = io_backend_toFtq_redirect_bits_cfiUpdate_pd_isCall; // @[Frontend.scala 144:22]
  assign ftq_io_fromBackend_redirect_bits_cfiUpdate_pd_isRet = io_backend_toFtq_redirect_bits_cfiUpdate_pd_isRet; // @[Frontend.scala 144:22]
  assign ftq_io_fromBackend_redirect_bits_cfiUpdate_target = io_backend_toFtq_redirect_bits_cfiUpdate_target; // @[Frontend.scala 144:22]
  assign ftq_io_fromBackend_redirect_bits_cfiUpdate_taken = io_backend_toFtq_redirect_bits_cfiUpdate_taken; // @[Frontend.scala 144:22]
  assign ftq_io_fromBackend_redirect_bits_cfiUpdate_isMisPred = io_backend_toFtq_redirect_bits_cfiUpdate_isMisPred; // @[Frontend.scala 144:22]
  assign ftq_io_toIfu_req_ready = ifu_io_ftqInter_fromFtq_req_ready & icache_io_fetch_req_ready; // @[Frontend.scala 117:64]
  assign ftq_io_mmioCommitRead_mmioFtqPtr_flag = ifu_io_mmioCommitRead_mmioFtqPtr_flag; // @[Frontend.scala 123:27]
  assign ftq_io_mmioCommitRead_mmioFtqPtr_value = ifu_io_mmioCommitRead_mmioFtqPtr_value; // @[Frontend.scala 123:27]
  assign tlbCsr_delay_clock = clock;
  assign tlbCsr_delay_io_in_satp_mode = io_tlbCsr_satp_mode; // @[Hold.scala 98:17]
  assign tlbCsr_delay_io_in_satp_asid = io_tlbCsr_satp_asid; // @[Hold.scala 98:17]
  assign tlbCsr_delay_io_in_satp_ppn = io_tlbCsr_satp_ppn; // @[Hold.scala 98:17]
  assign tlbCsr_delay_io_in_satp_changed = io_tlbCsr_satp_changed; // @[Hold.scala 98:17]
  assign tlbCsr_delay_io_in_priv_mxr = io_tlbCsr_priv_mxr; // @[Hold.scala 98:17]
  assign tlbCsr_delay_io_in_priv_sum = io_tlbCsr_priv_sum; // @[Hold.scala 98:17]
  assign tlbCsr_delay_io_in_priv_imode = io_tlbCsr_priv_imode; // @[Hold.scala 98:17]
  assign tlbCsr_delay_io_in_priv_dmode = io_tlbCsr_priv_dmode; // @[Hold.scala 98:17]
  assign csrCtrl_delay_clock = clock;
  assign csrCtrl_delay_io_in_icache_parity_enable = io_csrCtrl_icache_parity_enable; // @[Hold.scala 98:17]
  assign csrCtrl_delay_io_in_lvpred_disable = io_csrCtrl_lvpred_disable; // @[Hold.scala 98:17]
  assign csrCtrl_delay_io_in_no_spec_load = io_csrCtrl_no_spec_load; // @[Hold.scala 98:17]
  assign csrCtrl_delay_io_in_storeset_wait_store = io_csrCtrl_storeset_wait_store; // @[Hold.scala 98:17]
  assign csrCtrl_delay_io_in_lvpred_timeout = io_csrCtrl_lvpred_timeout; // @[Hold.scala 98:17]
  assign csrCtrl_delay_io_in_bp_ctrl_ubtb_enable = io_csrCtrl_bp_ctrl_ubtb_enable; // @[Hold.scala 98:17]
  assign csrCtrl_delay_io_in_bp_ctrl_btb_enable = io_csrCtrl_bp_ctrl_btb_enable; // @[Hold.scala 98:17]
  assign csrCtrl_delay_io_in_bp_ctrl_tage_enable = io_csrCtrl_bp_ctrl_tage_enable; // @[Hold.scala 98:17]
  assign csrCtrl_delay_io_in_bp_ctrl_sc_enable = io_csrCtrl_bp_ctrl_sc_enable; // @[Hold.scala 98:17]
  assign csrCtrl_delay_io_in_bp_ctrl_ras_enable = io_csrCtrl_bp_ctrl_ras_enable; // @[Hold.scala 98:17]
  assign csrCtrl_delay_io_in_sbuffer_threshold = io_csrCtrl_sbuffer_threshold; // @[Hold.scala 98:17]
  assign csrCtrl_delay_io_in_ldld_vio_check_enable = io_csrCtrl_ldld_vio_check_enable; // @[Hold.scala 98:17]
  assign csrCtrl_delay_io_in_cache_error_enable = io_csrCtrl_cache_error_enable; // @[Hold.scala 98:17]
  assign csrCtrl_delay_io_in_uncache_write_outstanding_enable = io_csrCtrl_uncache_write_outstanding_enable; // @[Hold.scala 98:17]
  assign csrCtrl_delay_io_in_fusion_enable = io_csrCtrl_fusion_enable; // @[Hold.scala 98:17]
  assign csrCtrl_delay_io_in_wfi_enable = io_csrCtrl_wfi_enable; // @[Hold.scala 98:17]
  assign csrCtrl_delay_io_in_svinval_enable = io_csrCtrl_svinval_enable; // @[Hold.scala 98:17]
  assign csrCtrl_delay_io_in_distribute_csr_wvalid = io_csrCtrl_distribute_csr_wvalid; // @[Hold.scala 98:17]
  assign csrCtrl_delay_io_in_distribute_csr_waddr = io_csrCtrl_distribute_csr_waddr; // @[Hold.scala 98:17]
  assign csrCtrl_delay_io_in_distribute_csr_wdata = io_csrCtrl_distribute_csr_wdata; // @[Hold.scala 98:17]
  assign csrCtrl_delay_io_in_singlestep = io_csrCtrl_singlestep; // @[Hold.scala 98:17]
  assign csrCtrl_delay_io_in_frontend_trigger_t_valid = io_csrCtrl_frontend_trigger_t_valid; // @[Hold.scala 98:17]
  assign csrCtrl_delay_io_in_frontend_trigger_t_bits_addr = io_csrCtrl_frontend_trigger_t_bits_addr; // @[Hold.scala 98:17]
  assign csrCtrl_delay_io_in_frontend_trigger_t_bits_tdata_matchType =
    io_csrCtrl_frontend_trigger_t_bits_tdata_matchType; // @[Hold.scala 98:17]
  assign csrCtrl_delay_io_in_frontend_trigger_t_bits_tdata_select = io_csrCtrl_frontend_trigger_t_bits_tdata_select; // @[Hold.scala 98:17]
  assign csrCtrl_delay_io_in_frontend_trigger_t_bits_tdata_timing = io_csrCtrl_frontend_trigger_t_bits_tdata_timing; // @[Hold.scala 98:17]
  assign csrCtrl_delay_io_in_frontend_trigger_t_bits_tdata_chain = io_csrCtrl_frontend_trigger_t_bits_tdata_chain; // @[Hold.scala 98:17]
  assign csrCtrl_delay_io_in_frontend_trigger_t_bits_tdata_tdata2 = io_csrCtrl_frontend_trigger_t_bits_tdata_tdata2; // @[Hold.scala 98:17]
  assign csrCtrl_delay_io_in_mem_trigger_t_valid = io_csrCtrl_mem_trigger_t_valid; // @[Hold.scala 98:17]
  assign csrCtrl_delay_io_in_mem_trigger_t_bits_addr = io_csrCtrl_mem_trigger_t_bits_addr; // @[Hold.scala 98:17]
  assign csrCtrl_delay_io_in_mem_trigger_t_bits_tdata_matchType = io_csrCtrl_mem_trigger_t_bits_tdata_matchType; // @[Hold.scala 98:17]
  assign csrCtrl_delay_io_in_mem_trigger_t_bits_tdata_select = io_csrCtrl_mem_trigger_t_bits_tdata_select; // @[Hold.scala 98:17]
  assign csrCtrl_delay_io_in_mem_trigger_t_bits_tdata_chain = io_csrCtrl_mem_trigger_t_bits_tdata_chain; // @[Hold.scala 98:17]
  assign csrCtrl_delay_io_in_mem_trigger_t_bits_tdata_tdata2 = io_csrCtrl_mem_trigger_t_bits_tdata_tdata2; // @[Hold.scala 98:17]
  assign csrCtrl_delay_io_in_trigger_enable_0 = io_csrCtrl_trigger_enable_0; // @[Hold.scala 98:17]
  assign csrCtrl_delay_io_in_trigger_enable_1 = io_csrCtrl_trigger_enable_1; // @[Hold.scala 98:17]
  assign csrCtrl_delay_io_in_trigger_enable_2 = io_csrCtrl_trigger_enable_2; // @[Hold.scala 98:17]
  assign csrCtrl_delay_io_in_trigger_enable_3 = io_csrCtrl_trigger_enable_3; // @[Hold.scala 98:17]
  assign csrCtrl_delay_io_in_trigger_enable_4 = io_csrCtrl_trigger_enable_4; // @[Hold.scala 98:17]
  assign csrCtrl_delay_io_in_trigger_enable_5 = io_csrCtrl_trigger_enable_5; // @[Hold.scala 98:17]
  assign csrCtrl_delay_io_in_trigger_enable_6 = io_csrCtrl_trigger_enable_6; // @[Hold.scala 98:17]
  assign csrCtrl_delay_io_in_trigger_enable_7 = io_csrCtrl_trigger_enable_7; // @[Hold.scala 98:17]
  assign csrCtrl_delay_io_in_trigger_enable_8 = io_csrCtrl_trigger_enable_8; // @[Hold.scala 98:17]
  assign csrCtrl_delay_io_in_trigger_enable_9 = io_csrCtrl_trigger_enable_9; // @[Hold.scala 98:17]
  assign pmp_clock = clock;
  assign pmp_reset = reset;
  assign pmp_io_distribute_csr_wvalid = csrCtrl_delay_io_out_distribute_csr_wvalid; // @[Frontend.scala 89:25]
  assign pmp_io_distribute_csr_waddr = csrCtrl_delay_io_out_distribute_csr_waddr; // @[Frontend.scala 89:25]
  assign pmp_io_distribute_csr_wdata = csrCtrl_delay_io_out_distribute_csr_wdata; // @[Frontend.scala 89:25]
  assign PMPChecker_io_check_env_mode = tlbCsr_delay_io_out_priv_imode; // @[Frontend.scala 88:26 PMP.scala 465:15]
  assign PMPChecker_io_check_env_pmp_0_cfg_l = pmp_io_pmp_0_cfg_l; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_0_cfg_a = pmp_io_pmp_0_cfg_a; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_0_cfg_x = pmp_io_pmp_0_cfg_x; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_0_cfg_w = pmp_io_pmp_0_cfg_w; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_0_cfg_r = pmp_io_pmp_0_cfg_r; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_0_addr = pmp_io_pmp_0_addr; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_0_mask = pmp_io_pmp_0_mask; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_1_cfg_l = pmp_io_pmp_1_cfg_l; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_1_cfg_a = pmp_io_pmp_1_cfg_a; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_1_cfg_x = pmp_io_pmp_1_cfg_x; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_1_cfg_w = pmp_io_pmp_1_cfg_w; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_1_cfg_r = pmp_io_pmp_1_cfg_r; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_1_addr = pmp_io_pmp_1_addr; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_1_mask = pmp_io_pmp_1_mask; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_2_cfg_l = pmp_io_pmp_2_cfg_l; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_2_cfg_a = pmp_io_pmp_2_cfg_a; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_2_cfg_x = pmp_io_pmp_2_cfg_x; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_2_cfg_w = pmp_io_pmp_2_cfg_w; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_2_cfg_r = pmp_io_pmp_2_cfg_r; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_2_addr = pmp_io_pmp_2_addr; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_2_mask = pmp_io_pmp_2_mask; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_3_cfg_l = pmp_io_pmp_3_cfg_l; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_3_cfg_a = pmp_io_pmp_3_cfg_a; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_3_cfg_x = pmp_io_pmp_3_cfg_x; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_3_cfg_w = pmp_io_pmp_3_cfg_w; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_3_cfg_r = pmp_io_pmp_3_cfg_r; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_3_addr = pmp_io_pmp_3_addr; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_3_mask = pmp_io_pmp_3_mask; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_4_cfg_l = pmp_io_pmp_4_cfg_l; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_4_cfg_a = pmp_io_pmp_4_cfg_a; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_4_cfg_x = pmp_io_pmp_4_cfg_x; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_4_cfg_w = pmp_io_pmp_4_cfg_w; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_4_cfg_r = pmp_io_pmp_4_cfg_r; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_4_addr = pmp_io_pmp_4_addr; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_4_mask = pmp_io_pmp_4_mask; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_5_cfg_l = pmp_io_pmp_5_cfg_l; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_5_cfg_a = pmp_io_pmp_5_cfg_a; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_5_cfg_x = pmp_io_pmp_5_cfg_x; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_5_cfg_w = pmp_io_pmp_5_cfg_w; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_5_cfg_r = pmp_io_pmp_5_cfg_r; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_5_addr = pmp_io_pmp_5_addr; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_5_mask = pmp_io_pmp_5_mask; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_6_cfg_l = pmp_io_pmp_6_cfg_l; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_6_cfg_a = pmp_io_pmp_6_cfg_a; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_6_cfg_x = pmp_io_pmp_6_cfg_x; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_6_cfg_w = pmp_io_pmp_6_cfg_w; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_6_cfg_r = pmp_io_pmp_6_cfg_r; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_6_addr = pmp_io_pmp_6_addr; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_6_mask = pmp_io_pmp_6_mask; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_7_cfg_l = pmp_io_pmp_7_cfg_l; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_7_cfg_a = pmp_io_pmp_7_cfg_a; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_7_cfg_x = pmp_io_pmp_7_cfg_x; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_7_cfg_w = pmp_io_pmp_7_cfg_w; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_7_cfg_r = pmp_io_pmp_7_cfg_r; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_7_addr = pmp_io_pmp_7_addr; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_7_mask = pmp_io_pmp_7_mask; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_8_cfg_l = pmp_io_pmp_8_cfg_l; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_8_cfg_a = pmp_io_pmp_8_cfg_a; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_8_cfg_x = pmp_io_pmp_8_cfg_x; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_8_cfg_w = pmp_io_pmp_8_cfg_w; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_8_cfg_r = pmp_io_pmp_8_cfg_r; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_8_addr = pmp_io_pmp_8_addr; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_8_mask = pmp_io_pmp_8_mask; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_9_cfg_l = pmp_io_pmp_9_cfg_l; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_9_cfg_a = pmp_io_pmp_9_cfg_a; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_9_cfg_x = pmp_io_pmp_9_cfg_x; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_9_cfg_w = pmp_io_pmp_9_cfg_w; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_9_cfg_r = pmp_io_pmp_9_cfg_r; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_9_addr = pmp_io_pmp_9_addr; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_9_mask = pmp_io_pmp_9_mask; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_10_cfg_l = pmp_io_pmp_10_cfg_l; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_10_cfg_a = pmp_io_pmp_10_cfg_a; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_10_cfg_x = pmp_io_pmp_10_cfg_x; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_10_cfg_w = pmp_io_pmp_10_cfg_w; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_10_cfg_r = pmp_io_pmp_10_cfg_r; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_10_addr = pmp_io_pmp_10_addr; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_10_mask = pmp_io_pmp_10_mask; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_11_cfg_l = pmp_io_pmp_11_cfg_l; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_11_cfg_a = pmp_io_pmp_11_cfg_a; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_11_cfg_x = pmp_io_pmp_11_cfg_x; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_11_cfg_w = pmp_io_pmp_11_cfg_w; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_11_cfg_r = pmp_io_pmp_11_cfg_r; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_11_addr = pmp_io_pmp_11_addr; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_11_mask = pmp_io_pmp_11_mask; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_12_cfg_l = pmp_io_pmp_12_cfg_l; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_12_cfg_a = pmp_io_pmp_12_cfg_a; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_12_cfg_x = pmp_io_pmp_12_cfg_x; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_12_cfg_w = pmp_io_pmp_12_cfg_w; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_12_cfg_r = pmp_io_pmp_12_cfg_r; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_12_addr = pmp_io_pmp_12_addr; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_12_mask = pmp_io_pmp_12_mask; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_13_cfg_l = pmp_io_pmp_13_cfg_l; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_13_cfg_a = pmp_io_pmp_13_cfg_a; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_13_cfg_x = pmp_io_pmp_13_cfg_x; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_13_cfg_w = pmp_io_pmp_13_cfg_w; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_13_cfg_r = pmp_io_pmp_13_cfg_r; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_13_addr = pmp_io_pmp_13_addr; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_13_mask = pmp_io_pmp_13_mask; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_14_cfg_l = pmp_io_pmp_14_cfg_l; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_14_cfg_a = pmp_io_pmp_14_cfg_a; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_14_cfg_x = pmp_io_pmp_14_cfg_x; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_14_cfg_w = pmp_io_pmp_14_cfg_w; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_14_cfg_r = pmp_io_pmp_14_cfg_r; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_14_addr = pmp_io_pmp_14_addr; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_14_mask = pmp_io_pmp_14_mask; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_15_cfg_l = pmp_io_pmp_15_cfg_l; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_15_cfg_a = pmp_io_pmp_15_cfg_a; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_15_cfg_x = pmp_io_pmp_15_cfg_x; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_15_cfg_w = pmp_io_pmp_15_cfg_w; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_15_cfg_r = pmp_io_pmp_15_cfg_r; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_15_addr = pmp_io_pmp_15_addr; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_15_mask = pmp_io_pmp_15_mask; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pma_0_cfg_c = pmp_io_pma_0_cfg_c; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_0_cfg_atomic = pmp_io_pma_0_cfg_atomic; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_0_cfg_a = pmp_io_pma_0_cfg_a; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_0_cfg_x = pmp_io_pma_0_cfg_x; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_0_cfg_w = pmp_io_pma_0_cfg_w; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_0_cfg_r = pmp_io_pma_0_cfg_r; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_0_addr = pmp_io_pma_0_addr; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_0_mask = pmp_io_pma_0_mask; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_1_cfg_c = pmp_io_pma_1_cfg_c; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_1_cfg_atomic = pmp_io_pma_1_cfg_atomic; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_1_cfg_a = pmp_io_pma_1_cfg_a; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_1_cfg_x = pmp_io_pma_1_cfg_x; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_1_cfg_w = pmp_io_pma_1_cfg_w; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_1_cfg_r = pmp_io_pma_1_cfg_r; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_1_addr = pmp_io_pma_1_addr; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_1_mask = pmp_io_pma_1_mask; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_2_cfg_c = pmp_io_pma_2_cfg_c; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_2_cfg_atomic = pmp_io_pma_2_cfg_atomic; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_2_cfg_a = pmp_io_pma_2_cfg_a; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_2_cfg_x = pmp_io_pma_2_cfg_x; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_2_cfg_w = pmp_io_pma_2_cfg_w; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_2_cfg_r = pmp_io_pma_2_cfg_r; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_2_addr = pmp_io_pma_2_addr; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_2_mask = pmp_io_pma_2_mask; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_3_cfg_c = pmp_io_pma_3_cfg_c; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_3_cfg_atomic = pmp_io_pma_3_cfg_atomic; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_3_cfg_a = pmp_io_pma_3_cfg_a; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_3_cfg_x = pmp_io_pma_3_cfg_x; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_3_cfg_w = pmp_io_pma_3_cfg_w; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_3_cfg_r = pmp_io_pma_3_cfg_r; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_3_addr = pmp_io_pma_3_addr; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_3_mask = pmp_io_pma_3_mask; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_4_cfg_c = pmp_io_pma_4_cfg_c; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_4_cfg_atomic = pmp_io_pma_4_cfg_atomic; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_4_cfg_a = pmp_io_pma_4_cfg_a; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_4_cfg_x = pmp_io_pma_4_cfg_x; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_4_cfg_w = pmp_io_pma_4_cfg_w; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_4_cfg_r = pmp_io_pma_4_cfg_r; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_4_addr = pmp_io_pma_4_addr; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_4_mask = pmp_io_pma_4_mask; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_5_cfg_c = pmp_io_pma_5_cfg_c; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_5_cfg_atomic = pmp_io_pma_5_cfg_atomic; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_5_cfg_a = pmp_io_pma_5_cfg_a; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_5_cfg_x = pmp_io_pma_5_cfg_x; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_5_cfg_w = pmp_io_pma_5_cfg_w; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_5_cfg_r = pmp_io_pma_5_cfg_r; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_5_addr = pmp_io_pma_5_addr; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_5_mask = pmp_io_pma_5_mask; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_6_cfg_c = pmp_io_pma_6_cfg_c; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_6_cfg_atomic = pmp_io_pma_6_cfg_atomic; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_6_cfg_a = pmp_io_pma_6_cfg_a; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_6_cfg_x = pmp_io_pma_6_cfg_x; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_6_cfg_w = pmp_io_pma_6_cfg_w; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_6_cfg_r = pmp_io_pma_6_cfg_r; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_6_addr = pmp_io_pma_6_addr; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_6_mask = pmp_io_pma_6_mask; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_7_cfg_c = pmp_io_pma_7_cfg_c; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_7_cfg_atomic = pmp_io_pma_7_cfg_atomic; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_7_cfg_a = pmp_io_pma_7_cfg_a; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_7_cfg_x = pmp_io_pma_7_cfg_x; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_7_cfg_w = pmp_io_pma_7_cfg_w; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_7_cfg_r = pmp_io_pma_7_cfg_r; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_7_addr = pmp_io_pma_7_addr; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_7_mask = pmp_io_pma_7_mask; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_8_cfg_c = pmp_io_pma_8_cfg_c; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_8_cfg_atomic = pmp_io_pma_8_cfg_atomic; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_8_cfg_a = pmp_io_pma_8_cfg_a; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_8_cfg_x = pmp_io_pma_8_cfg_x; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_8_cfg_w = pmp_io_pma_8_cfg_w; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_8_cfg_r = pmp_io_pma_8_cfg_r; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_8_addr = pmp_io_pma_8_addr; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_8_mask = pmp_io_pma_8_mask; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_9_cfg_c = pmp_io_pma_9_cfg_c; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_9_cfg_atomic = pmp_io_pma_9_cfg_atomic; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_9_cfg_a = pmp_io_pma_9_cfg_a; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_9_cfg_x = pmp_io_pma_9_cfg_x; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_9_cfg_w = pmp_io_pma_9_cfg_w; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_9_cfg_r = pmp_io_pma_9_cfg_r; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_9_addr = pmp_io_pma_9_addr; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_9_mask = pmp_io_pma_9_mask; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_10_cfg_c = pmp_io_pma_10_cfg_c; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_10_cfg_atomic = pmp_io_pma_10_cfg_atomic; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_10_cfg_a = pmp_io_pma_10_cfg_a; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_10_cfg_x = pmp_io_pma_10_cfg_x; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_10_cfg_w = pmp_io_pma_10_cfg_w; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_10_cfg_r = pmp_io_pma_10_cfg_r; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_10_addr = pmp_io_pma_10_addr; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_10_mask = pmp_io_pma_10_mask; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_11_cfg_c = pmp_io_pma_11_cfg_c; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_11_cfg_atomic = pmp_io_pma_11_cfg_atomic; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_11_cfg_a = pmp_io_pma_11_cfg_a; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_11_cfg_x = pmp_io_pma_11_cfg_x; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_11_cfg_w = pmp_io_pma_11_cfg_w; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_11_cfg_r = pmp_io_pma_11_cfg_r; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_11_addr = pmp_io_pma_11_addr; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_11_mask = pmp_io_pma_11_mask; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_12_cfg_c = pmp_io_pma_12_cfg_c; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_12_cfg_atomic = pmp_io_pma_12_cfg_atomic; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_12_cfg_a = pmp_io_pma_12_cfg_a; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_12_cfg_x = pmp_io_pma_12_cfg_x; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_12_cfg_w = pmp_io_pma_12_cfg_w; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_12_cfg_r = pmp_io_pma_12_cfg_r; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_12_addr = pmp_io_pma_12_addr; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_12_mask = pmp_io_pma_12_mask; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_13_cfg_c = pmp_io_pma_13_cfg_c; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_13_cfg_atomic = pmp_io_pma_13_cfg_atomic; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_13_cfg_a = pmp_io_pma_13_cfg_a; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_13_cfg_x = pmp_io_pma_13_cfg_x; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_13_cfg_w = pmp_io_pma_13_cfg_w; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_13_cfg_r = pmp_io_pma_13_cfg_r; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_13_addr = pmp_io_pma_13_addr; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_13_mask = pmp_io_pma_13_mask; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_14_cfg_c = pmp_io_pma_14_cfg_c; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_14_cfg_atomic = pmp_io_pma_14_cfg_atomic; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_14_cfg_a = pmp_io_pma_14_cfg_a; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_14_cfg_x = pmp_io_pma_14_cfg_x; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_14_cfg_w = pmp_io_pma_14_cfg_w; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_14_cfg_r = pmp_io_pma_14_cfg_r; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_14_addr = pmp_io_pma_14_addr; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_14_mask = pmp_io_pma_14_mask; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_15_cfg_c = pmp_io_pma_15_cfg_c; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_15_cfg_atomic = pmp_io_pma_15_cfg_atomic; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_15_cfg_a = pmp_io_pma_15_cfg_a; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_15_cfg_x = pmp_io_pma_15_cfg_x; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_15_cfg_w = pmp_io_pma_15_cfg_w; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_15_cfg_r = pmp_io_pma_15_cfg_r; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_15_addr = pmp_io_pma_15_addr; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_15_mask = pmp_io_pma_15_mask; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_io_req_bits_addr = icache_io_pmp_0_req_bits_addr; // @[Frontend.scala 90:29 91:18]
  assign PMPChecker_io_req_bits_cmd = 3'h2; // @[Frontend.scala 90:29 91:18]
  assign PMPChecker_1_io_check_env_mode = tlbCsr_delay_io_out_priv_imode; // @[Frontend.scala 88:26 PMP.scala 465:15]
  assign PMPChecker_1_io_check_env_pmp_0_cfg_l = pmp_io_pmp_0_cfg_l; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_0_cfg_a = pmp_io_pmp_0_cfg_a; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_0_cfg_x = pmp_io_pmp_0_cfg_x; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_0_cfg_w = pmp_io_pmp_0_cfg_w; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_0_cfg_r = pmp_io_pmp_0_cfg_r; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_0_addr = pmp_io_pmp_0_addr; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_0_mask = pmp_io_pmp_0_mask; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_1_cfg_l = pmp_io_pmp_1_cfg_l; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_1_cfg_a = pmp_io_pmp_1_cfg_a; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_1_cfg_x = pmp_io_pmp_1_cfg_x; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_1_cfg_w = pmp_io_pmp_1_cfg_w; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_1_cfg_r = pmp_io_pmp_1_cfg_r; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_1_addr = pmp_io_pmp_1_addr; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_1_mask = pmp_io_pmp_1_mask; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_2_cfg_l = pmp_io_pmp_2_cfg_l; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_2_cfg_a = pmp_io_pmp_2_cfg_a; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_2_cfg_x = pmp_io_pmp_2_cfg_x; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_2_cfg_w = pmp_io_pmp_2_cfg_w; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_2_cfg_r = pmp_io_pmp_2_cfg_r; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_2_addr = pmp_io_pmp_2_addr; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_2_mask = pmp_io_pmp_2_mask; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_3_cfg_l = pmp_io_pmp_3_cfg_l; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_3_cfg_a = pmp_io_pmp_3_cfg_a; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_3_cfg_x = pmp_io_pmp_3_cfg_x; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_3_cfg_w = pmp_io_pmp_3_cfg_w; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_3_cfg_r = pmp_io_pmp_3_cfg_r; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_3_addr = pmp_io_pmp_3_addr; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_3_mask = pmp_io_pmp_3_mask; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_4_cfg_l = pmp_io_pmp_4_cfg_l; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_4_cfg_a = pmp_io_pmp_4_cfg_a; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_4_cfg_x = pmp_io_pmp_4_cfg_x; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_4_cfg_w = pmp_io_pmp_4_cfg_w; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_4_cfg_r = pmp_io_pmp_4_cfg_r; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_4_addr = pmp_io_pmp_4_addr; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_4_mask = pmp_io_pmp_4_mask; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_5_cfg_l = pmp_io_pmp_5_cfg_l; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_5_cfg_a = pmp_io_pmp_5_cfg_a; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_5_cfg_x = pmp_io_pmp_5_cfg_x; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_5_cfg_w = pmp_io_pmp_5_cfg_w; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_5_cfg_r = pmp_io_pmp_5_cfg_r; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_5_addr = pmp_io_pmp_5_addr; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_5_mask = pmp_io_pmp_5_mask; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_6_cfg_l = pmp_io_pmp_6_cfg_l; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_6_cfg_a = pmp_io_pmp_6_cfg_a; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_6_cfg_x = pmp_io_pmp_6_cfg_x; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_6_cfg_w = pmp_io_pmp_6_cfg_w; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_6_cfg_r = pmp_io_pmp_6_cfg_r; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_6_addr = pmp_io_pmp_6_addr; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_6_mask = pmp_io_pmp_6_mask; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_7_cfg_l = pmp_io_pmp_7_cfg_l; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_7_cfg_a = pmp_io_pmp_7_cfg_a; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_7_cfg_x = pmp_io_pmp_7_cfg_x; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_7_cfg_w = pmp_io_pmp_7_cfg_w; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_7_cfg_r = pmp_io_pmp_7_cfg_r; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_7_addr = pmp_io_pmp_7_addr; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_7_mask = pmp_io_pmp_7_mask; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_8_cfg_l = pmp_io_pmp_8_cfg_l; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_8_cfg_a = pmp_io_pmp_8_cfg_a; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_8_cfg_x = pmp_io_pmp_8_cfg_x; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_8_cfg_w = pmp_io_pmp_8_cfg_w; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_8_cfg_r = pmp_io_pmp_8_cfg_r; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_8_addr = pmp_io_pmp_8_addr; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_8_mask = pmp_io_pmp_8_mask; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_9_cfg_l = pmp_io_pmp_9_cfg_l; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_9_cfg_a = pmp_io_pmp_9_cfg_a; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_9_cfg_x = pmp_io_pmp_9_cfg_x; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_9_cfg_w = pmp_io_pmp_9_cfg_w; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_9_cfg_r = pmp_io_pmp_9_cfg_r; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_9_addr = pmp_io_pmp_9_addr; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_9_mask = pmp_io_pmp_9_mask; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_10_cfg_l = pmp_io_pmp_10_cfg_l; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_10_cfg_a = pmp_io_pmp_10_cfg_a; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_10_cfg_x = pmp_io_pmp_10_cfg_x; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_10_cfg_w = pmp_io_pmp_10_cfg_w; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_10_cfg_r = pmp_io_pmp_10_cfg_r; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_10_addr = pmp_io_pmp_10_addr; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_10_mask = pmp_io_pmp_10_mask; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_11_cfg_l = pmp_io_pmp_11_cfg_l; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_11_cfg_a = pmp_io_pmp_11_cfg_a; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_11_cfg_x = pmp_io_pmp_11_cfg_x; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_11_cfg_w = pmp_io_pmp_11_cfg_w; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_11_cfg_r = pmp_io_pmp_11_cfg_r; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_11_addr = pmp_io_pmp_11_addr; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_11_mask = pmp_io_pmp_11_mask; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_12_cfg_l = pmp_io_pmp_12_cfg_l; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_12_cfg_a = pmp_io_pmp_12_cfg_a; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_12_cfg_x = pmp_io_pmp_12_cfg_x; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_12_cfg_w = pmp_io_pmp_12_cfg_w; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_12_cfg_r = pmp_io_pmp_12_cfg_r; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_12_addr = pmp_io_pmp_12_addr; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_12_mask = pmp_io_pmp_12_mask; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_13_cfg_l = pmp_io_pmp_13_cfg_l; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_13_cfg_a = pmp_io_pmp_13_cfg_a; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_13_cfg_x = pmp_io_pmp_13_cfg_x; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_13_cfg_w = pmp_io_pmp_13_cfg_w; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_13_cfg_r = pmp_io_pmp_13_cfg_r; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_13_addr = pmp_io_pmp_13_addr; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_13_mask = pmp_io_pmp_13_mask; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_14_cfg_l = pmp_io_pmp_14_cfg_l; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_14_cfg_a = pmp_io_pmp_14_cfg_a; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_14_cfg_x = pmp_io_pmp_14_cfg_x; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_14_cfg_w = pmp_io_pmp_14_cfg_w; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_14_cfg_r = pmp_io_pmp_14_cfg_r; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_14_addr = pmp_io_pmp_14_addr; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_14_mask = pmp_io_pmp_14_mask; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_15_cfg_l = pmp_io_pmp_15_cfg_l; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_15_cfg_a = pmp_io_pmp_15_cfg_a; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_15_cfg_x = pmp_io_pmp_15_cfg_x; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_15_cfg_w = pmp_io_pmp_15_cfg_w; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_15_cfg_r = pmp_io_pmp_15_cfg_r; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_15_addr = pmp_io_pmp_15_addr; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_15_mask = pmp_io_pmp_15_mask; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pma_0_cfg_c = pmp_io_pma_0_cfg_c; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_0_cfg_atomic = pmp_io_pma_0_cfg_atomic; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_0_cfg_a = pmp_io_pma_0_cfg_a; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_0_cfg_x = pmp_io_pma_0_cfg_x; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_0_cfg_w = pmp_io_pma_0_cfg_w; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_0_cfg_r = pmp_io_pma_0_cfg_r; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_0_addr = pmp_io_pma_0_addr; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_0_mask = pmp_io_pma_0_mask; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_1_cfg_c = pmp_io_pma_1_cfg_c; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_1_cfg_atomic = pmp_io_pma_1_cfg_atomic; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_1_cfg_a = pmp_io_pma_1_cfg_a; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_1_cfg_x = pmp_io_pma_1_cfg_x; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_1_cfg_w = pmp_io_pma_1_cfg_w; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_1_cfg_r = pmp_io_pma_1_cfg_r; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_1_addr = pmp_io_pma_1_addr; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_1_mask = pmp_io_pma_1_mask; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_2_cfg_c = pmp_io_pma_2_cfg_c; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_2_cfg_atomic = pmp_io_pma_2_cfg_atomic; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_2_cfg_a = pmp_io_pma_2_cfg_a; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_2_cfg_x = pmp_io_pma_2_cfg_x; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_2_cfg_w = pmp_io_pma_2_cfg_w; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_2_cfg_r = pmp_io_pma_2_cfg_r; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_2_addr = pmp_io_pma_2_addr; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_2_mask = pmp_io_pma_2_mask; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_3_cfg_c = pmp_io_pma_3_cfg_c; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_3_cfg_atomic = pmp_io_pma_3_cfg_atomic; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_3_cfg_a = pmp_io_pma_3_cfg_a; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_3_cfg_x = pmp_io_pma_3_cfg_x; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_3_cfg_w = pmp_io_pma_3_cfg_w; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_3_cfg_r = pmp_io_pma_3_cfg_r; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_3_addr = pmp_io_pma_3_addr; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_3_mask = pmp_io_pma_3_mask; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_4_cfg_c = pmp_io_pma_4_cfg_c; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_4_cfg_atomic = pmp_io_pma_4_cfg_atomic; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_4_cfg_a = pmp_io_pma_4_cfg_a; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_4_cfg_x = pmp_io_pma_4_cfg_x; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_4_cfg_w = pmp_io_pma_4_cfg_w; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_4_cfg_r = pmp_io_pma_4_cfg_r; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_4_addr = pmp_io_pma_4_addr; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_4_mask = pmp_io_pma_4_mask; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_5_cfg_c = pmp_io_pma_5_cfg_c; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_5_cfg_atomic = pmp_io_pma_5_cfg_atomic; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_5_cfg_a = pmp_io_pma_5_cfg_a; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_5_cfg_x = pmp_io_pma_5_cfg_x; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_5_cfg_w = pmp_io_pma_5_cfg_w; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_5_cfg_r = pmp_io_pma_5_cfg_r; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_5_addr = pmp_io_pma_5_addr; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_5_mask = pmp_io_pma_5_mask; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_6_cfg_c = pmp_io_pma_6_cfg_c; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_6_cfg_atomic = pmp_io_pma_6_cfg_atomic; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_6_cfg_a = pmp_io_pma_6_cfg_a; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_6_cfg_x = pmp_io_pma_6_cfg_x; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_6_cfg_w = pmp_io_pma_6_cfg_w; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_6_cfg_r = pmp_io_pma_6_cfg_r; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_6_addr = pmp_io_pma_6_addr; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_6_mask = pmp_io_pma_6_mask; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_7_cfg_c = pmp_io_pma_7_cfg_c; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_7_cfg_atomic = pmp_io_pma_7_cfg_atomic; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_7_cfg_a = pmp_io_pma_7_cfg_a; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_7_cfg_x = pmp_io_pma_7_cfg_x; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_7_cfg_w = pmp_io_pma_7_cfg_w; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_7_cfg_r = pmp_io_pma_7_cfg_r; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_7_addr = pmp_io_pma_7_addr; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_7_mask = pmp_io_pma_7_mask; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_8_cfg_c = pmp_io_pma_8_cfg_c; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_8_cfg_atomic = pmp_io_pma_8_cfg_atomic; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_8_cfg_a = pmp_io_pma_8_cfg_a; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_8_cfg_x = pmp_io_pma_8_cfg_x; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_8_cfg_w = pmp_io_pma_8_cfg_w; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_8_cfg_r = pmp_io_pma_8_cfg_r; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_8_addr = pmp_io_pma_8_addr; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_8_mask = pmp_io_pma_8_mask; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_9_cfg_c = pmp_io_pma_9_cfg_c; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_9_cfg_atomic = pmp_io_pma_9_cfg_atomic; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_9_cfg_a = pmp_io_pma_9_cfg_a; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_9_cfg_x = pmp_io_pma_9_cfg_x; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_9_cfg_w = pmp_io_pma_9_cfg_w; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_9_cfg_r = pmp_io_pma_9_cfg_r; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_9_addr = pmp_io_pma_9_addr; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_9_mask = pmp_io_pma_9_mask; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_10_cfg_c = pmp_io_pma_10_cfg_c; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_10_cfg_atomic = pmp_io_pma_10_cfg_atomic; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_10_cfg_a = pmp_io_pma_10_cfg_a; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_10_cfg_x = pmp_io_pma_10_cfg_x; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_10_cfg_w = pmp_io_pma_10_cfg_w; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_10_cfg_r = pmp_io_pma_10_cfg_r; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_10_addr = pmp_io_pma_10_addr; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_10_mask = pmp_io_pma_10_mask; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_11_cfg_c = pmp_io_pma_11_cfg_c; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_11_cfg_atomic = pmp_io_pma_11_cfg_atomic; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_11_cfg_a = pmp_io_pma_11_cfg_a; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_11_cfg_x = pmp_io_pma_11_cfg_x; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_11_cfg_w = pmp_io_pma_11_cfg_w; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_11_cfg_r = pmp_io_pma_11_cfg_r; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_11_addr = pmp_io_pma_11_addr; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_11_mask = pmp_io_pma_11_mask; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_12_cfg_c = pmp_io_pma_12_cfg_c; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_12_cfg_atomic = pmp_io_pma_12_cfg_atomic; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_12_cfg_a = pmp_io_pma_12_cfg_a; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_12_cfg_x = pmp_io_pma_12_cfg_x; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_12_cfg_w = pmp_io_pma_12_cfg_w; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_12_cfg_r = pmp_io_pma_12_cfg_r; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_12_addr = pmp_io_pma_12_addr; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_12_mask = pmp_io_pma_12_mask; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_13_cfg_c = pmp_io_pma_13_cfg_c; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_13_cfg_atomic = pmp_io_pma_13_cfg_atomic; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_13_cfg_a = pmp_io_pma_13_cfg_a; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_13_cfg_x = pmp_io_pma_13_cfg_x; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_13_cfg_w = pmp_io_pma_13_cfg_w; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_13_cfg_r = pmp_io_pma_13_cfg_r; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_13_addr = pmp_io_pma_13_addr; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_13_mask = pmp_io_pma_13_mask; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_14_cfg_c = pmp_io_pma_14_cfg_c; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_14_cfg_atomic = pmp_io_pma_14_cfg_atomic; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_14_cfg_a = pmp_io_pma_14_cfg_a; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_14_cfg_x = pmp_io_pma_14_cfg_x; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_14_cfg_w = pmp_io_pma_14_cfg_w; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_14_cfg_r = pmp_io_pma_14_cfg_r; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_14_addr = pmp_io_pma_14_addr; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_14_mask = pmp_io_pma_14_mask; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_15_cfg_c = pmp_io_pma_15_cfg_c; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_15_cfg_atomic = pmp_io_pma_15_cfg_atomic; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_15_cfg_a = pmp_io_pma_15_cfg_a; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_15_cfg_x = pmp_io_pma_15_cfg_x; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_15_cfg_w = pmp_io_pma_15_cfg_w; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_15_cfg_r = pmp_io_pma_15_cfg_r; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_15_addr = pmp_io_pma_15_addr; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_15_mask = pmp_io_pma_15_mask; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_1_io_req_bits_addr = icache_io_pmp_1_req_bits_addr; // @[Frontend.scala 90:29 92:18]
  assign PMPChecker_1_io_req_bits_cmd = 3'h2; // @[Frontend.scala 90:29 92:18]
  assign PMPChecker_2_io_check_env_mode = tlbCsr_delay_io_out_priv_imode; // @[Frontend.scala 88:26 PMP.scala 465:15]
  assign PMPChecker_2_io_check_env_pmp_0_cfg_l = pmp_io_pmp_0_cfg_l; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_0_cfg_a = pmp_io_pmp_0_cfg_a; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_0_cfg_x = pmp_io_pmp_0_cfg_x; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_0_cfg_w = pmp_io_pmp_0_cfg_w; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_0_cfg_r = pmp_io_pmp_0_cfg_r; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_0_addr = pmp_io_pmp_0_addr; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_0_mask = pmp_io_pmp_0_mask; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_1_cfg_l = pmp_io_pmp_1_cfg_l; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_1_cfg_a = pmp_io_pmp_1_cfg_a; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_1_cfg_x = pmp_io_pmp_1_cfg_x; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_1_cfg_w = pmp_io_pmp_1_cfg_w; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_1_cfg_r = pmp_io_pmp_1_cfg_r; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_1_addr = pmp_io_pmp_1_addr; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_1_mask = pmp_io_pmp_1_mask; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_2_cfg_l = pmp_io_pmp_2_cfg_l; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_2_cfg_a = pmp_io_pmp_2_cfg_a; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_2_cfg_x = pmp_io_pmp_2_cfg_x; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_2_cfg_w = pmp_io_pmp_2_cfg_w; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_2_cfg_r = pmp_io_pmp_2_cfg_r; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_2_addr = pmp_io_pmp_2_addr; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_2_mask = pmp_io_pmp_2_mask; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_3_cfg_l = pmp_io_pmp_3_cfg_l; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_3_cfg_a = pmp_io_pmp_3_cfg_a; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_3_cfg_x = pmp_io_pmp_3_cfg_x; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_3_cfg_w = pmp_io_pmp_3_cfg_w; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_3_cfg_r = pmp_io_pmp_3_cfg_r; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_3_addr = pmp_io_pmp_3_addr; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_3_mask = pmp_io_pmp_3_mask; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_4_cfg_l = pmp_io_pmp_4_cfg_l; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_4_cfg_a = pmp_io_pmp_4_cfg_a; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_4_cfg_x = pmp_io_pmp_4_cfg_x; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_4_cfg_w = pmp_io_pmp_4_cfg_w; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_4_cfg_r = pmp_io_pmp_4_cfg_r; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_4_addr = pmp_io_pmp_4_addr; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_4_mask = pmp_io_pmp_4_mask; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_5_cfg_l = pmp_io_pmp_5_cfg_l; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_5_cfg_a = pmp_io_pmp_5_cfg_a; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_5_cfg_x = pmp_io_pmp_5_cfg_x; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_5_cfg_w = pmp_io_pmp_5_cfg_w; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_5_cfg_r = pmp_io_pmp_5_cfg_r; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_5_addr = pmp_io_pmp_5_addr; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_5_mask = pmp_io_pmp_5_mask; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_6_cfg_l = pmp_io_pmp_6_cfg_l; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_6_cfg_a = pmp_io_pmp_6_cfg_a; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_6_cfg_x = pmp_io_pmp_6_cfg_x; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_6_cfg_w = pmp_io_pmp_6_cfg_w; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_6_cfg_r = pmp_io_pmp_6_cfg_r; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_6_addr = pmp_io_pmp_6_addr; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_6_mask = pmp_io_pmp_6_mask; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_7_cfg_l = pmp_io_pmp_7_cfg_l; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_7_cfg_a = pmp_io_pmp_7_cfg_a; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_7_cfg_x = pmp_io_pmp_7_cfg_x; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_7_cfg_w = pmp_io_pmp_7_cfg_w; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_7_cfg_r = pmp_io_pmp_7_cfg_r; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_7_addr = pmp_io_pmp_7_addr; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_7_mask = pmp_io_pmp_7_mask; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_8_cfg_l = pmp_io_pmp_8_cfg_l; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_8_cfg_a = pmp_io_pmp_8_cfg_a; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_8_cfg_x = pmp_io_pmp_8_cfg_x; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_8_cfg_w = pmp_io_pmp_8_cfg_w; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_8_cfg_r = pmp_io_pmp_8_cfg_r; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_8_addr = pmp_io_pmp_8_addr; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_8_mask = pmp_io_pmp_8_mask; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_9_cfg_l = pmp_io_pmp_9_cfg_l; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_9_cfg_a = pmp_io_pmp_9_cfg_a; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_9_cfg_x = pmp_io_pmp_9_cfg_x; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_9_cfg_w = pmp_io_pmp_9_cfg_w; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_9_cfg_r = pmp_io_pmp_9_cfg_r; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_9_addr = pmp_io_pmp_9_addr; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_9_mask = pmp_io_pmp_9_mask; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_10_cfg_l = pmp_io_pmp_10_cfg_l; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_10_cfg_a = pmp_io_pmp_10_cfg_a; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_10_cfg_x = pmp_io_pmp_10_cfg_x; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_10_cfg_w = pmp_io_pmp_10_cfg_w; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_10_cfg_r = pmp_io_pmp_10_cfg_r; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_10_addr = pmp_io_pmp_10_addr; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_10_mask = pmp_io_pmp_10_mask; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_11_cfg_l = pmp_io_pmp_11_cfg_l; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_11_cfg_a = pmp_io_pmp_11_cfg_a; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_11_cfg_x = pmp_io_pmp_11_cfg_x; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_11_cfg_w = pmp_io_pmp_11_cfg_w; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_11_cfg_r = pmp_io_pmp_11_cfg_r; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_11_addr = pmp_io_pmp_11_addr; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_11_mask = pmp_io_pmp_11_mask; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_12_cfg_l = pmp_io_pmp_12_cfg_l; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_12_cfg_a = pmp_io_pmp_12_cfg_a; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_12_cfg_x = pmp_io_pmp_12_cfg_x; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_12_cfg_w = pmp_io_pmp_12_cfg_w; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_12_cfg_r = pmp_io_pmp_12_cfg_r; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_12_addr = pmp_io_pmp_12_addr; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_12_mask = pmp_io_pmp_12_mask; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_13_cfg_l = pmp_io_pmp_13_cfg_l; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_13_cfg_a = pmp_io_pmp_13_cfg_a; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_13_cfg_x = pmp_io_pmp_13_cfg_x; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_13_cfg_w = pmp_io_pmp_13_cfg_w; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_13_cfg_r = pmp_io_pmp_13_cfg_r; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_13_addr = pmp_io_pmp_13_addr; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_13_mask = pmp_io_pmp_13_mask; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_14_cfg_l = pmp_io_pmp_14_cfg_l; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_14_cfg_a = pmp_io_pmp_14_cfg_a; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_14_cfg_x = pmp_io_pmp_14_cfg_x; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_14_cfg_w = pmp_io_pmp_14_cfg_w; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_14_cfg_r = pmp_io_pmp_14_cfg_r; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_14_addr = pmp_io_pmp_14_addr; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_14_mask = pmp_io_pmp_14_mask; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_15_cfg_l = pmp_io_pmp_15_cfg_l; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_15_cfg_a = pmp_io_pmp_15_cfg_a; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_15_cfg_x = pmp_io_pmp_15_cfg_x; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_15_cfg_w = pmp_io_pmp_15_cfg_w; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_15_cfg_r = pmp_io_pmp_15_cfg_r; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_15_addr = pmp_io_pmp_15_addr; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_15_mask = pmp_io_pmp_15_mask; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pma_0_cfg_c = pmp_io_pma_0_cfg_c; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_0_cfg_atomic = pmp_io_pma_0_cfg_atomic; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_0_cfg_a = pmp_io_pma_0_cfg_a; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_0_cfg_x = pmp_io_pma_0_cfg_x; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_0_cfg_w = pmp_io_pma_0_cfg_w; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_0_cfg_r = pmp_io_pma_0_cfg_r; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_0_addr = pmp_io_pma_0_addr; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_0_mask = pmp_io_pma_0_mask; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_1_cfg_c = pmp_io_pma_1_cfg_c; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_1_cfg_atomic = pmp_io_pma_1_cfg_atomic; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_1_cfg_a = pmp_io_pma_1_cfg_a; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_1_cfg_x = pmp_io_pma_1_cfg_x; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_1_cfg_w = pmp_io_pma_1_cfg_w; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_1_cfg_r = pmp_io_pma_1_cfg_r; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_1_addr = pmp_io_pma_1_addr; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_1_mask = pmp_io_pma_1_mask; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_2_cfg_c = pmp_io_pma_2_cfg_c; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_2_cfg_atomic = pmp_io_pma_2_cfg_atomic; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_2_cfg_a = pmp_io_pma_2_cfg_a; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_2_cfg_x = pmp_io_pma_2_cfg_x; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_2_cfg_w = pmp_io_pma_2_cfg_w; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_2_cfg_r = pmp_io_pma_2_cfg_r; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_2_addr = pmp_io_pma_2_addr; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_2_mask = pmp_io_pma_2_mask; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_3_cfg_c = pmp_io_pma_3_cfg_c; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_3_cfg_atomic = pmp_io_pma_3_cfg_atomic; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_3_cfg_a = pmp_io_pma_3_cfg_a; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_3_cfg_x = pmp_io_pma_3_cfg_x; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_3_cfg_w = pmp_io_pma_3_cfg_w; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_3_cfg_r = pmp_io_pma_3_cfg_r; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_3_addr = pmp_io_pma_3_addr; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_3_mask = pmp_io_pma_3_mask; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_4_cfg_c = pmp_io_pma_4_cfg_c; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_4_cfg_atomic = pmp_io_pma_4_cfg_atomic; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_4_cfg_a = pmp_io_pma_4_cfg_a; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_4_cfg_x = pmp_io_pma_4_cfg_x; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_4_cfg_w = pmp_io_pma_4_cfg_w; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_4_cfg_r = pmp_io_pma_4_cfg_r; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_4_addr = pmp_io_pma_4_addr; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_4_mask = pmp_io_pma_4_mask; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_5_cfg_c = pmp_io_pma_5_cfg_c; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_5_cfg_atomic = pmp_io_pma_5_cfg_atomic; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_5_cfg_a = pmp_io_pma_5_cfg_a; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_5_cfg_x = pmp_io_pma_5_cfg_x; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_5_cfg_w = pmp_io_pma_5_cfg_w; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_5_cfg_r = pmp_io_pma_5_cfg_r; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_5_addr = pmp_io_pma_5_addr; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_5_mask = pmp_io_pma_5_mask; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_6_cfg_c = pmp_io_pma_6_cfg_c; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_6_cfg_atomic = pmp_io_pma_6_cfg_atomic; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_6_cfg_a = pmp_io_pma_6_cfg_a; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_6_cfg_x = pmp_io_pma_6_cfg_x; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_6_cfg_w = pmp_io_pma_6_cfg_w; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_6_cfg_r = pmp_io_pma_6_cfg_r; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_6_addr = pmp_io_pma_6_addr; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_6_mask = pmp_io_pma_6_mask; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_7_cfg_c = pmp_io_pma_7_cfg_c; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_7_cfg_atomic = pmp_io_pma_7_cfg_atomic; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_7_cfg_a = pmp_io_pma_7_cfg_a; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_7_cfg_x = pmp_io_pma_7_cfg_x; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_7_cfg_w = pmp_io_pma_7_cfg_w; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_7_cfg_r = pmp_io_pma_7_cfg_r; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_7_addr = pmp_io_pma_7_addr; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_7_mask = pmp_io_pma_7_mask; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_8_cfg_c = pmp_io_pma_8_cfg_c; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_8_cfg_atomic = pmp_io_pma_8_cfg_atomic; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_8_cfg_a = pmp_io_pma_8_cfg_a; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_8_cfg_x = pmp_io_pma_8_cfg_x; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_8_cfg_w = pmp_io_pma_8_cfg_w; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_8_cfg_r = pmp_io_pma_8_cfg_r; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_8_addr = pmp_io_pma_8_addr; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_8_mask = pmp_io_pma_8_mask; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_9_cfg_c = pmp_io_pma_9_cfg_c; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_9_cfg_atomic = pmp_io_pma_9_cfg_atomic; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_9_cfg_a = pmp_io_pma_9_cfg_a; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_9_cfg_x = pmp_io_pma_9_cfg_x; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_9_cfg_w = pmp_io_pma_9_cfg_w; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_9_cfg_r = pmp_io_pma_9_cfg_r; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_9_addr = pmp_io_pma_9_addr; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_9_mask = pmp_io_pma_9_mask; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_10_cfg_c = pmp_io_pma_10_cfg_c; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_10_cfg_atomic = pmp_io_pma_10_cfg_atomic; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_10_cfg_a = pmp_io_pma_10_cfg_a; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_10_cfg_x = pmp_io_pma_10_cfg_x; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_10_cfg_w = pmp_io_pma_10_cfg_w; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_10_cfg_r = pmp_io_pma_10_cfg_r; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_10_addr = pmp_io_pma_10_addr; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_10_mask = pmp_io_pma_10_mask; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_11_cfg_c = pmp_io_pma_11_cfg_c; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_11_cfg_atomic = pmp_io_pma_11_cfg_atomic; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_11_cfg_a = pmp_io_pma_11_cfg_a; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_11_cfg_x = pmp_io_pma_11_cfg_x; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_11_cfg_w = pmp_io_pma_11_cfg_w; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_11_cfg_r = pmp_io_pma_11_cfg_r; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_11_addr = pmp_io_pma_11_addr; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_11_mask = pmp_io_pma_11_mask; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_12_cfg_c = pmp_io_pma_12_cfg_c; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_12_cfg_atomic = pmp_io_pma_12_cfg_atomic; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_12_cfg_a = pmp_io_pma_12_cfg_a; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_12_cfg_x = pmp_io_pma_12_cfg_x; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_12_cfg_w = pmp_io_pma_12_cfg_w; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_12_cfg_r = pmp_io_pma_12_cfg_r; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_12_addr = pmp_io_pma_12_addr; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_12_mask = pmp_io_pma_12_mask; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_13_cfg_c = pmp_io_pma_13_cfg_c; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_13_cfg_atomic = pmp_io_pma_13_cfg_atomic; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_13_cfg_a = pmp_io_pma_13_cfg_a; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_13_cfg_x = pmp_io_pma_13_cfg_x; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_13_cfg_w = pmp_io_pma_13_cfg_w; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_13_cfg_r = pmp_io_pma_13_cfg_r; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_13_addr = pmp_io_pma_13_addr; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_13_mask = pmp_io_pma_13_mask; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_14_cfg_c = pmp_io_pma_14_cfg_c; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_14_cfg_atomic = pmp_io_pma_14_cfg_atomic; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_14_cfg_a = pmp_io_pma_14_cfg_a; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_14_cfg_x = pmp_io_pma_14_cfg_x; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_14_cfg_w = pmp_io_pma_14_cfg_w; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_14_cfg_r = pmp_io_pma_14_cfg_r; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_14_addr = pmp_io_pma_14_addr; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_14_mask = pmp_io_pma_14_mask; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_15_cfg_c = pmp_io_pma_15_cfg_c; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_15_cfg_atomic = pmp_io_pma_15_cfg_atomic; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_15_cfg_a = pmp_io_pma_15_cfg_a; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_15_cfg_x = pmp_io_pma_15_cfg_x; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_15_cfg_w = pmp_io_pma_15_cfg_w; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_15_cfg_r = pmp_io_pma_15_cfg_r; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_15_addr = pmp_io_pma_15_addr; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_15_mask = pmp_io_pma_15_mask; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_2_io_req_bits_addr = 36'h0; // @[Frontend.scala 90:29 93:18]
  assign PMPChecker_2_io_req_bits_cmd = 3'h2; // @[Frontend.scala 90:29 93:18]
  assign PMPChecker_3_io_check_env_mode = tlbCsr_delay_io_out_priv_imode; // @[Frontend.scala 88:26 PMP.scala 465:15]
  assign PMPChecker_3_io_check_env_pmp_0_cfg_l = pmp_io_pmp_0_cfg_l; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_0_cfg_a = pmp_io_pmp_0_cfg_a; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_0_cfg_x = pmp_io_pmp_0_cfg_x; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_0_cfg_w = pmp_io_pmp_0_cfg_w; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_0_cfg_r = pmp_io_pmp_0_cfg_r; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_0_addr = pmp_io_pmp_0_addr; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_0_mask = pmp_io_pmp_0_mask; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_1_cfg_l = pmp_io_pmp_1_cfg_l; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_1_cfg_a = pmp_io_pmp_1_cfg_a; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_1_cfg_x = pmp_io_pmp_1_cfg_x; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_1_cfg_w = pmp_io_pmp_1_cfg_w; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_1_cfg_r = pmp_io_pmp_1_cfg_r; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_1_addr = pmp_io_pmp_1_addr; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_1_mask = pmp_io_pmp_1_mask; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_2_cfg_l = pmp_io_pmp_2_cfg_l; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_2_cfg_a = pmp_io_pmp_2_cfg_a; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_2_cfg_x = pmp_io_pmp_2_cfg_x; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_2_cfg_w = pmp_io_pmp_2_cfg_w; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_2_cfg_r = pmp_io_pmp_2_cfg_r; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_2_addr = pmp_io_pmp_2_addr; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_2_mask = pmp_io_pmp_2_mask; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_3_cfg_l = pmp_io_pmp_3_cfg_l; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_3_cfg_a = pmp_io_pmp_3_cfg_a; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_3_cfg_x = pmp_io_pmp_3_cfg_x; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_3_cfg_w = pmp_io_pmp_3_cfg_w; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_3_cfg_r = pmp_io_pmp_3_cfg_r; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_3_addr = pmp_io_pmp_3_addr; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_3_mask = pmp_io_pmp_3_mask; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_4_cfg_l = pmp_io_pmp_4_cfg_l; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_4_cfg_a = pmp_io_pmp_4_cfg_a; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_4_cfg_x = pmp_io_pmp_4_cfg_x; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_4_cfg_w = pmp_io_pmp_4_cfg_w; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_4_cfg_r = pmp_io_pmp_4_cfg_r; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_4_addr = pmp_io_pmp_4_addr; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_4_mask = pmp_io_pmp_4_mask; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_5_cfg_l = pmp_io_pmp_5_cfg_l; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_5_cfg_a = pmp_io_pmp_5_cfg_a; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_5_cfg_x = pmp_io_pmp_5_cfg_x; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_5_cfg_w = pmp_io_pmp_5_cfg_w; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_5_cfg_r = pmp_io_pmp_5_cfg_r; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_5_addr = pmp_io_pmp_5_addr; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_5_mask = pmp_io_pmp_5_mask; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_6_cfg_l = pmp_io_pmp_6_cfg_l; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_6_cfg_a = pmp_io_pmp_6_cfg_a; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_6_cfg_x = pmp_io_pmp_6_cfg_x; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_6_cfg_w = pmp_io_pmp_6_cfg_w; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_6_cfg_r = pmp_io_pmp_6_cfg_r; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_6_addr = pmp_io_pmp_6_addr; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_6_mask = pmp_io_pmp_6_mask; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_7_cfg_l = pmp_io_pmp_7_cfg_l; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_7_cfg_a = pmp_io_pmp_7_cfg_a; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_7_cfg_x = pmp_io_pmp_7_cfg_x; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_7_cfg_w = pmp_io_pmp_7_cfg_w; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_7_cfg_r = pmp_io_pmp_7_cfg_r; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_7_addr = pmp_io_pmp_7_addr; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_7_mask = pmp_io_pmp_7_mask; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_8_cfg_l = pmp_io_pmp_8_cfg_l; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_8_cfg_a = pmp_io_pmp_8_cfg_a; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_8_cfg_x = pmp_io_pmp_8_cfg_x; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_8_cfg_w = pmp_io_pmp_8_cfg_w; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_8_cfg_r = pmp_io_pmp_8_cfg_r; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_8_addr = pmp_io_pmp_8_addr; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_8_mask = pmp_io_pmp_8_mask; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_9_cfg_l = pmp_io_pmp_9_cfg_l; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_9_cfg_a = pmp_io_pmp_9_cfg_a; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_9_cfg_x = pmp_io_pmp_9_cfg_x; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_9_cfg_w = pmp_io_pmp_9_cfg_w; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_9_cfg_r = pmp_io_pmp_9_cfg_r; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_9_addr = pmp_io_pmp_9_addr; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_9_mask = pmp_io_pmp_9_mask; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_10_cfg_l = pmp_io_pmp_10_cfg_l; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_10_cfg_a = pmp_io_pmp_10_cfg_a; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_10_cfg_x = pmp_io_pmp_10_cfg_x; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_10_cfg_w = pmp_io_pmp_10_cfg_w; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_10_cfg_r = pmp_io_pmp_10_cfg_r; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_10_addr = pmp_io_pmp_10_addr; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_10_mask = pmp_io_pmp_10_mask; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_11_cfg_l = pmp_io_pmp_11_cfg_l; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_11_cfg_a = pmp_io_pmp_11_cfg_a; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_11_cfg_x = pmp_io_pmp_11_cfg_x; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_11_cfg_w = pmp_io_pmp_11_cfg_w; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_11_cfg_r = pmp_io_pmp_11_cfg_r; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_11_addr = pmp_io_pmp_11_addr; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_11_mask = pmp_io_pmp_11_mask; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_12_cfg_l = pmp_io_pmp_12_cfg_l; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_12_cfg_a = pmp_io_pmp_12_cfg_a; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_12_cfg_x = pmp_io_pmp_12_cfg_x; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_12_cfg_w = pmp_io_pmp_12_cfg_w; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_12_cfg_r = pmp_io_pmp_12_cfg_r; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_12_addr = pmp_io_pmp_12_addr; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_12_mask = pmp_io_pmp_12_mask; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_13_cfg_l = pmp_io_pmp_13_cfg_l; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_13_cfg_a = pmp_io_pmp_13_cfg_a; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_13_cfg_x = pmp_io_pmp_13_cfg_x; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_13_cfg_w = pmp_io_pmp_13_cfg_w; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_13_cfg_r = pmp_io_pmp_13_cfg_r; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_13_addr = pmp_io_pmp_13_addr; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_13_mask = pmp_io_pmp_13_mask; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_14_cfg_l = pmp_io_pmp_14_cfg_l; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_14_cfg_a = pmp_io_pmp_14_cfg_a; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_14_cfg_x = pmp_io_pmp_14_cfg_x; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_14_cfg_w = pmp_io_pmp_14_cfg_w; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_14_cfg_r = pmp_io_pmp_14_cfg_r; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_14_addr = pmp_io_pmp_14_addr; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_14_mask = pmp_io_pmp_14_mask; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_15_cfg_l = pmp_io_pmp_15_cfg_l; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_15_cfg_a = pmp_io_pmp_15_cfg_a; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_15_cfg_x = pmp_io_pmp_15_cfg_x; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_15_cfg_w = pmp_io_pmp_15_cfg_w; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_15_cfg_r = pmp_io_pmp_15_cfg_r; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_15_addr = pmp_io_pmp_15_addr; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_15_mask = pmp_io_pmp_15_mask; // @[Frontend.scala 88:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pma_0_cfg_c = pmp_io_pma_0_cfg_c; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_0_cfg_atomic = pmp_io_pma_0_cfg_atomic; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_0_cfg_a = pmp_io_pma_0_cfg_a; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_0_cfg_x = pmp_io_pma_0_cfg_x; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_0_cfg_w = pmp_io_pma_0_cfg_w; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_0_cfg_r = pmp_io_pma_0_cfg_r; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_0_addr = pmp_io_pma_0_addr; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_0_mask = pmp_io_pma_0_mask; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_1_cfg_c = pmp_io_pma_1_cfg_c; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_1_cfg_atomic = pmp_io_pma_1_cfg_atomic; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_1_cfg_a = pmp_io_pma_1_cfg_a; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_1_cfg_x = pmp_io_pma_1_cfg_x; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_1_cfg_w = pmp_io_pma_1_cfg_w; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_1_cfg_r = pmp_io_pma_1_cfg_r; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_1_addr = pmp_io_pma_1_addr; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_1_mask = pmp_io_pma_1_mask; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_2_cfg_c = pmp_io_pma_2_cfg_c; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_2_cfg_atomic = pmp_io_pma_2_cfg_atomic; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_2_cfg_a = pmp_io_pma_2_cfg_a; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_2_cfg_x = pmp_io_pma_2_cfg_x; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_2_cfg_w = pmp_io_pma_2_cfg_w; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_2_cfg_r = pmp_io_pma_2_cfg_r; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_2_addr = pmp_io_pma_2_addr; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_2_mask = pmp_io_pma_2_mask; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_3_cfg_c = pmp_io_pma_3_cfg_c; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_3_cfg_atomic = pmp_io_pma_3_cfg_atomic; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_3_cfg_a = pmp_io_pma_3_cfg_a; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_3_cfg_x = pmp_io_pma_3_cfg_x; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_3_cfg_w = pmp_io_pma_3_cfg_w; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_3_cfg_r = pmp_io_pma_3_cfg_r; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_3_addr = pmp_io_pma_3_addr; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_3_mask = pmp_io_pma_3_mask; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_4_cfg_c = pmp_io_pma_4_cfg_c; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_4_cfg_atomic = pmp_io_pma_4_cfg_atomic; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_4_cfg_a = pmp_io_pma_4_cfg_a; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_4_cfg_x = pmp_io_pma_4_cfg_x; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_4_cfg_w = pmp_io_pma_4_cfg_w; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_4_cfg_r = pmp_io_pma_4_cfg_r; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_4_addr = pmp_io_pma_4_addr; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_4_mask = pmp_io_pma_4_mask; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_5_cfg_c = pmp_io_pma_5_cfg_c; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_5_cfg_atomic = pmp_io_pma_5_cfg_atomic; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_5_cfg_a = pmp_io_pma_5_cfg_a; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_5_cfg_x = pmp_io_pma_5_cfg_x; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_5_cfg_w = pmp_io_pma_5_cfg_w; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_5_cfg_r = pmp_io_pma_5_cfg_r; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_5_addr = pmp_io_pma_5_addr; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_5_mask = pmp_io_pma_5_mask; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_6_cfg_c = pmp_io_pma_6_cfg_c; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_6_cfg_atomic = pmp_io_pma_6_cfg_atomic; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_6_cfg_a = pmp_io_pma_6_cfg_a; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_6_cfg_x = pmp_io_pma_6_cfg_x; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_6_cfg_w = pmp_io_pma_6_cfg_w; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_6_cfg_r = pmp_io_pma_6_cfg_r; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_6_addr = pmp_io_pma_6_addr; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_6_mask = pmp_io_pma_6_mask; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_7_cfg_c = pmp_io_pma_7_cfg_c; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_7_cfg_atomic = pmp_io_pma_7_cfg_atomic; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_7_cfg_a = pmp_io_pma_7_cfg_a; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_7_cfg_x = pmp_io_pma_7_cfg_x; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_7_cfg_w = pmp_io_pma_7_cfg_w; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_7_cfg_r = pmp_io_pma_7_cfg_r; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_7_addr = pmp_io_pma_7_addr; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_7_mask = pmp_io_pma_7_mask; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_8_cfg_c = pmp_io_pma_8_cfg_c; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_8_cfg_atomic = pmp_io_pma_8_cfg_atomic; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_8_cfg_a = pmp_io_pma_8_cfg_a; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_8_cfg_x = pmp_io_pma_8_cfg_x; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_8_cfg_w = pmp_io_pma_8_cfg_w; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_8_cfg_r = pmp_io_pma_8_cfg_r; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_8_addr = pmp_io_pma_8_addr; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_8_mask = pmp_io_pma_8_mask; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_9_cfg_c = pmp_io_pma_9_cfg_c; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_9_cfg_atomic = pmp_io_pma_9_cfg_atomic; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_9_cfg_a = pmp_io_pma_9_cfg_a; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_9_cfg_x = pmp_io_pma_9_cfg_x; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_9_cfg_w = pmp_io_pma_9_cfg_w; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_9_cfg_r = pmp_io_pma_9_cfg_r; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_9_addr = pmp_io_pma_9_addr; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_9_mask = pmp_io_pma_9_mask; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_10_cfg_c = pmp_io_pma_10_cfg_c; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_10_cfg_atomic = pmp_io_pma_10_cfg_atomic; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_10_cfg_a = pmp_io_pma_10_cfg_a; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_10_cfg_x = pmp_io_pma_10_cfg_x; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_10_cfg_w = pmp_io_pma_10_cfg_w; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_10_cfg_r = pmp_io_pma_10_cfg_r; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_10_addr = pmp_io_pma_10_addr; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_10_mask = pmp_io_pma_10_mask; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_11_cfg_c = pmp_io_pma_11_cfg_c; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_11_cfg_atomic = pmp_io_pma_11_cfg_atomic; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_11_cfg_a = pmp_io_pma_11_cfg_a; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_11_cfg_x = pmp_io_pma_11_cfg_x; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_11_cfg_w = pmp_io_pma_11_cfg_w; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_11_cfg_r = pmp_io_pma_11_cfg_r; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_11_addr = pmp_io_pma_11_addr; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_11_mask = pmp_io_pma_11_mask; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_12_cfg_c = pmp_io_pma_12_cfg_c; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_12_cfg_atomic = pmp_io_pma_12_cfg_atomic; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_12_cfg_a = pmp_io_pma_12_cfg_a; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_12_cfg_x = pmp_io_pma_12_cfg_x; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_12_cfg_w = pmp_io_pma_12_cfg_w; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_12_cfg_r = pmp_io_pma_12_cfg_r; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_12_addr = pmp_io_pma_12_addr; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_12_mask = pmp_io_pma_12_mask; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_13_cfg_c = pmp_io_pma_13_cfg_c; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_13_cfg_atomic = pmp_io_pma_13_cfg_atomic; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_13_cfg_a = pmp_io_pma_13_cfg_a; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_13_cfg_x = pmp_io_pma_13_cfg_x; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_13_cfg_w = pmp_io_pma_13_cfg_w; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_13_cfg_r = pmp_io_pma_13_cfg_r; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_13_addr = pmp_io_pma_13_addr; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_13_mask = pmp_io_pma_13_mask; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_14_cfg_c = pmp_io_pma_14_cfg_c; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_14_cfg_atomic = pmp_io_pma_14_cfg_atomic; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_14_cfg_a = pmp_io_pma_14_cfg_a; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_14_cfg_x = pmp_io_pma_14_cfg_x; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_14_cfg_w = pmp_io_pma_14_cfg_w; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_14_cfg_r = pmp_io_pma_14_cfg_r; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_14_addr = pmp_io_pma_14_addr; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_14_mask = pmp_io_pma_14_mask; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_15_cfg_c = pmp_io_pma_15_cfg_c; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_15_cfg_atomic = pmp_io_pma_15_cfg_atomic; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_15_cfg_a = pmp_io_pma_15_cfg_a; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_15_cfg_x = pmp_io_pma_15_cfg_x; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_15_cfg_w = pmp_io_pma_15_cfg_w; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_15_cfg_r = pmp_io_pma_15_cfg_r; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_15_addr = pmp_io_pma_15_addr; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_15_mask = pmp_io_pma_15_mask; // @[Frontend.scala 88:26 PMP.scala 467:14]
  assign PMPChecker_3_io_req_bits_addr = ifu_io_pmp_req_bits_addr; // @[Frontend.scala 90:29 94:18]
  assign PMPChecker_3_io_req_bits_cmd = 3'h2; // @[Frontend.scala 90:29 94:18]
  assign itlb_clock = clock;
  assign itlb_reset = reset;
  assign itlb_io_sfence_valid = io_sfence_valid; // @[MMUBundle.scala 448:17]
  assign itlb_io_sfence_bits_rs1 = io_sfence_bits_rs1; // @[MMUBundle.scala 448:17]
  assign itlb_io_sfence_bits_rs2 = io_sfence_bits_rs2; // @[MMUBundle.scala 448:17]
  assign itlb_io_sfence_bits_addr = io_sfence_bits_addr; // @[MMUBundle.scala 448:17]
  assign itlb_io_sfence_bits_asid = io_sfence_bits_asid; // @[MMUBundle.scala 448:17]
  assign itlb_io_csr_satp_mode = tlbCsr_delay_io_out_satp_mode; // @[MMUBundle.scala 449:14]
  assign itlb_io_csr_satp_asid = tlbCsr_delay_io_out_satp_asid; // @[MMUBundle.scala 449:14]
  assign itlb_io_csr_satp_changed = tlbCsr_delay_io_out_satp_changed; // @[MMUBundle.scala 449:14]
  assign itlb_io_csr_priv_imode = tlbCsr_delay_io_out_priv_imode; // @[MMUBundle.scala 449:14]
  assign itlb_io_requestor_0_req_valid = icache_io_itlb_0_req_valid; // @[Frontend.scala 105:73]
  assign itlb_io_requestor_0_req_bits_vaddr = icache_io_itlb_0_req_bits_vaddr; // @[Frontend.scala 105:73]
  assign itlb_io_requestor_0_req_bits_kill = icache_io_itlb_0_req_bits_kill; // @[Frontend.scala 105:73]
  assign itlb_io_requestor_0_resp_ready = icache_io_itlb_0_resp_ready; // @[Frontend.scala 105:73]
  assign itlb_io_requestor_1_req_valid = icache_io_itlb_1_req_valid; // @[Frontend.scala 105:73]
  assign itlb_io_requestor_1_req_bits_vaddr = icache_io_itlb_1_req_bits_vaddr; // @[Frontend.scala 105:73]
  assign itlb_io_requestor_1_req_bits_kill = icache_io_itlb_1_req_bits_kill; // @[Frontend.scala 105:73]
  assign itlb_io_requestor_1_resp_ready = icache_io_itlb_1_resp_ready; // @[Frontend.scala 105:73]
  assign itlb_io_requestor_3_req_valid = ifu_io_iTLBInter_req_valid; // @[Frontend.scala 106:24]
  assign itlb_io_requestor_3_req_bits_vaddr = ifu_io_iTLBInter_req_bits_vaddr; // @[Frontend.scala 106:24]
  assign itlb_io_flushPipe_0 = needFlush; // @[Frontend.scala 110:27]
  assign itlb_io_flushPipe_1 = needFlush; // @[Frontend.scala 110:27]
  assign itlb_io_flushPipe_3 = needFlush; // @[Frontend.scala 110:27]
  assign itlb_io_ptw_req_0_ready = io_ptw_req_0_ready; // @[MMUBundle.scala 487:9]
  assign itlb_io_ptw_req_1_ready = io_ptw_req_1_ready; // @[MMUBundle.scala 487:9]
  assign itlb_io_ptw_req_3_ready = io_ptw_req_3_ready; // @[MMUBundle.scala 487:9]
  assign itlb_io_ptw_resp_valid = io_ptw_resp_valid; // @[MMUBundle.scala 490:23]
  assign itlb_io_ptw_resp_bits_entry_tag = io_ptw_resp_bits_data_entry_tag; // @[MMUBundle.scala 489:22]
  assign itlb_io_ptw_resp_bits_entry_asid = io_ptw_resp_bits_data_entry_asid; // @[MMUBundle.scala 489:22]
  assign itlb_io_ptw_resp_bits_entry_ppn = io_ptw_resp_bits_data_entry_ppn; // @[MMUBundle.scala 489:22]
  assign itlb_io_ptw_resp_bits_entry_perm_d = io_ptw_resp_bits_data_entry_perm_d; // @[MMUBundle.scala 489:22]
  assign itlb_io_ptw_resp_bits_entry_perm_a = io_ptw_resp_bits_data_entry_perm_a; // @[MMUBundle.scala 489:22]
  assign itlb_io_ptw_resp_bits_entry_perm_g = io_ptw_resp_bits_data_entry_perm_g; // @[MMUBundle.scala 489:22]
  assign itlb_io_ptw_resp_bits_entry_perm_u = io_ptw_resp_bits_data_entry_perm_u; // @[MMUBundle.scala 489:22]
  assign itlb_io_ptw_resp_bits_entry_perm_x = io_ptw_resp_bits_data_entry_perm_x; // @[MMUBundle.scala 489:22]
  assign itlb_io_ptw_resp_bits_entry_perm_w = io_ptw_resp_bits_data_entry_perm_w; // @[MMUBundle.scala 489:22]
  assign itlb_io_ptw_resp_bits_entry_perm_r = io_ptw_resp_bits_data_entry_perm_r; // @[MMUBundle.scala 489:22]
  assign itlb_io_ptw_resp_bits_entry_level = io_ptw_resp_bits_data_entry_level; // @[MMUBundle.scala 489:22]
  assign itlb_io_ptw_resp_bits_pf = io_ptw_resp_bits_data_pf; // @[MMUBundle.scala 489:22]
  assign itlb_io_ptw_resp_bits_af = io_ptw_resp_bits_data_af; // @[MMUBundle.scala 489:22]
  assign pfevent_clock = clock;
  assign pfevent_reset = reset;
  assign pfevent_io_distribute_csr_wvalid = io_csrCtrl_distribute_csr_wvalid; // @[Frontend.scala 166:29]
  assign pfevent_io_distribute_csr_waddr = io_csrCtrl_distribute_csr_waddr; // @[Frontend.scala 166:29]
  assign pfevent_io_distribute_csr_wdata = io_csrCtrl_distribute_csr_wdata; // @[Frontend.scala 166:29]
  assign hpm_clock = clock;
  assign hpm_io_hpm_event_0 = pfevent_io_hpmevent_0; // @[PerfCounterUtils.scala 256:22]
  assign hpm_io_hpm_event_1 = pfevent_io_hpmevent_1; // @[PerfCounterUtils.scala 256:22]
  assign hpm_io_hpm_event_2 = pfevent_io_hpmevent_2; // @[PerfCounterUtils.scala 256:22]
  assign hpm_io_hpm_event_3 = pfevent_io_hpmevent_3; // @[PerfCounterUtils.scala 256:22]
  assign hpm_io_hpm_event_4 = pfevent_io_hpmevent_4; // @[PerfCounterUtils.scala 256:22]
  assign hpm_io_hpm_event_5 = pfevent_io_hpmevent_5; // @[PerfCounterUtils.scala 256:22]
  assign hpm_io_hpm_event_6 = pfevent_io_hpmevent_6; // @[PerfCounterUtils.scala 256:22]
  assign hpm_io_hpm_event_7 = pfevent_io_hpmevent_7; // @[PerfCounterUtils.scala 256:22]
  assign hpm_io_events_sets_0_value = ifu_io_perf_0_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_1_value = ifu_io_perf_1_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_2_value = ifu_io_perf_2_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_3_value = ifu_io_perf_3_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_4_value = ifu_io_perf_4_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_5_value = ifu_io_perf_5_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_6_value = ifu_io_perf_6_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_7_value = ifu_io_perf_7_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_8_value = ifu_io_perf_8_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_9_value = ifu_io_perf_9_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_10_value = ifu_io_perf_10_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_11_value = ifu_io_perf_11_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_12_value = ifu_io_perf_12_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_13_value = ibuffer_io_perf_0_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_14_value = ibuffer_io_perf_1_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_15_value = ibuffer_io_perf_2_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_16_value = ibuffer_io_perf_3_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_17_value = ibuffer_io_perf_4_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_18_value = ibuffer_io_perf_5_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_19_value = ibuffer_io_perf_6_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_20_value = ibuffer_io_perf_7_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_23_value = ftq_io_perf_0_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_24_value = ftq_io_perf_1_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_25_value = ftq_io_perf_2_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_26_value = ftq_io_perf_3_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_27_value = ftq_io_perf_4_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_28_value = ftq_io_perf_5_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_29_value = ftq_io_perf_6_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_30_value = ftq_io_perf_7_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_31_value = ftq_io_perf_8_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_32_value = ftq_io_perf_9_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_33_value = ftq_io_perf_10_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_34_value = ftq_io_perf_11_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_35_value = ftq_io_perf_12_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_36_value = ftq_io_perf_13_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_37_value = ftq_io_perf_14_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_38_value = ftq_io_perf_15_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_39_value = ftq_io_perf_16_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_40_value = ftq_io_perf_17_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_41_value = ftq_io_perf_18_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_42_value = ftq_io_perf_19_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_43_value = ftq_io_perf_20_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_44_value = ftq_io_perf_21_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_45_value = ftq_io_perf_22_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_46_value = ftq_io_perf_23_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_47_value = bpu_io_perf_0_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_48_value = bpu_io_perf_1_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_49_value = bpu_io_perf_2_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_50_value = bpu_io_perf_3_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_51_value = bpu_io_perf_4_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_52_value = bpu_io_perf_5_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_53_value = bpu_io_perf_6_value; // @[PerfCounterUtils.scala 257:24]
  always @(posedge clock) begin
    needFlush <= io_backend_toFtq_redirect_valid; // @[Frontend.scala 71:26]
    io_csrUpdate_REG_wvalid <= icache_io_csr_update_wvalid; // @[Frontend.scala 136:26]
    io_csrUpdate_REG_waddr <= icache_io_csr_update_waddr; // @[Frontend.scala 136:26]
    io_csrUpdate_REG_wdata <= icache_io_csr_update_wdata; // @[Frontend.scala 136:26]
    icache_io_csr_parity_enable_REG <= csrCtrl_delay_io_out_icache_parity_enable; // @[Frontend.scala 139:41]
    io_error_REG_paddr <= icache_io_error_paddr; // @[Frontend.scala 156:30]
    io_error_REG_report_to_beu <= icache_io_error_report_to_beu; // @[Frontend.scala 156:30]
    io_error_REG_1_paddr <= io_error_REG_paddr; // @[Frontend.scala 156:22]
    io_error_REG_1_report_to_beu <= io_error_REG_report_to_beu; // @[Frontend.scala 156:22]
    io_perf_0_value_REG <= hpm_io_perf_0_value; // @[PerfCounterUtils.scala 188:35]
    io_perf_0_value_REG_1 <= io_perf_0_value_REG; // @[PerfCounterUtils.scala 188:27]
    io_perf_1_value_REG <= hpm_io_perf_1_value; // @[PerfCounterUtils.scala 188:35]
    io_perf_1_value_REG_1 <= io_perf_1_value_REG; // @[PerfCounterUtils.scala 188:27]
    io_perf_2_value_REG <= hpm_io_perf_2_value; // @[PerfCounterUtils.scala 188:35]
    io_perf_2_value_REG_1 <= io_perf_2_value_REG; // @[PerfCounterUtils.scala 188:27]
    io_perf_3_value_REG <= hpm_io_perf_3_value; // @[PerfCounterUtils.scala 188:35]
    io_perf_3_value_REG_1 <= io_perf_3_value_REG; // @[PerfCounterUtils.scala 188:27]
    io_perf_4_value_REG <= hpm_io_perf_4_value; // @[PerfCounterUtils.scala 188:35]
    io_perf_4_value_REG_1 <= io_perf_4_value_REG; // @[PerfCounterUtils.scala 188:27]
    io_perf_5_value_REG <= hpm_io_perf_5_value; // @[PerfCounterUtils.scala 188:35]
    io_perf_5_value_REG_1 <= io_perf_5_value_REG; // @[PerfCounterUtils.scala 188:27]
    io_perf_6_value_REG <= hpm_io_perf_6_value; // @[PerfCounterUtils.scala 188:35]
    io_perf_6_value_REG_1 <= io_perf_6_value_REG; // @[PerfCounterUtils.scala 188:27]
    io_perf_7_value_REG <= hpm_io_perf_7_value; // @[PerfCounterUtils.scala 188:35]
    io_perf_7_value_REG_1 <= io_perf_7_value_REG; // @[PerfCounterUtils.scala 188:27]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  needFlush = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  io_csrUpdate_REG_wvalid = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  io_csrUpdate_REG_waddr = _RAND_2[11:0];
  _RAND_3 = {2{`RANDOM}};
  io_csrUpdate_REG_wdata = _RAND_3[63:0];
  _RAND_4 = {1{`RANDOM}};
  icache_io_csr_parity_enable_REG = _RAND_4[0:0];
  _RAND_5 = {2{`RANDOM}};
  io_error_REG_paddr = _RAND_5[35:0];
  _RAND_6 = {1{`RANDOM}};
  io_error_REG_report_to_beu = _RAND_6[0:0];
  _RAND_7 = {2{`RANDOM}};
  io_error_REG_1_paddr = _RAND_7[35:0];
  _RAND_8 = {1{`RANDOM}};
  io_error_REG_1_report_to_beu = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  io_perf_0_value_REG = _RAND_9[5:0];
  _RAND_10 = {1{`RANDOM}};
  io_perf_0_value_REG_1 = _RAND_10[5:0];
  _RAND_11 = {1{`RANDOM}};
  io_perf_1_value_REG = _RAND_11[5:0];
  _RAND_12 = {1{`RANDOM}};
  io_perf_1_value_REG_1 = _RAND_12[5:0];
  _RAND_13 = {1{`RANDOM}};
  io_perf_2_value_REG = _RAND_13[5:0];
  _RAND_14 = {1{`RANDOM}};
  io_perf_2_value_REG_1 = _RAND_14[5:0];
  _RAND_15 = {1{`RANDOM}};
  io_perf_3_value_REG = _RAND_15[5:0];
  _RAND_16 = {1{`RANDOM}};
  io_perf_3_value_REG_1 = _RAND_16[5:0];
  _RAND_17 = {1{`RANDOM}};
  io_perf_4_value_REG = _RAND_17[5:0];
  _RAND_18 = {1{`RANDOM}};
  io_perf_4_value_REG_1 = _RAND_18[5:0];
  _RAND_19 = {1{`RANDOM}};
  io_perf_5_value_REG = _RAND_19[5:0];
  _RAND_20 = {1{`RANDOM}};
  io_perf_5_value_REG_1 = _RAND_20[5:0];
  _RAND_21 = {1{`RANDOM}};
  io_perf_6_value_REG = _RAND_21[5:0];
  _RAND_22 = {1{`RANDOM}};
  io_perf_6_value_REG_1 = _RAND_22[5:0];
  _RAND_23 = {1{`RANDOM}};
  io_perf_7_value_REG = _RAND_23[5:0];
  _RAND_24 = {1{`RANDOM}};
  io_perf_7_value_REG_1 = _RAND_24[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule

