module DelayN_94(
  input  [7:0] io_in,
  output [7:0] io_out
);
  assign io_out = io_in; // @[Hold.scala 92:10]
endmodule

