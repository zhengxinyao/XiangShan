module bosc_mbist_controller_L3_dfx_top(
  input          io_mbist_ijtag_tck,
  input          io_mbist_ijtag_reset,
  input          io_mbist_ijtag_ce,
  input          io_mbist_ijtag_se,
  input          io_mbist_ijtag_ue,
  input          io_mbist_ijtag_sel,
  input          io_mbist_ijtag_si,
  output         io_mbist_ijtag_so,
  output         io_mbist_ijtag_diag_done,
  output [10:0]  io_hd2prf_out_trim_fuse,
  output [1:0]   io_hd2prf_out_sleep_fuse,
  output [19:0]  io_hsuspsr_out_trim_fuse,
  output [1:0]   io_hsuspsr_out_sleep_fuse,
  output [19:0]  io_uhdusplr_out_trim_fuse,
  output [1:0]   io_uhdusplr_out_sleep_fuse,
  output [19:0]  io_hduspsr_out_trim_fuse,
  output [1:0]   io_hduspsr_out_sleep_fuse,
  input  [10:0]  io_hd2prf_in_trim_fuse,
  input  [1:0]   io_hd2prf_in_sleep_fuse,
  input  [19:0]  io_hsuspsr_in_trim_fuse,
  input  [1:0]   io_hsuspsr_in_sleep_fuse,
  input  [19:0]  io_uhdusplr_in_trim_fuse,
  input  [1:0]   io_uhdusplr_in_sleep_fuse,
  input  [19:0]  io_hduspsr_in_trim_fuse,
  input  [1:0]   io_hduspsr_in_sleep_fuse,
  input          io_xsx_fscan_in_bypsel,
  input          io_xsx_fscan_in_wdis_b,
  input          io_xsx_fscan_in_rdis_b,
  input          io_xsx_fscan_in_init_en,
  input          io_xsx_fscan_in_init_val,
  input          io_xsl2_fscan_in_bypsel,
  input          io_xsl2_fscan_in_wdis_b,
  input          io_xsl2_fscan_in_rdis_b,
  input          io_xsl2_fscan_in_init_en,
  input          io_xsl2_fscan_in_init_val,
  input          io_fscan_clkungate,
  input          io_clock,
  input          io_bisr_shift_en,
  input          io_bisr_clock,
  input          io_bisr_reset,
  input          io_bisr_scan_in,
  output         io_bisr_scan_out,
  input          io_bisr_mem_chain_select,
  output         io_L3_bisr_shift_en,
  output         io_L3_bisr_clock,
  output         io_L3_bisr_reset,
  output         io_L3_bisr_scan_in,
  input          io_L3_bisr_scan_out,
  output [25:0]  slice_bankedData0_bank0_rowRepair,
  output [12:0]  slice_bankedData0_bank0_colRepair,
  output [25:0]  slice_bankedData0_bank1_rowRepair,
  output [12:0]  slice_bankedData0_bank1_colRepair,
  output [25:0]  slice_bankedData0_bank2_rowRepair,
  output [12:0]  slice_bankedData0_bank2_colRepair,
  output [25:0]  slice_bankedData0_bank3_rowRepair,
  output [12:0]  slice_bankedData0_bank3_colRepair,
  output [25:0]  slice_bankedData1_bank0_rowRepair,
  output [12:0]  slice_bankedData1_bank0_colRepair,
  output [25:0]  slice_bankedData1_bank1_rowRepair,
  output [12:0]  slice_bankedData1_bank1_colRepair,
  output [25:0]  slice_bankedData1_bank2_rowRepair,
  output [12:0]  slice_bankedData1_bank2_colRepair,
  output [25:0]  slice_bankedData1_bank3_rowRepair,
  output [12:0]  slice_bankedData1_bank3_colRepair,
  output [25:0]  slice_bankedData2_bank0_rowRepair,
  output [12:0]  slice_bankedData2_bank0_colRepair,
  output [25:0]  slice_bankedData2_bank1_rowRepair,
  output [12:0]  slice_bankedData2_bank1_colRepair,
  output [25:0]  slice_bankedData2_bank2_rowRepair,
  output [12:0]  slice_bankedData2_bank2_colRepair,
  output [25:0]  slice_bankedData2_bank3_rowRepair,
  output [12:0]  slice_bankedData2_bank3_colRepair,
  output [25:0]  slice_bankedData3_bank0_rowRepair,
  output [12:0]  slice_bankedData3_bank0_colRepair,
  output [25:0]  slice_bankedData3_bank1_rowRepair,
  output [12:0]  slice_bankedData3_bank1_colRepair,
  output [25:0]  slice_bankedData3_bank2_rowRepair,
  output [12:0]  slice_bankedData3_bank2_colRepair,
  output [25:0]  slice_bankedData3_bank3_rowRepair,
  output [12:0]  slice_bankedData3_bank3_colRepair,
  output [25:0]  slice_bankedData4_bank0_rowRepair,
  output [12:0]  slice_bankedData4_bank0_colRepair,
  output [25:0]  slice_bankedData4_bank1_rowRepair,
  output [12:0]  slice_bankedData4_bank1_colRepair,
  output [25:0]  slice_bankedData4_bank2_rowRepair,
  output [12:0]  slice_bankedData4_bank2_colRepair,
  output [25:0]  slice_bankedData4_bank3_rowRepair,
  output [12:0]  slice_bankedData4_bank3_colRepair,
  output [25:0]  slice_bankedData5_bank0_rowRepair,
  output [12:0]  slice_bankedData5_bank0_colRepair,
  output [25:0]  slice_bankedData5_bank1_rowRepair,
  output [12:0]  slice_bankedData5_bank1_colRepair,
  output [25:0]  slice_bankedData5_bank2_rowRepair,
  output [12:0]  slice_bankedData5_bank2_colRepair,
  output [25:0]  slice_bankedData5_bank3_rowRepair,
  output [12:0]  slice_bankedData5_bank3_colRepair,
  output [25:0]  slice_bankedData6_bank0_rowRepair,
  output [12:0]  slice_bankedData6_bank0_colRepair,
  output [25:0]  slice_bankedData6_bank1_rowRepair,
  output [12:0]  slice_bankedData6_bank1_colRepair,
  output [25:0]  slice_bankedData6_bank2_rowRepair,
  output [12:0]  slice_bankedData6_bank2_colRepair,
  output [25:0]  slice_bankedData6_bank3_rowRepair,
  output [12:0]  slice_bankedData6_bank3_colRepair,
  output [25:0]  slice_bankedData7_bank0_rowRepair,
  output [12:0]  slice_bankedData7_bank0_colRepair,
  output [25:0]  slice_bankedData7_bank1_rowRepair,
  output [12:0]  slice_bankedData7_bank1_colRepair,
  output [25:0]  slice_bankedData7_bank2_rowRepair,
  output [12:0]  slice_bankedData7_bank2_colRepair,
  output [25:0]  slice_bankedData7_bank3_rowRepair,
  output [12:0]  slice_bankedData7_bank3_colRepair,
  output [25:0]  slice_dataEcc0_bank0_rowRepair,
  output [12:0]  slice_dataEcc0_bank0_colRepair,
  output [25:0]  slice_dataEcc0_bank1_rowRepair,
  output [12:0]  slice_dataEcc0_bank1_colRepair,
  output [25:0]  slice_dataEcc0_bank2_rowRepair,
  output [12:0]  slice_dataEcc0_bank2_colRepair,
  output [25:0]  slice_dataEcc0_bank3_rowRepair,
  output [12:0]  slice_dataEcc0_bank3_colRepair,
  output [25:0]  slice_dataEcc1_bank0_rowRepair,
  output [12:0]  slice_dataEcc1_bank0_colRepair,
  output [25:0]  slice_dataEcc1_bank1_rowRepair,
  output [12:0]  slice_dataEcc1_bank1_colRepair,
  output [25:0]  slice_dataEcc1_bank2_rowRepair,
  output [12:0]  slice_dataEcc1_bank2_colRepair,
  output [25:0]  slice_dataEcc1_bank3_rowRepair,
  output [12:0]  slice_dataEcc1_bank3_colRepair,
  output [5:0]   io_L3_SRAM_array,
  output         io_L3_SRAM_all,
  output         io_L3_SRAM_req,
  input          io_L3_SRAM_ack,
  output         io_L3_SRAM_writeen,
  output [7:0]   io_L3_SRAM_be,
  output [11:0]  io_L3_SRAM_addr,
  output [167:0] io_L3_SRAM_indata,
  output         io_L3_SRAM_readen,
  input  [167:0] io_L3_SRAM_outdata,
  output         io_fscan_ram_L3_bypsel,
  output         io_fscan_ram_L3_wdis_b,
  output         io_fscan_ram_L3_rdis_b,
  output         io_fscan_ram_L3_init_en,
  output         io_fscan_ram_L3_init_val,
  output         io_fscan_ram_L3_clkungate
);
  mbist_controller_L3_dfx_wrap mbistControllers_l3 ( // @[HuanCun.scala 461:28]
    .i_L3_mbist_ijtag_tck(io_mbist_ijtag_tck),
    .i_L3_mbist_ijtag_reset(io_mbist_ijtag_reset),
    .i_L3_mbist_ijtag_ce(io_mbist_ijtag_ce),
    .i_L3_mbist_ijtag_se(io_mbist_ijtag_se),
    .i_L3_mbist_ijtag_ue(io_mbist_ijtag_ue),
    .i_L3_mbist_ijtag_sel(io_mbist_ijtag_sel),
    .i_L3_mbist_ijtag_si(io_mbist_ijtag_si),
    .o_L3_mbist_ijtag_so(io_mbist_ijtag_so),
    .o_L3_aary_mbist_diag_done(io_mbist_ijtag_diag_done),
    .o_L3_hsuspsr_trim_fuse_out(io_hsuspsr_out_trim_fuse),
    .o_L3_hsuspsr_sleep_fuse_out(io_hsuspsr_out_sleep_fuse),
    .o_L3_uhdusplr_trim_fuse_out(io_uhdusplr_out_trim_fuse),
    .o_L3_uhdusplr_sleep_fuse_out(io_uhdusplr_out_sleep_fuse),
    .i_L3_hsuspsr_trim_fuse_in(io_hsuspsr_in_trim_fuse),
    .i_L3_hsuspsr_sleep_fuse_in(io_hsuspsr_in_sleep_fuse),
    .i_L3_uhdusplr_trim_fuse_in(io_uhdusplr_in_trim_fuse),
    .i_L3_uhdusplr_sleep_fuse_in(io_uhdusplr_in_sleep_fuse),
    .i_xsx_fscan_ram_bypsel(io_xsx_fscan_in_bypsel),
    .i_xsx_fscan_ram_wdis_b(io_xsx_fscan_in_wdis_b),
    .i_xsx_fscan_ram_rdis_b(io_xsx_fscan_in_rdis_b),
    .i_xsx_fscan_ram_init_en(io_xsx_fscan_in_init_en),
    .i_xsx_fscan_ram_init_val(io_xsx_fscan_in_init_val),
    .i_xsl2_fscan_ram_bypsel(io_xsl2_fscan_in_bypsel),
    .i_xsl2_fscan_ram_wdis_b(io_xsl2_fscan_in_wdis_b),
    .i_xsl2_fscan_ram_rdis_b(io_xsl2_fscan_in_rdis_b),
    .i_xsl2_fscan_ram_init_en(io_xsl2_fscan_in_init_en),
    .i_xsl2_fscan_ram_init_val(io_xsl2_fscan_in_init_val),
    .i_fscan_clkungate(io_fscan_clkungate),
    .l3cacheOpt_clock(io_clock),
    .i_L3_mbist_bisr_mem_chain_select(io_bisr_mem_chain_select),
    .i_L3_mbist_bisr_shift_en(io_bisr_shift_en),
    .i_L3_mbist_bisr_clock(io_bisr_clock),
    .i_L3_mbist_bisr_reset(io_bisr_reset),
    .i_L3_mbist_bisr_scan_in(io_bisr_scan_in),
    .o_L3_mbist_bisr_scan_out(io_bisr_scan_out),
    .o_L3_bisr_shift_en(io_L3_bisr_shift_en),
    .o_L3_bisr_clock(io_L3_bisr_clock),
    .o_L3_bisr_reset(io_L3_bisr_reset),
    .o_L3_bisr_scan_in(io_L3_bisr_scan_in),
    .i_L3_bisr_scan_out(io_L3_bisr_scan_out),
    .slice_bankedData0_bank0_rowRepair(slice_bankedData0_bank0_rowRepair),
    .slice_bankedData0_bank0_colRepair(slice_bankedData0_bank0_colRepair),
    .slice_bankedData0_bank1_rowRepair(slice_bankedData0_bank1_rowRepair),
    .slice_bankedData0_bank1_colRepair(slice_bankedData0_bank1_colRepair),
    .slice_bankedData0_bank2_rowRepair(slice_bankedData0_bank2_rowRepair),
    .slice_bankedData0_bank2_colRepair(slice_bankedData0_bank2_colRepair),
    .slice_bankedData0_bank3_rowRepair(slice_bankedData0_bank3_rowRepair),
    .slice_bankedData0_bank3_colRepair(slice_bankedData0_bank3_colRepair),
    .slice_bankedData1_bank0_rowRepair(slice_bankedData1_bank0_rowRepair),
    .slice_bankedData1_bank0_colRepair(slice_bankedData1_bank0_colRepair),
    .slice_bankedData1_bank1_rowRepair(slice_bankedData1_bank1_rowRepair),
    .slice_bankedData1_bank1_colRepair(slice_bankedData1_bank1_colRepair),
    .slice_bankedData1_bank2_rowRepair(slice_bankedData1_bank2_rowRepair),
    .slice_bankedData1_bank2_colRepair(slice_bankedData1_bank2_colRepair),
    .slice_bankedData1_bank3_rowRepair(slice_bankedData1_bank3_rowRepair),
    .slice_bankedData1_bank3_colRepair(slice_bankedData1_bank3_colRepair),
    .slice_bankedData2_bank0_rowRepair(slice_bankedData2_bank0_rowRepair),
    .slice_bankedData2_bank0_colRepair(slice_bankedData2_bank0_colRepair),
    .slice_bankedData2_bank1_rowRepair(slice_bankedData2_bank1_rowRepair),
    .slice_bankedData2_bank1_colRepair(slice_bankedData2_bank1_colRepair),
    .slice_bankedData2_bank2_rowRepair(slice_bankedData2_bank2_rowRepair),
    .slice_bankedData2_bank2_colRepair(slice_bankedData2_bank2_colRepair),
    .slice_bankedData2_bank3_rowRepair(slice_bankedData2_bank3_rowRepair),
    .slice_bankedData2_bank3_colRepair(slice_bankedData2_bank3_colRepair),
    .slice_bankedData3_bank0_rowRepair(slice_bankedData3_bank0_rowRepair),
    .slice_bankedData3_bank0_colRepair(slice_bankedData3_bank0_colRepair),
    .slice_bankedData3_bank1_rowRepair(slice_bankedData3_bank1_rowRepair),
    .slice_bankedData3_bank1_colRepair(slice_bankedData3_bank1_colRepair),
    .slice_bankedData3_bank2_rowRepair(slice_bankedData3_bank2_rowRepair),
    .slice_bankedData3_bank2_colRepair(slice_bankedData3_bank2_colRepair),
    .slice_bankedData3_bank3_rowRepair(slice_bankedData3_bank3_rowRepair),
    .slice_bankedData3_bank3_colRepair(slice_bankedData3_bank3_colRepair),
    .slice_bankedData4_bank0_rowRepair(slice_bankedData4_bank0_rowRepair),
    .slice_bankedData4_bank0_colRepair(slice_bankedData4_bank0_colRepair),
    .slice_bankedData4_bank1_rowRepair(slice_bankedData4_bank1_rowRepair),
    .slice_bankedData4_bank1_colRepair(slice_bankedData4_bank1_colRepair),
    .slice_bankedData4_bank2_rowRepair(slice_bankedData4_bank2_rowRepair),
    .slice_bankedData4_bank2_colRepair(slice_bankedData4_bank2_colRepair),
    .slice_bankedData4_bank3_rowRepair(slice_bankedData4_bank3_rowRepair),
    .slice_bankedData4_bank3_colRepair(slice_bankedData4_bank3_colRepair),
    .slice_bankedData5_bank0_rowRepair(slice_bankedData5_bank0_rowRepair),
    .slice_bankedData5_bank0_colRepair(slice_bankedData5_bank0_colRepair),
    .slice_bankedData5_bank1_rowRepair(slice_bankedData5_bank1_rowRepair),
    .slice_bankedData5_bank1_colRepair(slice_bankedData5_bank1_colRepair),
    .slice_bankedData5_bank2_rowRepair(slice_bankedData5_bank2_rowRepair),
    .slice_bankedData5_bank2_colRepair(slice_bankedData5_bank2_colRepair),
    .slice_bankedData5_bank3_rowRepair(slice_bankedData5_bank3_rowRepair),
    .slice_bankedData5_bank3_colRepair(slice_bankedData5_bank3_colRepair),
    .slice_bankedData6_bank0_rowRepair(slice_bankedData6_bank0_rowRepair),
    .slice_bankedData6_bank0_colRepair(slice_bankedData6_bank0_colRepair),
    .slice_bankedData6_bank1_rowRepair(slice_bankedData6_bank1_rowRepair),
    .slice_bankedData6_bank1_colRepair(slice_bankedData6_bank1_colRepair),
    .slice_bankedData6_bank2_rowRepair(slice_bankedData6_bank2_rowRepair),
    .slice_bankedData6_bank2_colRepair(slice_bankedData6_bank2_colRepair),
    .slice_bankedData6_bank3_rowRepair(slice_bankedData6_bank3_rowRepair),
    .slice_bankedData6_bank3_colRepair(slice_bankedData6_bank3_colRepair),
    .slice_bankedData7_bank0_rowRepair(slice_bankedData7_bank0_rowRepair),
    .slice_bankedData7_bank0_colRepair(slice_bankedData7_bank0_colRepair),
    .slice_bankedData7_bank1_rowRepair(slice_bankedData7_bank1_rowRepair),
    .slice_bankedData7_bank1_colRepair(slice_bankedData7_bank1_colRepair),
    .slice_bankedData7_bank2_rowRepair(slice_bankedData7_bank2_rowRepair),
    .slice_bankedData7_bank2_colRepair(slice_bankedData7_bank2_colRepair),
    .slice_bankedData7_bank3_rowRepair(slice_bankedData7_bank3_rowRepair),
    .slice_bankedData7_bank3_colRepair(slice_bankedData7_bank3_colRepair),
    .slice_dataEccArray0_bank0_rowRepair(slice_dataEcc0_bank0_rowRepair),
    .slice_dataEccArray0_bank0_colRepair(slice_dataEcc0_bank0_colRepair),
    .slice_dataEccArray0_bank1_rowRepair(slice_dataEcc0_bank1_rowRepair),
    .slice_dataEccArray0_bank1_colRepair(slice_dataEcc0_bank1_colRepair),
    .slice_dataEccArray0_bank2_rowRepair(slice_dataEcc0_bank2_rowRepair),
    .slice_dataEccArray0_bank2_colRepair(slice_dataEcc0_bank2_colRepair),
    .slice_dataEccArray0_bank3_rowRepair(slice_dataEcc0_bank3_rowRepair),
    .slice_dataEccArray0_bank3_colRepair(slice_dataEcc0_bank3_colRepair),
    .slice_dataEccArray1_bank0_rowRepair(slice_dataEcc1_bank0_rowRepair),
    .slice_dataEccArray1_bank0_colRepair(slice_dataEcc1_bank0_colRepair),
    .slice_dataEccArray1_bank1_rowRepair(slice_dataEcc1_bank1_rowRepair),
    .slice_dataEccArray1_bank1_colRepair(slice_dataEcc1_bank1_colRepair),
    .slice_dataEccArray1_bank2_rowRepair(slice_dataEcc1_bank2_rowRepair),
    .slice_dataEccArray1_bank2_colRepair(slice_dataEcc1_bank2_colRepair),
    .slice_dataEccArray1_bank3_rowRepair(slice_dataEcc1_bank3_rowRepair),
    .slice_dataEccArray1_bank3_colRepair(slice_dataEcc1_bank3_colRepair),
    .o_L3_mbist_array(io_L3_SRAM_array),
    .o_L3_mbist_all(io_L3_SRAM_all),
    .o_L3_mbist_req(io_L3_SRAM_req),
    .i_L3_mbist_ack(io_L3_SRAM_ack),
    .o_L3_mbist_writeen(io_L3_SRAM_writeen),
    .o_L3_mbist_be(io_L3_SRAM_be),
    .o_L3_mbist_addr(io_L3_SRAM_addr),
    .o_L3_mbist_indata(io_L3_SRAM_indata),
    .o_L3_mbist_readen(io_L3_SRAM_readen),
    .i_L3_mbist_outdata(io_L3_SRAM_outdata),
    .o_L3_fscan_ram_bypsel(io_fscan_ram_L3_bypsel),
    .o_L3_fscan_ram_wdis_b(io_fscan_ram_L3_wdis_b),
    .o_L3_fscan_ram_rdis_b(io_fscan_ram_L3_rdis_b),
    .o_L3_fscan_ram_init_en(io_fscan_ram_L3_init_en),
    .o_L3_fscan_ram_init_val(io_fscan_ram_L3_init_val),
    .o_L3_fscan_clkungate(io_fscan_ram_L3_clkungate)
  );
  assign io_hd2prf_out_trim_fuse = 11'h0;
  assign io_hd2prf_out_sleep_fuse = 2'h0;
  assign io_hduspsr_out_trim_fuse = 20'h0;
  assign io_hduspsr_out_sleep_fuse = 2'h0;
endmodule

