module LoadQueueFlag(
  input         clock,
  input         reset,
  input         io_redirect_valid,
  input         io_redirect_bits_robIdx_flag,
  input  [4:0]  io_redirect_bits_robIdx_value,
  input         io_redirect_bits_level,
  output        io_enq_canAccept,
  input         io_enq_sqCanAccept,
  input         io_enq_req_0_valid,
  input         io_enq_req_0_bits_cf_trigger_backendEn_1,
  input  [6:0]  io_enq_req_0_bits_ctrl_fuOpType,
  input         io_enq_req_0_bits_ctrl_rfWen,
  input         io_enq_req_0_bits_ctrl_fpWen,
  input         io_enq_req_0_bits_ctrl_flushPipe,
  input         io_enq_req_0_bits_ctrl_replayInst,
  input  [5:0]  io_enq_req_0_bits_pdest,
  input         io_enq_req_0_bits_robIdx_flag,
  input  [4:0]  io_enq_req_0_bits_robIdx_value,
  input  [3:0]  io_enq_req_0_bits_lqIdx_value,
  input         io_enq_req_1_valid,
  input         io_enq_req_1_bits_cf_trigger_backendEn_1,
  input  [6:0]  io_enq_req_1_bits_ctrl_fuOpType,
  input         io_enq_req_1_bits_ctrl_rfWen,
  input         io_enq_req_1_bits_ctrl_fpWen,
  input         io_enq_req_1_bits_ctrl_flushPipe,
  input         io_enq_req_1_bits_ctrl_replayInst,
  input  [5:0]  io_enq_req_1_bits_pdest,
  input         io_enq_req_1_bits_robIdx_flag,
  input  [4:0]  io_enq_req_1_bits_robIdx_value,
  input  [3:0]  io_enq_req_1_bits_lqIdx_value,
  input         io_enq_req_2_valid,
  input         io_enq_req_2_bits_cf_trigger_backendEn_1,
  input  [6:0]  io_enq_req_2_bits_ctrl_fuOpType,
  input         io_enq_req_2_bits_ctrl_rfWen,
  input         io_enq_req_2_bits_ctrl_fpWen,
  input         io_enq_req_2_bits_ctrl_flushPipe,
  input         io_enq_req_2_bits_ctrl_replayInst,
  input  [5:0]  io_enq_req_2_bits_pdest,
  input         io_enq_req_2_bits_robIdx_flag,
  input  [4:0]  io_enq_req_2_bits_robIdx_value,
  input  [3:0]  io_enq_req_2_bits_lqIdx_value,
  input         io_enq_req_3_valid,
  input         io_enq_req_3_bits_cf_trigger_backendEn_1,
  input  [6:0]  io_enq_req_3_bits_ctrl_fuOpType,
  input         io_enq_req_3_bits_ctrl_rfWen,
  input         io_enq_req_3_bits_ctrl_fpWen,
  input         io_enq_req_3_bits_ctrl_flushPipe,
  input         io_enq_req_3_bits_ctrl_replayInst,
  input  [5:0]  io_enq_req_3_bits_pdest,
  input         io_enq_req_3_bits_robIdx_flag,
  input  [4:0]  io_enq_req_3_bits_robIdx_value,
  input  [3:0]  io_enq_req_3_bits_lqIdx_value,
  input         io_loadIn_0_valid,
  input         io_loadIn_0_bits_uop_cf_exceptionVec_4,
  input         io_loadIn_0_bits_uop_cf_exceptionVec_5,
  input         io_loadIn_0_bits_uop_cf_exceptionVec_13,
  input         io_loadIn_0_bits_uop_cf_trigger_backendEn_1,
  input         io_loadIn_0_bits_uop_cf_trigger_backendHit_0,
  input         io_loadIn_0_bits_uop_cf_trigger_backendHit_1,
  input         io_loadIn_0_bits_uop_cf_trigger_backendHit_4,
  input  [6:0]  io_loadIn_0_bits_uop_ctrl_fuOpType,
  input         io_loadIn_0_bits_uop_ctrl_rfWen,
  input         io_loadIn_0_bits_uop_ctrl_fpWen,
  input         io_loadIn_0_bits_uop_ctrl_replayInst,
  input  [5:0]  io_loadIn_0_bits_uop_pdest,
  input  [4:0]  io_loadIn_0_bits_uop_robIdx_value,
  input  [3:0]  io_loadIn_0_bits_uop_lqIdx_value,
  input  [38:0] io_loadIn_0_bits_vaddr,
  input  [35:0] io_loadIn_0_bits_paddr,
  input  [15:0] io_loadIn_0_bits_mask,
  input         io_loadIn_0_bits_miss,
  input         io_loadIn_0_bits_tlbMiss,
  input         io_loadIn_0_bits_mmio,
  input         io_loadIn_0_bits_replayInfo_cause_0,
  input         io_loadIn_0_bits_replayInfo_cause_1,
  input         io_loadIn_0_bits_replayInfo_cause_2,
  input         io_loadIn_0_bits_replayInfo_cause_3,
  input         io_loadIn_0_bits_replayInfo_cause_4,
  input         io_loadIn_0_bits_replayInfo_cause_5,
  input         io_loadIn_0_bits_replayInfo_cause_6,
  input         io_loadIn_0_bits_replayInfo_cause_7,
  input         io_loadIn_0_bits_lqDataWenDup_1,
  input         io_loadIn_0_bits_lqDataWenDup_2,
  input         io_loadIn_0_bits_lqDataWenDup_3,
  input         io_loadIn_0_bits_lqDataWenDup_5,
  input         io_loadIn_1_valid,
  input         io_loadIn_1_bits_uop_cf_exceptionVec_4,
  input         io_loadIn_1_bits_uop_cf_exceptionVec_5,
  input         io_loadIn_1_bits_uop_cf_exceptionVec_13,
  input         io_loadIn_1_bits_uop_cf_trigger_backendEn_1,
  input         io_loadIn_1_bits_uop_cf_trigger_backendHit_0,
  input         io_loadIn_1_bits_uop_cf_trigger_backendHit_1,
  input         io_loadIn_1_bits_uop_cf_trigger_backendHit_4,
  input  [6:0]  io_loadIn_1_bits_uop_ctrl_fuOpType,
  input         io_loadIn_1_bits_uop_ctrl_rfWen,
  input         io_loadIn_1_bits_uop_ctrl_fpWen,
  input         io_loadIn_1_bits_uop_ctrl_replayInst,
  input  [5:0]  io_loadIn_1_bits_uop_pdest,
  input  [4:0]  io_loadIn_1_bits_uop_robIdx_value,
  input  [3:0]  io_loadIn_1_bits_uop_lqIdx_value,
  input  [38:0] io_loadIn_1_bits_vaddr,
  input  [35:0] io_loadIn_1_bits_paddr,
  input  [15:0] io_loadIn_1_bits_mask,
  input         io_loadIn_1_bits_miss,
  input         io_loadIn_1_bits_tlbMiss,
  input         io_loadIn_1_bits_mmio,
  input         io_loadIn_1_bits_replayInfo_cause_0,
  input         io_loadIn_1_bits_replayInfo_cause_1,
  input         io_loadIn_1_bits_replayInfo_cause_2,
  input         io_loadIn_1_bits_replayInfo_cause_3,
  input         io_loadIn_1_bits_replayInfo_cause_4,
  input         io_loadIn_1_bits_replayInfo_cause_5,
  input         io_loadIn_1_bits_replayInfo_cause_6,
  input         io_loadIn_1_bits_replayInfo_cause_7,
  input         io_loadIn_1_bits_lqDataWenDup_1,
  input         io_loadIn_1_bits_lqDataWenDup_2,
  input         io_loadIn_1_bits_lqDataWenDup_3,
  input         io_loadIn_1_bits_lqDataWenDup_5,
  input         io_loadOut_0_ready,
  output        io_loadOut_0_valid,
  output        io_loadOut_0_bits_uop_cf_exceptionVec_4,
  output        io_loadOut_0_bits_uop_cf_exceptionVec_5,
  output        io_loadOut_0_bits_uop_cf_exceptionVec_13,
  output        io_loadOut_0_bits_uop_cf_trigger_backendEn_1,
  output        io_loadOut_0_bits_uop_cf_trigger_backendHit_0,
  output        io_loadOut_0_bits_uop_cf_trigger_backendHit_1,
  output        io_loadOut_0_bits_uop_cf_trigger_backendHit_4,
  output [6:0]  io_loadOut_0_bits_uop_ctrl_fuOpType,
  output        io_loadOut_0_bits_uop_ctrl_rfWen,
  output        io_loadOut_0_bits_uop_ctrl_fpWen,
  output        io_loadOut_0_bits_uop_ctrl_flushPipe,
  output        io_loadOut_0_bits_uop_ctrl_replayInst,
  output [5:0]  io_loadOut_0_bits_uop_pdest,
  output        io_loadOut_0_bits_uop_robIdx_flag,
  output [4:0]  io_loadOut_0_bits_uop_robIdx_value,
  output [63:0] io_ldRawDataOut_0_lqData,
  output [6:0]  io_ldRawDataOut_0_uop_ctrl_fuOpType,
  output        io_ldRawDataOut_0_uop_ctrl_fpWen,
  output [2:0]  io_ldRawDataOut_0_addrOffset,
  input         io_rob_pendingld,
  input         io_rob_commit,
  output        io_rob_isMMIO_0,
  output        io_rob_isMMIO_1,
  output [4:0]  io_rob_uop_0_robIdx_value,
  output [4:0]  io_rob_uop_1_robIdx_value,
  input         io_uncache_req_ready,
  output        io_uncache_req_valid,
  output [35:0] io_uncache_req_bits_addr,
  output [7:0]  io_uncache_req_bits_mask,
  output        io_uncache_resp_ready,
  input         io_uncache_resp_valid,
  input  [63:0] io_uncache_resp_bits_data,
  input         io_trigger_0_hitLoadAddrTriggerHitVec_0,
  input         io_trigger_0_hitLoadAddrTriggerHitVec_1,
  input         io_trigger_0_hitLoadAddrTriggerHitVec_2,
  output        io_trigger_0_lqLoadAddrTriggerHitVec_0,
  output        io_trigger_0_lqLoadAddrTriggerHitVec_1,
  output        io_trigger_0_lqLoadAddrTriggerHitVec_2,
  input         io_trigger_1_hitLoadAddrTriggerHitVec_0,
  input         io_trigger_1_hitLoadAddrTriggerHitVec_1,
  input         io_trigger_1_hitLoadAddrTriggerHitVec_2,
  output [38:0] io_exceptionAddr_vaddr,
  output        io_ldIssuePtr_flag,
  output [3:0]  io_ldIssuePtr_value,
  output [1:0]  io_lqDeq,
  output [4:0]  io_lqCancelCnt,
  output [5:0]  io_perf_0_value,
  output [5:0]  io_perf_1_value,
  output [5:0]  io_perf_2_value,
  output [5:0]  io_perf_3_value
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [63:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
`endif // RANDOMIZE_REG_INIT
  wire  vaddrModule_clock; // @[LoadQueueFlag.scala 63:27]
  wire [3:0] vaddrModule_io_raddr_1; // @[LoadQueueFlag.scala 63:27]
  wire [38:0] vaddrModule_io_rdata_1; // @[LoadQueueFlag.scala 63:27]
  wire  vaddrModule_io_wen_0; // @[LoadQueueFlag.scala 63:27]
  wire  vaddrModule_io_wen_1; // @[LoadQueueFlag.scala 63:27]
  wire [3:0] vaddrModule_io_waddr_0; // @[LoadQueueFlag.scala 63:27]
  wire [3:0] vaddrModule_io_waddr_1; // @[LoadQueueFlag.scala 63:27]
  wire [38:0] vaddrModule_io_wdata_0; // @[LoadQueueFlag.scala 63:27]
  wire [38:0] vaddrModule_io_wdata_1; // @[LoadQueueFlag.scala 63:27]
  wire  paddrModule_clock; // @[LoadQueueFlag.scala 72:27]
  wire [3:0] paddrModule_io_raddr_0; // @[LoadQueueFlag.scala 72:27]
  wire [35:0] paddrModule_io_rdata_0; // @[LoadQueueFlag.scala 72:27]
  wire  paddrModule_io_wen_0; // @[LoadQueueFlag.scala 72:27]
  wire  paddrModule_io_wen_1; // @[LoadQueueFlag.scala 72:27]
  wire [3:0] paddrModule_io_waddr_0; // @[LoadQueueFlag.scala 72:27]
  wire [3:0] paddrModule_io_waddr_1; // @[LoadQueueFlag.scala 72:27]
  wire [35:0] paddrModule_io_wdata_0; // @[LoadQueueFlag.scala 72:27]
  wire [35:0] paddrModule_io_wdata_1; // @[LoadQueueFlag.scala 72:27]
  wire  maskModule_clock; // @[LoadQueueFlag.scala 81:26]
  wire [3:0] maskModule_io_raddr_0; // @[LoadQueueFlag.scala 81:26]
  wire [7:0] maskModule_io_rdata_0; // @[LoadQueueFlag.scala 81:26]
  wire  maskModule_io_wen_0; // @[LoadQueueFlag.scala 81:26]
  wire  maskModule_io_wen_1; // @[LoadQueueFlag.scala 81:26]
  wire [3:0] maskModule_io_waddr_0; // @[LoadQueueFlag.scala 81:26]
  wire [3:0] maskModule_io_waddr_1; // @[LoadQueueFlag.scala 81:26]
  wire [7:0] maskModule_io_wdata_0; // @[LoadQueueFlag.scala 81:26]
  wire [7:0] maskModule_io_wdata_1; // @[LoadQueueFlag.scala 81:26]
  wire  vaddrTriggerResultModule_clock; // @[LoadQueueFlag.scala 105:40]
  wire [3:0] vaddrTriggerResultModule_io_raddr_0; // @[LoadQueueFlag.scala 105:40]
  wire  vaddrTriggerResultModule_io_rdata_0_0; // @[LoadQueueFlag.scala 105:40]
  wire  vaddrTriggerResultModule_io_rdata_0_1; // @[LoadQueueFlag.scala 105:40]
  wire  vaddrTriggerResultModule_io_rdata_0_2; // @[LoadQueueFlag.scala 105:40]
  wire  vaddrTriggerResultModule_io_wen_0; // @[LoadQueueFlag.scala 105:40]
  wire  vaddrTriggerResultModule_io_wen_1; // @[LoadQueueFlag.scala 105:40]
  wire [3:0] vaddrTriggerResultModule_io_waddr_0; // @[LoadQueueFlag.scala 105:40]
  wire [3:0] vaddrTriggerResultModule_io_waddr_1; // @[LoadQueueFlag.scala 105:40]
  wire  vaddrTriggerResultModule_io_wdata_0_0; // @[LoadQueueFlag.scala 105:40]
  wire  vaddrTriggerResultModule_io_wdata_0_1; // @[LoadQueueFlag.scala 105:40]
  wire  vaddrTriggerResultModule_io_wdata_0_2; // @[LoadQueueFlag.scala 105:40]
  wire  vaddrTriggerResultModule_io_wdata_1_0; // @[LoadQueueFlag.scala 105:40]
  wire  vaddrTriggerResultModule_io_wdata_1_1; // @[LoadQueueFlag.scala 105:40]
  wire  vaddrTriggerResultModule_io_wdata_1_2; // @[LoadQueueFlag.scala 105:40]
  reg  allocated_0; // @[LoadQueueFlag.scala 61:26]
  reg  allocated_1; // @[LoadQueueFlag.scala 61:26]
  reg  allocated_2; // @[LoadQueueFlag.scala 61:26]
  reg  allocated_3; // @[LoadQueueFlag.scala 61:26]
  reg  allocated_4; // @[LoadQueueFlag.scala 61:26]
  reg  allocated_5; // @[LoadQueueFlag.scala 61:26]
  reg  allocated_6; // @[LoadQueueFlag.scala 61:26]
  reg  allocated_7; // @[LoadQueueFlag.scala 61:26]
  reg  allocated_8; // @[LoadQueueFlag.scala 61:26]
  reg  allocated_9; // @[LoadQueueFlag.scala 61:26]
  reg  allocated_10; // @[LoadQueueFlag.scala 61:26]
  reg  allocated_11; // @[LoadQueueFlag.scala 61:26]
  reg  allocated_12; // @[LoadQueueFlag.scala 61:26]
  reg  allocated_13; // @[LoadQueueFlag.scala 61:26]
  reg  allocated_14; // @[LoadQueueFlag.scala 61:26]
  reg  allocated_15; // @[LoadQueueFlag.scala 61:26]
  reg  uop_0_cf_exceptionVec_4; // @[LoadQueueFlag.scala 62:16]
  reg  uop_0_cf_exceptionVec_5; // @[LoadQueueFlag.scala 62:16]
  reg  uop_0_cf_exceptionVec_13; // @[LoadQueueFlag.scala 62:16]
  reg  uop_0_cf_trigger_backendEn_1; // @[LoadQueueFlag.scala 62:16]
  reg  uop_0_cf_trigger_backendHit_0; // @[LoadQueueFlag.scala 62:16]
  reg  uop_0_cf_trigger_backendHit_1; // @[LoadQueueFlag.scala 62:16]
  reg  uop_0_cf_trigger_backendHit_4; // @[LoadQueueFlag.scala 62:16]
  reg [6:0] uop_0_ctrl_fuOpType; // @[LoadQueueFlag.scala 62:16]
  reg  uop_0_ctrl_rfWen; // @[LoadQueueFlag.scala 62:16]
  reg  uop_0_ctrl_fpWen; // @[LoadQueueFlag.scala 62:16]
  reg  uop_0_ctrl_flushPipe; // @[LoadQueueFlag.scala 62:16]
  reg  uop_0_ctrl_replayInst; // @[LoadQueueFlag.scala 62:16]
  reg [5:0] uop_0_pdest; // @[LoadQueueFlag.scala 62:16]
  reg  uop_0_robIdx_flag; // @[LoadQueueFlag.scala 62:16]
  reg [4:0] uop_0_robIdx_value; // @[LoadQueueFlag.scala 62:16]
  reg  uop_1_cf_exceptionVec_4; // @[LoadQueueFlag.scala 62:16]
  reg  uop_1_cf_exceptionVec_5; // @[LoadQueueFlag.scala 62:16]
  reg  uop_1_cf_exceptionVec_13; // @[LoadQueueFlag.scala 62:16]
  reg  uop_1_cf_trigger_backendEn_1; // @[LoadQueueFlag.scala 62:16]
  reg  uop_1_cf_trigger_backendHit_0; // @[LoadQueueFlag.scala 62:16]
  reg  uop_1_cf_trigger_backendHit_1; // @[LoadQueueFlag.scala 62:16]
  reg  uop_1_cf_trigger_backendHit_4; // @[LoadQueueFlag.scala 62:16]
  reg [6:0] uop_1_ctrl_fuOpType; // @[LoadQueueFlag.scala 62:16]
  reg  uop_1_ctrl_rfWen; // @[LoadQueueFlag.scala 62:16]
  reg  uop_1_ctrl_fpWen; // @[LoadQueueFlag.scala 62:16]
  reg  uop_1_ctrl_flushPipe; // @[LoadQueueFlag.scala 62:16]
  reg  uop_1_ctrl_replayInst; // @[LoadQueueFlag.scala 62:16]
  reg [5:0] uop_1_pdest; // @[LoadQueueFlag.scala 62:16]
  reg  uop_1_robIdx_flag; // @[LoadQueueFlag.scala 62:16]
  reg [4:0] uop_1_robIdx_value; // @[LoadQueueFlag.scala 62:16]
  reg  uop_2_cf_exceptionVec_4; // @[LoadQueueFlag.scala 62:16]
  reg  uop_2_cf_exceptionVec_5; // @[LoadQueueFlag.scala 62:16]
  reg  uop_2_cf_exceptionVec_13; // @[LoadQueueFlag.scala 62:16]
  reg  uop_2_cf_trigger_backendEn_1; // @[LoadQueueFlag.scala 62:16]
  reg  uop_2_cf_trigger_backendHit_0; // @[LoadQueueFlag.scala 62:16]
  reg  uop_2_cf_trigger_backendHit_1; // @[LoadQueueFlag.scala 62:16]
  reg  uop_2_cf_trigger_backendHit_4; // @[LoadQueueFlag.scala 62:16]
  reg [6:0] uop_2_ctrl_fuOpType; // @[LoadQueueFlag.scala 62:16]
  reg  uop_2_ctrl_rfWen; // @[LoadQueueFlag.scala 62:16]
  reg  uop_2_ctrl_fpWen; // @[LoadQueueFlag.scala 62:16]
  reg  uop_2_ctrl_flushPipe; // @[LoadQueueFlag.scala 62:16]
  reg  uop_2_ctrl_replayInst; // @[LoadQueueFlag.scala 62:16]
  reg [5:0] uop_2_pdest; // @[LoadQueueFlag.scala 62:16]
  reg  uop_2_robIdx_flag; // @[LoadQueueFlag.scala 62:16]
  reg [4:0] uop_2_robIdx_value; // @[LoadQueueFlag.scala 62:16]
  reg  uop_3_cf_exceptionVec_4; // @[LoadQueueFlag.scala 62:16]
  reg  uop_3_cf_exceptionVec_5; // @[LoadQueueFlag.scala 62:16]
  reg  uop_3_cf_exceptionVec_13; // @[LoadQueueFlag.scala 62:16]
  reg  uop_3_cf_trigger_backendEn_1; // @[LoadQueueFlag.scala 62:16]
  reg  uop_3_cf_trigger_backendHit_0; // @[LoadQueueFlag.scala 62:16]
  reg  uop_3_cf_trigger_backendHit_1; // @[LoadQueueFlag.scala 62:16]
  reg  uop_3_cf_trigger_backendHit_4; // @[LoadQueueFlag.scala 62:16]
  reg [6:0] uop_3_ctrl_fuOpType; // @[LoadQueueFlag.scala 62:16]
  reg  uop_3_ctrl_rfWen; // @[LoadQueueFlag.scala 62:16]
  reg  uop_3_ctrl_fpWen; // @[LoadQueueFlag.scala 62:16]
  reg  uop_3_ctrl_flushPipe; // @[LoadQueueFlag.scala 62:16]
  reg  uop_3_ctrl_replayInst; // @[LoadQueueFlag.scala 62:16]
  reg [5:0] uop_3_pdest; // @[LoadQueueFlag.scala 62:16]
  reg  uop_3_robIdx_flag; // @[LoadQueueFlag.scala 62:16]
  reg [4:0] uop_3_robIdx_value; // @[LoadQueueFlag.scala 62:16]
  reg  uop_4_cf_exceptionVec_4; // @[LoadQueueFlag.scala 62:16]
  reg  uop_4_cf_exceptionVec_5; // @[LoadQueueFlag.scala 62:16]
  reg  uop_4_cf_exceptionVec_13; // @[LoadQueueFlag.scala 62:16]
  reg  uop_4_cf_trigger_backendEn_1; // @[LoadQueueFlag.scala 62:16]
  reg  uop_4_cf_trigger_backendHit_0; // @[LoadQueueFlag.scala 62:16]
  reg  uop_4_cf_trigger_backendHit_1; // @[LoadQueueFlag.scala 62:16]
  reg  uop_4_cf_trigger_backendHit_4; // @[LoadQueueFlag.scala 62:16]
  reg [6:0] uop_4_ctrl_fuOpType; // @[LoadQueueFlag.scala 62:16]
  reg  uop_4_ctrl_rfWen; // @[LoadQueueFlag.scala 62:16]
  reg  uop_4_ctrl_fpWen; // @[LoadQueueFlag.scala 62:16]
  reg  uop_4_ctrl_flushPipe; // @[LoadQueueFlag.scala 62:16]
  reg  uop_4_ctrl_replayInst; // @[LoadQueueFlag.scala 62:16]
  reg [5:0] uop_4_pdest; // @[LoadQueueFlag.scala 62:16]
  reg  uop_4_robIdx_flag; // @[LoadQueueFlag.scala 62:16]
  reg [4:0] uop_4_robIdx_value; // @[LoadQueueFlag.scala 62:16]
  reg  uop_5_cf_exceptionVec_4; // @[LoadQueueFlag.scala 62:16]
  reg  uop_5_cf_exceptionVec_5; // @[LoadQueueFlag.scala 62:16]
  reg  uop_5_cf_exceptionVec_13; // @[LoadQueueFlag.scala 62:16]
  reg  uop_5_cf_trigger_backendEn_1; // @[LoadQueueFlag.scala 62:16]
  reg  uop_5_cf_trigger_backendHit_0; // @[LoadQueueFlag.scala 62:16]
  reg  uop_5_cf_trigger_backendHit_1; // @[LoadQueueFlag.scala 62:16]
  reg  uop_5_cf_trigger_backendHit_4; // @[LoadQueueFlag.scala 62:16]
  reg [6:0] uop_5_ctrl_fuOpType; // @[LoadQueueFlag.scala 62:16]
  reg  uop_5_ctrl_rfWen; // @[LoadQueueFlag.scala 62:16]
  reg  uop_5_ctrl_fpWen; // @[LoadQueueFlag.scala 62:16]
  reg  uop_5_ctrl_flushPipe; // @[LoadQueueFlag.scala 62:16]
  reg  uop_5_ctrl_replayInst; // @[LoadQueueFlag.scala 62:16]
  reg [5:0] uop_5_pdest; // @[LoadQueueFlag.scala 62:16]
  reg  uop_5_robIdx_flag; // @[LoadQueueFlag.scala 62:16]
  reg [4:0] uop_5_robIdx_value; // @[LoadQueueFlag.scala 62:16]
  reg  uop_6_cf_exceptionVec_4; // @[LoadQueueFlag.scala 62:16]
  reg  uop_6_cf_exceptionVec_5; // @[LoadQueueFlag.scala 62:16]
  reg  uop_6_cf_exceptionVec_13; // @[LoadQueueFlag.scala 62:16]
  reg  uop_6_cf_trigger_backendEn_1; // @[LoadQueueFlag.scala 62:16]
  reg  uop_6_cf_trigger_backendHit_0; // @[LoadQueueFlag.scala 62:16]
  reg  uop_6_cf_trigger_backendHit_1; // @[LoadQueueFlag.scala 62:16]
  reg  uop_6_cf_trigger_backendHit_4; // @[LoadQueueFlag.scala 62:16]
  reg [6:0] uop_6_ctrl_fuOpType; // @[LoadQueueFlag.scala 62:16]
  reg  uop_6_ctrl_rfWen; // @[LoadQueueFlag.scala 62:16]
  reg  uop_6_ctrl_fpWen; // @[LoadQueueFlag.scala 62:16]
  reg  uop_6_ctrl_flushPipe; // @[LoadQueueFlag.scala 62:16]
  reg  uop_6_ctrl_replayInst; // @[LoadQueueFlag.scala 62:16]
  reg [5:0] uop_6_pdest; // @[LoadQueueFlag.scala 62:16]
  reg  uop_6_robIdx_flag; // @[LoadQueueFlag.scala 62:16]
  reg [4:0] uop_6_robIdx_value; // @[LoadQueueFlag.scala 62:16]
  reg  uop_7_cf_exceptionVec_4; // @[LoadQueueFlag.scala 62:16]
  reg  uop_7_cf_exceptionVec_5; // @[LoadQueueFlag.scala 62:16]
  reg  uop_7_cf_exceptionVec_13; // @[LoadQueueFlag.scala 62:16]
  reg  uop_7_cf_trigger_backendEn_1; // @[LoadQueueFlag.scala 62:16]
  reg  uop_7_cf_trigger_backendHit_0; // @[LoadQueueFlag.scala 62:16]
  reg  uop_7_cf_trigger_backendHit_1; // @[LoadQueueFlag.scala 62:16]
  reg  uop_7_cf_trigger_backendHit_4; // @[LoadQueueFlag.scala 62:16]
  reg [6:0] uop_7_ctrl_fuOpType; // @[LoadQueueFlag.scala 62:16]
  reg  uop_7_ctrl_rfWen; // @[LoadQueueFlag.scala 62:16]
  reg  uop_7_ctrl_fpWen; // @[LoadQueueFlag.scala 62:16]
  reg  uop_7_ctrl_flushPipe; // @[LoadQueueFlag.scala 62:16]
  reg  uop_7_ctrl_replayInst; // @[LoadQueueFlag.scala 62:16]
  reg [5:0] uop_7_pdest; // @[LoadQueueFlag.scala 62:16]
  reg  uop_7_robIdx_flag; // @[LoadQueueFlag.scala 62:16]
  reg [4:0] uop_7_robIdx_value; // @[LoadQueueFlag.scala 62:16]
  reg  uop_8_cf_exceptionVec_4; // @[LoadQueueFlag.scala 62:16]
  reg  uop_8_cf_exceptionVec_5; // @[LoadQueueFlag.scala 62:16]
  reg  uop_8_cf_exceptionVec_13; // @[LoadQueueFlag.scala 62:16]
  reg  uop_8_cf_trigger_backendEn_1; // @[LoadQueueFlag.scala 62:16]
  reg  uop_8_cf_trigger_backendHit_0; // @[LoadQueueFlag.scala 62:16]
  reg  uop_8_cf_trigger_backendHit_1; // @[LoadQueueFlag.scala 62:16]
  reg  uop_8_cf_trigger_backendHit_4; // @[LoadQueueFlag.scala 62:16]
  reg [6:0] uop_8_ctrl_fuOpType; // @[LoadQueueFlag.scala 62:16]
  reg  uop_8_ctrl_rfWen; // @[LoadQueueFlag.scala 62:16]
  reg  uop_8_ctrl_fpWen; // @[LoadQueueFlag.scala 62:16]
  reg  uop_8_ctrl_flushPipe; // @[LoadQueueFlag.scala 62:16]
  reg  uop_8_ctrl_replayInst; // @[LoadQueueFlag.scala 62:16]
  reg [5:0] uop_8_pdest; // @[LoadQueueFlag.scala 62:16]
  reg  uop_8_robIdx_flag; // @[LoadQueueFlag.scala 62:16]
  reg [4:0] uop_8_robIdx_value; // @[LoadQueueFlag.scala 62:16]
  reg  uop_9_cf_exceptionVec_4; // @[LoadQueueFlag.scala 62:16]
  reg  uop_9_cf_exceptionVec_5; // @[LoadQueueFlag.scala 62:16]
  reg  uop_9_cf_exceptionVec_13; // @[LoadQueueFlag.scala 62:16]
  reg  uop_9_cf_trigger_backendEn_1; // @[LoadQueueFlag.scala 62:16]
  reg  uop_9_cf_trigger_backendHit_0; // @[LoadQueueFlag.scala 62:16]
  reg  uop_9_cf_trigger_backendHit_1; // @[LoadQueueFlag.scala 62:16]
  reg  uop_9_cf_trigger_backendHit_4; // @[LoadQueueFlag.scala 62:16]
  reg [6:0] uop_9_ctrl_fuOpType; // @[LoadQueueFlag.scala 62:16]
  reg  uop_9_ctrl_rfWen; // @[LoadQueueFlag.scala 62:16]
  reg  uop_9_ctrl_fpWen; // @[LoadQueueFlag.scala 62:16]
  reg  uop_9_ctrl_flushPipe; // @[LoadQueueFlag.scala 62:16]
  reg  uop_9_ctrl_replayInst; // @[LoadQueueFlag.scala 62:16]
  reg [5:0] uop_9_pdest; // @[LoadQueueFlag.scala 62:16]
  reg  uop_9_robIdx_flag; // @[LoadQueueFlag.scala 62:16]
  reg [4:0] uop_9_robIdx_value; // @[LoadQueueFlag.scala 62:16]
  reg  uop_10_cf_exceptionVec_4; // @[LoadQueueFlag.scala 62:16]
  reg  uop_10_cf_exceptionVec_5; // @[LoadQueueFlag.scala 62:16]
  reg  uop_10_cf_exceptionVec_13; // @[LoadQueueFlag.scala 62:16]
  reg  uop_10_cf_trigger_backendEn_1; // @[LoadQueueFlag.scala 62:16]
  reg  uop_10_cf_trigger_backendHit_0; // @[LoadQueueFlag.scala 62:16]
  reg  uop_10_cf_trigger_backendHit_1; // @[LoadQueueFlag.scala 62:16]
  reg  uop_10_cf_trigger_backendHit_4; // @[LoadQueueFlag.scala 62:16]
  reg [6:0] uop_10_ctrl_fuOpType; // @[LoadQueueFlag.scala 62:16]
  reg  uop_10_ctrl_rfWen; // @[LoadQueueFlag.scala 62:16]
  reg  uop_10_ctrl_fpWen; // @[LoadQueueFlag.scala 62:16]
  reg  uop_10_ctrl_flushPipe; // @[LoadQueueFlag.scala 62:16]
  reg  uop_10_ctrl_replayInst; // @[LoadQueueFlag.scala 62:16]
  reg [5:0] uop_10_pdest; // @[LoadQueueFlag.scala 62:16]
  reg  uop_10_robIdx_flag; // @[LoadQueueFlag.scala 62:16]
  reg [4:0] uop_10_robIdx_value; // @[LoadQueueFlag.scala 62:16]
  reg  uop_11_cf_exceptionVec_4; // @[LoadQueueFlag.scala 62:16]
  reg  uop_11_cf_exceptionVec_5; // @[LoadQueueFlag.scala 62:16]
  reg  uop_11_cf_exceptionVec_13; // @[LoadQueueFlag.scala 62:16]
  reg  uop_11_cf_trigger_backendEn_1; // @[LoadQueueFlag.scala 62:16]
  reg  uop_11_cf_trigger_backendHit_0; // @[LoadQueueFlag.scala 62:16]
  reg  uop_11_cf_trigger_backendHit_1; // @[LoadQueueFlag.scala 62:16]
  reg  uop_11_cf_trigger_backendHit_4; // @[LoadQueueFlag.scala 62:16]
  reg [6:0] uop_11_ctrl_fuOpType; // @[LoadQueueFlag.scala 62:16]
  reg  uop_11_ctrl_rfWen; // @[LoadQueueFlag.scala 62:16]
  reg  uop_11_ctrl_fpWen; // @[LoadQueueFlag.scala 62:16]
  reg  uop_11_ctrl_flushPipe; // @[LoadQueueFlag.scala 62:16]
  reg  uop_11_ctrl_replayInst; // @[LoadQueueFlag.scala 62:16]
  reg [5:0] uop_11_pdest; // @[LoadQueueFlag.scala 62:16]
  reg  uop_11_robIdx_flag; // @[LoadQueueFlag.scala 62:16]
  reg [4:0] uop_11_robIdx_value; // @[LoadQueueFlag.scala 62:16]
  reg  uop_12_cf_exceptionVec_4; // @[LoadQueueFlag.scala 62:16]
  reg  uop_12_cf_exceptionVec_5; // @[LoadQueueFlag.scala 62:16]
  reg  uop_12_cf_exceptionVec_13; // @[LoadQueueFlag.scala 62:16]
  reg  uop_12_cf_trigger_backendEn_1; // @[LoadQueueFlag.scala 62:16]
  reg  uop_12_cf_trigger_backendHit_0; // @[LoadQueueFlag.scala 62:16]
  reg  uop_12_cf_trigger_backendHit_1; // @[LoadQueueFlag.scala 62:16]
  reg  uop_12_cf_trigger_backendHit_4; // @[LoadQueueFlag.scala 62:16]
  reg [6:0] uop_12_ctrl_fuOpType; // @[LoadQueueFlag.scala 62:16]
  reg  uop_12_ctrl_rfWen; // @[LoadQueueFlag.scala 62:16]
  reg  uop_12_ctrl_fpWen; // @[LoadQueueFlag.scala 62:16]
  reg  uop_12_ctrl_flushPipe; // @[LoadQueueFlag.scala 62:16]
  reg  uop_12_ctrl_replayInst; // @[LoadQueueFlag.scala 62:16]
  reg [5:0] uop_12_pdest; // @[LoadQueueFlag.scala 62:16]
  reg  uop_12_robIdx_flag; // @[LoadQueueFlag.scala 62:16]
  reg [4:0] uop_12_robIdx_value; // @[LoadQueueFlag.scala 62:16]
  reg  uop_13_cf_exceptionVec_4; // @[LoadQueueFlag.scala 62:16]
  reg  uop_13_cf_exceptionVec_5; // @[LoadQueueFlag.scala 62:16]
  reg  uop_13_cf_exceptionVec_13; // @[LoadQueueFlag.scala 62:16]
  reg  uop_13_cf_trigger_backendEn_1; // @[LoadQueueFlag.scala 62:16]
  reg  uop_13_cf_trigger_backendHit_0; // @[LoadQueueFlag.scala 62:16]
  reg  uop_13_cf_trigger_backendHit_1; // @[LoadQueueFlag.scala 62:16]
  reg  uop_13_cf_trigger_backendHit_4; // @[LoadQueueFlag.scala 62:16]
  reg [6:0] uop_13_ctrl_fuOpType; // @[LoadQueueFlag.scala 62:16]
  reg  uop_13_ctrl_rfWen; // @[LoadQueueFlag.scala 62:16]
  reg  uop_13_ctrl_fpWen; // @[LoadQueueFlag.scala 62:16]
  reg  uop_13_ctrl_flushPipe; // @[LoadQueueFlag.scala 62:16]
  reg  uop_13_ctrl_replayInst; // @[LoadQueueFlag.scala 62:16]
  reg [5:0] uop_13_pdest; // @[LoadQueueFlag.scala 62:16]
  reg  uop_13_robIdx_flag; // @[LoadQueueFlag.scala 62:16]
  reg [4:0] uop_13_robIdx_value; // @[LoadQueueFlag.scala 62:16]
  reg  uop_14_cf_exceptionVec_4; // @[LoadQueueFlag.scala 62:16]
  reg  uop_14_cf_exceptionVec_5; // @[LoadQueueFlag.scala 62:16]
  reg  uop_14_cf_exceptionVec_13; // @[LoadQueueFlag.scala 62:16]
  reg  uop_14_cf_trigger_backendEn_1; // @[LoadQueueFlag.scala 62:16]
  reg  uop_14_cf_trigger_backendHit_0; // @[LoadQueueFlag.scala 62:16]
  reg  uop_14_cf_trigger_backendHit_1; // @[LoadQueueFlag.scala 62:16]
  reg  uop_14_cf_trigger_backendHit_4; // @[LoadQueueFlag.scala 62:16]
  reg [6:0] uop_14_ctrl_fuOpType; // @[LoadQueueFlag.scala 62:16]
  reg  uop_14_ctrl_rfWen; // @[LoadQueueFlag.scala 62:16]
  reg  uop_14_ctrl_fpWen; // @[LoadQueueFlag.scala 62:16]
  reg  uop_14_ctrl_flushPipe; // @[LoadQueueFlag.scala 62:16]
  reg  uop_14_ctrl_replayInst; // @[LoadQueueFlag.scala 62:16]
  reg [5:0] uop_14_pdest; // @[LoadQueueFlag.scala 62:16]
  reg  uop_14_robIdx_flag; // @[LoadQueueFlag.scala 62:16]
  reg [4:0] uop_14_robIdx_value; // @[LoadQueueFlag.scala 62:16]
  reg  uop_15_cf_exceptionVec_4; // @[LoadQueueFlag.scala 62:16]
  reg  uop_15_cf_exceptionVec_5; // @[LoadQueueFlag.scala 62:16]
  reg  uop_15_cf_exceptionVec_13; // @[LoadQueueFlag.scala 62:16]
  reg  uop_15_cf_trigger_backendEn_1; // @[LoadQueueFlag.scala 62:16]
  reg  uop_15_cf_trigger_backendHit_0; // @[LoadQueueFlag.scala 62:16]
  reg  uop_15_cf_trigger_backendHit_1; // @[LoadQueueFlag.scala 62:16]
  reg  uop_15_cf_trigger_backendHit_4; // @[LoadQueueFlag.scala 62:16]
  reg [6:0] uop_15_ctrl_fuOpType; // @[LoadQueueFlag.scala 62:16]
  reg  uop_15_ctrl_rfWen; // @[LoadQueueFlag.scala 62:16]
  reg  uop_15_ctrl_fpWen; // @[LoadQueueFlag.scala 62:16]
  reg  uop_15_ctrl_flushPipe; // @[LoadQueueFlag.scala 62:16]
  reg  uop_15_ctrl_replayInst; // @[LoadQueueFlag.scala 62:16]
  reg [5:0] uop_15_pdest; // @[LoadQueueFlag.scala 62:16]
  reg  uop_15_robIdx_flag; // @[LoadQueueFlag.scala 62:16]
  reg [4:0] uop_15_robIdx_value; // @[LoadQueueFlag.scala 62:16]
  reg  addrvalid_0; // @[LoadQueueFlag.scala 90:26]
  reg  addrvalid_1; // @[LoadQueueFlag.scala 90:26]
  reg  addrvalid_2; // @[LoadQueueFlag.scala 90:26]
  reg  addrvalid_3; // @[LoadQueueFlag.scala 90:26]
  reg  addrvalid_4; // @[LoadQueueFlag.scala 90:26]
  reg  addrvalid_5; // @[LoadQueueFlag.scala 90:26]
  reg  addrvalid_6; // @[LoadQueueFlag.scala 90:26]
  reg  addrvalid_7; // @[LoadQueueFlag.scala 90:26]
  reg  addrvalid_8; // @[LoadQueueFlag.scala 90:26]
  reg  addrvalid_9; // @[LoadQueueFlag.scala 90:26]
  reg  addrvalid_10; // @[LoadQueueFlag.scala 90:26]
  reg  addrvalid_11; // @[LoadQueueFlag.scala 90:26]
  reg  addrvalid_12; // @[LoadQueueFlag.scala 90:26]
  reg  addrvalid_13; // @[LoadQueueFlag.scala 90:26]
  reg  addrvalid_14; // @[LoadQueueFlag.scala 90:26]
  reg  addrvalid_15; // @[LoadQueueFlag.scala 90:26]
  reg  datavalid_0; // @[LoadQueueFlag.scala 91:26]
  reg  datavalid_1; // @[LoadQueueFlag.scala 91:26]
  reg  datavalid_2; // @[LoadQueueFlag.scala 91:26]
  reg  datavalid_3; // @[LoadQueueFlag.scala 91:26]
  reg  datavalid_4; // @[LoadQueueFlag.scala 91:26]
  reg  datavalid_5; // @[LoadQueueFlag.scala 91:26]
  reg  datavalid_6; // @[LoadQueueFlag.scala 91:26]
  reg  datavalid_7; // @[LoadQueueFlag.scala 91:26]
  reg  datavalid_8; // @[LoadQueueFlag.scala 91:26]
  reg  datavalid_9; // @[LoadQueueFlag.scala 91:26]
  reg  datavalid_10; // @[LoadQueueFlag.scala 91:26]
  reg  datavalid_11; // @[LoadQueueFlag.scala 91:26]
  reg  datavalid_12; // @[LoadQueueFlag.scala 91:26]
  reg  datavalid_13; // @[LoadQueueFlag.scala 91:26]
  reg  datavalid_14; // @[LoadQueueFlag.scala 91:26]
  reg  datavalid_15; // @[LoadQueueFlag.scala 91:26]
  reg  pending_0; // @[LoadQueueFlag.scala 92:24]
  reg  pending_1; // @[LoadQueueFlag.scala 92:24]
  reg  pending_2; // @[LoadQueueFlag.scala 92:24]
  reg  pending_3; // @[LoadQueueFlag.scala 92:24]
  reg  pending_4; // @[LoadQueueFlag.scala 92:24]
  reg  pending_5; // @[LoadQueueFlag.scala 92:24]
  reg  pending_6; // @[LoadQueueFlag.scala 92:24]
  reg  pending_7; // @[LoadQueueFlag.scala 92:24]
  reg  pending_8; // @[LoadQueueFlag.scala 92:24]
  reg  pending_9; // @[LoadQueueFlag.scala 92:24]
  reg  pending_10; // @[LoadQueueFlag.scala 92:24]
  reg  pending_11; // @[LoadQueueFlag.scala 92:24]
  reg  pending_12; // @[LoadQueueFlag.scala 92:24]
  reg  pending_13; // @[LoadQueueFlag.scala 92:24]
  reg  pending_14; // @[LoadQueueFlag.scala 92:24]
  reg  pending_15; // @[LoadQueueFlag.scala 92:24]
  reg  writebacked_0; // @[LoadQueueFlag.scala 93:28]
  reg  writebacked_1; // @[LoadQueueFlag.scala 93:28]
  reg  writebacked_2; // @[LoadQueueFlag.scala 93:28]
  reg  writebacked_3; // @[LoadQueueFlag.scala 93:28]
  reg  writebacked_4; // @[LoadQueueFlag.scala 93:28]
  reg  writebacked_5; // @[LoadQueueFlag.scala 93:28]
  reg  writebacked_6; // @[LoadQueueFlag.scala 93:28]
  reg  writebacked_7; // @[LoadQueueFlag.scala 93:28]
  reg  writebacked_8; // @[LoadQueueFlag.scala 93:28]
  reg  writebacked_9; // @[LoadQueueFlag.scala 93:28]
  reg  writebacked_10; // @[LoadQueueFlag.scala 93:28]
  reg  writebacked_11; // @[LoadQueueFlag.scala 93:28]
  reg  writebacked_12; // @[LoadQueueFlag.scala 93:28]
  reg  writebacked_13; // @[LoadQueueFlag.scala 93:28]
  reg  writebacked_14; // @[LoadQueueFlag.scala 93:28]
  reg  writebacked_15; // @[LoadQueueFlag.scala 93:28]
  reg  enqPtrExt_0_flag; // @[LoadQueueFlag.scala 116:26]
  reg [3:0] enqPtrExt_0_value; // @[LoadQueueFlag.scala 116:26]
  reg  lastCycleRedirect_valid; // @[LoadQueueFlag.scala 126:34]
  reg  deqPtrExt_rflag; // @[Reg.scala 28:20]
  reg [3:0] deqPtrExt_rvalue; // @[Reg.scala 28:20]
  wire [3:0] _validCount_T_2 = enqPtrExt_0_value - deqPtrExt_rvalue; // @[CircularQueuePtr.scala 81:21]
  wire [4:0] _GEN_31427 = {{1'd0}, enqPtrExt_0_value}; // @[CircularQueuePtr.scala 82:25]
  wire [4:0] _validCount_T_4 = 5'h10 + _GEN_31427; // @[CircularQueuePtr.scala 82:25]
  wire [4:0] _GEN_31428 = {{1'd0}, deqPtrExt_rvalue}; // @[CircularQueuePtr.scala 82:41]
  wire [4:0] _validCount_T_6 = _validCount_T_4 - _GEN_31428; // @[CircularQueuePtr.scala 82:41]
  wire [4:0] validCount = enqPtrExt_0_flag == deqPtrExt_rflag ? {{1'd0}, _validCount_T_2} : _validCount_T_6; // @[CircularQueuePtr.scala 80:8]
  wire [5:0] _needCancel_flushItself_T_1 = {uop_0_robIdx_flag,uop_0_robIdx_value}; // @[CircularQueuePtr.scala 61:50]
  wire [5:0] _needCancel_flushItself_T_2 = {io_redirect_bits_robIdx_flag,io_redirect_bits_robIdx_value}; // @[CircularQueuePtr.scala 61:70]
  wire  _needCancel_flushItself_T_3 = _needCancel_flushItself_T_1 == _needCancel_flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  needCancel_flushItself = io_redirect_bits_level & _needCancel_flushItself_T_3; // @[Rob.scala 122:51]
  wire  needCancel_differentFlag = uop_0_robIdx_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  needCancel_compare = uop_0_robIdx_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _needCancel_T = needCancel_differentFlag ^ needCancel_compare; // @[CircularQueuePtr.scala 88:19]
  wire  _needCancel_T_2 = io_redirect_valid & (needCancel_flushItself | _needCancel_T); // @[Rob.scala 123:20]
  wire  needCancel_0 = _needCancel_T_2 & allocated_0; // @[LoadQueueFlag.scala 133:42]
  wire [5:0] _needCancel_flushItself_T_5 = {uop_1_robIdx_flag,uop_1_robIdx_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _needCancel_flushItself_T_7 = _needCancel_flushItself_T_5 == _needCancel_flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  needCancel_flushItself_1 = io_redirect_bits_level & _needCancel_flushItself_T_7; // @[Rob.scala 122:51]
  wire  needCancel_differentFlag_1 = uop_1_robIdx_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  needCancel_compare_1 = uop_1_robIdx_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _needCancel_T_4 = needCancel_differentFlag_1 ^ needCancel_compare_1; // @[CircularQueuePtr.scala 88:19]
  wire  _needCancel_T_6 = io_redirect_valid & (needCancel_flushItself_1 | _needCancel_T_4); // @[Rob.scala 123:20]
  wire  needCancel_1 = _needCancel_T_6 & allocated_1; // @[LoadQueueFlag.scala 133:42]
  wire [5:0] _needCancel_flushItself_T_9 = {uop_2_robIdx_flag,uop_2_robIdx_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _needCancel_flushItself_T_11 = _needCancel_flushItself_T_9 == _needCancel_flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  needCancel_flushItself_2 = io_redirect_bits_level & _needCancel_flushItself_T_11; // @[Rob.scala 122:51]
  wire  needCancel_differentFlag_2 = uop_2_robIdx_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  needCancel_compare_2 = uop_2_robIdx_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _needCancel_T_8 = needCancel_differentFlag_2 ^ needCancel_compare_2; // @[CircularQueuePtr.scala 88:19]
  wire  _needCancel_T_10 = io_redirect_valid & (needCancel_flushItself_2 | _needCancel_T_8); // @[Rob.scala 123:20]
  wire  needCancel_2 = _needCancel_T_10 & allocated_2; // @[LoadQueueFlag.scala 133:42]
  wire [5:0] _needCancel_flushItself_T_13 = {uop_3_robIdx_flag,uop_3_robIdx_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _needCancel_flushItself_T_15 = _needCancel_flushItself_T_13 == _needCancel_flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  needCancel_flushItself_3 = io_redirect_bits_level & _needCancel_flushItself_T_15; // @[Rob.scala 122:51]
  wire  needCancel_differentFlag_3 = uop_3_robIdx_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  needCancel_compare_3 = uop_3_robIdx_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _needCancel_T_12 = needCancel_differentFlag_3 ^ needCancel_compare_3; // @[CircularQueuePtr.scala 88:19]
  wire  _needCancel_T_14 = io_redirect_valid & (needCancel_flushItself_3 | _needCancel_T_12); // @[Rob.scala 123:20]
  wire  needCancel_3 = _needCancel_T_14 & allocated_3; // @[LoadQueueFlag.scala 133:42]
  wire [5:0] _needCancel_flushItself_T_17 = {uop_4_robIdx_flag,uop_4_robIdx_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _needCancel_flushItself_T_19 = _needCancel_flushItself_T_17 == _needCancel_flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  needCancel_flushItself_4 = io_redirect_bits_level & _needCancel_flushItself_T_19; // @[Rob.scala 122:51]
  wire  needCancel_differentFlag_4 = uop_4_robIdx_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  needCancel_compare_4 = uop_4_robIdx_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _needCancel_T_16 = needCancel_differentFlag_4 ^ needCancel_compare_4; // @[CircularQueuePtr.scala 88:19]
  wire  _needCancel_T_18 = io_redirect_valid & (needCancel_flushItself_4 | _needCancel_T_16); // @[Rob.scala 123:20]
  wire  needCancel_4 = _needCancel_T_18 & allocated_4; // @[LoadQueueFlag.scala 133:42]
  wire [5:0] _needCancel_flushItself_T_21 = {uop_5_robIdx_flag,uop_5_robIdx_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _needCancel_flushItself_T_23 = _needCancel_flushItself_T_21 == _needCancel_flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  needCancel_flushItself_5 = io_redirect_bits_level & _needCancel_flushItself_T_23; // @[Rob.scala 122:51]
  wire  needCancel_differentFlag_5 = uop_5_robIdx_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  needCancel_compare_5 = uop_5_robIdx_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _needCancel_T_20 = needCancel_differentFlag_5 ^ needCancel_compare_5; // @[CircularQueuePtr.scala 88:19]
  wire  _needCancel_T_22 = io_redirect_valid & (needCancel_flushItself_5 | _needCancel_T_20); // @[Rob.scala 123:20]
  wire  needCancel_5 = _needCancel_T_22 & allocated_5; // @[LoadQueueFlag.scala 133:42]
  wire [5:0] _needCancel_flushItself_T_25 = {uop_6_robIdx_flag,uop_6_robIdx_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _needCancel_flushItself_T_27 = _needCancel_flushItself_T_25 == _needCancel_flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  needCancel_flushItself_6 = io_redirect_bits_level & _needCancel_flushItself_T_27; // @[Rob.scala 122:51]
  wire  needCancel_differentFlag_6 = uop_6_robIdx_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  needCancel_compare_6 = uop_6_robIdx_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _needCancel_T_24 = needCancel_differentFlag_6 ^ needCancel_compare_6; // @[CircularQueuePtr.scala 88:19]
  wire  _needCancel_T_26 = io_redirect_valid & (needCancel_flushItself_6 | _needCancel_T_24); // @[Rob.scala 123:20]
  wire  needCancel_6 = _needCancel_T_26 & allocated_6; // @[LoadQueueFlag.scala 133:42]
  wire [5:0] _needCancel_flushItself_T_29 = {uop_7_robIdx_flag,uop_7_robIdx_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _needCancel_flushItself_T_31 = _needCancel_flushItself_T_29 == _needCancel_flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  needCancel_flushItself_7 = io_redirect_bits_level & _needCancel_flushItself_T_31; // @[Rob.scala 122:51]
  wire  needCancel_differentFlag_7 = uop_7_robIdx_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  needCancel_compare_7 = uop_7_robIdx_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _needCancel_T_28 = needCancel_differentFlag_7 ^ needCancel_compare_7; // @[CircularQueuePtr.scala 88:19]
  wire  _needCancel_T_30 = io_redirect_valid & (needCancel_flushItself_7 | _needCancel_T_28); // @[Rob.scala 123:20]
  wire  needCancel_7 = _needCancel_T_30 & allocated_7; // @[LoadQueueFlag.scala 133:42]
  wire [5:0] _needCancel_flushItself_T_33 = {uop_8_robIdx_flag,uop_8_robIdx_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _needCancel_flushItself_T_35 = _needCancel_flushItself_T_33 == _needCancel_flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  needCancel_flushItself_8 = io_redirect_bits_level & _needCancel_flushItself_T_35; // @[Rob.scala 122:51]
  wire  needCancel_differentFlag_8 = uop_8_robIdx_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  needCancel_compare_8 = uop_8_robIdx_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _needCancel_T_32 = needCancel_differentFlag_8 ^ needCancel_compare_8; // @[CircularQueuePtr.scala 88:19]
  wire  _needCancel_T_34 = io_redirect_valid & (needCancel_flushItself_8 | _needCancel_T_32); // @[Rob.scala 123:20]
  wire  needCancel_8 = _needCancel_T_34 & allocated_8; // @[LoadQueueFlag.scala 133:42]
  wire [5:0] _needCancel_flushItself_T_37 = {uop_9_robIdx_flag,uop_9_robIdx_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _needCancel_flushItself_T_39 = _needCancel_flushItself_T_37 == _needCancel_flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  needCancel_flushItself_9 = io_redirect_bits_level & _needCancel_flushItself_T_39; // @[Rob.scala 122:51]
  wire  needCancel_differentFlag_9 = uop_9_robIdx_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  needCancel_compare_9 = uop_9_robIdx_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _needCancel_T_36 = needCancel_differentFlag_9 ^ needCancel_compare_9; // @[CircularQueuePtr.scala 88:19]
  wire  _needCancel_T_38 = io_redirect_valid & (needCancel_flushItself_9 | _needCancel_T_36); // @[Rob.scala 123:20]
  wire  needCancel_9 = _needCancel_T_38 & allocated_9; // @[LoadQueueFlag.scala 133:42]
  wire [5:0] _needCancel_flushItself_T_41 = {uop_10_robIdx_flag,uop_10_robIdx_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _needCancel_flushItself_T_43 = _needCancel_flushItself_T_41 == _needCancel_flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  needCancel_flushItself_10 = io_redirect_bits_level & _needCancel_flushItself_T_43; // @[Rob.scala 122:51]
  wire  needCancel_differentFlag_10 = uop_10_robIdx_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  needCancel_compare_10 = uop_10_robIdx_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _needCancel_T_40 = needCancel_differentFlag_10 ^ needCancel_compare_10; // @[CircularQueuePtr.scala 88:19]
  wire  _needCancel_T_42 = io_redirect_valid & (needCancel_flushItself_10 | _needCancel_T_40); // @[Rob.scala 123:20]
  wire  needCancel_10 = _needCancel_T_42 & allocated_10; // @[LoadQueueFlag.scala 133:42]
  wire [5:0] _needCancel_flushItself_T_45 = {uop_11_robIdx_flag,uop_11_robIdx_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _needCancel_flushItself_T_47 = _needCancel_flushItself_T_45 == _needCancel_flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  needCancel_flushItself_11 = io_redirect_bits_level & _needCancel_flushItself_T_47; // @[Rob.scala 122:51]
  wire  needCancel_differentFlag_11 = uop_11_robIdx_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  needCancel_compare_11 = uop_11_robIdx_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _needCancel_T_44 = needCancel_differentFlag_11 ^ needCancel_compare_11; // @[CircularQueuePtr.scala 88:19]
  wire  _needCancel_T_46 = io_redirect_valid & (needCancel_flushItself_11 | _needCancel_T_44); // @[Rob.scala 123:20]
  wire  needCancel_11 = _needCancel_T_46 & allocated_11; // @[LoadQueueFlag.scala 133:42]
  wire [5:0] _needCancel_flushItself_T_49 = {uop_12_robIdx_flag,uop_12_robIdx_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _needCancel_flushItself_T_51 = _needCancel_flushItself_T_49 == _needCancel_flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  needCancel_flushItself_12 = io_redirect_bits_level & _needCancel_flushItself_T_51; // @[Rob.scala 122:51]
  wire  needCancel_differentFlag_12 = uop_12_robIdx_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  needCancel_compare_12 = uop_12_robIdx_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _needCancel_T_48 = needCancel_differentFlag_12 ^ needCancel_compare_12; // @[CircularQueuePtr.scala 88:19]
  wire  _needCancel_T_50 = io_redirect_valid & (needCancel_flushItself_12 | _needCancel_T_48); // @[Rob.scala 123:20]
  wire  needCancel_12 = _needCancel_T_50 & allocated_12; // @[LoadQueueFlag.scala 133:42]
  wire [5:0] _needCancel_flushItself_T_53 = {uop_13_robIdx_flag,uop_13_robIdx_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _needCancel_flushItself_T_55 = _needCancel_flushItself_T_53 == _needCancel_flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  needCancel_flushItself_13 = io_redirect_bits_level & _needCancel_flushItself_T_55; // @[Rob.scala 122:51]
  wire  needCancel_differentFlag_13 = uop_13_robIdx_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  needCancel_compare_13 = uop_13_robIdx_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _needCancel_T_52 = needCancel_differentFlag_13 ^ needCancel_compare_13; // @[CircularQueuePtr.scala 88:19]
  wire  _needCancel_T_54 = io_redirect_valid & (needCancel_flushItself_13 | _needCancel_T_52); // @[Rob.scala 123:20]
  wire  needCancel_13 = _needCancel_T_54 & allocated_13; // @[LoadQueueFlag.scala 133:42]
  wire [5:0] _needCancel_flushItself_T_57 = {uop_14_robIdx_flag,uop_14_robIdx_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _needCancel_flushItself_T_59 = _needCancel_flushItself_T_57 == _needCancel_flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  needCancel_flushItself_14 = io_redirect_bits_level & _needCancel_flushItself_T_59; // @[Rob.scala 122:51]
  wire  needCancel_differentFlag_14 = uop_14_robIdx_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  needCancel_compare_14 = uop_14_robIdx_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _needCancel_T_56 = needCancel_differentFlag_14 ^ needCancel_compare_14; // @[CircularQueuePtr.scala 88:19]
  wire  _needCancel_T_58 = io_redirect_valid & (needCancel_flushItself_14 | _needCancel_T_56); // @[Rob.scala 123:20]
  wire  needCancel_14 = _needCancel_T_58 & allocated_14; // @[LoadQueueFlag.scala 133:42]
  wire [5:0] _needCancel_flushItself_T_61 = {uop_15_robIdx_flag,uop_15_robIdx_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _needCancel_flushItself_T_63 = _needCancel_flushItself_T_61 == _needCancel_flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  needCancel_flushItself_15 = io_redirect_bits_level & _needCancel_flushItself_T_63; // @[Rob.scala 122:51]
  wire  needCancel_differentFlag_15 = uop_15_robIdx_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  needCancel_compare_15 = uop_15_robIdx_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _needCancel_T_60 = needCancel_differentFlag_15 ^ needCancel_compare_15; // @[CircularQueuePtr.scala 88:19]
  wire  _needCancel_T_62 = io_redirect_valid & (needCancel_flushItself_15 | _needCancel_T_60); // @[Rob.scala 123:20]
  wire  needCancel_15 = _needCancel_T_62 & allocated_15; // @[LoadQueueFlag.scala 133:42]
  reg  lastNeedCancel_0; // @[LoadQueueFlag.scala 135:31]
  reg  lastNeedCancel_1; // @[LoadQueueFlag.scala 135:31]
  reg  lastNeedCancel_2; // @[LoadQueueFlag.scala 135:31]
  reg  lastNeedCancel_3; // @[LoadQueueFlag.scala 135:31]
  reg  lastNeedCancel_4; // @[LoadQueueFlag.scala 135:31]
  reg  lastNeedCancel_5; // @[LoadQueueFlag.scala 135:31]
  reg  lastNeedCancel_6; // @[LoadQueueFlag.scala 135:31]
  reg  lastNeedCancel_7; // @[LoadQueueFlag.scala 135:31]
  reg  lastNeedCancel_8; // @[LoadQueueFlag.scala 135:31]
  reg  lastNeedCancel_9; // @[LoadQueueFlag.scala 135:31]
  reg  lastNeedCancel_10; // @[LoadQueueFlag.scala 135:31]
  reg  lastNeedCancel_11; // @[LoadQueueFlag.scala 135:31]
  reg  lastNeedCancel_12; // @[LoadQueueFlag.scala 135:31]
  reg  lastNeedCancel_13; // @[LoadQueueFlag.scala 135:31]
  reg  lastNeedCancel_14; // @[LoadQueueFlag.scala 135:31]
  reg  lastNeedCancel_15; // @[LoadQueueFlag.scala 135:31]
  wire [5:0] _enqCancel_flushItself_T_1 = {io_enq_req_0_bits_robIdx_flag,io_enq_req_0_bits_robIdx_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _enqCancel_flushItself_T_3 = _enqCancel_flushItself_T_1 == _needCancel_flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  enqCancel_flushItself = io_redirect_bits_level & _enqCancel_flushItself_T_3; // @[Rob.scala 122:51]
  wire  enqCancel_differentFlag = io_enq_req_0_bits_robIdx_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  enqCancel_compare = io_enq_req_0_bits_robIdx_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _enqCancel_T = enqCancel_differentFlag ^ enqCancel_compare; // @[CircularQueuePtr.scala 88:19]
  wire  enqCancel_0 = io_redirect_valid & (enqCancel_flushItself | _enqCancel_T); // @[Rob.scala 123:20]
  wire [5:0] _enqCancel_flushItself_T_5 = {io_enq_req_1_bits_robIdx_flag,io_enq_req_1_bits_robIdx_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _enqCancel_flushItself_T_7 = _enqCancel_flushItself_T_5 == _needCancel_flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  enqCancel_flushItself_1 = io_redirect_bits_level & _enqCancel_flushItself_T_7; // @[Rob.scala 122:51]
  wire  enqCancel_differentFlag_1 = io_enq_req_1_bits_robIdx_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  enqCancel_compare_1 = io_enq_req_1_bits_robIdx_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _enqCancel_T_2 = enqCancel_differentFlag_1 ^ enqCancel_compare_1; // @[CircularQueuePtr.scala 88:19]
  wire  enqCancel_1 = io_redirect_valid & (enqCancel_flushItself_1 | _enqCancel_T_2); // @[Rob.scala 123:20]
  wire [5:0] _enqCancel_flushItself_T_9 = {io_enq_req_2_bits_robIdx_flag,io_enq_req_2_bits_robIdx_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _enqCancel_flushItself_T_11 = _enqCancel_flushItself_T_9 == _needCancel_flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  enqCancel_flushItself_2 = io_redirect_bits_level & _enqCancel_flushItself_T_11; // @[Rob.scala 122:51]
  wire  enqCancel_differentFlag_2 = io_enq_req_2_bits_robIdx_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  enqCancel_compare_2 = io_enq_req_2_bits_robIdx_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _enqCancel_T_4 = enqCancel_differentFlag_2 ^ enqCancel_compare_2; // @[CircularQueuePtr.scala 88:19]
  wire  enqCancel_2 = io_redirect_valid & (enqCancel_flushItself_2 | _enqCancel_T_4); // @[Rob.scala 123:20]
  wire [5:0] _enqCancel_flushItself_T_13 = {io_enq_req_3_bits_robIdx_flag,io_enq_req_3_bits_robIdx_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _enqCancel_flushItself_T_15 = _enqCancel_flushItself_T_13 == _needCancel_flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  enqCancel_flushItself_3 = io_redirect_bits_level & _enqCancel_flushItself_T_15; // @[Rob.scala 122:51]
  wire  enqCancel_differentFlag_3 = io_enq_req_3_bits_robIdx_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  enqCancel_compare_3 = io_enq_req_3_bits_robIdx_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _enqCancel_T_6 = enqCancel_differentFlag_3 ^ enqCancel_compare_3; // @[CircularQueuePtr.scala 88:19]
  wire  enqCancel_3 = io_redirect_valid & (enqCancel_flushItself_3 | _enqCancel_T_6); // @[Rob.scala 123:20]
  reg  lastEnqCancel_REG_0; // @[LoadQueueFlag.scala 137:39]
  reg  lastEnqCancel_REG_1; // @[LoadQueueFlag.scala 137:39]
  reg  lastEnqCancel_REG_2; // @[LoadQueueFlag.scala 137:39]
  reg  lastEnqCancel_REG_3; // @[LoadQueueFlag.scala 137:39]
  wire [1:0] _lastEnqCancel_T_4 = lastEnqCancel_REG_0 + lastEnqCancel_REG_1; // @[Bitwise.scala 48:55]
  wire [1:0] _lastEnqCancel_T_6 = lastEnqCancel_REG_2 + lastEnqCancel_REG_3; // @[Bitwise.scala 48:55]
  wire [2:0] lastEnqCancel = _lastEnqCancel_T_4 + _lastEnqCancel_T_6; // @[Bitwise.scala 48:55]
  wire [1:0] _lastCycleCancelCount_T = lastNeedCancel_0 + lastNeedCancel_1; // @[Bitwise.scala 48:55]
  wire [1:0] _lastCycleCancelCount_T_2 = lastNeedCancel_2 + lastNeedCancel_3; // @[Bitwise.scala 48:55]
  wire [2:0] _lastCycleCancelCount_T_4 = _lastCycleCancelCount_T + _lastCycleCancelCount_T_2; // @[Bitwise.scala 48:55]
  wire [1:0] _lastCycleCancelCount_T_6 = lastNeedCancel_4 + lastNeedCancel_5; // @[Bitwise.scala 48:55]
  wire [1:0] _lastCycleCancelCount_T_8 = lastNeedCancel_6 + lastNeedCancel_7; // @[Bitwise.scala 48:55]
  wire [2:0] _lastCycleCancelCount_T_10 = _lastCycleCancelCount_T_6 + _lastCycleCancelCount_T_8; // @[Bitwise.scala 48:55]
  wire [3:0] _lastCycleCancelCount_T_12 = _lastCycleCancelCount_T_4 + _lastCycleCancelCount_T_10; // @[Bitwise.scala 48:55]
  wire [1:0] _lastCycleCancelCount_T_14 = lastNeedCancel_8 + lastNeedCancel_9; // @[Bitwise.scala 48:55]
  wire [1:0] _lastCycleCancelCount_T_16 = lastNeedCancel_10 + lastNeedCancel_11; // @[Bitwise.scala 48:55]
  wire [2:0] _lastCycleCancelCount_T_18 = _lastCycleCancelCount_T_14 + _lastCycleCancelCount_T_16; // @[Bitwise.scala 48:55]
  wire [1:0] _lastCycleCancelCount_T_20 = lastNeedCancel_12 + lastNeedCancel_13; // @[Bitwise.scala 48:55]
  wire [1:0] _lastCycleCancelCount_T_22 = lastNeedCancel_14 + lastNeedCancel_15; // @[Bitwise.scala 48:55]
  wire [2:0] _lastCycleCancelCount_T_24 = _lastCycleCancelCount_T_20 + _lastCycleCancelCount_T_22; // @[Bitwise.scala 48:55]
  wire [3:0] _lastCycleCancelCount_T_26 = _lastCycleCancelCount_T_18 + _lastCycleCancelCount_T_24; // @[Bitwise.scala 48:55]
  wire [4:0] lastCycleCancelCount = _lastCycleCancelCount_T_12 + _lastCycleCancelCount_T_26; // @[Bitwise.scala 48:55]
  wire [1:0] _enqCount_T_1 = io_enq_req_0_valid + io_enq_req_1_valid; // @[Bitwise.scala 48:55]
  wire [1:0] _enqCount_T_3 = io_enq_req_2_valid + io_enq_req_3_valid; // @[Bitwise.scala 48:55]
  wire [2:0] _enqCount_T_5 = _enqCount_T_1 + _enqCount_T_3; // @[Bitwise.scala 48:55]
  wire [2:0] enqCount = io_enq_canAccept & io_enq_sqCanAccept ? _enqCount_T_5 : 3'h0; // @[LoadQueueFlag.scala 139:21]
  wire [4:0] _GEN_31429 = {{2'd0}, lastEnqCancel}; // @[LoadQueueFlag.scala 143:70]
  wire [4:0] _T_1 = lastCycleCancelCount + _GEN_31429; // @[LoadQueueFlag.scala 143:70]
  wire [4:0] _flipped_new_ptr_T_1 = 5'h10 - _T_1; // @[CircularQueuePtr.scala 54:50]
  wire [4:0] _flipped_new_ptr_new_ptr_T = {enqPtrExt_0_flag,enqPtrExt_0_value}; // @[Cat.scala 31:58]
  wire [4:0] _flipped_new_ptr_new_ptr_T_2 = _flipped_new_ptr_new_ptr_T + _flipped_new_ptr_T_1; // @[CircularQueuePtr.scala 39:46]
  wire [3:0] flipped_new_ptr_value = _flipped_new_ptr_new_ptr_T_2[3:0]; // @[CircularQueuePtr.scala 39:59]
  wire  flipped_new_ptr_flag = _flipped_new_ptr_new_ptr_T_2[4]; // @[CircularQueuePtr.scala 39:59]
  wire  new_ptr_flag = ~flipped_new_ptr_flag; // @[CircularQueuePtr.scala 56:21]
  wire [4:0] _GEN_31433 = {{2'd0}, enqCount}; // @[CircularQueuePtr.scala 39:46]
  wire [4:0] _new_ptr_T_2 = _flipped_new_ptr_new_ptr_T + _GEN_31433; // @[CircularQueuePtr.scala 39:46]
  wire [3:0] new_ptr_4_value = _new_ptr_T_2[3:0]; // @[CircularQueuePtr.scala 39:59]
  wire  new_ptr_4_flag = _new_ptr_T_2[4]; // @[CircularQueuePtr.scala 39:59]
  wire [4:0] _deqLookupVec_new_ptr_T = {deqPtrExt_rflag,deqPtrExt_rvalue}; // @[Cat.scala 31:58]
  wire [5:0] _deqLookupVec_new_ptr_T_1 = {{1'd0}, _deqLookupVec_new_ptr_T}; // @[CircularQueuePtr.scala 39:46]
  wire [3:0] deqLookupVec_new_ptr_value = _deqLookupVec_new_ptr_T_1[3:0]; // @[CircularQueuePtr.scala 39:59]
  wire  deqLookupVec_new_ptr_flag = _deqLookupVec_new_ptr_T_1[4]; // @[CircularQueuePtr.scala 39:59]
  wire [4:0] _deqLookupVec_new_ptr_T_7 = _deqLookupVec_new_ptr_T + 5'h1; // @[CircularQueuePtr.scala 39:46]
  wire [3:0] deqLookupVec_new_ptr_1_value = _deqLookupVec_new_ptr_T_7[3:0]; // @[CircularQueuePtr.scala 39:59]
  wire  deqLookupVec_new_ptr_1_flag = _deqLookupVec_new_ptr_T_7[4]; // @[CircularQueuePtr.scala 39:59]
  wire  _GEN_9 = 4'h1 == deqLookupVec_new_ptr_value ? allocated_1 : allocated_0; // @[LoadQueueFlag.scala 153:{72,72}]
  wire  _GEN_10 = 4'h2 == deqLookupVec_new_ptr_value ? allocated_2 : _GEN_9; // @[LoadQueueFlag.scala 153:{72,72}]
  wire  _GEN_11 = 4'h3 == deqLookupVec_new_ptr_value ? allocated_3 : _GEN_10; // @[LoadQueueFlag.scala 153:{72,72}]
  wire  _GEN_12 = 4'h4 == deqLookupVec_new_ptr_value ? allocated_4 : _GEN_11; // @[LoadQueueFlag.scala 153:{72,72}]
  wire  _GEN_13 = 4'h5 == deqLookupVec_new_ptr_value ? allocated_5 : _GEN_12; // @[LoadQueueFlag.scala 153:{72,72}]
  wire  _GEN_14 = 4'h6 == deqLookupVec_new_ptr_value ? allocated_6 : _GEN_13; // @[LoadQueueFlag.scala 153:{72,72}]
  wire  _GEN_15 = 4'h7 == deqLookupVec_new_ptr_value ? allocated_7 : _GEN_14; // @[LoadQueueFlag.scala 153:{72,72}]
  wire  _GEN_16 = 4'h8 == deqLookupVec_new_ptr_value ? allocated_8 : _GEN_15; // @[LoadQueueFlag.scala 153:{72,72}]
  wire  _GEN_17 = 4'h9 == deqLookupVec_new_ptr_value ? allocated_9 : _GEN_16; // @[LoadQueueFlag.scala 153:{72,72}]
  wire  _GEN_18 = 4'ha == deqLookupVec_new_ptr_value ? allocated_10 : _GEN_17; // @[LoadQueueFlag.scala 153:{72,72}]
  wire  _GEN_19 = 4'hb == deqLookupVec_new_ptr_value ? allocated_11 : _GEN_18; // @[LoadQueueFlag.scala 153:{72,72}]
  wire  _GEN_20 = 4'hc == deqLookupVec_new_ptr_value ? allocated_12 : _GEN_19; // @[LoadQueueFlag.scala 153:{72,72}]
  wire  _GEN_21 = 4'hd == deqLookupVec_new_ptr_value ? allocated_13 : _GEN_20; // @[LoadQueueFlag.scala 153:{72,72}]
  wire  _GEN_22 = 4'he == deqLookupVec_new_ptr_value ? allocated_14 : _GEN_21; // @[LoadQueueFlag.scala 153:{72,72}]
  wire  _GEN_23 = 4'hf == deqLookupVec_new_ptr_value ? allocated_15 : _GEN_22; // @[LoadQueueFlag.scala 153:{72,72}]
  wire  _GEN_25 = 4'h1 == deqLookupVec_new_ptr_value ? datavalid_1 : datavalid_0; // @[LoadQueueFlag.scala 153:{72,72}]
  wire  _GEN_26 = 4'h2 == deqLookupVec_new_ptr_value ? datavalid_2 : _GEN_25; // @[LoadQueueFlag.scala 153:{72,72}]
  wire  _GEN_27 = 4'h3 == deqLookupVec_new_ptr_value ? datavalid_3 : _GEN_26; // @[LoadQueueFlag.scala 153:{72,72}]
  wire  _GEN_28 = 4'h4 == deqLookupVec_new_ptr_value ? datavalid_4 : _GEN_27; // @[LoadQueueFlag.scala 153:{72,72}]
  wire  _GEN_29 = 4'h5 == deqLookupVec_new_ptr_value ? datavalid_5 : _GEN_28; // @[LoadQueueFlag.scala 153:{72,72}]
  wire  _GEN_30 = 4'h6 == deqLookupVec_new_ptr_value ? datavalid_6 : _GEN_29; // @[LoadQueueFlag.scala 153:{72,72}]
  wire  _GEN_31 = 4'h7 == deqLookupVec_new_ptr_value ? datavalid_7 : _GEN_30; // @[LoadQueueFlag.scala 153:{72,72}]
  wire  _GEN_32 = 4'h8 == deqLookupVec_new_ptr_value ? datavalid_8 : _GEN_31; // @[LoadQueueFlag.scala 153:{72,72}]
  wire  _GEN_33 = 4'h9 == deqLookupVec_new_ptr_value ? datavalid_9 : _GEN_32; // @[LoadQueueFlag.scala 153:{72,72}]
  wire  _GEN_34 = 4'ha == deqLookupVec_new_ptr_value ? datavalid_10 : _GEN_33; // @[LoadQueueFlag.scala 153:{72,72}]
  wire  _GEN_35 = 4'hb == deqLookupVec_new_ptr_value ? datavalid_11 : _GEN_34; // @[LoadQueueFlag.scala 153:{72,72}]
  wire  _GEN_36 = 4'hc == deqLookupVec_new_ptr_value ? datavalid_12 : _GEN_35; // @[LoadQueueFlag.scala 153:{72,72}]
  wire  _GEN_37 = 4'hd == deqLookupVec_new_ptr_value ? datavalid_13 : _GEN_36; // @[LoadQueueFlag.scala 153:{72,72}]
  wire  _GEN_38 = 4'he == deqLookupVec_new_ptr_value ? datavalid_14 : _GEN_37; // @[LoadQueueFlag.scala 153:{72,72}]
  wire  _GEN_39 = 4'hf == deqLookupVec_new_ptr_value ? datavalid_15 : _GEN_38; // @[LoadQueueFlag.scala 153:{72,72}]
  wire  _GEN_41 = 4'h1 == deqLookupVec_new_ptr_value ? addrvalid_1 : addrvalid_0; // @[LoadQueueFlag.scala 153:{96,96}]
  wire  _GEN_42 = 4'h2 == deqLookupVec_new_ptr_value ? addrvalid_2 : _GEN_41; // @[LoadQueueFlag.scala 153:{96,96}]
  wire  _GEN_43 = 4'h3 == deqLookupVec_new_ptr_value ? addrvalid_3 : _GEN_42; // @[LoadQueueFlag.scala 153:{96,96}]
  wire  _GEN_44 = 4'h4 == deqLookupVec_new_ptr_value ? addrvalid_4 : _GEN_43; // @[LoadQueueFlag.scala 153:{96,96}]
  wire  _GEN_45 = 4'h5 == deqLookupVec_new_ptr_value ? addrvalid_5 : _GEN_44; // @[LoadQueueFlag.scala 153:{96,96}]
  wire  _GEN_46 = 4'h6 == deqLookupVec_new_ptr_value ? addrvalid_6 : _GEN_45; // @[LoadQueueFlag.scala 153:{96,96}]
  wire  _GEN_47 = 4'h7 == deqLookupVec_new_ptr_value ? addrvalid_7 : _GEN_46; // @[LoadQueueFlag.scala 153:{96,96}]
  wire  _GEN_48 = 4'h8 == deqLookupVec_new_ptr_value ? addrvalid_8 : _GEN_47; // @[LoadQueueFlag.scala 153:{96,96}]
  wire  _GEN_49 = 4'h9 == deqLookupVec_new_ptr_value ? addrvalid_9 : _GEN_48; // @[LoadQueueFlag.scala 153:{96,96}]
  wire  _GEN_50 = 4'ha == deqLookupVec_new_ptr_value ? addrvalid_10 : _GEN_49; // @[LoadQueueFlag.scala 153:{96,96}]
  wire  _GEN_51 = 4'hb == deqLookupVec_new_ptr_value ? addrvalid_11 : _GEN_50; // @[LoadQueueFlag.scala 153:{96,96}]
  wire  _GEN_52 = 4'hc == deqLookupVec_new_ptr_value ? addrvalid_12 : _GEN_51; // @[LoadQueueFlag.scala 153:{96,96}]
  wire  _GEN_53 = 4'hd == deqLookupVec_new_ptr_value ? addrvalid_13 : _GEN_52; // @[LoadQueueFlag.scala 153:{96,96}]
  wire  _GEN_54 = 4'he == deqLookupVec_new_ptr_value ? addrvalid_14 : _GEN_53; // @[LoadQueueFlag.scala 153:{96,96}]
  wire  _GEN_55 = 4'hf == deqLookupVec_new_ptr_value ? addrvalid_15 : _GEN_54; // @[LoadQueueFlag.scala 153:{96,96}]
  wire  _GEN_57 = 4'h1 == deqLookupVec_new_ptr_value ? writebacked_1 : writebacked_0; // @[LoadQueueFlag.scala 153:{121,121}]
  wire  _GEN_58 = 4'h2 == deqLookupVec_new_ptr_value ? writebacked_2 : _GEN_57; // @[LoadQueueFlag.scala 153:{121,121}]
  wire  _GEN_59 = 4'h3 == deqLookupVec_new_ptr_value ? writebacked_3 : _GEN_58; // @[LoadQueueFlag.scala 153:{121,121}]
  wire  _GEN_60 = 4'h4 == deqLookupVec_new_ptr_value ? writebacked_4 : _GEN_59; // @[LoadQueueFlag.scala 153:{121,121}]
  wire  _GEN_61 = 4'h5 == deqLookupVec_new_ptr_value ? writebacked_5 : _GEN_60; // @[LoadQueueFlag.scala 153:{121,121}]
  wire  _GEN_62 = 4'h6 == deqLookupVec_new_ptr_value ? writebacked_6 : _GEN_61; // @[LoadQueueFlag.scala 153:{121,121}]
  wire  _GEN_63 = 4'h7 == deqLookupVec_new_ptr_value ? writebacked_7 : _GEN_62; // @[LoadQueueFlag.scala 153:{121,121}]
  wire  _GEN_64 = 4'h8 == deqLookupVec_new_ptr_value ? writebacked_8 : _GEN_63; // @[LoadQueueFlag.scala 153:{121,121}]
  wire  _GEN_65 = 4'h9 == deqLookupVec_new_ptr_value ? writebacked_9 : _GEN_64; // @[LoadQueueFlag.scala 153:{121,121}]
  wire  _GEN_66 = 4'ha == deqLookupVec_new_ptr_value ? writebacked_10 : _GEN_65; // @[LoadQueueFlag.scala 153:{121,121}]
  wire  _GEN_67 = 4'hb == deqLookupVec_new_ptr_value ? writebacked_11 : _GEN_66; // @[LoadQueueFlag.scala 153:{121,121}]
  wire  _GEN_68 = 4'hc == deqLookupVec_new_ptr_value ? writebacked_12 : _GEN_67; // @[LoadQueueFlag.scala 153:{121,121}]
  wire  _GEN_69 = 4'hd == deqLookupVec_new_ptr_value ? writebacked_13 : _GEN_68; // @[LoadQueueFlag.scala 153:{121,121}]
  wire  _GEN_70 = 4'he == deqLookupVec_new_ptr_value ? writebacked_14 : _GEN_69; // @[LoadQueueFlag.scala 153:{121,121}]
  wire  _GEN_71 = 4'hf == deqLookupVec_new_ptr_value ? writebacked_15 : _GEN_70; // @[LoadQueueFlag.scala 153:{121,121}]
  wire [4:0] _deqLookup_T_3 = {deqLookupVec_new_ptr_flag,deqLookupVec_new_ptr_value}; // @[CircularQueuePtr.scala 63:50]
  wire  _deqLookup_T_5 = _deqLookup_T_3 != _flipped_new_ptr_new_ptr_T; // @[CircularQueuePtr.scala 63:52]
  wire  deqLookup_0 = _GEN_23 & _GEN_39 & _GEN_55 & _GEN_71 & _deqLookup_T_5; // @[LoadQueueFlag.scala 153:147]
  wire  _GEN_73 = 4'h1 == deqLookupVec_new_ptr_1_value ? allocated_1 : allocated_0; // @[LoadQueueFlag.scala 153:{72,72}]
  wire  _GEN_74 = 4'h2 == deqLookupVec_new_ptr_1_value ? allocated_2 : _GEN_73; // @[LoadQueueFlag.scala 153:{72,72}]
  wire  _GEN_75 = 4'h3 == deqLookupVec_new_ptr_1_value ? allocated_3 : _GEN_74; // @[LoadQueueFlag.scala 153:{72,72}]
  wire  _GEN_76 = 4'h4 == deqLookupVec_new_ptr_1_value ? allocated_4 : _GEN_75; // @[LoadQueueFlag.scala 153:{72,72}]
  wire  _GEN_77 = 4'h5 == deqLookupVec_new_ptr_1_value ? allocated_5 : _GEN_76; // @[LoadQueueFlag.scala 153:{72,72}]
  wire  _GEN_78 = 4'h6 == deqLookupVec_new_ptr_1_value ? allocated_6 : _GEN_77; // @[LoadQueueFlag.scala 153:{72,72}]
  wire  _GEN_79 = 4'h7 == deqLookupVec_new_ptr_1_value ? allocated_7 : _GEN_78; // @[LoadQueueFlag.scala 153:{72,72}]
  wire  _GEN_80 = 4'h8 == deqLookupVec_new_ptr_1_value ? allocated_8 : _GEN_79; // @[LoadQueueFlag.scala 153:{72,72}]
  wire  _GEN_81 = 4'h9 == deqLookupVec_new_ptr_1_value ? allocated_9 : _GEN_80; // @[LoadQueueFlag.scala 153:{72,72}]
  wire  _GEN_82 = 4'ha == deqLookupVec_new_ptr_1_value ? allocated_10 : _GEN_81; // @[LoadQueueFlag.scala 153:{72,72}]
  wire  _GEN_83 = 4'hb == deqLookupVec_new_ptr_1_value ? allocated_11 : _GEN_82; // @[LoadQueueFlag.scala 153:{72,72}]
  wire  _GEN_84 = 4'hc == deqLookupVec_new_ptr_1_value ? allocated_12 : _GEN_83; // @[LoadQueueFlag.scala 153:{72,72}]
  wire  _GEN_85 = 4'hd == deqLookupVec_new_ptr_1_value ? allocated_13 : _GEN_84; // @[LoadQueueFlag.scala 153:{72,72}]
  wire  _GEN_86 = 4'he == deqLookupVec_new_ptr_1_value ? allocated_14 : _GEN_85; // @[LoadQueueFlag.scala 153:{72,72}]
  wire  _GEN_87 = 4'hf == deqLookupVec_new_ptr_1_value ? allocated_15 : _GEN_86; // @[LoadQueueFlag.scala 153:{72,72}]
  wire  _GEN_89 = 4'h1 == deqLookupVec_new_ptr_1_value ? datavalid_1 : datavalid_0; // @[LoadQueueFlag.scala 153:{72,72}]
  wire  _GEN_90 = 4'h2 == deqLookupVec_new_ptr_1_value ? datavalid_2 : _GEN_89; // @[LoadQueueFlag.scala 153:{72,72}]
  wire  _GEN_91 = 4'h3 == deqLookupVec_new_ptr_1_value ? datavalid_3 : _GEN_90; // @[LoadQueueFlag.scala 153:{72,72}]
  wire  _GEN_92 = 4'h4 == deqLookupVec_new_ptr_1_value ? datavalid_4 : _GEN_91; // @[LoadQueueFlag.scala 153:{72,72}]
  wire  _GEN_93 = 4'h5 == deqLookupVec_new_ptr_1_value ? datavalid_5 : _GEN_92; // @[LoadQueueFlag.scala 153:{72,72}]
  wire  _GEN_94 = 4'h6 == deqLookupVec_new_ptr_1_value ? datavalid_6 : _GEN_93; // @[LoadQueueFlag.scala 153:{72,72}]
  wire  _GEN_95 = 4'h7 == deqLookupVec_new_ptr_1_value ? datavalid_7 : _GEN_94; // @[LoadQueueFlag.scala 153:{72,72}]
  wire  _GEN_96 = 4'h8 == deqLookupVec_new_ptr_1_value ? datavalid_8 : _GEN_95; // @[LoadQueueFlag.scala 153:{72,72}]
  wire  _GEN_97 = 4'h9 == deqLookupVec_new_ptr_1_value ? datavalid_9 : _GEN_96; // @[LoadQueueFlag.scala 153:{72,72}]
  wire  _GEN_98 = 4'ha == deqLookupVec_new_ptr_1_value ? datavalid_10 : _GEN_97; // @[LoadQueueFlag.scala 153:{72,72}]
  wire  _GEN_99 = 4'hb == deqLookupVec_new_ptr_1_value ? datavalid_11 : _GEN_98; // @[LoadQueueFlag.scala 153:{72,72}]
  wire  _GEN_100 = 4'hc == deqLookupVec_new_ptr_1_value ? datavalid_12 : _GEN_99; // @[LoadQueueFlag.scala 153:{72,72}]
  wire  _GEN_101 = 4'hd == deqLookupVec_new_ptr_1_value ? datavalid_13 : _GEN_100; // @[LoadQueueFlag.scala 153:{72,72}]
  wire  _GEN_102 = 4'he == deqLookupVec_new_ptr_1_value ? datavalid_14 : _GEN_101; // @[LoadQueueFlag.scala 153:{72,72}]
  wire  _GEN_103 = 4'hf == deqLookupVec_new_ptr_1_value ? datavalid_15 : _GEN_102; // @[LoadQueueFlag.scala 153:{72,72}]
  wire  _GEN_105 = 4'h1 == deqLookupVec_new_ptr_1_value ? addrvalid_1 : addrvalid_0; // @[LoadQueueFlag.scala 153:{96,96}]
  wire  _GEN_106 = 4'h2 == deqLookupVec_new_ptr_1_value ? addrvalid_2 : _GEN_105; // @[LoadQueueFlag.scala 153:{96,96}]
  wire  _GEN_107 = 4'h3 == deqLookupVec_new_ptr_1_value ? addrvalid_3 : _GEN_106; // @[LoadQueueFlag.scala 153:{96,96}]
  wire  _GEN_108 = 4'h4 == deqLookupVec_new_ptr_1_value ? addrvalid_4 : _GEN_107; // @[LoadQueueFlag.scala 153:{96,96}]
  wire  _GEN_109 = 4'h5 == deqLookupVec_new_ptr_1_value ? addrvalid_5 : _GEN_108; // @[LoadQueueFlag.scala 153:{96,96}]
  wire  _GEN_110 = 4'h6 == deqLookupVec_new_ptr_1_value ? addrvalid_6 : _GEN_109; // @[LoadQueueFlag.scala 153:{96,96}]
  wire  _GEN_111 = 4'h7 == deqLookupVec_new_ptr_1_value ? addrvalid_7 : _GEN_110; // @[LoadQueueFlag.scala 153:{96,96}]
  wire  _GEN_112 = 4'h8 == deqLookupVec_new_ptr_1_value ? addrvalid_8 : _GEN_111; // @[LoadQueueFlag.scala 153:{96,96}]
  wire  _GEN_113 = 4'h9 == deqLookupVec_new_ptr_1_value ? addrvalid_9 : _GEN_112; // @[LoadQueueFlag.scala 153:{96,96}]
  wire  _GEN_114 = 4'ha == deqLookupVec_new_ptr_1_value ? addrvalid_10 : _GEN_113; // @[LoadQueueFlag.scala 153:{96,96}]
  wire  _GEN_115 = 4'hb == deqLookupVec_new_ptr_1_value ? addrvalid_11 : _GEN_114; // @[LoadQueueFlag.scala 153:{96,96}]
  wire  _GEN_116 = 4'hc == deqLookupVec_new_ptr_1_value ? addrvalid_12 : _GEN_115; // @[LoadQueueFlag.scala 153:{96,96}]
  wire  _GEN_117 = 4'hd == deqLookupVec_new_ptr_1_value ? addrvalid_13 : _GEN_116; // @[LoadQueueFlag.scala 153:{96,96}]
  wire  _GEN_118 = 4'he == deqLookupVec_new_ptr_1_value ? addrvalid_14 : _GEN_117; // @[LoadQueueFlag.scala 153:{96,96}]
  wire  _GEN_119 = 4'hf == deqLookupVec_new_ptr_1_value ? addrvalid_15 : _GEN_118; // @[LoadQueueFlag.scala 153:{96,96}]
  wire  _GEN_121 = 4'h1 == deqLookupVec_new_ptr_1_value ? writebacked_1 : writebacked_0; // @[LoadQueueFlag.scala 153:{121,121}]
  wire  _GEN_122 = 4'h2 == deqLookupVec_new_ptr_1_value ? writebacked_2 : _GEN_121; // @[LoadQueueFlag.scala 153:{121,121}]
  wire  _GEN_123 = 4'h3 == deqLookupVec_new_ptr_1_value ? writebacked_3 : _GEN_122; // @[LoadQueueFlag.scala 153:{121,121}]
  wire  _GEN_124 = 4'h4 == deqLookupVec_new_ptr_1_value ? writebacked_4 : _GEN_123; // @[LoadQueueFlag.scala 153:{121,121}]
  wire  _GEN_125 = 4'h5 == deqLookupVec_new_ptr_1_value ? writebacked_5 : _GEN_124; // @[LoadQueueFlag.scala 153:{121,121}]
  wire  _GEN_126 = 4'h6 == deqLookupVec_new_ptr_1_value ? writebacked_6 : _GEN_125; // @[LoadQueueFlag.scala 153:{121,121}]
  wire  _GEN_127 = 4'h7 == deqLookupVec_new_ptr_1_value ? writebacked_7 : _GEN_126; // @[LoadQueueFlag.scala 153:{121,121}]
  wire  _GEN_128 = 4'h8 == deqLookupVec_new_ptr_1_value ? writebacked_8 : _GEN_127; // @[LoadQueueFlag.scala 153:{121,121}]
  wire  _GEN_129 = 4'h9 == deqLookupVec_new_ptr_1_value ? writebacked_9 : _GEN_128; // @[LoadQueueFlag.scala 153:{121,121}]
  wire  _GEN_130 = 4'ha == deqLookupVec_new_ptr_1_value ? writebacked_10 : _GEN_129; // @[LoadQueueFlag.scala 153:{121,121}]
  wire  _GEN_131 = 4'hb == deqLookupVec_new_ptr_1_value ? writebacked_11 : _GEN_130; // @[LoadQueueFlag.scala 153:{121,121}]
  wire  _GEN_132 = 4'hc == deqLookupVec_new_ptr_1_value ? writebacked_12 : _GEN_131; // @[LoadQueueFlag.scala 153:{121,121}]
  wire  _GEN_133 = 4'hd == deqLookupVec_new_ptr_1_value ? writebacked_13 : _GEN_132; // @[LoadQueueFlag.scala 153:{121,121}]
  wire  _GEN_134 = 4'he == deqLookupVec_new_ptr_1_value ? writebacked_14 : _GEN_133; // @[LoadQueueFlag.scala 153:{121,121}]
  wire  _GEN_135 = 4'hf == deqLookupVec_new_ptr_1_value ? writebacked_15 : _GEN_134; // @[LoadQueueFlag.scala 153:{121,121}]
  wire [4:0] _deqLookup_T_10 = {deqLookupVec_new_ptr_1_flag,deqLookupVec_new_ptr_1_value}; // @[CircularQueuePtr.scala 63:50]
  wire  _deqLookup_T_12 = _deqLookup_T_10 != _flipped_new_ptr_new_ptr_T; // @[CircularQueuePtr.scala 63:52]
  wire  deqLookup_1 = _GEN_87 & _GEN_103 & _GEN_119 & _GEN_135 & _deqLookup_T_12; // @[LoadQueueFlag.scala 153:147]
  wire  _GEN_137 = 4'h1 == deqLookupVec_new_ptr_value ? needCancel_1 : needCancel_0; // @[LoadQueueFlag.scala 154:{39,39}]
  wire  _GEN_138 = 4'h2 == deqLookupVec_new_ptr_value ? needCancel_2 : _GEN_137; // @[LoadQueueFlag.scala 154:{39,39}]
  wire  _GEN_139 = 4'h3 == deqLookupVec_new_ptr_value ? needCancel_3 : _GEN_138; // @[LoadQueueFlag.scala 154:{39,39}]
  wire  _GEN_140 = 4'h4 == deqLookupVec_new_ptr_value ? needCancel_4 : _GEN_139; // @[LoadQueueFlag.scala 154:{39,39}]
  wire  _GEN_141 = 4'h5 == deqLookupVec_new_ptr_value ? needCancel_5 : _GEN_140; // @[LoadQueueFlag.scala 154:{39,39}]
  wire  _GEN_142 = 4'h6 == deqLookupVec_new_ptr_value ? needCancel_6 : _GEN_141; // @[LoadQueueFlag.scala 154:{39,39}]
  wire  _GEN_143 = 4'h7 == deqLookupVec_new_ptr_value ? needCancel_7 : _GEN_142; // @[LoadQueueFlag.scala 154:{39,39}]
  wire  _GEN_144 = 4'h8 == deqLookupVec_new_ptr_value ? needCancel_8 : _GEN_143; // @[LoadQueueFlag.scala 154:{39,39}]
  wire  _GEN_145 = 4'h9 == deqLookupVec_new_ptr_value ? needCancel_9 : _GEN_144; // @[LoadQueueFlag.scala 154:{39,39}]
  wire  _GEN_146 = 4'ha == deqLookupVec_new_ptr_value ? needCancel_10 : _GEN_145; // @[LoadQueueFlag.scala 154:{39,39}]
  wire  _GEN_147 = 4'hb == deqLookupVec_new_ptr_value ? needCancel_11 : _GEN_146; // @[LoadQueueFlag.scala 154:{39,39}]
  wire  _GEN_148 = 4'hc == deqLookupVec_new_ptr_value ? needCancel_12 : _GEN_147; // @[LoadQueueFlag.scala 154:{39,39}]
  wire  _GEN_149 = 4'hd == deqLookupVec_new_ptr_value ? needCancel_13 : _GEN_148; // @[LoadQueueFlag.scala 154:{39,39}]
  wire  _GEN_150 = 4'he == deqLookupVec_new_ptr_value ? needCancel_14 : _GEN_149; // @[LoadQueueFlag.scala 154:{39,39}]
  wire  deqInSameRedirectCycle_0 = 4'hf == deqLookupVec_new_ptr_value ? needCancel_15 : _GEN_150; // @[LoadQueueFlag.scala 154:{39,39}]
  wire  _GEN_153 = 4'h1 == deqLookupVec_new_ptr_1_value ? needCancel_1 : needCancel_0; // @[LoadQueueFlag.scala 154:{39,39}]
  wire  _GEN_154 = 4'h2 == deqLookupVec_new_ptr_1_value ? needCancel_2 : _GEN_153; // @[LoadQueueFlag.scala 154:{39,39}]
  wire  _GEN_155 = 4'h3 == deqLookupVec_new_ptr_1_value ? needCancel_3 : _GEN_154; // @[LoadQueueFlag.scala 154:{39,39}]
  wire  _GEN_156 = 4'h4 == deqLookupVec_new_ptr_1_value ? needCancel_4 : _GEN_155; // @[LoadQueueFlag.scala 154:{39,39}]
  wire  _GEN_157 = 4'h5 == deqLookupVec_new_ptr_1_value ? needCancel_5 : _GEN_156; // @[LoadQueueFlag.scala 154:{39,39}]
  wire  _GEN_158 = 4'h6 == deqLookupVec_new_ptr_1_value ? needCancel_6 : _GEN_157; // @[LoadQueueFlag.scala 154:{39,39}]
  wire  _GEN_159 = 4'h7 == deqLookupVec_new_ptr_1_value ? needCancel_7 : _GEN_158; // @[LoadQueueFlag.scala 154:{39,39}]
  wire  _GEN_160 = 4'h8 == deqLookupVec_new_ptr_1_value ? needCancel_8 : _GEN_159; // @[LoadQueueFlag.scala 154:{39,39}]
  wire  _GEN_161 = 4'h9 == deqLookupVec_new_ptr_1_value ? needCancel_9 : _GEN_160; // @[LoadQueueFlag.scala 154:{39,39}]
  wire  _GEN_162 = 4'ha == deqLookupVec_new_ptr_1_value ? needCancel_10 : _GEN_161; // @[LoadQueueFlag.scala 154:{39,39}]
  wire  _GEN_163 = 4'hb == deqLookupVec_new_ptr_1_value ? needCancel_11 : _GEN_162; // @[LoadQueueFlag.scala 154:{39,39}]
  wire  _GEN_164 = 4'hc == deqLookupVec_new_ptr_1_value ? needCancel_12 : _GEN_163; // @[LoadQueueFlag.scala 154:{39,39}]
  wire  _GEN_165 = 4'hd == deqLookupVec_new_ptr_1_value ? needCancel_13 : _GEN_164; // @[LoadQueueFlag.scala 154:{39,39}]
  wire  _GEN_166 = 4'he == deqLookupVec_new_ptr_1_value ? needCancel_14 : _GEN_165; // @[LoadQueueFlag.scala 154:{39,39}]
  wire  deqInSameRedirectCycle_1 = 4'hf == deqLookupVec_new_ptr_1_value ? needCancel_15 : _GEN_166; // @[LoadQueueFlag.scala 154:{39,39}]
  wire [1:0] _deqCountMask_T = {deqLookup_1,deqLookup_0}; // @[LoadQueueFlag.scala 157:29]
  wire [1:0] _deqCountMask_T_1 = {deqInSameRedirectCycle_1,deqInSameRedirectCycle_0}; // @[LoadQueueFlag.scala 157:62]
  wire [1:0] _deqCountMask_T_2 = ~_deqCountMask_T_1; // @[LoadQueueFlag.scala 157:38]
  wire [1:0] deqCountMask = _deqCountMask_T & _deqCountMask_T_2; // @[LoadQueueFlag.scala 157:36]
  wire [1:0] _commitCount_T = ~deqCountMask; // @[LoadQueueFlag.scala 158:48]
  wire [1:0] _commitCount_T_3 = _commitCount_T[1] ? 2'h2 : 2'h0; // @[Mux.scala 47:70]
  wire [1:0] _commitCount_T_4 = _commitCount_T[0] ? 2'h1 : _commitCount_T_3; // @[Mux.scala 47:70]
  wire [1:0] _commitCount_T_6 = _commitCount_T_4 - 2'h1; // @[LoadQueueFlag.scala 158:63]
  wire [1:0] commitCount = _commitCount_T_6[0] + _commitCount_T_6[1]; // @[Bitwise.scala 48:55]
  reg [1:0] lastCommitCount; // @[LoadQueueFlag.scala 159:32]
  wire  deqPtrUpdateEna = lastCommitCount != 2'h0; // @[LoadQueueFlag.scala 164:41]
  wire [4:0] _GEN_31437 = {{3'd0}, lastCommitCount}; // @[CircularQueuePtr.scala 39:46]
  wire [4:0] _deqPtrExtNext_new_ptr_T_2 = _deqLookupVec_new_ptr_T + _GEN_31437; // @[CircularQueuePtr.scala 39:46]
  wire [3:0] deqPtrExtNext_new_ptr_value = _deqPtrExtNext_new_ptr_T_2[3:0]; // @[CircularQueuePtr.scala 39:59]
  wire  deqPtrExtNext_new_ptr_flag = _deqPtrExtNext_new_ptr_T_2[4]; // @[CircularQueuePtr.scala 39:59]
  reg [1:0] io_lqDeq_REG; // @[LoadQueueFlag.scala 168:22]
  reg [4:0] io_lqCancelCnt_REG; // @[LoadQueueFlag.scala 169:28]
  wire  _GEN_270 = 4'h0 == io_enq_req_0_bits_lqIdx_value | allocated_0; // @[LoadQueueFlag.scala 205:{24,24} 61:26]
  wire  _GEN_271 = 4'h1 == io_enq_req_0_bits_lqIdx_value | allocated_1; // @[LoadQueueFlag.scala 205:{24,24} 61:26]
  wire  _GEN_272 = 4'h2 == io_enq_req_0_bits_lqIdx_value | allocated_2; // @[LoadQueueFlag.scala 205:{24,24} 61:26]
  wire  _GEN_273 = 4'h3 == io_enq_req_0_bits_lqIdx_value | allocated_3; // @[LoadQueueFlag.scala 205:{24,24} 61:26]
  wire  _GEN_274 = 4'h4 == io_enq_req_0_bits_lqIdx_value | allocated_4; // @[LoadQueueFlag.scala 205:{24,24} 61:26]
  wire  _GEN_275 = 4'h5 == io_enq_req_0_bits_lqIdx_value | allocated_5; // @[LoadQueueFlag.scala 205:{24,24} 61:26]
  wire  _GEN_276 = 4'h6 == io_enq_req_0_bits_lqIdx_value | allocated_6; // @[LoadQueueFlag.scala 205:{24,24} 61:26]
  wire  _GEN_277 = 4'h7 == io_enq_req_0_bits_lqIdx_value | allocated_7; // @[LoadQueueFlag.scala 205:{24,24} 61:26]
  wire  _GEN_278 = 4'h8 == io_enq_req_0_bits_lqIdx_value | allocated_8; // @[LoadQueueFlag.scala 205:{24,24} 61:26]
  wire  _GEN_279 = 4'h9 == io_enq_req_0_bits_lqIdx_value | allocated_9; // @[LoadQueueFlag.scala 205:{24,24} 61:26]
  wire  _GEN_280 = 4'ha == io_enq_req_0_bits_lqIdx_value | allocated_10; // @[LoadQueueFlag.scala 205:{24,24} 61:26]
  wire  _GEN_281 = 4'hb == io_enq_req_0_bits_lqIdx_value | allocated_11; // @[LoadQueueFlag.scala 205:{24,24} 61:26]
  wire  _GEN_282 = 4'hc == io_enq_req_0_bits_lqIdx_value | allocated_12; // @[LoadQueueFlag.scala 205:{24,24} 61:26]
  wire  _GEN_283 = 4'hd == io_enq_req_0_bits_lqIdx_value | allocated_13; // @[LoadQueueFlag.scala 205:{24,24} 61:26]
  wire  _GEN_284 = 4'he == io_enq_req_0_bits_lqIdx_value | allocated_14; // @[LoadQueueFlag.scala 205:{24,24} 61:26]
  wire  _GEN_285 = 4'hf == io_enq_req_0_bits_lqIdx_value | allocated_15; // @[LoadQueueFlag.scala 205:{24,24} 61:26]
  wire  _GEN_398 = 4'h0 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_0_cf_exceptionVec_4; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_399 = 4'h1 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_1_cf_exceptionVec_4; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_400 = 4'h2 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_2_cf_exceptionVec_4; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_401 = 4'h3 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_3_cf_exceptionVec_4; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_402 = 4'h4 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_4_cf_exceptionVec_4; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_403 = 4'h5 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_5_cf_exceptionVec_4; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_404 = 4'h6 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_6_cf_exceptionVec_4; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_405 = 4'h7 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_7_cf_exceptionVec_4; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_406 = 4'h8 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_8_cf_exceptionVec_4; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_407 = 4'h9 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_9_cf_exceptionVec_4; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_408 = 4'ha == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_10_cf_exceptionVec_4; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_409 = 4'hb == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_11_cf_exceptionVec_4; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_410 = 4'hc == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_12_cf_exceptionVec_4; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_411 = 4'hd == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_13_cf_exceptionVec_4; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_412 = 4'he == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_14_cf_exceptionVec_4; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_413 = 4'hf == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_15_cf_exceptionVec_4; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_414 = 4'h0 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_0_cf_exceptionVec_5; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_415 = 4'h1 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_1_cf_exceptionVec_5; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_416 = 4'h2 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_2_cf_exceptionVec_5; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_417 = 4'h3 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_3_cf_exceptionVec_5; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_418 = 4'h4 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_4_cf_exceptionVec_5; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_419 = 4'h5 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_5_cf_exceptionVec_5; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_420 = 4'h6 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_6_cf_exceptionVec_5; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_421 = 4'h7 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_7_cf_exceptionVec_5; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_422 = 4'h8 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_8_cf_exceptionVec_5; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_423 = 4'h9 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_9_cf_exceptionVec_5; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_424 = 4'ha == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_10_cf_exceptionVec_5; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_425 = 4'hb == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_11_cf_exceptionVec_5; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_426 = 4'hc == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_12_cf_exceptionVec_5; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_427 = 4'hd == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_13_cf_exceptionVec_5; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_428 = 4'he == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_14_cf_exceptionVec_5; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_429 = 4'hf == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_15_cf_exceptionVec_5; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_542 = 4'h0 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_0_cf_exceptionVec_13; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_543 = 4'h1 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_1_cf_exceptionVec_13; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_544 = 4'h2 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_2_cf_exceptionVec_13; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_545 = 4'h3 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_3_cf_exceptionVec_13; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_546 = 4'h4 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_4_cf_exceptionVec_13; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_547 = 4'h5 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_5_cf_exceptionVec_13; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_548 = 4'h6 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_6_cf_exceptionVec_13; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_549 = 4'h7 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_7_cf_exceptionVec_13; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_550 = 4'h8 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_8_cf_exceptionVec_13; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_551 = 4'h9 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_9_cf_exceptionVec_13; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_552 = 4'ha == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_10_cf_exceptionVec_13; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_553 = 4'hb == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_11_cf_exceptionVec_13; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_554 = 4'hc == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_12_cf_exceptionVec_13; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_555 = 4'hd == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_13_cf_exceptionVec_13; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_556 = 4'he == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_14_cf_exceptionVec_13; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_557 = 4'hf == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_15_cf_exceptionVec_13; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_670 = 4'h0 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_cf_trigger_backendEn_1 :
    uop_0_cf_trigger_backendEn_1; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_671 = 4'h1 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_cf_trigger_backendEn_1 :
    uop_1_cf_trigger_backendEn_1; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_672 = 4'h2 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_cf_trigger_backendEn_1 :
    uop_2_cf_trigger_backendEn_1; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_673 = 4'h3 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_cf_trigger_backendEn_1 :
    uop_3_cf_trigger_backendEn_1; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_674 = 4'h4 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_cf_trigger_backendEn_1 :
    uop_4_cf_trigger_backendEn_1; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_675 = 4'h5 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_cf_trigger_backendEn_1 :
    uop_5_cf_trigger_backendEn_1; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_676 = 4'h6 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_cf_trigger_backendEn_1 :
    uop_6_cf_trigger_backendEn_1; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_677 = 4'h7 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_cf_trigger_backendEn_1 :
    uop_7_cf_trigger_backendEn_1; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_678 = 4'h8 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_cf_trigger_backendEn_1 :
    uop_8_cf_trigger_backendEn_1; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_679 = 4'h9 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_cf_trigger_backendEn_1 :
    uop_9_cf_trigger_backendEn_1; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_680 = 4'ha == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_cf_trigger_backendEn_1 :
    uop_10_cf_trigger_backendEn_1; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_681 = 4'hb == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_cf_trigger_backendEn_1 :
    uop_11_cf_trigger_backendEn_1; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_682 = 4'hc == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_cf_trigger_backendEn_1 :
    uop_12_cf_trigger_backendEn_1; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_683 = 4'hd == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_cf_trigger_backendEn_1 :
    uop_13_cf_trigger_backendEn_1; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_684 = 4'he == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_cf_trigger_backendEn_1 :
    uop_14_cf_trigger_backendEn_1; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_685 = 4'hf == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_cf_trigger_backendEn_1 :
    uop_15_cf_trigger_backendEn_1; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_686 = 4'h0 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_0_cf_trigger_backendHit_0; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_687 = 4'h1 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_1_cf_trigger_backendHit_0; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_688 = 4'h2 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_2_cf_trigger_backendHit_0; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_689 = 4'h3 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_3_cf_trigger_backendHit_0; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_690 = 4'h4 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_4_cf_trigger_backendHit_0; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_691 = 4'h5 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_5_cf_trigger_backendHit_0; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_692 = 4'h6 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_6_cf_trigger_backendHit_0; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_693 = 4'h7 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_7_cf_trigger_backendHit_0; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_694 = 4'h8 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_8_cf_trigger_backendHit_0; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_695 = 4'h9 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_9_cf_trigger_backendHit_0; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_696 = 4'ha == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_10_cf_trigger_backendHit_0; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_697 = 4'hb == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_11_cf_trigger_backendHit_0; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_698 = 4'hc == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_12_cf_trigger_backendHit_0; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_699 = 4'hd == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_13_cf_trigger_backendHit_0; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_700 = 4'he == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_14_cf_trigger_backendHit_0; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_701 = 4'hf == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_15_cf_trigger_backendHit_0; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_702 = 4'h0 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_0_cf_trigger_backendHit_1; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_703 = 4'h1 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_1_cf_trigger_backendHit_1; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_704 = 4'h2 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_2_cf_trigger_backendHit_1; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_705 = 4'h3 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_3_cf_trigger_backendHit_1; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_706 = 4'h4 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_4_cf_trigger_backendHit_1; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_707 = 4'h5 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_5_cf_trigger_backendHit_1; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_708 = 4'h6 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_6_cf_trigger_backendHit_1; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_709 = 4'h7 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_7_cf_trigger_backendHit_1; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_710 = 4'h8 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_8_cf_trigger_backendHit_1; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_711 = 4'h9 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_9_cf_trigger_backendHit_1; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_712 = 4'ha == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_10_cf_trigger_backendHit_1; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_713 = 4'hb == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_11_cf_trigger_backendHit_1; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_714 = 4'hc == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_12_cf_trigger_backendHit_1; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_715 = 4'hd == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_13_cf_trigger_backendHit_1; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_716 = 4'he == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_14_cf_trigger_backendHit_1; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_717 = 4'hf == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_15_cf_trigger_backendHit_1; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_750 = 4'h0 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_0_cf_trigger_backendHit_4; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_751 = 4'h1 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_1_cf_trigger_backendHit_4; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_752 = 4'h2 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_2_cf_trigger_backendHit_4; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_753 = 4'h3 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_3_cf_trigger_backendHit_4; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_754 = 4'h4 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_4_cf_trigger_backendHit_4; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_755 = 4'h5 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_5_cf_trigger_backendHit_4; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_756 = 4'h6 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_6_cf_trigger_backendHit_4; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_757 = 4'h7 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_7_cf_trigger_backendHit_4; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_758 = 4'h8 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_8_cf_trigger_backendHit_4; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_759 = 4'h9 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_9_cf_trigger_backendHit_4; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_760 = 4'ha == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_10_cf_trigger_backendHit_4; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_761 = 4'hb == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_11_cf_trigger_backendHit_4; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_762 = 4'hc == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_12_cf_trigger_backendHit_4; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_763 = 4'hd == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_13_cf_trigger_backendHit_4; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_764 = 4'he == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_14_cf_trigger_backendHit_4; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_765 = 4'hf == io_enq_req_0_bits_lqIdx_value ? 1'h0 : uop_15_cf_trigger_backendHit_4; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire [6:0] _GEN_1182 = 4'h0 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_ctrl_fuOpType : uop_0_ctrl_fuOpType; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire [6:0] _GEN_1183 = 4'h1 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_ctrl_fuOpType : uop_1_ctrl_fuOpType; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire [6:0] _GEN_1184 = 4'h2 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_ctrl_fuOpType : uop_2_ctrl_fuOpType; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire [6:0] _GEN_1185 = 4'h3 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_ctrl_fuOpType : uop_3_ctrl_fuOpType; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire [6:0] _GEN_1186 = 4'h4 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_ctrl_fuOpType : uop_4_ctrl_fuOpType; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire [6:0] _GEN_1187 = 4'h5 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_ctrl_fuOpType : uop_5_ctrl_fuOpType; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire [6:0] _GEN_1188 = 4'h6 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_ctrl_fuOpType : uop_6_ctrl_fuOpType; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire [6:0] _GEN_1189 = 4'h7 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_ctrl_fuOpType : uop_7_ctrl_fuOpType; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire [6:0] _GEN_1190 = 4'h8 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_ctrl_fuOpType : uop_8_ctrl_fuOpType; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire [6:0] _GEN_1191 = 4'h9 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_ctrl_fuOpType : uop_9_ctrl_fuOpType; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire [6:0] _GEN_1192 = 4'ha == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_ctrl_fuOpType : uop_10_ctrl_fuOpType; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire [6:0] _GEN_1193 = 4'hb == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_ctrl_fuOpType : uop_11_ctrl_fuOpType; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire [6:0] _GEN_1194 = 4'hc == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_ctrl_fuOpType : uop_12_ctrl_fuOpType; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire [6:0] _GEN_1195 = 4'hd == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_ctrl_fuOpType : uop_13_ctrl_fuOpType; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire [6:0] _GEN_1196 = 4'he == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_ctrl_fuOpType : uop_14_ctrl_fuOpType; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire [6:0] _GEN_1197 = 4'hf == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_ctrl_fuOpType : uop_15_ctrl_fuOpType; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_1198 = 4'h0 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_ctrl_rfWen : uop_0_ctrl_rfWen; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_1199 = 4'h1 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_ctrl_rfWen : uop_1_ctrl_rfWen; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_1200 = 4'h2 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_ctrl_rfWen : uop_2_ctrl_rfWen; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_1201 = 4'h3 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_ctrl_rfWen : uop_3_ctrl_rfWen; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_1202 = 4'h4 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_ctrl_rfWen : uop_4_ctrl_rfWen; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_1203 = 4'h5 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_ctrl_rfWen : uop_5_ctrl_rfWen; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_1204 = 4'h6 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_ctrl_rfWen : uop_6_ctrl_rfWen; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_1205 = 4'h7 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_ctrl_rfWen : uop_7_ctrl_rfWen; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_1206 = 4'h8 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_ctrl_rfWen : uop_8_ctrl_rfWen; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_1207 = 4'h9 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_ctrl_rfWen : uop_9_ctrl_rfWen; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_1208 = 4'ha == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_ctrl_rfWen : uop_10_ctrl_rfWen; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_1209 = 4'hb == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_ctrl_rfWen : uop_11_ctrl_rfWen; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_1210 = 4'hc == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_ctrl_rfWen : uop_12_ctrl_rfWen; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_1211 = 4'hd == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_ctrl_rfWen : uop_13_ctrl_rfWen; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_1212 = 4'he == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_ctrl_rfWen : uop_14_ctrl_rfWen; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_1213 = 4'hf == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_ctrl_rfWen : uop_15_ctrl_rfWen; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_1214 = 4'h0 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_ctrl_fpWen : uop_0_ctrl_fpWen; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_1215 = 4'h1 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_ctrl_fpWen : uop_1_ctrl_fpWen; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_1216 = 4'h2 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_ctrl_fpWen : uop_2_ctrl_fpWen; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_1217 = 4'h3 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_ctrl_fpWen : uop_3_ctrl_fpWen; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_1218 = 4'h4 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_ctrl_fpWen : uop_4_ctrl_fpWen; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_1219 = 4'h5 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_ctrl_fpWen : uop_5_ctrl_fpWen; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_1220 = 4'h6 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_ctrl_fpWen : uop_6_ctrl_fpWen; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_1221 = 4'h7 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_ctrl_fpWen : uop_7_ctrl_fpWen; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_1222 = 4'h8 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_ctrl_fpWen : uop_8_ctrl_fpWen; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_1223 = 4'h9 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_ctrl_fpWen : uop_9_ctrl_fpWen; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_1224 = 4'ha == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_ctrl_fpWen : uop_10_ctrl_fpWen; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_1225 = 4'hb == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_ctrl_fpWen : uop_11_ctrl_fpWen; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_1226 = 4'hc == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_ctrl_fpWen : uop_12_ctrl_fpWen; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_1227 = 4'hd == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_ctrl_fpWen : uop_13_ctrl_fpWen; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_1228 = 4'he == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_ctrl_fpWen : uop_14_ctrl_fpWen; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_1229 = 4'hf == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_ctrl_fpWen : uop_15_ctrl_fpWen; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_1278 = 4'h0 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_ctrl_flushPipe : uop_0_ctrl_flushPipe; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_1279 = 4'h1 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_ctrl_flushPipe : uop_1_ctrl_flushPipe; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_1280 = 4'h2 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_ctrl_flushPipe : uop_2_ctrl_flushPipe; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_1281 = 4'h3 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_ctrl_flushPipe : uop_3_ctrl_flushPipe; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_1282 = 4'h4 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_ctrl_flushPipe : uop_4_ctrl_flushPipe; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_1283 = 4'h5 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_ctrl_flushPipe : uop_5_ctrl_flushPipe; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_1284 = 4'h6 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_ctrl_flushPipe : uop_6_ctrl_flushPipe; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_1285 = 4'h7 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_ctrl_flushPipe : uop_7_ctrl_flushPipe; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_1286 = 4'h8 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_ctrl_flushPipe : uop_8_ctrl_flushPipe; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_1287 = 4'h9 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_ctrl_flushPipe : uop_9_ctrl_flushPipe; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_1288 = 4'ha == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_ctrl_flushPipe : uop_10_ctrl_flushPipe; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_1289 = 4'hb == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_ctrl_flushPipe : uop_11_ctrl_flushPipe; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_1290 = 4'hc == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_ctrl_flushPipe : uop_12_ctrl_flushPipe; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_1291 = 4'hd == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_ctrl_flushPipe : uop_13_ctrl_flushPipe; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_1292 = 4'he == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_ctrl_flushPipe : uop_14_ctrl_flushPipe; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_1293 = 4'hf == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_ctrl_flushPipe : uop_15_ctrl_flushPipe; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_1598 = 4'h0 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_ctrl_replayInst : uop_0_ctrl_replayInst; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_1599 = 4'h1 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_ctrl_replayInst : uop_1_ctrl_replayInst; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_1600 = 4'h2 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_ctrl_replayInst : uop_2_ctrl_replayInst; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_1601 = 4'h3 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_ctrl_replayInst : uop_3_ctrl_replayInst; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_1602 = 4'h4 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_ctrl_replayInst : uop_4_ctrl_replayInst; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_1603 = 4'h5 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_ctrl_replayInst : uop_5_ctrl_replayInst; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_1604 = 4'h6 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_ctrl_replayInst : uop_6_ctrl_replayInst; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_1605 = 4'h7 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_ctrl_replayInst : uop_7_ctrl_replayInst; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_1606 = 4'h8 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_ctrl_replayInst : uop_8_ctrl_replayInst; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_1607 = 4'h9 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_ctrl_replayInst : uop_9_ctrl_replayInst; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_1608 = 4'ha == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_ctrl_replayInst : uop_10_ctrl_replayInst; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_1609 = 4'hb == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_ctrl_replayInst : uop_11_ctrl_replayInst; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_1610 = 4'hc == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_ctrl_replayInst : uop_12_ctrl_replayInst; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_1611 = 4'hd == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_ctrl_replayInst : uop_13_ctrl_replayInst; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_1612 = 4'he == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_ctrl_replayInst : uop_14_ctrl_replayInst; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_1613 = 4'hf == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_ctrl_replayInst : uop_15_ctrl_replayInst; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire [5:0] _GEN_1710 = 4'h0 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_pdest : uop_0_pdest; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire [5:0] _GEN_1711 = 4'h1 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_pdest : uop_1_pdest; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire [5:0] _GEN_1712 = 4'h2 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_pdest : uop_2_pdest; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire [5:0] _GEN_1713 = 4'h3 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_pdest : uop_3_pdest; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire [5:0] _GEN_1714 = 4'h4 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_pdest : uop_4_pdest; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire [5:0] _GEN_1715 = 4'h5 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_pdest : uop_5_pdest; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire [5:0] _GEN_1716 = 4'h6 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_pdest : uop_6_pdest; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire [5:0] _GEN_1717 = 4'h7 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_pdest : uop_7_pdest; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire [5:0] _GEN_1718 = 4'h8 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_pdest : uop_8_pdest; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire [5:0] _GEN_1719 = 4'h9 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_pdest : uop_9_pdest; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire [5:0] _GEN_1720 = 4'ha == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_pdest : uop_10_pdest; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire [5:0] _GEN_1721 = 4'hb == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_pdest : uop_11_pdest; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire [5:0] _GEN_1722 = 4'hc == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_pdest : uop_12_pdest; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire [5:0] _GEN_1723 = 4'hd == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_pdest : uop_13_pdest; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire [5:0] _GEN_1724 = 4'he == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_pdest : uop_14_pdest; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire [5:0] _GEN_1725 = 4'hf == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_pdest : uop_15_pdest; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_1742 = 4'h0 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_robIdx_flag : uop_0_robIdx_flag; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_1743 = 4'h1 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_robIdx_flag : uop_1_robIdx_flag; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_1744 = 4'h2 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_robIdx_flag : uop_2_robIdx_flag; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_1745 = 4'h3 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_robIdx_flag : uop_3_robIdx_flag; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_1746 = 4'h4 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_robIdx_flag : uop_4_robIdx_flag; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_1747 = 4'h5 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_robIdx_flag : uop_5_robIdx_flag; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_1748 = 4'h6 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_robIdx_flag : uop_6_robIdx_flag; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_1749 = 4'h7 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_robIdx_flag : uop_7_robIdx_flag; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_1750 = 4'h8 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_robIdx_flag : uop_8_robIdx_flag; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_1751 = 4'h9 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_robIdx_flag : uop_9_robIdx_flag; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_1752 = 4'ha == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_robIdx_flag : uop_10_robIdx_flag; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_1753 = 4'hb == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_robIdx_flag : uop_11_robIdx_flag; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_1754 = 4'hc == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_robIdx_flag : uop_12_robIdx_flag; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_1755 = 4'hd == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_robIdx_flag : uop_13_robIdx_flag; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_1756 = 4'he == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_robIdx_flag : uop_14_robIdx_flag; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_1757 = 4'hf == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_robIdx_flag : uop_15_robIdx_flag; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire [4:0] _GEN_1758 = 4'h0 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_robIdx_value : uop_0_robIdx_value; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire [4:0] _GEN_1759 = 4'h1 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_robIdx_value : uop_1_robIdx_value; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire [4:0] _GEN_1760 = 4'h2 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_robIdx_value : uop_2_robIdx_value; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire [4:0] _GEN_1761 = 4'h3 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_robIdx_value : uop_3_robIdx_value; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire [4:0] _GEN_1762 = 4'h4 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_robIdx_value : uop_4_robIdx_value; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire [4:0] _GEN_1763 = 4'h5 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_robIdx_value : uop_5_robIdx_value; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire [4:0] _GEN_1764 = 4'h6 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_robIdx_value : uop_6_robIdx_value; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire [4:0] _GEN_1765 = 4'h7 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_robIdx_value : uop_7_robIdx_value; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire [4:0] _GEN_1766 = 4'h8 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_robIdx_value : uop_8_robIdx_value; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire [4:0] _GEN_1767 = 4'h9 == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_robIdx_value : uop_9_robIdx_value; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire [4:0] _GEN_1768 = 4'ha == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_robIdx_value : uop_10_robIdx_value; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire [4:0] _GEN_1769 = 4'hb == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_robIdx_value : uop_11_robIdx_value; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire [4:0] _GEN_1770 = 4'hc == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_robIdx_value : uop_12_robIdx_value; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire [4:0] _GEN_1771 = 4'hd == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_robIdx_value : uop_13_robIdx_value; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire [4:0] _GEN_1772 = 4'he == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_robIdx_value : uop_14_robIdx_value; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire [4:0] _GEN_1773 = 4'hf == io_enq_req_0_bits_lqIdx_value ? io_enq_req_0_bits_robIdx_value : uop_15_robIdx_value; // @[LoadQueueFlag.scala 206:{18,18} 62:16]
  wire  _GEN_2110 = 4'h0 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : _GEN_398; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_2111 = 4'h1 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : _GEN_399; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_2112 = 4'h2 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : _GEN_400; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_2113 = 4'h3 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : _GEN_401; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_2114 = 4'h4 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : _GEN_402; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_2115 = 4'h5 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : _GEN_403; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_2116 = 4'h6 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : _GEN_404; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_2117 = 4'h7 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : _GEN_405; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_2118 = 4'h8 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : _GEN_406; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_2119 = 4'h9 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : _GEN_407; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_2120 = 4'ha == io_enq_req_0_bits_lqIdx_value ? 1'h0 : _GEN_408; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_2121 = 4'hb == io_enq_req_0_bits_lqIdx_value ? 1'h0 : _GEN_409; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_2122 = 4'hc == io_enq_req_0_bits_lqIdx_value ? 1'h0 : _GEN_410; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_2123 = 4'hd == io_enq_req_0_bits_lqIdx_value ? 1'h0 : _GEN_411; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_2124 = 4'he == io_enq_req_0_bits_lqIdx_value ? 1'h0 : _GEN_412; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_2125 = 4'hf == io_enq_req_0_bits_lqIdx_value ? 1'h0 : _GEN_413; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_2126 = 4'h0 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : _GEN_414; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_2127 = 4'h1 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : _GEN_415; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_2128 = 4'h2 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : _GEN_416; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_2129 = 4'h3 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : _GEN_417; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_2130 = 4'h4 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : _GEN_418; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_2131 = 4'h5 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : _GEN_419; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_2132 = 4'h6 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : _GEN_420; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_2133 = 4'h7 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : _GEN_421; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_2134 = 4'h8 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : _GEN_422; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_2135 = 4'h9 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : _GEN_423; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_2136 = 4'ha == io_enq_req_0_bits_lqIdx_value ? 1'h0 : _GEN_424; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_2137 = 4'hb == io_enq_req_0_bits_lqIdx_value ? 1'h0 : _GEN_425; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_2138 = 4'hc == io_enq_req_0_bits_lqIdx_value ? 1'h0 : _GEN_426; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_2139 = 4'hd == io_enq_req_0_bits_lqIdx_value ? 1'h0 : _GEN_427; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_2140 = 4'he == io_enq_req_0_bits_lqIdx_value ? 1'h0 : _GEN_428; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_2141 = 4'hf == io_enq_req_0_bits_lqIdx_value ? 1'h0 : _GEN_429; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_2254 = 4'h0 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : _GEN_542; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_2255 = 4'h1 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : _GEN_543; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_2256 = 4'h2 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : _GEN_544; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_2257 = 4'h3 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : _GEN_545; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_2258 = 4'h4 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : _GEN_546; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_2259 = 4'h5 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : _GEN_547; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_2260 = 4'h6 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : _GEN_548; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_2261 = 4'h7 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : _GEN_549; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_2262 = 4'h8 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : _GEN_550; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_2263 = 4'h9 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : _GEN_551; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_2264 = 4'ha == io_enq_req_0_bits_lqIdx_value ? 1'h0 : _GEN_552; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_2265 = 4'hb == io_enq_req_0_bits_lqIdx_value ? 1'h0 : _GEN_553; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_2266 = 4'hc == io_enq_req_0_bits_lqIdx_value ? 1'h0 : _GEN_554; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_2267 = 4'hd == io_enq_req_0_bits_lqIdx_value ? 1'h0 : _GEN_555; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_2268 = 4'he == io_enq_req_0_bits_lqIdx_value ? 1'h0 : _GEN_556; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_2269 = 4'hf == io_enq_req_0_bits_lqIdx_value ? 1'h0 : _GEN_557; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_2302 = 4'h0 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : addrvalid_0; // @[LoadQueueFlag.scala 211:{24,24} 90:26]
  wire  _GEN_2303 = 4'h1 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : addrvalid_1; // @[LoadQueueFlag.scala 211:{24,24} 90:26]
  wire  _GEN_2304 = 4'h2 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : addrvalid_2; // @[LoadQueueFlag.scala 211:{24,24} 90:26]
  wire  _GEN_2305 = 4'h3 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : addrvalid_3; // @[LoadQueueFlag.scala 211:{24,24} 90:26]
  wire  _GEN_2306 = 4'h4 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : addrvalid_4; // @[LoadQueueFlag.scala 211:{24,24} 90:26]
  wire  _GEN_2307 = 4'h5 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : addrvalid_5; // @[LoadQueueFlag.scala 211:{24,24} 90:26]
  wire  _GEN_2308 = 4'h6 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : addrvalid_6; // @[LoadQueueFlag.scala 211:{24,24} 90:26]
  wire  _GEN_2309 = 4'h7 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : addrvalid_7; // @[LoadQueueFlag.scala 211:{24,24} 90:26]
  wire  _GEN_2310 = 4'h8 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : addrvalid_8; // @[LoadQueueFlag.scala 211:{24,24} 90:26]
  wire  _GEN_2311 = 4'h9 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : addrvalid_9; // @[LoadQueueFlag.scala 211:{24,24} 90:26]
  wire  _GEN_2312 = 4'ha == io_enq_req_0_bits_lqIdx_value ? 1'h0 : addrvalid_10; // @[LoadQueueFlag.scala 211:{24,24} 90:26]
  wire  _GEN_2313 = 4'hb == io_enq_req_0_bits_lqIdx_value ? 1'h0 : addrvalid_11; // @[LoadQueueFlag.scala 211:{24,24} 90:26]
  wire  _GEN_2314 = 4'hc == io_enq_req_0_bits_lqIdx_value ? 1'h0 : addrvalid_12; // @[LoadQueueFlag.scala 211:{24,24} 90:26]
  wire  _GEN_2315 = 4'hd == io_enq_req_0_bits_lqIdx_value ? 1'h0 : addrvalid_13; // @[LoadQueueFlag.scala 211:{24,24} 90:26]
  wire  _GEN_2316 = 4'he == io_enq_req_0_bits_lqIdx_value ? 1'h0 : addrvalid_14; // @[LoadQueueFlag.scala 211:{24,24} 90:26]
  wire  _GEN_2317 = 4'hf == io_enq_req_0_bits_lqIdx_value ? 1'h0 : addrvalid_15; // @[LoadQueueFlag.scala 211:{24,24} 90:26]
  wire  _GEN_2318 = 4'h0 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : datavalid_0; // @[LoadQueueFlag.scala 212:{24,24} 91:26]
  wire  _GEN_2319 = 4'h1 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : datavalid_1; // @[LoadQueueFlag.scala 212:{24,24} 91:26]
  wire  _GEN_2320 = 4'h2 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : datavalid_2; // @[LoadQueueFlag.scala 212:{24,24} 91:26]
  wire  _GEN_2321 = 4'h3 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : datavalid_3; // @[LoadQueueFlag.scala 212:{24,24} 91:26]
  wire  _GEN_2322 = 4'h4 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : datavalid_4; // @[LoadQueueFlag.scala 212:{24,24} 91:26]
  wire  _GEN_2323 = 4'h5 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : datavalid_5; // @[LoadQueueFlag.scala 212:{24,24} 91:26]
  wire  _GEN_2324 = 4'h6 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : datavalid_6; // @[LoadQueueFlag.scala 212:{24,24} 91:26]
  wire  _GEN_2325 = 4'h7 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : datavalid_7; // @[LoadQueueFlag.scala 212:{24,24} 91:26]
  wire  _GEN_2326 = 4'h8 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : datavalid_8; // @[LoadQueueFlag.scala 212:{24,24} 91:26]
  wire  _GEN_2327 = 4'h9 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : datavalid_9; // @[LoadQueueFlag.scala 212:{24,24} 91:26]
  wire  _GEN_2328 = 4'ha == io_enq_req_0_bits_lqIdx_value ? 1'h0 : datavalid_10; // @[LoadQueueFlag.scala 212:{24,24} 91:26]
  wire  _GEN_2329 = 4'hb == io_enq_req_0_bits_lqIdx_value ? 1'h0 : datavalid_11; // @[LoadQueueFlag.scala 212:{24,24} 91:26]
  wire  _GEN_2330 = 4'hc == io_enq_req_0_bits_lqIdx_value ? 1'h0 : datavalid_12; // @[LoadQueueFlag.scala 212:{24,24} 91:26]
  wire  _GEN_2331 = 4'hd == io_enq_req_0_bits_lqIdx_value ? 1'h0 : datavalid_13; // @[LoadQueueFlag.scala 212:{24,24} 91:26]
  wire  _GEN_2332 = 4'he == io_enq_req_0_bits_lqIdx_value ? 1'h0 : datavalid_14; // @[LoadQueueFlag.scala 212:{24,24} 91:26]
  wire  _GEN_2333 = 4'hf == io_enq_req_0_bits_lqIdx_value ? 1'h0 : datavalid_15; // @[LoadQueueFlag.scala 212:{24,24} 91:26]
  wire  _GEN_2334 = 4'h0 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : pending_0; // @[LoadQueueFlag.scala 213:{22,22} 92:24]
  wire  _GEN_2335 = 4'h1 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : pending_1; // @[LoadQueueFlag.scala 213:{22,22} 92:24]
  wire  _GEN_2336 = 4'h2 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : pending_2; // @[LoadQueueFlag.scala 213:{22,22} 92:24]
  wire  _GEN_2337 = 4'h3 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : pending_3; // @[LoadQueueFlag.scala 213:{22,22} 92:24]
  wire  _GEN_2338 = 4'h4 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : pending_4; // @[LoadQueueFlag.scala 213:{22,22} 92:24]
  wire  _GEN_2339 = 4'h5 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : pending_5; // @[LoadQueueFlag.scala 213:{22,22} 92:24]
  wire  _GEN_2340 = 4'h6 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : pending_6; // @[LoadQueueFlag.scala 213:{22,22} 92:24]
  wire  _GEN_2341 = 4'h7 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : pending_7; // @[LoadQueueFlag.scala 213:{22,22} 92:24]
  wire  _GEN_2342 = 4'h8 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : pending_8; // @[LoadQueueFlag.scala 213:{22,22} 92:24]
  wire  _GEN_2343 = 4'h9 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : pending_9; // @[LoadQueueFlag.scala 213:{22,22} 92:24]
  wire  _GEN_2344 = 4'ha == io_enq_req_0_bits_lqIdx_value ? 1'h0 : pending_10; // @[LoadQueueFlag.scala 213:{22,22} 92:24]
  wire  _GEN_2345 = 4'hb == io_enq_req_0_bits_lqIdx_value ? 1'h0 : pending_11; // @[LoadQueueFlag.scala 213:{22,22} 92:24]
  wire  _GEN_2346 = 4'hc == io_enq_req_0_bits_lqIdx_value ? 1'h0 : pending_12; // @[LoadQueueFlag.scala 213:{22,22} 92:24]
  wire  _GEN_2347 = 4'hd == io_enq_req_0_bits_lqIdx_value ? 1'h0 : pending_13; // @[LoadQueueFlag.scala 213:{22,22} 92:24]
  wire  _GEN_2348 = 4'he == io_enq_req_0_bits_lqIdx_value ? 1'h0 : pending_14; // @[LoadQueueFlag.scala 213:{22,22} 92:24]
  wire  _GEN_2349 = 4'hf == io_enq_req_0_bits_lqIdx_value ? 1'h0 : pending_15; // @[LoadQueueFlag.scala 213:{22,22} 92:24]
  wire  _GEN_2350 = 4'h0 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : writebacked_0; // @[LoadQueueFlag.scala 214:{26,26} 93:28]
  wire  _GEN_2351 = 4'h1 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : writebacked_1; // @[LoadQueueFlag.scala 214:{26,26} 93:28]
  wire  _GEN_2352 = 4'h2 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : writebacked_2; // @[LoadQueueFlag.scala 214:{26,26} 93:28]
  wire  _GEN_2353 = 4'h3 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : writebacked_3; // @[LoadQueueFlag.scala 214:{26,26} 93:28]
  wire  _GEN_2354 = 4'h4 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : writebacked_4; // @[LoadQueueFlag.scala 214:{26,26} 93:28]
  wire  _GEN_2355 = 4'h5 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : writebacked_5; // @[LoadQueueFlag.scala 214:{26,26} 93:28]
  wire  _GEN_2356 = 4'h6 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : writebacked_6; // @[LoadQueueFlag.scala 214:{26,26} 93:28]
  wire  _GEN_2357 = 4'h7 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : writebacked_7; // @[LoadQueueFlag.scala 214:{26,26} 93:28]
  wire  _GEN_2358 = 4'h8 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : writebacked_8; // @[LoadQueueFlag.scala 214:{26,26} 93:28]
  wire  _GEN_2359 = 4'h9 == io_enq_req_0_bits_lqIdx_value ? 1'h0 : writebacked_9; // @[LoadQueueFlag.scala 214:{26,26} 93:28]
  wire  _GEN_2360 = 4'ha == io_enq_req_0_bits_lqIdx_value ? 1'h0 : writebacked_10; // @[LoadQueueFlag.scala 214:{26,26} 93:28]
  wire  _GEN_2361 = 4'hb == io_enq_req_0_bits_lqIdx_value ? 1'h0 : writebacked_11; // @[LoadQueueFlag.scala 214:{26,26} 93:28]
  wire  _GEN_2362 = 4'hc == io_enq_req_0_bits_lqIdx_value ? 1'h0 : writebacked_12; // @[LoadQueueFlag.scala 214:{26,26} 93:28]
  wire  _GEN_2363 = 4'hd == io_enq_req_0_bits_lqIdx_value ? 1'h0 : writebacked_13; // @[LoadQueueFlag.scala 214:{26,26} 93:28]
  wire  _GEN_2364 = 4'he == io_enq_req_0_bits_lqIdx_value ? 1'h0 : writebacked_14; // @[LoadQueueFlag.scala 214:{26,26} 93:28]
  wire  _GEN_2365 = 4'hf == io_enq_req_0_bits_lqIdx_value ? 1'h0 : writebacked_15; // @[LoadQueueFlag.scala 214:{26,26} 93:28]
  wire  _GEN_2414 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_270 : allocated_0; // @[LoadQueueFlag.scala 204:43 61:26]
  wire  _GEN_2415 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_271 : allocated_1; // @[LoadQueueFlag.scala 204:43 61:26]
  wire  _GEN_2416 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_272 : allocated_2; // @[LoadQueueFlag.scala 204:43 61:26]
  wire  _GEN_2417 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_273 : allocated_3; // @[LoadQueueFlag.scala 204:43 61:26]
  wire  _GEN_2418 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_274 : allocated_4; // @[LoadQueueFlag.scala 204:43 61:26]
  wire  _GEN_2419 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_275 : allocated_5; // @[LoadQueueFlag.scala 204:43 61:26]
  wire  _GEN_2420 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_276 : allocated_6; // @[LoadQueueFlag.scala 204:43 61:26]
  wire  _GEN_2421 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_277 : allocated_7; // @[LoadQueueFlag.scala 204:43 61:26]
  wire  _GEN_2422 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_278 : allocated_8; // @[LoadQueueFlag.scala 204:43 61:26]
  wire  _GEN_2423 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_279 : allocated_9; // @[LoadQueueFlag.scala 204:43 61:26]
  wire  _GEN_2424 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_280 : allocated_10; // @[LoadQueueFlag.scala 204:43 61:26]
  wire  _GEN_2425 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_281 : allocated_11; // @[LoadQueueFlag.scala 204:43 61:26]
  wire  _GEN_2426 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_282 : allocated_12; // @[LoadQueueFlag.scala 204:43 61:26]
  wire  _GEN_2427 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_283 : allocated_13; // @[LoadQueueFlag.scala 204:43 61:26]
  wire  _GEN_2428 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_284 : allocated_14; // @[LoadQueueFlag.scala 204:43 61:26]
  wire  _GEN_2429 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_285 : allocated_15; // @[LoadQueueFlag.scala 204:43 61:26]
  wire  _GEN_2542 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2110 : uop_0_cf_exceptionVec_4; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2543 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2111 : uop_1_cf_exceptionVec_4; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2544 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2112 : uop_2_cf_exceptionVec_4; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2545 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2113 : uop_3_cf_exceptionVec_4; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2546 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2114 : uop_4_cf_exceptionVec_4; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2547 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2115 : uop_5_cf_exceptionVec_4; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2548 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2116 : uop_6_cf_exceptionVec_4; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2549 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2117 : uop_7_cf_exceptionVec_4; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2550 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2118 : uop_8_cf_exceptionVec_4; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2551 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2119 : uop_9_cf_exceptionVec_4; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2552 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2120 : uop_10_cf_exceptionVec_4; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2553 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2121 : uop_11_cf_exceptionVec_4; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2554 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2122 : uop_12_cf_exceptionVec_4; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2555 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2123 : uop_13_cf_exceptionVec_4; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2556 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2124 : uop_14_cf_exceptionVec_4; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2557 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2125 : uop_15_cf_exceptionVec_4; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2558 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2126 : uop_0_cf_exceptionVec_5; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2559 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2127 : uop_1_cf_exceptionVec_5; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2560 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2128 : uop_2_cf_exceptionVec_5; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2561 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2129 : uop_3_cf_exceptionVec_5; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2562 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2130 : uop_4_cf_exceptionVec_5; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2563 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2131 : uop_5_cf_exceptionVec_5; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2564 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2132 : uop_6_cf_exceptionVec_5; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2565 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2133 : uop_7_cf_exceptionVec_5; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2566 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2134 : uop_8_cf_exceptionVec_5; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2567 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2135 : uop_9_cf_exceptionVec_5; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2568 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2136 : uop_10_cf_exceptionVec_5; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2569 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2137 : uop_11_cf_exceptionVec_5; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2570 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2138 : uop_12_cf_exceptionVec_5; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2571 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2139 : uop_13_cf_exceptionVec_5; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2572 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2140 : uop_14_cf_exceptionVec_5; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2573 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2141 : uop_15_cf_exceptionVec_5; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2686 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2254 : uop_0_cf_exceptionVec_13; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2687 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2255 : uop_1_cf_exceptionVec_13; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2688 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2256 : uop_2_cf_exceptionVec_13; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2689 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2257 : uop_3_cf_exceptionVec_13; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2690 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2258 : uop_4_cf_exceptionVec_13; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2691 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2259 : uop_5_cf_exceptionVec_13; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2692 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2260 : uop_6_cf_exceptionVec_13; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2693 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2261 : uop_7_cf_exceptionVec_13; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2694 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2262 : uop_8_cf_exceptionVec_13; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2695 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2263 : uop_9_cf_exceptionVec_13; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2696 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2264 : uop_10_cf_exceptionVec_13; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2697 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2265 : uop_11_cf_exceptionVec_13; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2698 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2266 : uop_12_cf_exceptionVec_13; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2699 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2267 : uop_13_cf_exceptionVec_13; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2700 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2268 : uop_14_cf_exceptionVec_13; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2701 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2269 : uop_15_cf_exceptionVec_13; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2814 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_670 : uop_0_cf_trigger_backendEn_1; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2815 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_671 : uop_1_cf_trigger_backendEn_1; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2816 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_672 : uop_2_cf_trigger_backendEn_1; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2817 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_673 : uop_3_cf_trigger_backendEn_1; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2818 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_674 : uop_4_cf_trigger_backendEn_1; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2819 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_675 : uop_5_cf_trigger_backendEn_1; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2820 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_676 : uop_6_cf_trigger_backendEn_1; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2821 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_677 : uop_7_cf_trigger_backendEn_1; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2822 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_678 : uop_8_cf_trigger_backendEn_1; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2823 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_679 : uop_9_cf_trigger_backendEn_1; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2824 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_680 : uop_10_cf_trigger_backendEn_1; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2825 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_681 : uop_11_cf_trigger_backendEn_1; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2826 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_682 : uop_12_cf_trigger_backendEn_1; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2827 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_683 : uop_13_cf_trigger_backendEn_1; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2828 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_684 : uop_14_cf_trigger_backendEn_1; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2829 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_685 : uop_15_cf_trigger_backendEn_1; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2830 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_686 : uop_0_cf_trigger_backendHit_0; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2831 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_687 : uop_1_cf_trigger_backendHit_0; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2832 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_688 : uop_2_cf_trigger_backendHit_0; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2833 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_689 : uop_3_cf_trigger_backendHit_0; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2834 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_690 : uop_4_cf_trigger_backendHit_0; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2835 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_691 : uop_5_cf_trigger_backendHit_0; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2836 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_692 : uop_6_cf_trigger_backendHit_0; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2837 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_693 : uop_7_cf_trigger_backendHit_0; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2838 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_694 : uop_8_cf_trigger_backendHit_0; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2839 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_695 : uop_9_cf_trigger_backendHit_0; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2840 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_696 : uop_10_cf_trigger_backendHit_0; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2841 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_697 : uop_11_cf_trigger_backendHit_0; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2842 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_698 : uop_12_cf_trigger_backendHit_0; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2843 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_699 : uop_13_cf_trigger_backendHit_0; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2844 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_700 : uop_14_cf_trigger_backendHit_0; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2845 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_701 : uop_15_cf_trigger_backendHit_0; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2846 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_702 : uop_0_cf_trigger_backendHit_1; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2847 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_703 : uop_1_cf_trigger_backendHit_1; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2848 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_704 : uop_2_cf_trigger_backendHit_1; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2849 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_705 : uop_3_cf_trigger_backendHit_1; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2850 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_706 : uop_4_cf_trigger_backendHit_1; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2851 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_707 : uop_5_cf_trigger_backendHit_1; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2852 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_708 : uop_6_cf_trigger_backendHit_1; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2853 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_709 : uop_7_cf_trigger_backendHit_1; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2854 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_710 : uop_8_cf_trigger_backendHit_1; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2855 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_711 : uop_9_cf_trigger_backendHit_1; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2856 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_712 : uop_10_cf_trigger_backendHit_1; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2857 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_713 : uop_11_cf_trigger_backendHit_1; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2858 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_714 : uop_12_cf_trigger_backendHit_1; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2859 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_715 : uop_13_cf_trigger_backendHit_1; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2860 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_716 : uop_14_cf_trigger_backendHit_1; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2861 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_717 : uop_15_cf_trigger_backendHit_1; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2894 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_750 : uop_0_cf_trigger_backendHit_4; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2895 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_751 : uop_1_cf_trigger_backendHit_4; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2896 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_752 : uop_2_cf_trigger_backendHit_4; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2897 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_753 : uop_3_cf_trigger_backendHit_4; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2898 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_754 : uop_4_cf_trigger_backendHit_4; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2899 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_755 : uop_5_cf_trigger_backendHit_4; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2900 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_756 : uop_6_cf_trigger_backendHit_4; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2901 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_757 : uop_7_cf_trigger_backendHit_4; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2902 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_758 : uop_8_cf_trigger_backendHit_4; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2903 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_759 : uop_9_cf_trigger_backendHit_4; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2904 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_760 : uop_10_cf_trigger_backendHit_4; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2905 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_761 : uop_11_cf_trigger_backendHit_4; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2906 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_762 : uop_12_cf_trigger_backendHit_4; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2907 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_763 : uop_13_cf_trigger_backendHit_4; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2908 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_764 : uop_14_cf_trigger_backendHit_4; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_2909 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_765 : uop_15_cf_trigger_backendHit_4; // @[LoadQueueFlag.scala 204:43 62:16]
  wire [6:0] _GEN_3326 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1182 : uop_0_ctrl_fuOpType; // @[LoadQueueFlag.scala 204:43 62:16]
  wire [6:0] _GEN_3327 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1183 : uop_1_ctrl_fuOpType; // @[LoadQueueFlag.scala 204:43 62:16]
  wire [6:0] _GEN_3328 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1184 : uop_2_ctrl_fuOpType; // @[LoadQueueFlag.scala 204:43 62:16]
  wire [6:0] _GEN_3329 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1185 : uop_3_ctrl_fuOpType; // @[LoadQueueFlag.scala 204:43 62:16]
  wire [6:0] _GEN_3330 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1186 : uop_4_ctrl_fuOpType; // @[LoadQueueFlag.scala 204:43 62:16]
  wire [6:0] _GEN_3331 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1187 : uop_5_ctrl_fuOpType; // @[LoadQueueFlag.scala 204:43 62:16]
  wire [6:0] _GEN_3332 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1188 : uop_6_ctrl_fuOpType; // @[LoadQueueFlag.scala 204:43 62:16]
  wire [6:0] _GEN_3333 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1189 : uop_7_ctrl_fuOpType; // @[LoadQueueFlag.scala 204:43 62:16]
  wire [6:0] _GEN_3334 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1190 : uop_8_ctrl_fuOpType; // @[LoadQueueFlag.scala 204:43 62:16]
  wire [6:0] _GEN_3335 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1191 : uop_9_ctrl_fuOpType; // @[LoadQueueFlag.scala 204:43 62:16]
  wire [6:0] _GEN_3336 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1192 : uop_10_ctrl_fuOpType; // @[LoadQueueFlag.scala 204:43 62:16]
  wire [6:0] _GEN_3337 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1193 : uop_11_ctrl_fuOpType; // @[LoadQueueFlag.scala 204:43 62:16]
  wire [6:0] _GEN_3338 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1194 : uop_12_ctrl_fuOpType; // @[LoadQueueFlag.scala 204:43 62:16]
  wire [6:0] _GEN_3339 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1195 : uop_13_ctrl_fuOpType; // @[LoadQueueFlag.scala 204:43 62:16]
  wire [6:0] _GEN_3340 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1196 : uop_14_ctrl_fuOpType; // @[LoadQueueFlag.scala 204:43 62:16]
  wire [6:0] _GEN_3341 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1197 : uop_15_ctrl_fuOpType; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_3342 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1198 : uop_0_ctrl_rfWen; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_3343 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1199 : uop_1_ctrl_rfWen; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_3344 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1200 : uop_2_ctrl_rfWen; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_3345 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1201 : uop_3_ctrl_rfWen; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_3346 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1202 : uop_4_ctrl_rfWen; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_3347 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1203 : uop_5_ctrl_rfWen; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_3348 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1204 : uop_6_ctrl_rfWen; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_3349 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1205 : uop_7_ctrl_rfWen; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_3350 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1206 : uop_8_ctrl_rfWen; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_3351 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1207 : uop_9_ctrl_rfWen; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_3352 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1208 : uop_10_ctrl_rfWen; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_3353 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1209 : uop_11_ctrl_rfWen; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_3354 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1210 : uop_12_ctrl_rfWen; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_3355 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1211 : uop_13_ctrl_rfWen; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_3356 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1212 : uop_14_ctrl_rfWen; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_3357 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1213 : uop_15_ctrl_rfWen; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_3358 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1214 : uop_0_ctrl_fpWen; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_3359 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1215 : uop_1_ctrl_fpWen; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_3360 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1216 : uop_2_ctrl_fpWen; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_3361 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1217 : uop_3_ctrl_fpWen; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_3362 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1218 : uop_4_ctrl_fpWen; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_3363 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1219 : uop_5_ctrl_fpWen; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_3364 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1220 : uop_6_ctrl_fpWen; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_3365 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1221 : uop_7_ctrl_fpWen; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_3366 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1222 : uop_8_ctrl_fpWen; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_3367 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1223 : uop_9_ctrl_fpWen; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_3368 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1224 : uop_10_ctrl_fpWen; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_3369 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1225 : uop_11_ctrl_fpWen; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_3370 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1226 : uop_12_ctrl_fpWen; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_3371 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1227 : uop_13_ctrl_fpWen; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_3372 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1228 : uop_14_ctrl_fpWen; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_3373 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1229 : uop_15_ctrl_fpWen; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_3422 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1278 : uop_0_ctrl_flushPipe; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_3423 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1279 : uop_1_ctrl_flushPipe; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_3424 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1280 : uop_2_ctrl_flushPipe; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_3425 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1281 : uop_3_ctrl_flushPipe; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_3426 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1282 : uop_4_ctrl_flushPipe; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_3427 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1283 : uop_5_ctrl_flushPipe; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_3428 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1284 : uop_6_ctrl_flushPipe; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_3429 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1285 : uop_7_ctrl_flushPipe; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_3430 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1286 : uop_8_ctrl_flushPipe; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_3431 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1287 : uop_9_ctrl_flushPipe; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_3432 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1288 : uop_10_ctrl_flushPipe; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_3433 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1289 : uop_11_ctrl_flushPipe; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_3434 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1290 : uop_12_ctrl_flushPipe; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_3435 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1291 : uop_13_ctrl_flushPipe; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_3436 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1292 : uop_14_ctrl_flushPipe; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_3437 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1293 : uop_15_ctrl_flushPipe; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_3742 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1598 : uop_0_ctrl_replayInst; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_3743 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1599 : uop_1_ctrl_replayInst; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_3744 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1600 : uop_2_ctrl_replayInst; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_3745 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1601 : uop_3_ctrl_replayInst; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_3746 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1602 : uop_4_ctrl_replayInst; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_3747 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1603 : uop_5_ctrl_replayInst; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_3748 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1604 : uop_6_ctrl_replayInst; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_3749 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1605 : uop_7_ctrl_replayInst; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_3750 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1606 : uop_8_ctrl_replayInst; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_3751 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1607 : uop_9_ctrl_replayInst; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_3752 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1608 : uop_10_ctrl_replayInst; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_3753 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1609 : uop_11_ctrl_replayInst; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_3754 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1610 : uop_12_ctrl_replayInst; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_3755 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1611 : uop_13_ctrl_replayInst; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_3756 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1612 : uop_14_ctrl_replayInst; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_3757 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1613 : uop_15_ctrl_replayInst; // @[LoadQueueFlag.scala 204:43 62:16]
  wire [5:0] _GEN_3854 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1710 : uop_0_pdest; // @[LoadQueueFlag.scala 204:43 62:16]
  wire [5:0] _GEN_3855 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1711 : uop_1_pdest; // @[LoadQueueFlag.scala 204:43 62:16]
  wire [5:0] _GEN_3856 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1712 : uop_2_pdest; // @[LoadQueueFlag.scala 204:43 62:16]
  wire [5:0] _GEN_3857 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1713 : uop_3_pdest; // @[LoadQueueFlag.scala 204:43 62:16]
  wire [5:0] _GEN_3858 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1714 : uop_4_pdest; // @[LoadQueueFlag.scala 204:43 62:16]
  wire [5:0] _GEN_3859 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1715 : uop_5_pdest; // @[LoadQueueFlag.scala 204:43 62:16]
  wire [5:0] _GEN_3860 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1716 : uop_6_pdest; // @[LoadQueueFlag.scala 204:43 62:16]
  wire [5:0] _GEN_3861 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1717 : uop_7_pdest; // @[LoadQueueFlag.scala 204:43 62:16]
  wire [5:0] _GEN_3862 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1718 : uop_8_pdest; // @[LoadQueueFlag.scala 204:43 62:16]
  wire [5:0] _GEN_3863 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1719 : uop_9_pdest; // @[LoadQueueFlag.scala 204:43 62:16]
  wire [5:0] _GEN_3864 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1720 : uop_10_pdest; // @[LoadQueueFlag.scala 204:43 62:16]
  wire [5:0] _GEN_3865 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1721 : uop_11_pdest; // @[LoadQueueFlag.scala 204:43 62:16]
  wire [5:0] _GEN_3866 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1722 : uop_12_pdest; // @[LoadQueueFlag.scala 204:43 62:16]
  wire [5:0] _GEN_3867 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1723 : uop_13_pdest; // @[LoadQueueFlag.scala 204:43 62:16]
  wire [5:0] _GEN_3868 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1724 : uop_14_pdest; // @[LoadQueueFlag.scala 204:43 62:16]
  wire [5:0] _GEN_3869 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1725 : uop_15_pdest; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_3886 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1742 : uop_0_robIdx_flag; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_3887 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1743 : uop_1_robIdx_flag; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_3888 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1744 : uop_2_robIdx_flag; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_3889 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1745 : uop_3_robIdx_flag; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_3890 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1746 : uop_4_robIdx_flag; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_3891 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1747 : uop_5_robIdx_flag; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_3892 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1748 : uop_6_robIdx_flag; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_3893 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1749 : uop_7_robIdx_flag; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_3894 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1750 : uop_8_robIdx_flag; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_3895 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1751 : uop_9_robIdx_flag; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_3896 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1752 : uop_10_robIdx_flag; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_3897 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1753 : uop_11_robIdx_flag; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_3898 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1754 : uop_12_robIdx_flag; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_3899 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1755 : uop_13_robIdx_flag; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_3900 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1756 : uop_14_robIdx_flag; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_3901 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1757 : uop_15_robIdx_flag; // @[LoadQueueFlag.scala 204:43 62:16]
  wire [4:0] _GEN_3902 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1758 : uop_0_robIdx_value; // @[LoadQueueFlag.scala 204:43 62:16]
  wire [4:0] _GEN_3903 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1759 : uop_1_robIdx_value; // @[LoadQueueFlag.scala 204:43 62:16]
  wire [4:0] _GEN_3904 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1760 : uop_2_robIdx_value; // @[LoadQueueFlag.scala 204:43 62:16]
  wire [4:0] _GEN_3905 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1761 : uop_3_robIdx_value; // @[LoadQueueFlag.scala 204:43 62:16]
  wire [4:0] _GEN_3906 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1762 : uop_4_robIdx_value; // @[LoadQueueFlag.scala 204:43 62:16]
  wire [4:0] _GEN_3907 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1763 : uop_5_robIdx_value; // @[LoadQueueFlag.scala 204:43 62:16]
  wire [4:0] _GEN_3908 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1764 : uop_6_robIdx_value; // @[LoadQueueFlag.scala 204:43 62:16]
  wire [4:0] _GEN_3909 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1765 : uop_7_robIdx_value; // @[LoadQueueFlag.scala 204:43 62:16]
  wire [4:0] _GEN_3910 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1766 : uop_8_robIdx_value; // @[LoadQueueFlag.scala 204:43 62:16]
  wire [4:0] _GEN_3911 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1767 : uop_9_robIdx_value; // @[LoadQueueFlag.scala 204:43 62:16]
  wire [4:0] _GEN_3912 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1768 : uop_10_robIdx_value; // @[LoadQueueFlag.scala 204:43 62:16]
  wire [4:0] _GEN_3913 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1769 : uop_11_robIdx_value; // @[LoadQueueFlag.scala 204:43 62:16]
  wire [4:0] _GEN_3914 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1770 : uop_12_robIdx_value; // @[LoadQueueFlag.scala 204:43 62:16]
  wire [4:0] _GEN_3915 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1771 : uop_13_robIdx_value; // @[LoadQueueFlag.scala 204:43 62:16]
  wire [4:0] _GEN_3916 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1772 : uop_14_robIdx_value; // @[LoadQueueFlag.scala 204:43 62:16]
  wire [4:0] _GEN_3917 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_1773 : uop_15_robIdx_value; // @[LoadQueueFlag.scala 204:43 62:16]
  wire  _GEN_4158 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2302 : addrvalid_0; // @[LoadQueueFlag.scala 204:43 90:26]
  wire  _GEN_4159 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2303 : addrvalid_1; // @[LoadQueueFlag.scala 204:43 90:26]
  wire  _GEN_4160 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2304 : addrvalid_2; // @[LoadQueueFlag.scala 204:43 90:26]
  wire  _GEN_4161 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2305 : addrvalid_3; // @[LoadQueueFlag.scala 204:43 90:26]
  wire  _GEN_4162 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2306 : addrvalid_4; // @[LoadQueueFlag.scala 204:43 90:26]
  wire  _GEN_4163 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2307 : addrvalid_5; // @[LoadQueueFlag.scala 204:43 90:26]
  wire  _GEN_4164 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2308 : addrvalid_6; // @[LoadQueueFlag.scala 204:43 90:26]
  wire  _GEN_4165 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2309 : addrvalid_7; // @[LoadQueueFlag.scala 204:43 90:26]
  wire  _GEN_4166 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2310 : addrvalid_8; // @[LoadQueueFlag.scala 204:43 90:26]
  wire  _GEN_4167 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2311 : addrvalid_9; // @[LoadQueueFlag.scala 204:43 90:26]
  wire  _GEN_4168 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2312 : addrvalid_10; // @[LoadQueueFlag.scala 204:43 90:26]
  wire  _GEN_4169 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2313 : addrvalid_11; // @[LoadQueueFlag.scala 204:43 90:26]
  wire  _GEN_4170 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2314 : addrvalid_12; // @[LoadQueueFlag.scala 204:43 90:26]
  wire  _GEN_4171 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2315 : addrvalid_13; // @[LoadQueueFlag.scala 204:43 90:26]
  wire  _GEN_4172 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2316 : addrvalid_14; // @[LoadQueueFlag.scala 204:43 90:26]
  wire  _GEN_4173 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2317 : addrvalid_15; // @[LoadQueueFlag.scala 204:43 90:26]
  wire  _GEN_4174 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2318 : datavalid_0; // @[LoadQueueFlag.scala 204:43 91:26]
  wire  _GEN_4175 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2319 : datavalid_1; // @[LoadQueueFlag.scala 204:43 91:26]
  wire  _GEN_4176 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2320 : datavalid_2; // @[LoadQueueFlag.scala 204:43 91:26]
  wire  _GEN_4177 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2321 : datavalid_3; // @[LoadQueueFlag.scala 204:43 91:26]
  wire  _GEN_4178 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2322 : datavalid_4; // @[LoadQueueFlag.scala 204:43 91:26]
  wire  _GEN_4179 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2323 : datavalid_5; // @[LoadQueueFlag.scala 204:43 91:26]
  wire  _GEN_4180 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2324 : datavalid_6; // @[LoadQueueFlag.scala 204:43 91:26]
  wire  _GEN_4181 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2325 : datavalid_7; // @[LoadQueueFlag.scala 204:43 91:26]
  wire  _GEN_4182 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2326 : datavalid_8; // @[LoadQueueFlag.scala 204:43 91:26]
  wire  _GEN_4183 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2327 : datavalid_9; // @[LoadQueueFlag.scala 204:43 91:26]
  wire  _GEN_4184 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2328 : datavalid_10; // @[LoadQueueFlag.scala 204:43 91:26]
  wire  _GEN_4185 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2329 : datavalid_11; // @[LoadQueueFlag.scala 204:43 91:26]
  wire  _GEN_4186 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2330 : datavalid_12; // @[LoadQueueFlag.scala 204:43 91:26]
  wire  _GEN_4187 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2331 : datavalid_13; // @[LoadQueueFlag.scala 204:43 91:26]
  wire  _GEN_4188 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2332 : datavalid_14; // @[LoadQueueFlag.scala 204:43 91:26]
  wire  _GEN_4189 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2333 : datavalid_15; // @[LoadQueueFlag.scala 204:43 91:26]
  wire  _GEN_4190 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2334 : pending_0; // @[LoadQueueFlag.scala 204:43 92:24]
  wire  _GEN_4191 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2335 : pending_1; // @[LoadQueueFlag.scala 204:43 92:24]
  wire  _GEN_4192 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2336 : pending_2; // @[LoadQueueFlag.scala 204:43 92:24]
  wire  _GEN_4193 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2337 : pending_3; // @[LoadQueueFlag.scala 204:43 92:24]
  wire  _GEN_4194 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2338 : pending_4; // @[LoadQueueFlag.scala 204:43 92:24]
  wire  _GEN_4195 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2339 : pending_5; // @[LoadQueueFlag.scala 204:43 92:24]
  wire  _GEN_4196 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2340 : pending_6; // @[LoadQueueFlag.scala 204:43 92:24]
  wire  _GEN_4197 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2341 : pending_7; // @[LoadQueueFlag.scala 204:43 92:24]
  wire  _GEN_4198 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2342 : pending_8; // @[LoadQueueFlag.scala 204:43 92:24]
  wire  _GEN_4199 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2343 : pending_9; // @[LoadQueueFlag.scala 204:43 92:24]
  wire  _GEN_4200 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2344 : pending_10; // @[LoadQueueFlag.scala 204:43 92:24]
  wire  _GEN_4201 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2345 : pending_11; // @[LoadQueueFlag.scala 204:43 92:24]
  wire  _GEN_4202 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2346 : pending_12; // @[LoadQueueFlag.scala 204:43 92:24]
  wire  _GEN_4203 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2347 : pending_13; // @[LoadQueueFlag.scala 204:43 92:24]
  wire  _GEN_4204 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2348 : pending_14; // @[LoadQueueFlag.scala 204:43 92:24]
  wire  _GEN_4205 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2349 : pending_15; // @[LoadQueueFlag.scala 204:43 92:24]
  wire  _GEN_4206 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2350 : writebacked_0; // @[LoadQueueFlag.scala 204:43 93:28]
  wire  _GEN_4207 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2351 : writebacked_1; // @[LoadQueueFlag.scala 204:43 93:28]
  wire  _GEN_4208 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2352 : writebacked_2; // @[LoadQueueFlag.scala 204:43 93:28]
  wire  _GEN_4209 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2353 : writebacked_3; // @[LoadQueueFlag.scala 204:43 93:28]
  wire  _GEN_4210 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2354 : writebacked_4; // @[LoadQueueFlag.scala 204:43 93:28]
  wire  _GEN_4211 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2355 : writebacked_5; // @[LoadQueueFlag.scala 204:43 93:28]
  wire  _GEN_4212 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2356 : writebacked_6; // @[LoadQueueFlag.scala 204:43 93:28]
  wire  _GEN_4213 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2357 : writebacked_7; // @[LoadQueueFlag.scala 204:43 93:28]
  wire  _GEN_4214 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2358 : writebacked_8; // @[LoadQueueFlag.scala 204:43 93:28]
  wire  _GEN_4215 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2359 : writebacked_9; // @[LoadQueueFlag.scala 204:43 93:28]
  wire  _GEN_4216 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2360 : writebacked_10; // @[LoadQueueFlag.scala 204:43 93:28]
  wire  _GEN_4217 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2361 : writebacked_11; // @[LoadQueueFlag.scala 204:43 93:28]
  wire  _GEN_4218 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2362 : writebacked_12; // @[LoadQueueFlag.scala 204:43 93:28]
  wire  _GEN_4219 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2363 : writebacked_13; // @[LoadQueueFlag.scala 204:43 93:28]
  wire  _GEN_4220 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2364 : writebacked_14; // @[LoadQueueFlag.scala 204:43 93:28]
  wire  _GEN_4221 = io_enq_req_0_valid & ~enqCancel_0 ? _GEN_2365 : writebacked_15; // @[LoadQueueFlag.scala 204:43 93:28]
  wire  _GEN_4270 = 4'h0 == io_enq_req_1_bits_lqIdx_value | _GEN_2414; // @[LoadQueueFlag.scala 205:{24,24}]
  wire  _GEN_4271 = 4'h1 == io_enq_req_1_bits_lqIdx_value | _GEN_2415; // @[LoadQueueFlag.scala 205:{24,24}]
  wire  _GEN_4272 = 4'h2 == io_enq_req_1_bits_lqIdx_value | _GEN_2416; // @[LoadQueueFlag.scala 205:{24,24}]
  wire  _GEN_4273 = 4'h3 == io_enq_req_1_bits_lqIdx_value | _GEN_2417; // @[LoadQueueFlag.scala 205:{24,24}]
  wire  _GEN_4274 = 4'h4 == io_enq_req_1_bits_lqIdx_value | _GEN_2418; // @[LoadQueueFlag.scala 205:{24,24}]
  wire  _GEN_4275 = 4'h5 == io_enq_req_1_bits_lqIdx_value | _GEN_2419; // @[LoadQueueFlag.scala 205:{24,24}]
  wire  _GEN_4276 = 4'h6 == io_enq_req_1_bits_lqIdx_value | _GEN_2420; // @[LoadQueueFlag.scala 205:{24,24}]
  wire  _GEN_4277 = 4'h7 == io_enq_req_1_bits_lqIdx_value | _GEN_2421; // @[LoadQueueFlag.scala 205:{24,24}]
  wire  _GEN_4278 = 4'h8 == io_enq_req_1_bits_lqIdx_value | _GEN_2422; // @[LoadQueueFlag.scala 205:{24,24}]
  wire  _GEN_4279 = 4'h9 == io_enq_req_1_bits_lqIdx_value | _GEN_2423; // @[LoadQueueFlag.scala 205:{24,24}]
  wire  _GEN_4280 = 4'ha == io_enq_req_1_bits_lqIdx_value | _GEN_2424; // @[LoadQueueFlag.scala 205:{24,24}]
  wire  _GEN_4281 = 4'hb == io_enq_req_1_bits_lqIdx_value | _GEN_2425; // @[LoadQueueFlag.scala 205:{24,24}]
  wire  _GEN_4282 = 4'hc == io_enq_req_1_bits_lqIdx_value | _GEN_2426; // @[LoadQueueFlag.scala 205:{24,24}]
  wire  _GEN_4283 = 4'hd == io_enq_req_1_bits_lqIdx_value | _GEN_2427; // @[LoadQueueFlag.scala 205:{24,24}]
  wire  _GEN_4284 = 4'he == io_enq_req_1_bits_lqIdx_value | _GEN_2428; // @[LoadQueueFlag.scala 205:{24,24}]
  wire  _GEN_4285 = 4'hf == io_enq_req_1_bits_lqIdx_value | _GEN_2429; // @[LoadQueueFlag.scala 205:{24,24}]
  wire  _GEN_4398 = 4'h0 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2542; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4399 = 4'h1 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2543; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4400 = 4'h2 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2544; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4401 = 4'h3 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2545; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4402 = 4'h4 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2546; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4403 = 4'h5 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2547; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4404 = 4'h6 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2548; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4405 = 4'h7 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2549; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4406 = 4'h8 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2550; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4407 = 4'h9 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2551; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4408 = 4'ha == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2552; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4409 = 4'hb == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2553; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4410 = 4'hc == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2554; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4411 = 4'hd == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2555; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4412 = 4'he == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2556; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4413 = 4'hf == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2557; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4414 = 4'h0 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2558; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4415 = 4'h1 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2559; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4416 = 4'h2 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2560; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4417 = 4'h3 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2561; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4418 = 4'h4 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2562; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4419 = 4'h5 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2563; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4420 = 4'h6 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2564; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4421 = 4'h7 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2565; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4422 = 4'h8 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2566; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4423 = 4'h9 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2567; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4424 = 4'ha == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2568; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4425 = 4'hb == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2569; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4426 = 4'hc == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2570; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4427 = 4'hd == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2571; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4428 = 4'he == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2572; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4429 = 4'hf == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2573; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4542 = 4'h0 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2686; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4543 = 4'h1 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2687; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4544 = 4'h2 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2688; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4545 = 4'h3 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2689; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4546 = 4'h4 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2690; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4547 = 4'h5 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2691; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4548 = 4'h6 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2692; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4549 = 4'h7 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2693; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4550 = 4'h8 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2694; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4551 = 4'h9 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2695; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4552 = 4'ha == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2696; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4553 = 4'hb == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2697; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4554 = 4'hc == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2698; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4555 = 4'hd == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2699; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4556 = 4'he == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2700; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4557 = 4'hf == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2701; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4670 = 4'h0 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_cf_trigger_backendEn_1 : _GEN_2814; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4671 = 4'h1 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_cf_trigger_backendEn_1 : _GEN_2815; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4672 = 4'h2 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_cf_trigger_backendEn_1 : _GEN_2816; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4673 = 4'h3 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_cf_trigger_backendEn_1 : _GEN_2817; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4674 = 4'h4 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_cf_trigger_backendEn_1 : _GEN_2818; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4675 = 4'h5 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_cf_trigger_backendEn_1 : _GEN_2819; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4676 = 4'h6 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_cf_trigger_backendEn_1 : _GEN_2820; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4677 = 4'h7 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_cf_trigger_backendEn_1 : _GEN_2821; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4678 = 4'h8 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_cf_trigger_backendEn_1 : _GEN_2822; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4679 = 4'h9 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_cf_trigger_backendEn_1 : _GEN_2823; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4680 = 4'ha == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_cf_trigger_backendEn_1 : _GEN_2824; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4681 = 4'hb == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_cf_trigger_backendEn_1 : _GEN_2825; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4682 = 4'hc == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_cf_trigger_backendEn_1 : _GEN_2826; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4683 = 4'hd == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_cf_trigger_backendEn_1 : _GEN_2827; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4684 = 4'he == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_cf_trigger_backendEn_1 : _GEN_2828; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4685 = 4'hf == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_cf_trigger_backendEn_1 : _GEN_2829; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4686 = 4'h0 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2830; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4687 = 4'h1 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2831; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4688 = 4'h2 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2832; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4689 = 4'h3 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2833; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4690 = 4'h4 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2834; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4691 = 4'h5 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2835; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4692 = 4'h6 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2836; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4693 = 4'h7 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2837; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4694 = 4'h8 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2838; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4695 = 4'h9 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2839; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4696 = 4'ha == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2840; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4697 = 4'hb == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2841; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4698 = 4'hc == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2842; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4699 = 4'hd == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2843; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4700 = 4'he == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2844; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4701 = 4'hf == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2845; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4702 = 4'h0 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2846; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4703 = 4'h1 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2847; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4704 = 4'h2 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2848; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4705 = 4'h3 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2849; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4706 = 4'h4 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2850; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4707 = 4'h5 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2851; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4708 = 4'h6 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2852; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4709 = 4'h7 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2853; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4710 = 4'h8 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2854; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4711 = 4'h9 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2855; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4712 = 4'ha == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2856; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4713 = 4'hb == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2857; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4714 = 4'hc == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2858; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4715 = 4'hd == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2859; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4716 = 4'he == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2860; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4717 = 4'hf == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2861; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4750 = 4'h0 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2894; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4751 = 4'h1 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2895; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4752 = 4'h2 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2896; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4753 = 4'h3 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2897; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4754 = 4'h4 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2898; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4755 = 4'h5 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2899; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4756 = 4'h6 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2900; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4757 = 4'h7 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2901; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4758 = 4'h8 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2902; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4759 = 4'h9 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2903; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4760 = 4'ha == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2904; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4761 = 4'hb == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2905; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4762 = 4'hc == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2906; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4763 = 4'hd == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2907; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4764 = 4'he == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2908; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_4765 = 4'hf == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_2909; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [6:0] _GEN_5182 = 4'h0 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_ctrl_fuOpType : _GEN_3326; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [6:0] _GEN_5183 = 4'h1 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_ctrl_fuOpType : _GEN_3327; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [6:0] _GEN_5184 = 4'h2 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_ctrl_fuOpType : _GEN_3328; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [6:0] _GEN_5185 = 4'h3 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_ctrl_fuOpType : _GEN_3329; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [6:0] _GEN_5186 = 4'h4 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_ctrl_fuOpType : _GEN_3330; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [6:0] _GEN_5187 = 4'h5 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_ctrl_fuOpType : _GEN_3331; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [6:0] _GEN_5188 = 4'h6 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_ctrl_fuOpType : _GEN_3332; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [6:0] _GEN_5189 = 4'h7 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_ctrl_fuOpType : _GEN_3333; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [6:0] _GEN_5190 = 4'h8 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_ctrl_fuOpType : _GEN_3334; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [6:0] _GEN_5191 = 4'h9 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_ctrl_fuOpType : _GEN_3335; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [6:0] _GEN_5192 = 4'ha == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_ctrl_fuOpType : _GEN_3336; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [6:0] _GEN_5193 = 4'hb == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_ctrl_fuOpType : _GEN_3337; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [6:0] _GEN_5194 = 4'hc == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_ctrl_fuOpType : _GEN_3338; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [6:0] _GEN_5195 = 4'hd == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_ctrl_fuOpType : _GEN_3339; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [6:0] _GEN_5196 = 4'he == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_ctrl_fuOpType : _GEN_3340; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [6:0] _GEN_5197 = 4'hf == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_ctrl_fuOpType : _GEN_3341; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_5198 = 4'h0 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_ctrl_rfWen : _GEN_3342; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_5199 = 4'h1 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_ctrl_rfWen : _GEN_3343; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_5200 = 4'h2 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_ctrl_rfWen : _GEN_3344; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_5201 = 4'h3 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_ctrl_rfWen : _GEN_3345; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_5202 = 4'h4 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_ctrl_rfWen : _GEN_3346; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_5203 = 4'h5 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_ctrl_rfWen : _GEN_3347; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_5204 = 4'h6 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_ctrl_rfWen : _GEN_3348; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_5205 = 4'h7 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_ctrl_rfWen : _GEN_3349; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_5206 = 4'h8 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_ctrl_rfWen : _GEN_3350; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_5207 = 4'h9 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_ctrl_rfWen : _GEN_3351; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_5208 = 4'ha == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_ctrl_rfWen : _GEN_3352; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_5209 = 4'hb == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_ctrl_rfWen : _GEN_3353; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_5210 = 4'hc == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_ctrl_rfWen : _GEN_3354; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_5211 = 4'hd == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_ctrl_rfWen : _GEN_3355; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_5212 = 4'he == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_ctrl_rfWen : _GEN_3356; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_5213 = 4'hf == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_ctrl_rfWen : _GEN_3357; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_5214 = 4'h0 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_ctrl_fpWen : _GEN_3358; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_5215 = 4'h1 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_ctrl_fpWen : _GEN_3359; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_5216 = 4'h2 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_ctrl_fpWen : _GEN_3360; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_5217 = 4'h3 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_ctrl_fpWen : _GEN_3361; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_5218 = 4'h4 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_ctrl_fpWen : _GEN_3362; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_5219 = 4'h5 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_ctrl_fpWen : _GEN_3363; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_5220 = 4'h6 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_ctrl_fpWen : _GEN_3364; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_5221 = 4'h7 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_ctrl_fpWen : _GEN_3365; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_5222 = 4'h8 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_ctrl_fpWen : _GEN_3366; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_5223 = 4'h9 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_ctrl_fpWen : _GEN_3367; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_5224 = 4'ha == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_ctrl_fpWen : _GEN_3368; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_5225 = 4'hb == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_ctrl_fpWen : _GEN_3369; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_5226 = 4'hc == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_ctrl_fpWen : _GEN_3370; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_5227 = 4'hd == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_ctrl_fpWen : _GEN_3371; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_5228 = 4'he == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_ctrl_fpWen : _GEN_3372; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_5229 = 4'hf == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_ctrl_fpWen : _GEN_3373; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_5278 = 4'h0 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_ctrl_flushPipe : _GEN_3422; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_5279 = 4'h1 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_ctrl_flushPipe : _GEN_3423; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_5280 = 4'h2 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_ctrl_flushPipe : _GEN_3424; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_5281 = 4'h3 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_ctrl_flushPipe : _GEN_3425; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_5282 = 4'h4 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_ctrl_flushPipe : _GEN_3426; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_5283 = 4'h5 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_ctrl_flushPipe : _GEN_3427; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_5284 = 4'h6 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_ctrl_flushPipe : _GEN_3428; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_5285 = 4'h7 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_ctrl_flushPipe : _GEN_3429; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_5286 = 4'h8 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_ctrl_flushPipe : _GEN_3430; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_5287 = 4'h9 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_ctrl_flushPipe : _GEN_3431; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_5288 = 4'ha == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_ctrl_flushPipe : _GEN_3432; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_5289 = 4'hb == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_ctrl_flushPipe : _GEN_3433; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_5290 = 4'hc == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_ctrl_flushPipe : _GEN_3434; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_5291 = 4'hd == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_ctrl_flushPipe : _GEN_3435; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_5292 = 4'he == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_ctrl_flushPipe : _GEN_3436; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_5293 = 4'hf == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_ctrl_flushPipe : _GEN_3437; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_5598 = 4'h0 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_ctrl_replayInst : _GEN_3742; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_5599 = 4'h1 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_ctrl_replayInst : _GEN_3743; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_5600 = 4'h2 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_ctrl_replayInst : _GEN_3744; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_5601 = 4'h3 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_ctrl_replayInst : _GEN_3745; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_5602 = 4'h4 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_ctrl_replayInst : _GEN_3746; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_5603 = 4'h5 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_ctrl_replayInst : _GEN_3747; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_5604 = 4'h6 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_ctrl_replayInst : _GEN_3748; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_5605 = 4'h7 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_ctrl_replayInst : _GEN_3749; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_5606 = 4'h8 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_ctrl_replayInst : _GEN_3750; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_5607 = 4'h9 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_ctrl_replayInst : _GEN_3751; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_5608 = 4'ha == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_ctrl_replayInst : _GEN_3752; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_5609 = 4'hb == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_ctrl_replayInst : _GEN_3753; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_5610 = 4'hc == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_ctrl_replayInst : _GEN_3754; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_5611 = 4'hd == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_ctrl_replayInst : _GEN_3755; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_5612 = 4'he == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_ctrl_replayInst : _GEN_3756; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_5613 = 4'hf == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_ctrl_replayInst : _GEN_3757; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [5:0] _GEN_5710 = 4'h0 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_pdest : _GEN_3854; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [5:0] _GEN_5711 = 4'h1 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_pdest : _GEN_3855; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [5:0] _GEN_5712 = 4'h2 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_pdest : _GEN_3856; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [5:0] _GEN_5713 = 4'h3 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_pdest : _GEN_3857; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [5:0] _GEN_5714 = 4'h4 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_pdest : _GEN_3858; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [5:0] _GEN_5715 = 4'h5 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_pdest : _GEN_3859; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [5:0] _GEN_5716 = 4'h6 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_pdest : _GEN_3860; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [5:0] _GEN_5717 = 4'h7 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_pdest : _GEN_3861; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [5:0] _GEN_5718 = 4'h8 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_pdest : _GEN_3862; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [5:0] _GEN_5719 = 4'h9 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_pdest : _GEN_3863; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [5:0] _GEN_5720 = 4'ha == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_pdest : _GEN_3864; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [5:0] _GEN_5721 = 4'hb == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_pdest : _GEN_3865; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [5:0] _GEN_5722 = 4'hc == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_pdest : _GEN_3866; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [5:0] _GEN_5723 = 4'hd == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_pdest : _GEN_3867; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [5:0] _GEN_5724 = 4'he == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_pdest : _GEN_3868; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [5:0] _GEN_5725 = 4'hf == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_pdest : _GEN_3869; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_5742 = 4'h0 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_robIdx_flag : _GEN_3886; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_5743 = 4'h1 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_robIdx_flag : _GEN_3887; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_5744 = 4'h2 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_robIdx_flag : _GEN_3888; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_5745 = 4'h3 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_robIdx_flag : _GEN_3889; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_5746 = 4'h4 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_robIdx_flag : _GEN_3890; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_5747 = 4'h5 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_robIdx_flag : _GEN_3891; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_5748 = 4'h6 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_robIdx_flag : _GEN_3892; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_5749 = 4'h7 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_robIdx_flag : _GEN_3893; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_5750 = 4'h8 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_robIdx_flag : _GEN_3894; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_5751 = 4'h9 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_robIdx_flag : _GEN_3895; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_5752 = 4'ha == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_robIdx_flag : _GEN_3896; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_5753 = 4'hb == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_robIdx_flag : _GEN_3897; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_5754 = 4'hc == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_robIdx_flag : _GEN_3898; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_5755 = 4'hd == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_robIdx_flag : _GEN_3899; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_5756 = 4'he == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_robIdx_flag : _GEN_3900; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_5757 = 4'hf == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_robIdx_flag : _GEN_3901; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [4:0] _GEN_5758 = 4'h0 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_robIdx_value : _GEN_3902; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [4:0] _GEN_5759 = 4'h1 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_robIdx_value : _GEN_3903; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [4:0] _GEN_5760 = 4'h2 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_robIdx_value : _GEN_3904; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [4:0] _GEN_5761 = 4'h3 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_robIdx_value : _GEN_3905; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [4:0] _GEN_5762 = 4'h4 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_robIdx_value : _GEN_3906; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [4:0] _GEN_5763 = 4'h5 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_robIdx_value : _GEN_3907; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [4:0] _GEN_5764 = 4'h6 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_robIdx_value : _GEN_3908; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [4:0] _GEN_5765 = 4'h7 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_robIdx_value : _GEN_3909; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [4:0] _GEN_5766 = 4'h8 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_robIdx_value : _GEN_3910; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [4:0] _GEN_5767 = 4'h9 == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_robIdx_value : _GEN_3911; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [4:0] _GEN_5768 = 4'ha == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_robIdx_value : _GEN_3912; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [4:0] _GEN_5769 = 4'hb == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_robIdx_value : _GEN_3913; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [4:0] _GEN_5770 = 4'hc == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_robIdx_value : _GEN_3914; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [4:0] _GEN_5771 = 4'hd == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_robIdx_value : _GEN_3915; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [4:0] _GEN_5772 = 4'he == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_robIdx_value : _GEN_3916; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [4:0] _GEN_5773 = 4'hf == io_enq_req_1_bits_lqIdx_value ? io_enq_req_1_bits_robIdx_value : _GEN_3917; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_6118 = 4'h0 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4398; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_6119 = 4'h1 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4399; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_6120 = 4'h2 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4400; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_6121 = 4'h3 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4401; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_6122 = 4'h4 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4402; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_6123 = 4'h5 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4403; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_6124 = 4'h6 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4404; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_6125 = 4'h7 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4405; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_6126 = 4'h8 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4406; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_6127 = 4'h9 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4407; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_6128 = 4'ha == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4408; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_6129 = 4'hb == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4409; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_6130 = 4'hc == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4410; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_6131 = 4'hd == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4411; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_6132 = 4'he == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4412; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_6133 = 4'hf == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4413; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_6134 = 4'h0 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4414; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_6135 = 4'h1 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4415; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_6136 = 4'h2 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4416; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_6137 = 4'h3 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4417; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_6138 = 4'h4 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4418; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_6139 = 4'h5 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4419; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_6140 = 4'h6 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4420; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_6141 = 4'h7 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4421; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_6142 = 4'h8 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4422; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_6143 = 4'h9 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4423; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_6144 = 4'ha == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4424; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_6145 = 4'hb == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4425; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_6146 = 4'hc == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4426; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_6147 = 4'hd == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4427; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_6148 = 4'he == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4428; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_6149 = 4'hf == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4429; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_6262 = 4'h0 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4542; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_6263 = 4'h1 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4543; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_6264 = 4'h2 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4544; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_6265 = 4'h3 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4545; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_6266 = 4'h4 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4546; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_6267 = 4'h5 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4547; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_6268 = 4'h6 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4548; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_6269 = 4'h7 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4549; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_6270 = 4'h8 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4550; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_6271 = 4'h9 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4551; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_6272 = 4'ha == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4552; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_6273 = 4'hb == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4553; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_6274 = 4'hc == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4554; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_6275 = 4'hd == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4555; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_6276 = 4'he == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4556; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_6277 = 4'hf == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4557; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_6310 = 4'h0 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4158; // @[LoadQueueFlag.scala 211:{24,24}]
  wire  _GEN_6311 = 4'h1 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4159; // @[LoadQueueFlag.scala 211:{24,24}]
  wire  _GEN_6312 = 4'h2 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4160; // @[LoadQueueFlag.scala 211:{24,24}]
  wire  _GEN_6313 = 4'h3 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4161; // @[LoadQueueFlag.scala 211:{24,24}]
  wire  _GEN_6314 = 4'h4 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4162; // @[LoadQueueFlag.scala 211:{24,24}]
  wire  _GEN_6315 = 4'h5 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4163; // @[LoadQueueFlag.scala 211:{24,24}]
  wire  _GEN_6316 = 4'h6 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4164; // @[LoadQueueFlag.scala 211:{24,24}]
  wire  _GEN_6317 = 4'h7 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4165; // @[LoadQueueFlag.scala 211:{24,24}]
  wire  _GEN_6318 = 4'h8 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4166; // @[LoadQueueFlag.scala 211:{24,24}]
  wire  _GEN_6319 = 4'h9 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4167; // @[LoadQueueFlag.scala 211:{24,24}]
  wire  _GEN_6320 = 4'ha == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4168; // @[LoadQueueFlag.scala 211:{24,24}]
  wire  _GEN_6321 = 4'hb == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4169; // @[LoadQueueFlag.scala 211:{24,24}]
  wire  _GEN_6322 = 4'hc == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4170; // @[LoadQueueFlag.scala 211:{24,24}]
  wire  _GEN_6323 = 4'hd == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4171; // @[LoadQueueFlag.scala 211:{24,24}]
  wire  _GEN_6324 = 4'he == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4172; // @[LoadQueueFlag.scala 211:{24,24}]
  wire  _GEN_6325 = 4'hf == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4173; // @[LoadQueueFlag.scala 211:{24,24}]
  wire  _GEN_6326 = 4'h0 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4174; // @[LoadQueueFlag.scala 212:{24,24}]
  wire  _GEN_6327 = 4'h1 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4175; // @[LoadQueueFlag.scala 212:{24,24}]
  wire  _GEN_6328 = 4'h2 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4176; // @[LoadQueueFlag.scala 212:{24,24}]
  wire  _GEN_6329 = 4'h3 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4177; // @[LoadQueueFlag.scala 212:{24,24}]
  wire  _GEN_6330 = 4'h4 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4178; // @[LoadQueueFlag.scala 212:{24,24}]
  wire  _GEN_6331 = 4'h5 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4179; // @[LoadQueueFlag.scala 212:{24,24}]
  wire  _GEN_6332 = 4'h6 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4180; // @[LoadQueueFlag.scala 212:{24,24}]
  wire  _GEN_6333 = 4'h7 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4181; // @[LoadQueueFlag.scala 212:{24,24}]
  wire  _GEN_6334 = 4'h8 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4182; // @[LoadQueueFlag.scala 212:{24,24}]
  wire  _GEN_6335 = 4'h9 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4183; // @[LoadQueueFlag.scala 212:{24,24}]
  wire  _GEN_6336 = 4'ha == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4184; // @[LoadQueueFlag.scala 212:{24,24}]
  wire  _GEN_6337 = 4'hb == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4185; // @[LoadQueueFlag.scala 212:{24,24}]
  wire  _GEN_6338 = 4'hc == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4186; // @[LoadQueueFlag.scala 212:{24,24}]
  wire  _GEN_6339 = 4'hd == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4187; // @[LoadQueueFlag.scala 212:{24,24}]
  wire  _GEN_6340 = 4'he == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4188; // @[LoadQueueFlag.scala 212:{24,24}]
  wire  _GEN_6341 = 4'hf == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4189; // @[LoadQueueFlag.scala 212:{24,24}]
  wire  _GEN_6342 = 4'h0 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4190; // @[LoadQueueFlag.scala 213:{22,22}]
  wire  _GEN_6343 = 4'h1 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4191; // @[LoadQueueFlag.scala 213:{22,22}]
  wire  _GEN_6344 = 4'h2 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4192; // @[LoadQueueFlag.scala 213:{22,22}]
  wire  _GEN_6345 = 4'h3 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4193; // @[LoadQueueFlag.scala 213:{22,22}]
  wire  _GEN_6346 = 4'h4 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4194; // @[LoadQueueFlag.scala 213:{22,22}]
  wire  _GEN_6347 = 4'h5 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4195; // @[LoadQueueFlag.scala 213:{22,22}]
  wire  _GEN_6348 = 4'h6 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4196; // @[LoadQueueFlag.scala 213:{22,22}]
  wire  _GEN_6349 = 4'h7 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4197; // @[LoadQueueFlag.scala 213:{22,22}]
  wire  _GEN_6350 = 4'h8 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4198; // @[LoadQueueFlag.scala 213:{22,22}]
  wire  _GEN_6351 = 4'h9 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4199; // @[LoadQueueFlag.scala 213:{22,22}]
  wire  _GEN_6352 = 4'ha == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4200; // @[LoadQueueFlag.scala 213:{22,22}]
  wire  _GEN_6353 = 4'hb == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4201; // @[LoadQueueFlag.scala 213:{22,22}]
  wire  _GEN_6354 = 4'hc == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4202; // @[LoadQueueFlag.scala 213:{22,22}]
  wire  _GEN_6355 = 4'hd == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4203; // @[LoadQueueFlag.scala 213:{22,22}]
  wire  _GEN_6356 = 4'he == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4204; // @[LoadQueueFlag.scala 213:{22,22}]
  wire  _GEN_6357 = 4'hf == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4205; // @[LoadQueueFlag.scala 213:{22,22}]
  wire  _GEN_6358 = 4'h0 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4206; // @[LoadQueueFlag.scala 214:{26,26}]
  wire  _GEN_6359 = 4'h1 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4207; // @[LoadQueueFlag.scala 214:{26,26}]
  wire  _GEN_6360 = 4'h2 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4208; // @[LoadQueueFlag.scala 214:{26,26}]
  wire  _GEN_6361 = 4'h3 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4209; // @[LoadQueueFlag.scala 214:{26,26}]
  wire  _GEN_6362 = 4'h4 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4210; // @[LoadQueueFlag.scala 214:{26,26}]
  wire  _GEN_6363 = 4'h5 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4211; // @[LoadQueueFlag.scala 214:{26,26}]
  wire  _GEN_6364 = 4'h6 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4212; // @[LoadQueueFlag.scala 214:{26,26}]
  wire  _GEN_6365 = 4'h7 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4213; // @[LoadQueueFlag.scala 214:{26,26}]
  wire  _GEN_6366 = 4'h8 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4214; // @[LoadQueueFlag.scala 214:{26,26}]
  wire  _GEN_6367 = 4'h9 == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4215; // @[LoadQueueFlag.scala 214:{26,26}]
  wire  _GEN_6368 = 4'ha == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4216; // @[LoadQueueFlag.scala 214:{26,26}]
  wire  _GEN_6369 = 4'hb == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4217; // @[LoadQueueFlag.scala 214:{26,26}]
  wire  _GEN_6370 = 4'hc == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4218; // @[LoadQueueFlag.scala 214:{26,26}]
  wire  _GEN_6371 = 4'hd == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4219; // @[LoadQueueFlag.scala 214:{26,26}]
  wire  _GEN_6372 = 4'he == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4220; // @[LoadQueueFlag.scala 214:{26,26}]
  wire  _GEN_6373 = 4'hf == io_enq_req_1_bits_lqIdx_value ? 1'h0 : _GEN_4221; // @[LoadQueueFlag.scala 214:{26,26}]
  wire  _GEN_6422 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_4270 : _GEN_2414; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6423 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_4271 : _GEN_2415; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6424 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_4272 : _GEN_2416; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6425 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_4273 : _GEN_2417; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6426 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_4274 : _GEN_2418; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6427 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_4275 : _GEN_2419; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6428 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_4276 : _GEN_2420; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6429 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_4277 : _GEN_2421; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6430 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_4278 : _GEN_2422; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6431 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_4279 : _GEN_2423; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6432 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_4280 : _GEN_2424; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6433 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_4281 : _GEN_2425; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6434 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_4282 : _GEN_2426; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6435 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_4283 : _GEN_2427; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6436 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_4284 : _GEN_2428; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6437 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_4285 : _GEN_2429; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6550 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6118 : _GEN_2542; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6551 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6119 : _GEN_2543; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6552 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6120 : _GEN_2544; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6553 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6121 : _GEN_2545; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6554 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6122 : _GEN_2546; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6555 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6123 : _GEN_2547; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6556 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6124 : _GEN_2548; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6557 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6125 : _GEN_2549; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6558 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6126 : _GEN_2550; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6559 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6127 : _GEN_2551; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6560 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6128 : _GEN_2552; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6561 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6129 : _GEN_2553; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6562 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6130 : _GEN_2554; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6563 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6131 : _GEN_2555; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6564 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6132 : _GEN_2556; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6565 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6133 : _GEN_2557; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6566 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6134 : _GEN_2558; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6567 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6135 : _GEN_2559; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6568 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6136 : _GEN_2560; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6569 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6137 : _GEN_2561; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6570 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6138 : _GEN_2562; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6571 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6139 : _GEN_2563; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6572 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6140 : _GEN_2564; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6573 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6141 : _GEN_2565; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6574 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6142 : _GEN_2566; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6575 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6143 : _GEN_2567; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6576 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6144 : _GEN_2568; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6577 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6145 : _GEN_2569; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6578 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6146 : _GEN_2570; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6579 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6147 : _GEN_2571; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6580 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6148 : _GEN_2572; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6581 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6149 : _GEN_2573; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6694 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6262 : _GEN_2686; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6695 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6263 : _GEN_2687; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6696 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6264 : _GEN_2688; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6697 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6265 : _GEN_2689; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6698 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6266 : _GEN_2690; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6699 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6267 : _GEN_2691; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6700 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6268 : _GEN_2692; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6701 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6269 : _GEN_2693; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6702 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6270 : _GEN_2694; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6703 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6271 : _GEN_2695; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6704 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6272 : _GEN_2696; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6705 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6273 : _GEN_2697; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6706 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6274 : _GEN_2698; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6707 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6275 : _GEN_2699; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6708 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6276 : _GEN_2700; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6709 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6277 : _GEN_2701; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6822 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_4670 : _GEN_2814; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6823 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_4671 : _GEN_2815; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6824 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_4672 : _GEN_2816; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6825 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_4673 : _GEN_2817; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6826 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_4674 : _GEN_2818; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6827 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_4675 : _GEN_2819; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6828 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_4676 : _GEN_2820; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6829 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_4677 : _GEN_2821; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6830 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_4678 : _GEN_2822; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6831 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_4679 : _GEN_2823; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6832 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_4680 : _GEN_2824; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6833 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_4681 : _GEN_2825; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6834 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_4682 : _GEN_2826; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6835 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_4683 : _GEN_2827; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6836 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_4684 : _GEN_2828; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6837 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_4685 : _GEN_2829; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6838 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_4686 : _GEN_2830; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6839 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_4687 : _GEN_2831; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6840 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_4688 : _GEN_2832; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6841 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_4689 : _GEN_2833; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6842 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_4690 : _GEN_2834; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6843 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_4691 : _GEN_2835; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6844 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_4692 : _GEN_2836; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6845 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_4693 : _GEN_2837; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6846 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_4694 : _GEN_2838; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6847 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_4695 : _GEN_2839; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6848 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_4696 : _GEN_2840; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6849 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_4697 : _GEN_2841; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6850 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_4698 : _GEN_2842; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6851 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_4699 : _GEN_2843; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6852 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_4700 : _GEN_2844; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6853 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_4701 : _GEN_2845; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6854 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_4702 : _GEN_2846; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6855 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_4703 : _GEN_2847; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6856 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_4704 : _GEN_2848; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6857 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_4705 : _GEN_2849; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6858 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_4706 : _GEN_2850; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6859 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_4707 : _GEN_2851; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6860 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_4708 : _GEN_2852; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6861 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_4709 : _GEN_2853; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6862 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_4710 : _GEN_2854; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6863 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_4711 : _GEN_2855; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6864 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_4712 : _GEN_2856; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6865 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_4713 : _GEN_2857; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6866 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_4714 : _GEN_2858; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6867 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_4715 : _GEN_2859; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6868 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_4716 : _GEN_2860; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6869 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_4717 : _GEN_2861; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6902 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_4750 : _GEN_2894; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6903 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_4751 : _GEN_2895; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6904 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_4752 : _GEN_2896; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6905 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_4753 : _GEN_2897; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6906 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_4754 : _GEN_2898; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6907 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_4755 : _GEN_2899; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6908 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_4756 : _GEN_2900; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6909 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_4757 : _GEN_2901; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6910 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_4758 : _GEN_2902; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6911 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_4759 : _GEN_2903; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6912 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_4760 : _GEN_2904; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6913 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_4761 : _GEN_2905; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6914 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_4762 : _GEN_2906; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6915 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_4763 : _GEN_2907; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6916 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_4764 : _GEN_2908; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_6917 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_4765 : _GEN_2909; // @[LoadQueueFlag.scala 204:43]
  wire [6:0] _GEN_7334 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5182 : _GEN_3326; // @[LoadQueueFlag.scala 204:43]
  wire [6:0] _GEN_7335 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5183 : _GEN_3327; // @[LoadQueueFlag.scala 204:43]
  wire [6:0] _GEN_7336 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5184 : _GEN_3328; // @[LoadQueueFlag.scala 204:43]
  wire [6:0] _GEN_7337 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5185 : _GEN_3329; // @[LoadQueueFlag.scala 204:43]
  wire [6:0] _GEN_7338 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5186 : _GEN_3330; // @[LoadQueueFlag.scala 204:43]
  wire [6:0] _GEN_7339 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5187 : _GEN_3331; // @[LoadQueueFlag.scala 204:43]
  wire [6:0] _GEN_7340 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5188 : _GEN_3332; // @[LoadQueueFlag.scala 204:43]
  wire [6:0] _GEN_7341 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5189 : _GEN_3333; // @[LoadQueueFlag.scala 204:43]
  wire [6:0] _GEN_7342 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5190 : _GEN_3334; // @[LoadQueueFlag.scala 204:43]
  wire [6:0] _GEN_7343 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5191 : _GEN_3335; // @[LoadQueueFlag.scala 204:43]
  wire [6:0] _GEN_7344 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5192 : _GEN_3336; // @[LoadQueueFlag.scala 204:43]
  wire [6:0] _GEN_7345 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5193 : _GEN_3337; // @[LoadQueueFlag.scala 204:43]
  wire [6:0] _GEN_7346 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5194 : _GEN_3338; // @[LoadQueueFlag.scala 204:43]
  wire [6:0] _GEN_7347 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5195 : _GEN_3339; // @[LoadQueueFlag.scala 204:43]
  wire [6:0] _GEN_7348 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5196 : _GEN_3340; // @[LoadQueueFlag.scala 204:43]
  wire [6:0] _GEN_7349 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5197 : _GEN_3341; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_7350 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5198 : _GEN_3342; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_7351 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5199 : _GEN_3343; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_7352 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5200 : _GEN_3344; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_7353 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5201 : _GEN_3345; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_7354 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5202 : _GEN_3346; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_7355 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5203 : _GEN_3347; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_7356 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5204 : _GEN_3348; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_7357 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5205 : _GEN_3349; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_7358 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5206 : _GEN_3350; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_7359 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5207 : _GEN_3351; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_7360 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5208 : _GEN_3352; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_7361 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5209 : _GEN_3353; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_7362 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5210 : _GEN_3354; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_7363 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5211 : _GEN_3355; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_7364 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5212 : _GEN_3356; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_7365 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5213 : _GEN_3357; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_7366 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5214 : _GEN_3358; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_7367 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5215 : _GEN_3359; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_7368 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5216 : _GEN_3360; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_7369 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5217 : _GEN_3361; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_7370 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5218 : _GEN_3362; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_7371 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5219 : _GEN_3363; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_7372 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5220 : _GEN_3364; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_7373 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5221 : _GEN_3365; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_7374 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5222 : _GEN_3366; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_7375 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5223 : _GEN_3367; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_7376 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5224 : _GEN_3368; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_7377 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5225 : _GEN_3369; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_7378 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5226 : _GEN_3370; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_7379 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5227 : _GEN_3371; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_7380 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5228 : _GEN_3372; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_7381 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5229 : _GEN_3373; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_7430 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5278 : _GEN_3422; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_7431 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5279 : _GEN_3423; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_7432 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5280 : _GEN_3424; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_7433 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5281 : _GEN_3425; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_7434 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5282 : _GEN_3426; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_7435 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5283 : _GEN_3427; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_7436 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5284 : _GEN_3428; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_7437 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5285 : _GEN_3429; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_7438 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5286 : _GEN_3430; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_7439 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5287 : _GEN_3431; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_7440 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5288 : _GEN_3432; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_7441 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5289 : _GEN_3433; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_7442 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5290 : _GEN_3434; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_7443 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5291 : _GEN_3435; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_7444 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5292 : _GEN_3436; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_7445 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5293 : _GEN_3437; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_7750 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5598 : _GEN_3742; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_7751 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5599 : _GEN_3743; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_7752 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5600 : _GEN_3744; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_7753 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5601 : _GEN_3745; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_7754 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5602 : _GEN_3746; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_7755 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5603 : _GEN_3747; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_7756 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5604 : _GEN_3748; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_7757 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5605 : _GEN_3749; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_7758 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5606 : _GEN_3750; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_7759 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5607 : _GEN_3751; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_7760 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5608 : _GEN_3752; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_7761 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5609 : _GEN_3753; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_7762 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5610 : _GEN_3754; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_7763 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5611 : _GEN_3755; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_7764 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5612 : _GEN_3756; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_7765 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5613 : _GEN_3757; // @[LoadQueueFlag.scala 204:43]
  wire [5:0] _GEN_7862 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5710 : _GEN_3854; // @[LoadQueueFlag.scala 204:43]
  wire [5:0] _GEN_7863 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5711 : _GEN_3855; // @[LoadQueueFlag.scala 204:43]
  wire [5:0] _GEN_7864 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5712 : _GEN_3856; // @[LoadQueueFlag.scala 204:43]
  wire [5:0] _GEN_7865 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5713 : _GEN_3857; // @[LoadQueueFlag.scala 204:43]
  wire [5:0] _GEN_7866 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5714 : _GEN_3858; // @[LoadQueueFlag.scala 204:43]
  wire [5:0] _GEN_7867 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5715 : _GEN_3859; // @[LoadQueueFlag.scala 204:43]
  wire [5:0] _GEN_7868 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5716 : _GEN_3860; // @[LoadQueueFlag.scala 204:43]
  wire [5:0] _GEN_7869 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5717 : _GEN_3861; // @[LoadQueueFlag.scala 204:43]
  wire [5:0] _GEN_7870 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5718 : _GEN_3862; // @[LoadQueueFlag.scala 204:43]
  wire [5:0] _GEN_7871 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5719 : _GEN_3863; // @[LoadQueueFlag.scala 204:43]
  wire [5:0] _GEN_7872 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5720 : _GEN_3864; // @[LoadQueueFlag.scala 204:43]
  wire [5:0] _GEN_7873 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5721 : _GEN_3865; // @[LoadQueueFlag.scala 204:43]
  wire [5:0] _GEN_7874 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5722 : _GEN_3866; // @[LoadQueueFlag.scala 204:43]
  wire [5:0] _GEN_7875 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5723 : _GEN_3867; // @[LoadQueueFlag.scala 204:43]
  wire [5:0] _GEN_7876 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5724 : _GEN_3868; // @[LoadQueueFlag.scala 204:43]
  wire [5:0] _GEN_7877 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5725 : _GEN_3869; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_7894 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5742 : _GEN_3886; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_7895 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5743 : _GEN_3887; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_7896 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5744 : _GEN_3888; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_7897 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5745 : _GEN_3889; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_7898 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5746 : _GEN_3890; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_7899 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5747 : _GEN_3891; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_7900 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5748 : _GEN_3892; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_7901 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5749 : _GEN_3893; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_7902 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5750 : _GEN_3894; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_7903 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5751 : _GEN_3895; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_7904 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5752 : _GEN_3896; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_7905 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5753 : _GEN_3897; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_7906 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5754 : _GEN_3898; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_7907 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5755 : _GEN_3899; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_7908 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5756 : _GEN_3900; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_7909 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5757 : _GEN_3901; // @[LoadQueueFlag.scala 204:43]
  wire [4:0] _GEN_7910 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5758 : _GEN_3902; // @[LoadQueueFlag.scala 204:43]
  wire [4:0] _GEN_7911 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5759 : _GEN_3903; // @[LoadQueueFlag.scala 204:43]
  wire [4:0] _GEN_7912 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5760 : _GEN_3904; // @[LoadQueueFlag.scala 204:43]
  wire [4:0] _GEN_7913 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5761 : _GEN_3905; // @[LoadQueueFlag.scala 204:43]
  wire [4:0] _GEN_7914 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5762 : _GEN_3906; // @[LoadQueueFlag.scala 204:43]
  wire [4:0] _GEN_7915 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5763 : _GEN_3907; // @[LoadQueueFlag.scala 204:43]
  wire [4:0] _GEN_7916 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5764 : _GEN_3908; // @[LoadQueueFlag.scala 204:43]
  wire [4:0] _GEN_7917 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5765 : _GEN_3909; // @[LoadQueueFlag.scala 204:43]
  wire [4:0] _GEN_7918 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5766 : _GEN_3910; // @[LoadQueueFlag.scala 204:43]
  wire [4:0] _GEN_7919 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5767 : _GEN_3911; // @[LoadQueueFlag.scala 204:43]
  wire [4:0] _GEN_7920 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5768 : _GEN_3912; // @[LoadQueueFlag.scala 204:43]
  wire [4:0] _GEN_7921 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5769 : _GEN_3913; // @[LoadQueueFlag.scala 204:43]
  wire [4:0] _GEN_7922 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5770 : _GEN_3914; // @[LoadQueueFlag.scala 204:43]
  wire [4:0] _GEN_7923 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5771 : _GEN_3915; // @[LoadQueueFlag.scala 204:43]
  wire [4:0] _GEN_7924 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5772 : _GEN_3916; // @[LoadQueueFlag.scala 204:43]
  wire [4:0] _GEN_7925 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_5773 : _GEN_3917; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_8166 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6310 : _GEN_4158; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_8167 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6311 : _GEN_4159; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_8168 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6312 : _GEN_4160; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_8169 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6313 : _GEN_4161; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_8170 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6314 : _GEN_4162; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_8171 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6315 : _GEN_4163; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_8172 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6316 : _GEN_4164; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_8173 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6317 : _GEN_4165; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_8174 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6318 : _GEN_4166; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_8175 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6319 : _GEN_4167; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_8176 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6320 : _GEN_4168; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_8177 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6321 : _GEN_4169; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_8178 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6322 : _GEN_4170; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_8179 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6323 : _GEN_4171; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_8180 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6324 : _GEN_4172; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_8181 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6325 : _GEN_4173; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_8182 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6326 : _GEN_4174; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_8183 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6327 : _GEN_4175; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_8184 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6328 : _GEN_4176; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_8185 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6329 : _GEN_4177; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_8186 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6330 : _GEN_4178; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_8187 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6331 : _GEN_4179; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_8188 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6332 : _GEN_4180; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_8189 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6333 : _GEN_4181; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_8190 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6334 : _GEN_4182; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_8191 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6335 : _GEN_4183; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_8192 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6336 : _GEN_4184; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_8193 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6337 : _GEN_4185; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_8194 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6338 : _GEN_4186; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_8195 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6339 : _GEN_4187; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_8196 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6340 : _GEN_4188; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_8197 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6341 : _GEN_4189; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_8198 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6342 : _GEN_4190; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_8199 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6343 : _GEN_4191; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_8200 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6344 : _GEN_4192; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_8201 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6345 : _GEN_4193; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_8202 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6346 : _GEN_4194; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_8203 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6347 : _GEN_4195; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_8204 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6348 : _GEN_4196; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_8205 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6349 : _GEN_4197; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_8206 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6350 : _GEN_4198; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_8207 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6351 : _GEN_4199; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_8208 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6352 : _GEN_4200; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_8209 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6353 : _GEN_4201; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_8210 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6354 : _GEN_4202; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_8211 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6355 : _GEN_4203; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_8212 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6356 : _GEN_4204; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_8213 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6357 : _GEN_4205; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_8214 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6358 : _GEN_4206; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_8215 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6359 : _GEN_4207; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_8216 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6360 : _GEN_4208; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_8217 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6361 : _GEN_4209; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_8218 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6362 : _GEN_4210; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_8219 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6363 : _GEN_4211; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_8220 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6364 : _GEN_4212; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_8221 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6365 : _GEN_4213; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_8222 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6366 : _GEN_4214; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_8223 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6367 : _GEN_4215; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_8224 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6368 : _GEN_4216; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_8225 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6369 : _GEN_4217; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_8226 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6370 : _GEN_4218; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_8227 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6371 : _GEN_4219; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_8228 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6372 : _GEN_4220; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_8229 = io_enq_req_1_valid & ~enqCancel_1 ? _GEN_6373 : _GEN_4221; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_8278 = 4'h0 == io_enq_req_2_bits_lqIdx_value | _GEN_6422; // @[LoadQueueFlag.scala 205:{24,24}]
  wire  _GEN_8279 = 4'h1 == io_enq_req_2_bits_lqIdx_value | _GEN_6423; // @[LoadQueueFlag.scala 205:{24,24}]
  wire  _GEN_8280 = 4'h2 == io_enq_req_2_bits_lqIdx_value | _GEN_6424; // @[LoadQueueFlag.scala 205:{24,24}]
  wire  _GEN_8281 = 4'h3 == io_enq_req_2_bits_lqIdx_value | _GEN_6425; // @[LoadQueueFlag.scala 205:{24,24}]
  wire  _GEN_8282 = 4'h4 == io_enq_req_2_bits_lqIdx_value | _GEN_6426; // @[LoadQueueFlag.scala 205:{24,24}]
  wire  _GEN_8283 = 4'h5 == io_enq_req_2_bits_lqIdx_value | _GEN_6427; // @[LoadQueueFlag.scala 205:{24,24}]
  wire  _GEN_8284 = 4'h6 == io_enq_req_2_bits_lqIdx_value | _GEN_6428; // @[LoadQueueFlag.scala 205:{24,24}]
  wire  _GEN_8285 = 4'h7 == io_enq_req_2_bits_lqIdx_value | _GEN_6429; // @[LoadQueueFlag.scala 205:{24,24}]
  wire  _GEN_8286 = 4'h8 == io_enq_req_2_bits_lqIdx_value | _GEN_6430; // @[LoadQueueFlag.scala 205:{24,24}]
  wire  _GEN_8287 = 4'h9 == io_enq_req_2_bits_lqIdx_value | _GEN_6431; // @[LoadQueueFlag.scala 205:{24,24}]
  wire  _GEN_8288 = 4'ha == io_enq_req_2_bits_lqIdx_value | _GEN_6432; // @[LoadQueueFlag.scala 205:{24,24}]
  wire  _GEN_8289 = 4'hb == io_enq_req_2_bits_lqIdx_value | _GEN_6433; // @[LoadQueueFlag.scala 205:{24,24}]
  wire  _GEN_8290 = 4'hc == io_enq_req_2_bits_lqIdx_value | _GEN_6434; // @[LoadQueueFlag.scala 205:{24,24}]
  wire  _GEN_8291 = 4'hd == io_enq_req_2_bits_lqIdx_value | _GEN_6435; // @[LoadQueueFlag.scala 205:{24,24}]
  wire  _GEN_8292 = 4'he == io_enq_req_2_bits_lqIdx_value | _GEN_6436; // @[LoadQueueFlag.scala 205:{24,24}]
  wire  _GEN_8293 = 4'hf == io_enq_req_2_bits_lqIdx_value | _GEN_6437; // @[LoadQueueFlag.scala 205:{24,24}]
  wire  _GEN_8406 = 4'h0 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6550; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8407 = 4'h1 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6551; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8408 = 4'h2 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6552; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8409 = 4'h3 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6553; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8410 = 4'h4 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6554; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8411 = 4'h5 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6555; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8412 = 4'h6 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6556; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8413 = 4'h7 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6557; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8414 = 4'h8 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6558; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8415 = 4'h9 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6559; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8416 = 4'ha == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6560; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8417 = 4'hb == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6561; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8418 = 4'hc == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6562; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8419 = 4'hd == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6563; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8420 = 4'he == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6564; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8421 = 4'hf == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6565; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8422 = 4'h0 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6566; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8423 = 4'h1 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6567; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8424 = 4'h2 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6568; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8425 = 4'h3 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6569; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8426 = 4'h4 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6570; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8427 = 4'h5 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6571; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8428 = 4'h6 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6572; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8429 = 4'h7 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6573; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8430 = 4'h8 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6574; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8431 = 4'h9 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6575; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8432 = 4'ha == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6576; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8433 = 4'hb == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6577; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8434 = 4'hc == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6578; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8435 = 4'hd == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6579; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8436 = 4'he == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6580; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8437 = 4'hf == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6581; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8550 = 4'h0 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6694; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8551 = 4'h1 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6695; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8552 = 4'h2 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6696; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8553 = 4'h3 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6697; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8554 = 4'h4 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6698; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8555 = 4'h5 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6699; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8556 = 4'h6 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6700; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8557 = 4'h7 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6701; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8558 = 4'h8 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6702; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8559 = 4'h9 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6703; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8560 = 4'ha == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6704; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8561 = 4'hb == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6705; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8562 = 4'hc == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6706; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8563 = 4'hd == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6707; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8564 = 4'he == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6708; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8565 = 4'hf == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6709; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8678 = 4'h0 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_cf_trigger_backendEn_1 : _GEN_6822; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8679 = 4'h1 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_cf_trigger_backendEn_1 : _GEN_6823; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8680 = 4'h2 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_cf_trigger_backendEn_1 : _GEN_6824; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8681 = 4'h3 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_cf_trigger_backendEn_1 : _GEN_6825; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8682 = 4'h4 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_cf_trigger_backendEn_1 : _GEN_6826; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8683 = 4'h5 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_cf_trigger_backendEn_1 : _GEN_6827; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8684 = 4'h6 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_cf_trigger_backendEn_1 : _GEN_6828; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8685 = 4'h7 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_cf_trigger_backendEn_1 : _GEN_6829; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8686 = 4'h8 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_cf_trigger_backendEn_1 : _GEN_6830; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8687 = 4'h9 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_cf_trigger_backendEn_1 : _GEN_6831; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8688 = 4'ha == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_cf_trigger_backendEn_1 : _GEN_6832; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8689 = 4'hb == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_cf_trigger_backendEn_1 : _GEN_6833; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8690 = 4'hc == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_cf_trigger_backendEn_1 : _GEN_6834; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8691 = 4'hd == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_cf_trigger_backendEn_1 : _GEN_6835; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8692 = 4'he == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_cf_trigger_backendEn_1 : _GEN_6836; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8693 = 4'hf == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_cf_trigger_backendEn_1 : _GEN_6837; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8694 = 4'h0 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6838; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8695 = 4'h1 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6839; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8696 = 4'h2 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6840; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8697 = 4'h3 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6841; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8698 = 4'h4 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6842; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8699 = 4'h5 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6843; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8700 = 4'h6 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6844; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8701 = 4'h7 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6845; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8702 = 4'h8 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6846; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8703 = 4'h9 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6847; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8704 = 4'ha == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6848; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8705 = 4'hb == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6849; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8706 = 4'hc == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6850; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8707 = 4'hd == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6851; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8708 = 4'he == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6852; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8709 = 4'hf == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6853; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8710 = 4'h0 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6854; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8711 = 4'h1 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6855; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8712 = 4'h2 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6856; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8713 = 4'h3 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6857; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8714 = 4'h4 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6858; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8715 = 4'h5 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6859; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8716 = 4'h6 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6860; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8717 = 4'h7 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6861; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8718 = 4'h8 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6862; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8719 = 4'h9 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6863; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8720 = 4'ha == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6864; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8721 = 4'hb == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6865; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8722 = 4'hc == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6866; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8723 = 4'hd == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6867; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8724 = 4'he == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6868; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8725 = 4'hf == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6869; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8758 = 4'h0 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6902; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8759 = 4'h1 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6903; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8760 = 4'h2 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6904; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8761 = 4'h3 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6905; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8762 = 4'h4 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6906; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8763 = 4'h5 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6907; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8764 = 4'h6 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6908; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8765 = 4'h7 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6909; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8766 = 4'h8 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6910; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8767 = 4'h9 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6911; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8768 = 4'ha == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6912; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8769 = 4'hb == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6913; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8770 = 4'hc == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6914; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8771 = 4'hd == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6915; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8772 = 4'he == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6916; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_8773 = 4'hf == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_6917; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [6:0] _GEN_9190 = 4'h0 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_ctrl_fuOpType : _GEN_7334; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [6:0] _GEN_9191 = 4'h1 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_ctrl_fuOpType : _GEN_7335; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [6:0] _GEN_9192 = 4'h2 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_ctrl_fuOpType : _GEN_7336; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [6:0] _GEN_9193 = 4'h3 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_ctrl_fuOpType : _GEN_7337; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [6:0] _GEN_9194 = 4'h4 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_ctrl_fuOpType : _GEN_7338; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [6:0] _GEN_9195 = 4'h5 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_ctrl_fuOpType : _GEN_7339; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [6:0] _GEN_9196 = 4'h6 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_ctrl_fuOpType : _GEN_7340; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [6:0] _GEN_9197 = 4'h7 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_ctrl_fuOpType : _GEN_7341; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [6:0] _GEN_9198 = 4'h8 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_ctrl_fuOpType : _GEN_7342; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [6:0] _GEN_9199 = 4'h9 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_ctrl_fuOpType : _GEN_7343; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [6:0] _GEN_9200 = 4'ha == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_ctrl_fuOpType : _GEN_7344; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [6:0] _GEN_9201 = 4'hb == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_ctrl_fuOpType : _GEN_7345; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [6:0] _GEN_9202 = 4'hc == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_ctrl_fuOpType : _GEN_7346; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [6:0] _GEN_9203 = 4'hd == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_ctrl_fuOpType : _GEN_7347; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [6:0] _GEN_9204 = 4'he == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_ctrl_fuOpType : _GEN_7348; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [6:0] _GEN_9205 = 4'hf == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_ctrl_fuOpType : _GEN_7349; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_9206 = 4'h0 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_ctrl_rfWen : _GEN_7350; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_9207 = 4'h1 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_ctrl_rfWen : _GEN_7351; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_9208 = 4'h2 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_ctrl_rfWen : _GEN_7352; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_9209 = 4'h3 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_ctrl_rfWen : _GEN_7353; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_9210 = 4'h4 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_ctrl_rfWen : _GEN_7354; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_9211 = 4'h5 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_ctrl_rfWen : _GEN_7355; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_9212 = 4'h6 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_ctrl_rfWen : _GEN_7356; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_9213 = 4'h7 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_ctrl_rfWen : _GEN_7357; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_9214 = 4'h8 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_ctrl_rfWen : _GEN_7358; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_9215 = 4'h9 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_ctrl_rfWen : _GEN_7359; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_9216 = 4'ha == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_ctrl_rfWen : _GEN_7360; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_9217 = 4'hb == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_ctrl_rfWen : _GEN_7361; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_9218 = 4'hc == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_ctrl_rfWen : _GEN_7362; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_9219 = 4'hd == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_ctrl_rfWen : _GEN_7363; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_9220 = 4'he == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_ctrl_rfWen : _GEN_7364; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_9221 = 4'hf == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_ctrl_rfWen : _GEN_7365; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_9222 = 4'h0 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_ctrl_fpWen : _GEN_7366; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_9223 = 4'h1 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_ctrl_fpWen : _GEN_7367; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_9224 = 4'h2 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_ctrl_fpWen : _GEN_7368; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_9225 = 4'h3 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_ctrl_fpWen : _GEN_7369; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_9226 = 4'h4 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_ctrl_fpWen : _GEN_7370; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_9227 = 4'h5 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_ctrl_fpWen : _GEN_7371; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_9228 = 4'h6 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_ctrl_fpWen : _GEN_7372; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_9229 = 4'h7 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_ctrl_fpWen : _GEN_7373; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_9230 = 4'h8 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_ctrl_fpWen : _GEN_7374; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_9231 = 4'h9 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_ctrl_fpWen : _GEN_7375; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_9232 = 4'ha == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_ctrl_fpWen : _GEN_7376; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_9233 = 4'hb == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_ctrl_fpWen : _GEN_7377; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_9234 = 4'hc == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_ctrl_fpWen : _GEN_7378; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_9235 = 4'hd == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_ctrl_fpWen : _GEN_7379; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_9236 = 4'he == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_ctrl_fpWen : _GEN_7380; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_9237 = 4'hf == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_ctrl_fpWen : _GEN_7381; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_9286 = 4'h0 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_ctrl_flushPipe : _GEN_7430; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_9287 = 4'h1 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_ctrl_flushPipe : _GEN_7431; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_9288 = 4'h2 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_ctrl_flushPipe : _GEN_7432; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_9289 = 4'h3 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_ctrl_flushPipe : _GEN_7433; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_9290 = 4'h4 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_ctrl_flushPipe : _GEN_7434; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_9291 = 4'h5 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_ctrl_flushPipe : _GEN_7435; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_9292 = 4'h6 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_ctrl_flushPipe : _GEN_7436; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_9293 = 4'h7 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_ctrl_flushPipe : _GEN_7437; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_9294 = 4'h8 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_ctrl_flushPipe : _GEN_7438; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_9295 = 4'h9 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_ctrl_flushPipe : _GEN_7439; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_9296 = 4'ha == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_ctrl_flushPipe : _GEN_7440; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_9297 = 4'hb == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_ctrl_flushPipe : _GEN_7441; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_9298 = 4'hc == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_ctrl_flushPipe : _GEN_7442; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_9299 = 4'hd == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_ctrl_flushPipe : _GEN_7443; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_9300 = 4'he == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_ctrl_flushPipe : _GEN_7444; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_9301 = 4'hf == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_ctrl_flushPipe : _GEN_7445; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_9606 = 4'h0 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_ctrl_replayInst : _GEN_7750; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_9607 = 4'h1 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_ctrl_replayInst : _GEN_7751; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_9608 = 4'h2 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_ctrl_replayInst : _GEN_7752; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_9609 = 4'h3 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_ctrl_replayInst : _GEN_7753; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_9610 = 4'h4 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_ctrl_replayInst : _GEN_7754; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_9611 = 4'h5 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_ctrl_replayInst : _GEN_7755; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_9612 = 4'h6 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_ctrl_replayInst : _GEN_7756; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_9613 = 4'h7 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_ctrl_replayInst : _GEN_7757; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_9614 = 4'h8 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_ctrl_replayInst : _GEN_7758; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_9615 = 4'h9 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_ctrl_replayInst : _GEN_7759; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_9616 = 4'ha == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_ctrl_replayInst : _GEN_7760; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_9617 = 4'hb == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_ctrl_replayInst : _GEN_7761; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_9618 = 4'hc == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_ctrl_replayInst : _GEN_7762; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_9619 = 4'hd == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_ctrl_replayInst : _GEN_7763; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_9620 = 4'he == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_ctrl_replayInst : _GEN_7764; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_9621 = 4'hf == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_ctrl_replayInst : _GEN_7765; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [5:0] _GEN_9718 = 4'h0 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_pdest : _GEN_7862; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [5:0] _GEN_9719 = 4'h1 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_pdest : _GEN_7863; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [5:0] _GEN_9720 = 4'h2 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_pdest : _GEN_7864; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [5:0] _GEN_9721 = 4'h3 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_pdest : _GEN_7865; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [5:0] _GEN_9722 = 4'h4 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_pdest : _GEN_7866; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [5:0] _GEN_9723 = 4'h5 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_pdest : _GEN_7867; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [5:0] _GEN_9724 = 4'h6 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_pdest : _GEN_7868; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [5:0] _GEN_9725 = 4'h7 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_pdest : _GEN_7869; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [5:0] _GEN_9726 = 4'h8 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_pdest : _GEN_7870; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [5:0] _GEN_9727 = 4'h9 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_pdest : _GEN_7871; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [5:0] _GEN_9728 = 4'ha == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_pdest : _GEN_7872; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [5:0] _GEN_9729 = 4'hb == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_pdest : _GEN_7873; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [5:0] _GEN_9730 = 4'hc == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_pdest : _GEN_7874; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [5:0] _GEN_9731 = 4'hd == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_pdest : _GEN_7875; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [5:0] _GEN_9732 = 4'he == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_pdest : _GEN_7876; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [5:0] _GEN_9733 = 4'hf == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_pdest : _GEN_7877; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_9750 = 4'h0 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_robIdx_flag : _GEN_7894; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_9751 = 4'h1 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_robIdx_flag : _GEN_7895; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_9752 = 4'h2 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_robIdx_flag : _GEN_7896; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_9753 = 4'h3 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_robIdx_flag : _GEN_7897; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_9754 = 4'h4 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_robIdx_flag : _GEN_7898; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_9755 = 4'h5 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_robIdx_flag : _GEN_7899; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_9756 = 4'h6 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_robIdx_flag : _GEN_7900; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_9757 = 4'h7 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_robIdx_flag : _GEN_7901; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_9758 = 4'h8 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_robIdx_flag : _GEN_7902; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_9759 = 4'h9 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_robIdx_flag : _GEN_7903; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_9760 = 4'ha == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_robIdx_flag : _GEN_7904; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_9761 = 4'hb == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_robIdx_flag : _GEN_7905; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_9762 = 4'hc == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_robIdx_flag : _GEN_7906; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_9763 = 4'hd == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_robIdx_flag : _GEN_7907; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_9764 = 4'he == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_robIdx_flag : _GEN_7908; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_9765 = 4'hf == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_robIdx_flag : _GEN_7909; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [4:0] _GEN_9766 = 4'h0 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_robIdx_value : _GEN_7910; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [4:0] _GEN_9767 = 4'h1 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_robIdx_value : _GEN_7911; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [4:0] _GEN_9768 = 4'h2 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_robIdx_value : _GEN_7912; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [4:0] _GEN_9769 = 4'h3 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_robIdx_value : _GEN_7913; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [4:0] _GEN_9770 = 4'h4 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_robIdx_value : _GEN_7914; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [4:0] _GEN_9771 = 4'h5 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_robIdx_value : _GEN_7915; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [4:0] _GEN_9772 = 4'h6 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_robIdx_value : _GEN_7916; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [4:0] _GEN_9773 = 4'h7 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_robIdx_value : _GEN_7917; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [4:0] _GEN_9774 = 4'h8 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_robIdx_value : _GEN_7918; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [4:0] _GEN_9775 = 4'h9 == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_robIdx_value : _GEN_7919; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [4:0] _GEN_9776 = 4'ha == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_robIdx_value : _GEN_7920; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [4:0] _GEN_9777 = 4'hb == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_robIdx_value : _GEN_7921; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [4:0] _GEN_9778 = 4'hc == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_robIdx_value : _GEN_7922; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [4:0] _GEN_9779 = 4'hd == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_robIdx_value : _GEN_7923; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [4:0] _GEN_9780 = 4'he == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_robIdx_value : _GEN_7924; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [4:0] _GEN_9781 = 4'hf == io_enq_req_2_bits_lqIdx_value ? io_enq_req_2_bits_robIdx_value : _GEN_7925; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_10126 = 4'h0 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8406; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_10127 = 4'h1 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8407; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_10128 = 4'h2 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8408; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_10129 = 4'h3 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8409; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_10130 = 4'h4 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8410; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_10131 = 4'h5 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8411; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_10132 = 4'h6 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8412; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_10133 = 4'h7 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8413; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_10134 = 4'h8 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8414; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_10135 = 4'h9 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8415; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_10136 = 4'ha == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8416; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_10137 = 4'hb == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8417; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_10138 = 4'hc == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8418; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_10139 = 4'hd == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8419; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_10140 = 4'he == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8420; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_10141 = 4'hf == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8421; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_10142 = 4'h0 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8422; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_10143 = 4'h1 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8423; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_10144 = 4'h2 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8424; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_10145 = 4'h3 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8425; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_10146 = 4'h4 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8426; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_10147 = 4'h5 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8427; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_10148 = 4'h6 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8428; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_10149 = 4'h7 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8429; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_10150 = 4'h8 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8430; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_10151 = 4'h9 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8431; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_10152 = 4'ha == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8432; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_10153 = 4'hb == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8433; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_10154 = 4'hc == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8434; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_10155 = 4'hd == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8435; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_10156 = 4'he == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8436; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_10157 = 4'hf == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8437; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_10270 = 4'h0 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8550; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_10271 = 4'h1 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8551; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_10272 = 4'h2 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8552; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_10273 = 4'h3 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8553; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_10274 = 4'h4 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8554; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_10275 = 4'h5 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8555; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_10276 = 4'h6 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8556; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_10277 = 4'h7 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8557; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_10278 = 4'h8 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8558; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_10279 = 4'h9 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8559; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_10280 = 4'ha == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8560; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_10281 = 4'hb == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8561; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_10282 = 4'hc == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8562; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_10283 = 4'hd == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8563; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_10284 = 4'he == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8564; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_10285 = 4'hf == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8565; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_10318 = 4'h0 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8166; // @[LoadQueueFlag.scala 211:{24,24}]
  wire  _GEN_10319 = 4'h1 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8167; // @[LoadQueueFlag.scala 211:{24,24}]
  wire  _GEN_10320 = 4'h2 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8168; // @[LoadQueueFlag.scala 211:{24,24}]
  wire  _GEN_10321 = 4'h3 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8169; // @[LoadQueueFlag.scala 211:{24,24}]
  wire  _GEN_10322 = 4'h4 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8170; // @[LoadQueueFlag.scala 211:{24,24}]
  wire  _GEN_10323 = 4'h5 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8171; // @[LoadQueueFlag.scala 211:{24,24}]
  wire  _GEN_10324 = 4'h6 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8172; // @[LoadQueueFlag.scala 211:{24,24}]
  wire  _GEN_10325 = 4'h7 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8173; // @[LoadQueueFlag.scala 211:{24,24}]
  wire  _GEN_10326 = 4'h8 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8174; // @[LoadQueueFlag.scala 211:{24,24}]
  wire  _GEN_10327 = 4'h9 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8175; // @[LoadQueueFlag.scala 211:{24,24}]
  wire  _GEN_10328 = 4'ha == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8176; // @[LoadQueueFlag.scala 211:{24,24}]
  wire  _GEN_10329 = 4'hb == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8177; // @[LoadQueueFlag.scala 211:{24,24}]
  wire  _GEN_10330 = 4'hc == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8178; // @[LoadQueueFlag.scala 211:{24,24}]
  wire  _GEN_10331 = 4'hd == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8179; // @[LoadQueueFlag.scala 211:{24,24}]
  wire  _GEN_10332 = 4'he == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8180; // @[LoadQueueFlag.scala 211:{24,24}]
  wire  _GEN_10333 = 4'hf == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8181; // @[LoadQueueFlag.scala 211:{24,24}]
  wire  _GEN_10334 = 4'h0 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8182; // @[LoadQueueFlag.scala 212:{24,24}]
  wire  _GEN_10335 = 4'h1 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8183; // @[LoadQueueFlag.scala 212:{24,24}]
  wire  _GEN_10336 = 4'h2 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8184; // @[LoadQueueFlag.scala 212:{24,24}]
  wire  _GEN_10337 = 4'h3 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8185; // @[LoadQueueFlag.scala 212:{24,24}]
  wire  _GEN_10338 = 4'h4 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8186; // @[LoadQueueFlag.scala 212:{24,24}]
  wire  _GEN_10339 = 4'h5 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8187; // @[LoadQueueFlag.scala 212:{24,24}]
  wire  _GEN_10340 = 4'h6 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8188; // @[LoadQueueFlag.scala 212:{24,24}]
  wire  _GEN_10341 = 4'h7 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8189; // @[LoadQueueFlag.scala 212:{24,24}]
  wire  _GEN_10342 = 4'h8 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8190; // @[LoadQueueFlag.scala 212:{24,24}]
  wire  _GEN_10343 = 4'h9 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8191; // @[LoadQueueFlag.scala 212:{24,24}]
  wire  _GEN_10344 = 4'ha == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8192; // @[LoadQueueFlag.scala 212:{24,24}]
  wire  _GEN_10345 = 4'hb == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8193; // @[LoadQueueFlag.scala 212:{24,24}]
  wire  _GEN_10346 = 4'hc == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8194; // @[LoadQueueFlag.scala 212:{24,24}]
  wire  _GEN_10347 = 4'hd == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8195; // @[LoadQueueFlag.scala 212:{24,24}]
  wire  _GEN_10348 = 4'he == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8196; // @[LoadQueueFlag.scala 212:{24,24}]
  wire  _GEN_10349 = 4'hf == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8197; // @[LoadQueueFlag.scala 212:{24,24}]
  wire  _GEN_10350 = 4'h0 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8198; // @[LoadQueueFlag.scala 213:{22,22}]
  wire  _GEN_10351 = 4'h1 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8199; // @[LoadQueueFlag.scala 213:{22,22}]
  wire  _GEN_10352 = 4'h2 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8200; // @[LoadQueueFlag.scala 213:{22,22}]
  wire  _GEN_10353 = 4'h3 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8201; // @[LoadQueueFlag.scala 213:{22,22}]
  wire  _GEN_10354 = 4'h4 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8202; // @[LoadQueueFlag.scala 213:{22,22}]
  wire  _GEN_10355 = 4'h5 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8203; // @[LoadQueueFlag.scala 213:{22,22}]
  wire  _GEN_10356 = 4'h6 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8204; // @[LoadQueueFlag.scala 213:{22,22}]
  wire  _GEN_10357 = 4'h7 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8205; // @[LoadQueueFlag.scala 213:{22,22}]
  wire  _GEN_10358 = 4'h8 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8206; // @[LoadQueueFlag.scala 213:{22,22}]
  wire  _GEN_10359 = 4'h9 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8207; // @[LoadQueueFlag.scala 213:{22,22}]
  wire  _GEN_10360 = 4'ha == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8208; // @[LoadQueueFlag.scala 213:{22,22}]
  wire  _GEN_10361 = 4'hb == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8209; // @[LoadQueueFlag.scala 213:{22,22}]
  wire  _GEN_10362 = 4'hc == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8210; // @[LoadQueueFlag.scala 213:{22,22}]
  wire  _GEN_10363 = 4'hd == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8211; // @[LoadQueueFlag.scala 213:{22,22}]
  wire  _GEN_10364 = 4'he == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8212; // @[LoadQueueFlag.scala 213:{22,22}]
  wire  _GEN_10365 = 4'hf == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8213; // @[LoadQueueFlag.scala 213:{22,22}]
  wire  _GEN_10366 = 4'h0 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8214; // @[LoadQueueFlag.scala 214:{26,26}]
  wire  _GEN_10367 = 4'h1 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8215; // @[LoadQueueFlag.scala 214:{26,26}]
  wire  _GEN_10368 = 4'h2 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8216; // @[LoadQueueFlag.scala 214:{26,26}]
  wire  _GEN_10369 = 4'h3 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8217; // @[LoadQueueFlag.scala 214:{26,26}]
  wire  _GEN_10370 = 4'h4 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8218; // @[LoadQueueFlag.scala 214:{26,26}]
  wire  _GEN_10371 = 4'h5 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8219; // @[LoadQueueFlag.scala 214:{26,26}]
  wire  _GEN_10372 = 4'h6 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8220; // @[LoadQueueFlag.scala 214:{26,26}]
  wire  _GEN_10373 = 4'h7 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8221; // @[LoadQueueFlag.scala 214:{26,26}]
  wire  _GEN_10374 = 4'h8 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8222; // @[LoadQueueFlag.scala 214:{26,26}]
  wire  _GEN_10375 = 4'h9 == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8223; // @[LoadQueueFlag.scala 214:{26,26}]
  wire  _GEN_10376 = 4'ha == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8224; // @[LoadQueueFlag.scala 214:{26,26}]
  wire  _GEN_10377 = 4'hb == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8225; // @[LoadQueueFlag.scala 214:{26,26}]
  wire  _GEN_10378 = 4'hc == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8226; // @[LoadQueueFlag.scala 214:{26,26}]
  wire  _GEN_10379 = 4'hd == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8227; // @[LoadQueueFlag.scala 214:{26,26}]
  wire  _GEN_10380 = 4'he == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8228; // @[LoadQueueFlag.scala 214:{26,26}]
  wire  _GEN_10381 = 4'hf == io_enq_req_2_bits_lqIdx_value ? 1'h0 : _GEN_8229; // @[LoadQueueFlag.scala 214:{26,26}]
  wire  _GEN_10430 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_8278 : _GEN_6422; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10431 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_8279 : _GEN_6423; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10432 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_8280 : _GEN_6424; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10433 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_8281 : _GEN_6425; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10434 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_8282 : _GEN_6426; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10435 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_8283 : _GEN_6427; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10436 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_8284 : _GEN_6428; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10437 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_8285 : _GEN_6429; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10438 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_8286 : _GEN_6430; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10439 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_8287 : _GEN_6431; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10440 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_8288 : _GEN_6432; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10441 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_8289 : _GEN_6433; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10442 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_8290 : _GEN_6434; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10443 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_8291 : _GEN_6435; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10444 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_8292 : _GEN_6436; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10445 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_8293 : _GEN_6437; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10558 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10126 : _GEN_6550; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10559 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10127 : _GEN_6551; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10560 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10128 : _GEN_6552; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10561 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10129 : _GEN_6553; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10562 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10130 : _GEN_6554; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10563 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10131 : _GEN_6555; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10564 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10132 : _GEN_6556; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10565 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10133 : _GEN_6557; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10566 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10134 : _GEN_6558; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10567 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10135 : _GEN_6559; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10568 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10136 : _GEN_6560; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10569 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10137 : _GEN_6561; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10570 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10138 : _GEN_6562; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10571 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10139 : _GEN_6563; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10572 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10140 : _GEN_6564; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10573 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10141 : _GEN_6565; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10574 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10142 : _GEN_6566; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10575 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10143 : _GEN_6567; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10576 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10144 : _GEN_6568; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10577 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10145 : _GEN_6569; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10578 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10146 : _GEN_6570; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10579 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10147 : _GEN_6571; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10580 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10148 : _GEN_6572; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10581 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10149 : _GEN_6573; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10582 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10150 : _GEN_6574; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10583 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10151 : _GEN_6575; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10584 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10152 : _GEN_6576; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10585 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10153 : _GEN_6577; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10586 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10154 : _GEN_6578; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10587 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10155 : _GEN_6579; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10588 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10156 : _GEN_6580; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10589 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10157 : _GEN_6581; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10702 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10270 : _GEN_6694; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10703 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10271 : _GEN_6695; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10704 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10272 : _GEN_6696; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10705 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10273 : _GEN_6697; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10706 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10274 : _GEN_6698; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10707 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10275 : _GEN_6699; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10708 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10276 : _GEN_6700; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10709 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10277 : _GEN_6701; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10710 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10278 : _GEN_6702; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10711 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10279 : _GEN_6703; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10712 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10280 : _GEN_6704; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10713 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10281 : _GEN_6705; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10714 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10282 : _GEN_6706; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10715 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10283 : _GEN_6707; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10716 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10284 : _GEN_6708; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10717 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10285 : _GEN_6709; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10830 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_8678 : _GEN_6822; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10831 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_8679 : _GEN_6823; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10832 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_8680 : _GEN_6824; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10833 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_8681 : _GEN_6825; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10834 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_8682 : _GEN_6826; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10835 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_8683 : _GEN_6827; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10836 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_8684 : _GEN_6828; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10837 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_8685 : _GEN_6829; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10838 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_8686 : _GEN_6830; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10839 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_8687 : _GEN_6831; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10840 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_8688 : _GEN_6832; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10841 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_8689 : _GEN_6833; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10842 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_8690 : _GEN_6834; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10843 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_8691 : _GEN_6835; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10844 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_8692 : _GEN_6836; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10845 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_8693 : _GEN_6837; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10846 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_8694 : _GEN_6838; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10847 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_8695 : _GEN_6839; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10848 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_8696 : _GEN_6840; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10849 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_8697 : _GEN_6841; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10850 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_8698 : _GEN_6842; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10851 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_8699 : _GEN_6843; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10852 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_8700 : _GEN_6844; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10853 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_8701 : _GEN_6845; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10854 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_8702 : _GEN_6846; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10855 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_8703 : _GEN_6847; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10856 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_8704 : _GEN_6848; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10857 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_8705 : _GEN_6849; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10858 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_8706 : _GEN_6850; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10859 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_8707 : _GEN_6851; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10860 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_8708 : _GEN_6852; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10861 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_8709 : _GEN_6853; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10862 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_8710 : _GEN_6854; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10863 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_8711 : _GEN_6855; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10864 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_8712 : _GEN_6856; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10865 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_8713 : _GEN_6857; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10866 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_8714 : _GEN_6858; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10867 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_8715 : _GEN_6859; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10868 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_8716 : _GEN_6860; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10869 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_8717 : _GEN_6861; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10870 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_8718 : _GEN_6862; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10871 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_8719 : _GEN_6863; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10872 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_8720 : _GEN_6864; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10873 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_8721 : _GEN_6865; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10874 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_8722 : _GEN_6866; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10875 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_8723 : _GEN_6867; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10876 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_8724 : _GEN_6868; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10877 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_8725 : _GEN_6869; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10910 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_8758 : _GEN_6902; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10911 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_8759 : _GEN_6903; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10912 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_8760 : _GEN_6904; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10913 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_8761 : _GEN_6905; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10914 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_8762 : _GEN_6906; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10915 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_8763 : _GEN_6907; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10916 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_8764 : _GEN_6908; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10917 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_8765 : _GEN_6909; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10918 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_8766 : _GEN_6910; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10919 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_8767 : _GEN_6911; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10920 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_8768 : _GEN_6912; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10921 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_8769 : _GEN_6913; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10922 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_8770 : _GEN_6914; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10923 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_8771 : _GEN_6915; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10924 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_8772 : _GEN_6916; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_10925 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_8773 : _GEN_6917; // @[LoadQueueFlag.scala 204:43]
  wire [6:0] _GEN_11342 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9190 : _GEN_7334; // @[LoadQueueFlag.scala 204:43]
  wire [6:0] _GEN_11343 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9191 : _GEN_7335; // @[LoadQueueFlag.scala 204:43]
  wire [6:0] _GEN_11344 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9192 : _GEN_7336; // @[LoadQueueFlag.scala 204:43]
  wire [6:0] _GEN_11345 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9193 : _GEN_7337; // @[LoadQueueFlag.scala 204:43]
  wire [6:0] _GEN_11346 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9194 : _GEN_7338; // @[LoadQueueFlag.scala 204:43]
  wire [6:0] _GEN_11347 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9195 : _GEN_7339; // @[LoadQueueFlag.scala 204:43]
  wire [6:0] _GEN_11348 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9196 : _GEN_7340; // @[LoadQueueFlag.scala 204:43]
  wire [6:0] _GEN_11349 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9197 : _GEN_7341; // @[LoadQueueFlag.scala 204:43]
  wire [6:0] _GEN_11350 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9198 : _GEN_7342; // @[LoadQueueFlag.scala 204:43]
  wire [6:0] _GEN_11351 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9199 : _GEN_7343; // @[LoadQueueFlag.scala 204:43]
  wire [6:0] _GEN_11352 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9200 : _GEN_7344; // @[LoadQueueFlag.scala 204:43]
  wire [6:0] _GEN_11353 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9201 : _GEN_7345; // @[LoadQueueFlag.scala 204:43]
  wire [6:0] _GEN_11354 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9202 : _GEN_7346; // @[LoadQueueFlag.scala 204:43]
  wire [6:0] _GEN_11355 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9203 : _GEN_7347; // @[LoadQueueFlag.scala 204:43]
  wire [6:0] _GEN_11356 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9204 : _GEN_7348; // @[LoadQueueFlag.scala 204:43]
  wire [6:0] _GEN_11357 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9205 : _GEN_7349; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_11358 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9206 : _GEN_7350; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_11359 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9207 : _GEN_7351; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_11360 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9208 : _GEN_7352; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_11361 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9209 : _GEN_7353; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_11362 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9210 : _GEN_7354; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_11363 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9211 : _GEN_7355; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_11364 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9212 : _GEN_7356; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_11365 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9213 : _GEN_7357; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_11366 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9214 : _GEN_7358; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_11367 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9215 : _GEN_7359; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_11368 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9216 : _GEN_7360; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_11369 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9217 : _GEN_7361; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_11370 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9218 : _GEN_7362; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_11371 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9219 : _GEN_7363; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_11372 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9220 : _GEN_7364; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_11373 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9221 : _GEN_7365; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_11374 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9222 : _GEN_7366; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_11375 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9223 : _GEN_7367; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_11376 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9224 : _GEN_7368; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_11377 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9225 : _GEN_7369; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_11378 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9226 : _GEN_7370; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_11379 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9227 : _GEN_7371; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_11380 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9228 : _GEN_7372; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_11381 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9229 : _GEN_7373; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_11382 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9230 : _GEN_7374; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_11383 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9231 : _GEN_7375; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_11384 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9232 : _GEN_7376; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_11385 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9233 : _GEN_7377; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_11386 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9234 : _GEN_7378; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_11387 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9235 : _GEN_7379; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_11388 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9236 : _GEN_7380; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_11389 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9237 : _GEN_7381; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_11438 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9286 : _GEN_7430; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_11439 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9287 : _GEN_7431; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_11440 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9288 : _GEN_7432; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_11441 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9289 : _GEN_7433; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_11442 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9290 : _GEN_7434; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_11443 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9291 : _GEN_7435; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_11444 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9292 : _GEN_7436; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_11445 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9293 : _GEN_7437; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_11446 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9294 : _GEN_7438; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_11447 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9295 : _GEN_7439; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_11448 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9296 : _GEN_7440; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_11449 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9297 : _GEN_7441; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_11450 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9298 : _GEN_7442; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_11451 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9299 : _GEN_7443; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_11452 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9300 : _GEN_7444; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_11453 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9301 : _GEN_7445; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_11758 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9606 : _GEN_7750; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_11759 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9607 : _GEN_7751; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_11760 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9608 : _GEN_7752; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_11761 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9609 : _GEN_7753; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_11762 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9610 : _GEN_7754; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_11763 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9611 : _GEN_7755; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_11764 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9612 : _GEN_7756; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_11765 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9613 : _GEN_7757; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_11766 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9614 : _GEN_7758; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_11767 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9615 : _GEN_7759; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_11768 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9616 : _GEN_7760; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_11769 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9617 : _GEN_7761; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_11770 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9618 : _GEN_7762; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_11771 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9619 : _GEN_7763; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_11772 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9620 : _GEN_7764; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_11773 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9621 : _GEN_7765; // @[LoadQueueFlag.scala 204:43]
  wire [5:0] _GEN_11870 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9718 : _GEN_7862; // @[LoadQueueFlag.scala 204:43]
  wire [5:0] _GEN_11871 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9719 : _GEN_7863; // @[LoadQueueFlag.scala 204:43]
  wire [5:0] _GEN_11872 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9720 : _GEN_7864; // @[LoadQueueFlag.scala 204:43]
  wire [5:0] _GEN_11873 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9721 : _GEN_7865; // @[LoadQueueFlag.scala 204:43]
  wire [5:0] _GEN_11874 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9722 : _GEN_7866; // @[LoadQueueFlag.scala 204:43]
  wire [5:0] _GEN_11875 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9723 : _GEN_7867; // @[LoadQueueFlag.scala 204:43]
  wire [5:0] _GEN_11876 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9724 : _GEN_7868; // @[LoadQueueFlag.scala 204:43]
  wire [5:0] _GEN_11877 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9725 : _GEN_7869; // @[LoadQueueFlag.scala 204:43]
  wire [5:0] _GEN_11878 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9726 : _GEN_7870; // @[LoadQueueFlag.scala 204:43]
  wire [5:0] _GEN_11879 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9727 : _GEN_7871; // @[LoadQueueFlag.scala 204:43]
  wire [5:0] _GEN_11880 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9728 : _GEN_7872; // @[LoadQueueFlag.scala 204:43]
  wire [5:0] _GEN_11881 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9729 : _GEN_7873; // @[LoadQueueFlag.scala 204:43]
  wire [5:0] _GEN_11882 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9730 : _GEN_7874; // @[LoadQueueFlag.scala 204:43]
  wire [5:0] _GEN_11883 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9731 : _GEN_7875; // @[LoadQueueFlag.scala 204:43]
  wire [5:0] _GEN_11884 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9732 : _GEN_7876; // @[LoadQueueFlag.scala 204:43]
  wire [5:0] _GEN_11885 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9733 : _GEN_7877; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_11902 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9750 : _GEN_7894; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_11903 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9751 : _GEN_7895; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_11904 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9752 : _GEN_7896; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_11905 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9753 : _GEN_7897; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_11906 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9754 : _GEN_7898; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_11907 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9755 : _GEN_7899; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_11908 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9756 : _GEN_7900; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_11909 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9757 : _GEN_7901; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_11910 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9758 : _GEN_7902; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_11911 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9759 : _GEN_7903; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_11912 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9760 : _GEN_7904; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_11913 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9761 : _GEN_7905; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_11914 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9762 : _GEN_7906; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_11915 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9763 : _GEN_7907; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_11916 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9764 : _GEN_7908; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_11917 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9765 : _GEN_7909; // @[LoadQueueFlag.scala 204:43]
  wire [4:0] _GEN_11918 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9766 : _GEN_7910; // @[LoadQueueFlag.scala 204:43]
  wire [4:0] _GEN_11919 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9767 : _GEN_7911; // @[LoadQueueFlag.scala 204:43]
  wire [4:0] _GEN_11920 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9768 : _GEN_7912; // @[LoadQueueFlag.scala 204:43]
  wire [4:0] _GEN_11921 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9769 : _GEN_7913; // @[LoadQueueFlag.scala 204:43]
  wire [4:0] _GEN_11922 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9770 : _GEN_7914; // @[LoadQueueFlag.scala 204:43]
  wire [4:0] _GEN_11923 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9771 : _GEN_7915; // @[LoadQueueFlag.scala 204:43]
  wire [4:0] _GEN_11924 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9772 : _GEN_7916; // @[LoadQueueFlag.scala 204:43]
  wire [4:0] _GEN_11925 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9773 : _GEN_7917; // @[LoadQueueFlag.scala 204:43]
  wire [4:0] _GEN_11926 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9774 : _GEN_7918; // @[LoadQueueFlag.scala 204:43]
  wire [4:0] _GEN_11927 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9775 : _GEN_7919; // @[LoadQueueFlag.scala 204:43]
  wire [4:0] _GEN_11928 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9776 : _GEN_7920; // @[LoadQueueFlag.scala 204:43]
  wire [4:0] _GEN_11929 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9777 : _GEN_7921; // @[LoadQueueFlag.scala 204:43]
  wire [4:0] _GEN_11930 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9778 : _GEN_7922; // @[LoadQueueFlag.scala 204:43]
  wire [4:0] _GEN_11931 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9779 : _GEN_7923; // @[LoadQueueFlag.scala 204:43]
  wire [4:0] _GEN_11932 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9780 : _GEN_7924; // @[LoadQueueFlag.scala 204:43]
  wire [4:0] _GEN_11933 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_9781 : _GEN_7925; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_12174 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10318 : _GEN_8166; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_12175 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10319 : _GEN_8167; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_12176 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10320 : _GEN_8168; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_12177 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10321 : _GEN_8169; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_12178 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10322 : _GEN_8170; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_12179 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10323 : _GEN_8171; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_12180 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10324 : _GEN_8172; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_12181 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10325 : _GEN_8173; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_12182 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10326 : _GEN_8174; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_12183 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10327 : _GEN_8175; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_12184 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10328 : _GEN_8176; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_12185 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10329 : _GEN_8177; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_12186 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10330 : _GEN_8178; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_12187 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10331 : _GEN_8179; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_12188 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10332 : _GEN_8180; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_12189 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10333 : _GEN_8181; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_12190 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10334 : _GEN_8182; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_12191 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10335 : _GEN_8183; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_12192 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10336 : _GEN_8184; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_12193 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10337 : _GEN_8185; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_12194 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10338 : _GEN_8186; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_12195 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10339 : _GEN_8187; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_12196 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10340 : _GEN_8188; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_12197 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10341 : _GEN_8189; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_12198 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10342 : _GEN_8190; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_12199 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10343 : _GEN_8191; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_12200 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10344 : _GEN_8192; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_12201 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10345 : _GEN_8193; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_12202 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10346 : _GEN_8194; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_12203 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10347 : _GEN_8195; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_12204 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10348 : _GEN_8196; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_12205 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10349 : _GEN_8197; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_12206 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10350 : _GEN_8198; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_12207 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10351 : _GEN_8199; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_12208 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10352 : _GEN_8200; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_12209 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10353 : _GEN_8201; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_12210 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10354 : _GEN_8202; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_12211 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10355 : _GEN_8203; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_12212 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10356 : _GEN_8204; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_12213 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10357 : _GEN_8205; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_12214 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10358 : _GEN_8206; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_12215 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10359 : _GEN_8207; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_12216 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10360 : _GEN_8208; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_12217 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10361 : _GEN_8209; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_12218 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10362 : _GEN_8210; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_12219 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10363 : _GEN_8211; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_12220 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10364 : _GEN_8212; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_12221 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10365 : _GEN_8213; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_12222 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10366 : _GEN_8214; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_12223 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10367 : _GEN_8215; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_12224 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10368 : _GEN_8216; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_12225 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10369 : _GEN_8217; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_12226 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10370 : _GEN_8218; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_12227 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10371 : _GEN_8219; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_12228 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10372 : _GEN_8220; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_12229 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10373 : _GEN_8221; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_12230 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10374 : _GEN_8222; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_12231 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10375 : _GEN_8223; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_12232 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10376 : _GEN_8224; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_12233 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10377 : _GEN_8225; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_12234 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10378 : _GEN_8226; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_12235 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10379 : _GEN_8227; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_12236 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10380 : _GEN_8228; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_12237 = io_enq_req_2_valid & ~enqCancel_2 ? _GEN_10381 : _GEN_8229; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_12286 = 4'h0 == io_enq_req_3_bits_lqIdx_value | _GEN_10430; // @[LoadQueueFlag.scala 205:{24,24}]
  wire  _GEN_12287 = 4'h1 == io_enq_req_3_bits_lqIdx_value | _GEN_10431; // @[LoadQueueFlag.scala 205:{24,24}]
  wire  _GEN_12288 = 4'h2 == io_enq_req_3_bits_lqIdx_value | _GEN_10432; // @[LoadQueueFlag.scala 205:{24,24}]
  wire  _GEN_12289 = 4'h3 == io_enq_req_3_bits_lqIdx_value | _GEN_10433; // @[LoadQueueFlag.scala 205:{24,24}]
  wire  _GEN_12290 = 4'h4 == io_enq_req_3_bits_lqIdx_value | _GEN_10434; // @[LoadQueueFlag.scala 205:{24,24}]
  wire  _GEN_12291 = 4'h5 == io_enq_req_3_bits_lqIdx_value | _GEN_10435; // @[LoadQueueFlag.scala 205:{24,24}]
  wire  _GEN_12292 = 4'h6 == io_enq_req_3_bits_lqIdx_value | _GEN_10436; // @[LoadQueueFlag.scala 205:{24,24}]
  wire  _GEN_12293 = 4'h7 == io_enq_req_3_bits_lqIdx_value | _GEN_10437; // @[LoadQueueFlag.scala 205:{24,24}]
  wire  _GEN_12294 = 4'h8 == io_enq_req_3_bits_lqIdx_value | _GEN_10438; // @[LoadQueueFlag.scala 205:{24,24}]
  wire  _GEN_12295 = 4'h9 == io_enq_req_3_bits_lqIdx_value | _GEN_10439; // @[LoadQueueFlag.scala 205:{24,24}]
  wire  _GEN_12296 = 4'ha == io_enq_req_3_bits_lqIdx_value | _GEN_10440; // @[LoadQueueFlag.scala 205:{24,24}]
  wire  _GEN_12297 = 4'hb == io_enq_req_3_bits_lqIdx_value | _GEN_10441; // @[LoadQueueFlag.scala 205:{24,24}]
  wire  _GEN_12298 = 4'hc == io_enq_req_3_bits_lqIdx_value | _GEN_10442; // @[LoadQueueFlag.scala 205:{24,24}]
  wire  _GEN_12299 = 4'hd == io_enq_req_3_bits_lqIdx_value | _GEN_10443; // @[LoadQueueFlag.scala 205:{24,24}]
  wire  _GEN_12300 = 4'he == io_enq_req_3_bits_lqIdx_value | _GEN_10444; // @[LoadQueueFlag.scala 205:{24,24}]
  wire  _GEN_12301 = 4'hf == io_enq_req_3_bits_lqIdx_value | _GEN_10445; // @[LoadQueueFlag.scala 205:{24,24}]
  wire  _GEN_12414 = 4'h0 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10558; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12415 = 4'h1 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10559; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12416 = 4'h2 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10560; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12417 = 4'h3 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10561; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12418 = 4'h4 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10562; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12419 = 4'h5 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10563; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12420 = 4'h6 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10564; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12421 = 4'h7 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10565; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12422 = 4'h8 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10566; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12423 = 4'h9 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10567; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12424 = 4'ha == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10568; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12425 = 4'hb == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10569; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12426 = 4'hc == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10570; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12427 = 4'hd == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10571; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12428 = 4'he == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10572; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12429 = 4'hf == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10573; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12430 = 4'h0 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10574; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12431 = 4'h1 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10575; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12432 = 4'h2 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10576; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12433 = 4'h3 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10577; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12434 = 4'h4 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10578; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12435 = 4'h5 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10579; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12436 = 4'h6 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10580; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12437 = 4'h7 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10581; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12438 = 4'h8 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10582; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12439 = 4'h9 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10583; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12440 = 4'ha == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10584; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12441 = 4'hb == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10585; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12442 = 4'hc == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10586; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12443 = 4'hd == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10587; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12444 = 4'he == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10588; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12445 = 4'hf == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10589; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12558 = 4'h0 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10702; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12559 = 4'h1 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10703; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12560 = 4'h2 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10704; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12561 = 4'h3 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10705; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12562 = 4'h4 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10706; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12563 = 4'h5 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10707; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12564 = 4'h6 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10708; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12565 = 4'h7 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10709; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12566 = 4'h8 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10710; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12567 = 4'h9 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10711; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12568 = 4'ha == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10712; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12569 = 4'hb == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10713; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12570 = 4'hc == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10714; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12571 = 4'hd == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10715; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12572 = 4'he == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10716; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12573 = 4'hf == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10717; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12686 = 4'h0 == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_cf_trigger_backendEn_1 : _GEN_10830; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12687 = 4'h1 == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_cf_trigger_backendEn_1 : _GEN_10831; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12688 = 4'h2 == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_cf_trigger_backendEn_1 : _GEN_10832; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12689 = 4'h3 == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_cf_trigger_backendEn_1 : _GEN_10833; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12690 = 4'h4 == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_cf_trigger_backendEn_1 : _GEN_10834; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12691 = 4'h5 == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_cf_trigger_backendEn_1 : _GEN_10835; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12692 = 4'h6 == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_cf_trigger_backendEn_1 : _GEN_10836; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12693 = 4'h7 == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_cf_trigger_backendEn_1 : _GEN_10837; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12694 = 4'h8 == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_cf_trigger_backendEn_1 : _GEN_10838; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12695 = 4'h9 == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_cf_trigger_backendEn_1 : _GEN_10839; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12696 = 4'ha == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_cf_trigger_backendEn_1 : _GEN_10840; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12697 = 4'hb == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_cf_trigger_backendEn_1 : _GEN_10841; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12698 = 4'hc == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_cf_trigger_backendEn_1 : _GEN_10842; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12699 = 4'hd == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_cf_trigger_backendEn_1 : _GEN_10843; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12700 = 4'he == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_cf_trigger_backendEn_1 : _GEN_10844; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12701 = 4'hf == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_cf_trigger_backendEn_1 : _GEN_10845; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12702 = 4'h0 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10846; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12703 = 4'h1 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10847; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12704 = 4'h2 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10848; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12705 = 4'h3 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10849; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12706 = 4'h4 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10850; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12707 = 4'h5 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10851; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12708 = 4'h6 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10852; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12709 = 4'h7 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10853; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12710 = 4'h8 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10854; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12711 = 4'h9 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10855; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12712 = 4'ha == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10856; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12713 = 4'hb == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10857; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12714 = 4'hc == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10858; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12715 = 4'hd == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10859; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12716 = 4'he == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10860; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12717 = 4'hf == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10861; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12718 = 4'h0 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10862; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12719 = 4'h1 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10863; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12720 = 4'h2 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10864; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12721 = 4'h3 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10865; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12722 = 4'h4 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10866; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12723 = 4'h5 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10867; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12724 = 4'h6 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10868; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12725 = 4'h7 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10869; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12726 = 4'h8 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10870; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12727 = 4'h9 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10871; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12728 = 4'ha == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10872; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12729 = 4'hb == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10873; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12730 = 4'hc == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10874; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12731 = 4'hd == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10875; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12732 = 4'he == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10876; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12733 = 4'hf == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10877; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12766 = 4'h0 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10910; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12767 = 4'h1 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10911; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12768 = 4'h2 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10912; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12769 = 4'h3 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10913; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12770 = 4'h4 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10914; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12771 = 4'h5 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10915; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12772 = 4'h6 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10916; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12773 = 4'h7 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10917; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12774 = 4'h8 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10918; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12775 = 4'h9 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10919; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12776 = 4'ha == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10920; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12777 = 4'hb == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10921; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12778 = 4'hc == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10922; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12779 = 4'hd == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10923; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12780 = 4'he == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10924; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_12781 = 4'hf == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_10925; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [6:0] _GEN_13198 = 4'h0 == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_ctrl_fuOpType : _GEN_11342; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [6:0] _GEN_13199 = 4'h1 == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_ctrl_fuOpType : _GEN_11343; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [6:0] _GEN_13200 = 4'h2 == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_ctrl_fuOpType : _GEN_11344; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [6:0] _GEN_13201 = 4'h3 == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_ctrl_fuOpType : _GEN_11345; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [6:0] _GEN_13202 = 4'h4 == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_ctrl_fuOpType : _GEN_11346; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [6:0] _GEN_13203 = 4'h5 == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_ctrl_fuOpType : _GEN_11347; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [6:0] _GEN_13204 = 4'h6 == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_ctrl_fuOpType : _GEN_11348; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [6:0] _GEN_13205 = 4'h7 == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_ctrl_fuOpType : _GEN_11349; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [6:0] _GEN_13206 = 4'h8 == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_ctrl_fuOpType : _GEN_11350; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [6:0] _GEN_13207 = 4'h9 == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_ctrl_fuOpType : _GEN_11351; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [6:0] _GEN_13208 = 4'ha == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_ctrl_fuOpType : _GEN_11352; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [6:0] _GEN_13209 = 4'hb == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_ctrl_fuOpType : _GEN_11353; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [6:0] _GEN_13210 = 4'hc == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_ctrl_fuOpType : _GEN_11354; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [6:0] _GEN_13211 = 4'hd == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_ctrl_fuOpType : _GEN_11355; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [6:0] _GEN_13212 = 4'he == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_ctrl_fuOpType : _GEN_11356; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [6:0] _GEN_13213 = 4'hf == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_ctrl_fuOpType : _GEN_11357; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_13214 = 4'h0 == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_ctrl_rfWen : _GEN_11358; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_13215 = 4'h1 == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_ctrl_rfWen : _GEN_11359; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_13216 = 4'h2 == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_ctrl_rfWen : _GEN_11360; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_13217 = 4'h3 == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_ctrl_rfWen : _GEN_11361; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_13218 = 4'h4 == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_ctrl_rfWen : _GEN_11362; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_13219 = 4'h5 == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_ctrl_rfWen : _GEN_11363; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_13220 = 4'h6 == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_ctrl_rfWen : _GEN_11364; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_13221 = 4'h7 == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_ctrl_rfWen : _GEN_11365; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_13222 = 4'h8 == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_ctrl_rfWen : _GEN_11366; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_13223 = 4'h9 == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_ctrl_rfWen : _GEN_11367; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_13224 = 4'ha == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_ctrl_rfWen : _GEN_11368; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_13225 = 4'hb == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_ctrl_rfWen : _GEN_11369; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_13226 = 4'hc == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_ctrl_rfWen : _GEN_11370; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_13227 = 4'hd == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_ctrl_rfWen : _GEN_11371; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_13228 = 4'he == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_ctrl_rfWen : _GEN_11372; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_13229 = 4'hf == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_ctrl_rfWen : _GEN_11373; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_13230 = 4'h0 == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_ctrl_fpWen : _GEN_11374; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_13231 = 4'h1 == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_ctrl_fpWen : _GEN_11375; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_13232 = 4'h2 == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_ctrl_fpWen : _GEN_11376; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_13233 = 4'h3 == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_ctrl_fpWen : _GEN_11377; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_13234 = 4'h4 == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_ctrl_fpWen : _GEN_11378; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_13235 = 4'h5 == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_ctrl_fpWen : _GEN_11379; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_13236 = 4'h6 == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_ctrl_fpWen : _GEN_11380; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_13237 = 4'h7 == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_ctrl_fpWen : _GEN_11381; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_13238 = 4'h8 == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_ctrl_fpWen : _GEN_11382; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_13239 = 4'h9 == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_ctrl_fpWen : _GEN_11383; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_13240 = 4'ha == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_ctrl_fpWen : _GEN_11384; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_13241 = 4'hb == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_ctrl_fpWen : _GEN_11385; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_13242 = 4'hc == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_ctrl_fpWen : _GEN_11386; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_13243 = 4'hd == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_ctrl_fpWen : _GEN_11387; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_13244 = 4'he == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_ctrl_fpWen : _GEN_11388; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_13245 = 4'hf == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_ctrl_fpWen : _GEN_11389; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_13294 = 4'h0 == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_ctrl_flushPipe : _GEN_11438; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_13295 = 4'h1 == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_ctrl_flushPipe : _GEN_11439; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_13296 = 4'h2 == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_ctrl_flushPipe : _GEN_11440; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_13297 = 4'h3 == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_ctrl_flushPipe : _GEN_11441; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_13298 = 4'h4 == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_ctrl_flushPipe : _GEN_11442; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_13299 = 4'h5 == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_ctrl_flushPipe : _GEN_11443; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_13300 = 4'h6 == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_ctrl_flushPipe : _GEN_11444; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_13301 = 4'h7 == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_ctrl_flushPipe : _GEN_11445; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_13302 = 4'h8 == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_ctrl_flushPipe : _GEN_11446; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_13303 = 4'h9 == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_ctrl_flushPipe : _GEN_11447; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_13304 = 4'ha == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_ctrl_flushPipe : _GEN_11448; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_13305 = 4'hb == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_ctrl_flushPipe : _GEN_11449; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_13306 = 4'hc == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_ctrl_flushPipe : _GEN_11450; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_13307 = 4'hd == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_ctrl_flushPipe : _GEN_11451; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_13308 = 4'he == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_ctrl_flushPipe : _GEN_11452; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_13309 = 4'hf == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_ctrl_flushPipe : _GEN_11453; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_13614 = 4'h0 == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_ctrl_replayInst : _GEN_11758; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_13615 = 4'h1 == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_ctrl_replayInst : _GEN_11759; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_13616 = 4'h2 == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_ctrl_replayInst : _GEN_11760; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_13617 = 4'h3 == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_ctrl_replayInst : _GEN_11761; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_13618 = 4'h4 == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_ctrl_replayInst : _GEN_11762; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_13619 = 4'h5 == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_ctrl_replayInst : _GEN_11763; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_13620 = 4'h6 == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_ctrl_replayInst : _GEN_11764; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_13621 = 4'h7 == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_ctrl_replayInst : _GEN_11765; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_13622 = 4'h8 == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_ctrl_replayInst : _GEN_11766; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_13623 = 4'h9 == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_ctrl_replayInst : _GEN_11767; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_13624 = 4'ha == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_ctrl_replayInst : _GEN_11768; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_13625 = 4'hb == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_ctrl_replayInst : _GEN_11769; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_13626 = 4'hc == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_ctrl_replayInst : _GEN_11770; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_13627 = 4'hd == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_ctrl_replayInst : _GEN_11771; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_13628 = 4'he == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_ctrl_replayInst : _GEN_11772; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_13629 = 4'hf == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_ctrl_replayInst : _GEN_11773; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [5:0] _GEN_13726 = 4'h0 == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_pdest : _GEN_11870; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [5:0] _GEN_13727 = 4'h1 == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_pdest : _GEN_11871; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [5:0] _GEN_13728 = 4'h2 == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_pdest : _GEN_11872; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [5:0] _GEN_13729 = 4'h3 == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_pdest : _GEN_11873; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [5:0] _GEN_13730 = 4'h4 == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_pdest : _GEN_11874; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [5:0] _GEN_13731 = 4'h5 == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_pdest : _GEN_11875; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [5:0] _GEN_13732 = 4'h6 == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_pdest : _GEN_11876; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [5:0] _GEN_13733 = 4'h7 == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_pdest : _GEN_11877; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [5:0] _GEN_13734 = 4'h8 == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_pdest : _GEN_11878; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [5:0] _GEN_13735 = 4'h9 == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_pdest : _GEN_11879; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [5:0] _GEN_13736 = 4'ha == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_pdest : _GEN_11880; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [5:0] _GEN_13737 = 4'hb == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_pdest : _GEN_11881; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [5:0] _GEN_13738 = 4'hc == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_pdest : _GEN_11882; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [5:0] _GEN_13739 = 4'hd == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_pdest : _GEN_11883; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [5:0] _GEN_13740 = 4'he == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_pdest : _GEN_11884; // @[LoadQueueFlag.scala 206:{18,18}]
  wire [5:0] _GEN_13741 = 4'hf == io_enq_req_3_bits_lqIdx_value ? io_enq_req_3_bits_pdest : _GEN_11885; // @[LoadQueueFlag.scala 206:{18,18}]
  wire  _GEN_14134 = 4'h0 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12414; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_14135 = 4'h1 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12415; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_14136 = 4'h2 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12416; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_14137 = 4'h3 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12417; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_14138 = 4'h4 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12418; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_14139 = 4'h5 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12419; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_14140 = 4'h6 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12420; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_14141 = 4'h7 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12421; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_14142 = 4'h8 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12422; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_14143 = 4'h9 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12423; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_14144 = 4'ha == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12424; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_14145 = 4'hb == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12425; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_14146 = 4'hc == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12426; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_14147 = 4'hd == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12427; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_14148 = 4'he == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12428; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_14149 = 4'hf == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12429; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_14150 = 4'h0 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12430; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_14151 = 4'h1 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12431; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_14152 = 4'h2 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12432; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_14153 = 4'h3 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12433; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_14154 = 4'h4 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12434; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_14155 = 4'h5 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12435; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_14156 = 4'h6 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12436; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_14157 = 4'h7 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12437; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_14158 = 4'h8 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12438; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_14159 = 4'h9 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12439; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_14160 = 4'ha == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12440; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_14161 = 4'hb == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12441; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_14162 = 4'hc == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12442; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_14163 = 4'hd == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12443; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_14164 = 4'he == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12444; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_14165 = 4'hf == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12445; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_14278 = 4'h0 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12558; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_14279 = 4'h1 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12559; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_14280 = 4'h2 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12560; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_14281 = 4'h3 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12561; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_14282 = 4'h4 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12562; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_14283 = 4'h5 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12563; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_14284 = 4'h6 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12564; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_14285 = 4'h7 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12565; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_14286 = 4'h8 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12566; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_14287 = 4'h9 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12567; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_14288 = 4'ha == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12568; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_14289 = 4'hb == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12569; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_14290 = 4'hc == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12570; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_14291 = 4'hd == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12571; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_14292 = 4'he == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12572; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_14293 = 4'hf == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12573; // @[LoadQueueFlag.scala 208:{34,34}]
  wire  _GEN_14326 = 4'h0 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12174; // @[LoadQueueFlag.scala 211:{24,24}]
  wire  _GEN_14327 = 4'h1 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12175; // @[LoadQueueFlag.scala 211:{24,24}]
  wire  _GEN_14328 = 4'h2 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12176; // @[LoadQueueFlag.scala 211:{24,24}]
  wire  _GEN_14329 = 4'h3 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12177; // @[LoadQueueFlag.scala 211:{24,24}]
  wire  _GEN_14330 = 4'h4 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12178; // @[LoadQueueFlag.scala 211:{24,24}]
  wire  _GEN_14331 = 4'h5 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12179; // @[LoadQueueFlag.scala 211:{24,24}]
  wire  _GEN_14332 = 4'h6 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12180; // @[LoadQueueFlag.scala 211:{24,24}]
  wire  _GEN_14333 = 4'h7 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12181; // @[LoadQueueFlag.scala 211:{24,24}]
  wire  _GEN_14334 = 4'h8 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12182; // @[LoadQueueFlag.scala 211:{24,24}]
  wire  _GEN_14335 = 4'h9 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12183; // @[LoadQueueFlag.scala 211:{24,24}]
  wire  _GEN_14336 = 4'ha == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12184; // @[LoadQueueFlag.scala 211:{24,24}]
  wire  _GEN_14337 = 4'hb == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12185; // @[LoadQueueFlag.scala 211:{24,24}]
  wire  _GEN_14338 = 4'hc == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12186; // @[LoadQueueFlag.scala 211:{24,24}]
  wire  _GEN_14339 = 4'hd == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12187; // @[LoadQueueFlag.scala 211:{24,24}]
  wire  _GEN_14340 = 4'he == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12188; // @[LoadQueueFlag.scala 211:{24,24}]
  wire  _GEN_14341 = 4'hf == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12189; // @[LoadQueueFlag.scala 211:{24,24}]
  wire  _GEN_14342 = 4'h0 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12190; // @[LoadQueueFlag.scala 212:{24,24}]
  wire  _GEN_14343 = 4'h1 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12191; // @[LoadQueueFlag.scala 212:{24,24}]
  wire  _GEN_14344 = 4'h2 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12192; // @[LoadQueueFlag.scala 212:{24,24}]
  wire  _GEN_14345 = 4'h3 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12193; // @[LoadQueueFlag.scala 212:{24,24}]
  wire  _GEN_14346 = 4'h4 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12194; // @[LoadQueueFlag.scala 212:{24,24}]
  wire  _GEN_14347 = 4'h5 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12195; // @[LoadQueueFlag.scala 212:{24,24}]
  wire  _GEN_14348 = 4'h6 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12196; // @[LoadQueueFlag.scala 212:{24,24}]
  wire  _GEN_14349 = 4'h7 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12197; // @[LoadQueueFlag.scala 212:{24,24}]
  wire  _GEN_14350 = 4'h8 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12198; // @[LoadQueueFlag.scala 212:{24,24}]
  wire  _GEN_14351 = 4'h9 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12199; // @[LoadQueueFlag.scala 212:{24,24}]
  wire  _GEN_14352 = 4'ha == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12200; // @[LoadQueueFlag.scala 212:{24,24}]
  wire  _GEN_14353 = 4'hb == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12201; // @[LoadQueueFlag.scala 212:{24,24}]
  wire  _GEN_14354 = 4'hc == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12202; // @[LoadQueueFlag.scala 212:{24,24}]
  wire  _GEN_14355 = 4'hd == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12203; // @[LoadQueueFlag.scala 212:{24,24}]
  wire  _GEN_14356 = 4'he == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12204; // @[LoadQueueFlag.scala 212:{24,24}]
  wire  _GEN_14357 = 4'hf == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12205; // @[LoadQueueFlag.scala 212:{24,24}]
  wire  _GEN_14358 = 4'h0 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12206; // @[LoadQueueFlag.scala 213:{22,22}]
  wire  _GEN_14359 = 4'h1 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12207; // @[LoadQueueFlag.scala 213:{22,22}]
  wire  _GEN_14360 = 4'h2 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12208; // @[LoadQueueFlag.scala 213:{22,22}]
  wire  _GEN_14361 = 4'h3 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12209; // @[LoadQueueFlag.scala 213:{22,22}]
  wire  _GEN_14362 = 4'h4 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12210; // @[LoadQueueFlag.scala 213:{22,22}]
  wire  _GEN_14363 = 4'h5 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12211; // @[LoadQueueFlag.scala 213:{22,22}]
  wire  _GEN_14364 = 4'h6 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12212; // @[LoadQueueFlag.scala 213:{22,22}]
  wire  _GEN_14365 = 4'h7 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12213; // @[LoadQueueFlag.scala 213:{22,22}]
  wire  _GEN_14366 = 4'h8 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12214; // @[LoadQueueFlag.scala 213:{22,22}]
  wire  _GEN_14367 = 4'h9 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12215; // @[LoadQueueFlag.scala 213:{22,22}]
  wire  _GEN_14368 = 4'ha == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12216; // @[LoadQueueFlag.scala 213:{22,22}]
  wire  _GEN_14369 = 4'hb == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12217; // @[LoadQueueFlag.scala 213:{22,22}]
  wire  _GEN_14370 = 4'hc == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12218; // @[LoadQueueFlag.scala 213:{22,22}]
  wire  _GEN_14371 = 4'hd == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12219; // @[LoadQueueFlag.scala 213:{22,22}]
  wire  _GEN_14372 = 4'he == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12220; // @[LoadQueueFlag.scala 213:{22,22}]
  wire  _GEN_14373 = 4'hf == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12221; // @[LoadQueueFlag.scala 213:{22,22}]
  wire  _GEN_14374 = 4'h0 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12222; // @[LoadQueueFlag.scala 214:{26,26}]
  wire  _GEN_14375 = 4'h1 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12223; // @[LoadQueueFlag.scala 214:{26,26}]
  wire  _GEN_14376 = 4'h2 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12224; // @[LoadQueueFlag.scala 214:{26,26}]
  wire  _GEN_14377 = 4'h3 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12225; // @[LoadQueueFlag.scala 214:{26,26}]
  wire  _GEN_14378 = 4'h4 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12226; // @[LoadQueueFlag.scala 214:{26,26}]
  wire  _GEN_14379 = 4'h5 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12227; // @[LoadQueueFlag.scala 214:{26,26}]
  wire  _GEN_14380 = 4'h6 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12228; // @[LoadQueueFlag.scala 214:{26,26}]
  wire  _GEN_14381 = 4'h7 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12229; // @[LoadQueueFlag.scala 214:{26,26}]
  wire  _GEN_14382 = 4'h8 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12230; // @[LoadQueueFlag.scala 214:{26,26}]
  wire  _GEN_14383 = 4'h9 == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12231; // @[LoadQueueFlag.scala 214:{26,26}]
  wire  _GEN_14384 = 4'ha == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12232; // @[LoadQueueFlag.scala 214:{26,26}]
  wire  _GEN_14385 = 4'hb == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12233; // @[LoadQueueFlag.scala 214:{26,26}]
  wire  _GEN_14386 = 4'hc == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12234; // @[LoadQueueFlag.scala 214:{26,26}]
  wire  _GEN_14387 = 4'hd == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12235; // @[LoadQueueFlag.scala 214:{26,26}]
  wire  _GEN_14388 = 4'he == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12236; // @[LoadQueueFlag.scala 214:{26,26}]
  wire  _GEN_14389 = 4'hf == io_enq_req_3_bits_lqIdx_value ? 1'h0 : _GEN_12237; // @[LoadQueueFlag.scala 214:{26,26}]
  wire  _GEN_14438 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_12286 : _GEN_10430; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14439 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_12287 : _GEN_10431; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14440 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_12288 : _GEN_10432; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14441 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_12289 : _GEN_10433; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14442 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_12290 : _GEN_10434; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14443 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_12291 : _GEN_10435; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14444 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_12292 : _GEN_10436; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14445 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_12293 : _GEN_10437; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14446 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_12294 : _GEN_10438; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14447 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_12295 : _GEN_10439; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14448 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_12296 : _GEN_10440; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14449 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_12297 : _GEN_10441; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14450 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_12298 : _GEN_10442; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14451 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_12299 : _GEN_10443; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14452 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_12300 : _GEN_10444; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14453 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_12301 : _GEN_10445; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14566 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14134 : _GEN_10558; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14567 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14135 : _GEN_10559; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14568 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14136 : _GEN_10560; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14569 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14137 : _GEN_10561; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14570 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14138 : _GEN_10562; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14571 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14139 : _GEN_10563; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14572 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14140 : _GEN_10564; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14573 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14141 : _GEN_10565; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14574 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14142 : _GEN_10566; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14575 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14143 : _GEN_10567; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14576 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14144 : _GEN_10568; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14577 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14145 : _GEN_10569; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14578 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14146 : _GEN_10570; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14579 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14147 : _GEN_10571; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14580 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14148 : _GEN_10572; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14581 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14149 : _GEN_10573; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14582 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14150 : _GEN_10574; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14583 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14151 : _GEN_10575; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14584 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14152 : _GEN_10576; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14585 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14153 : _GEN_10577; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14586 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14154 : _GEN_10578; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14587 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14155 : _GEN_10579; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14588 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14156 : _GEN_10580; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14589 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14157 : _GEN_10581; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14590 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14158 : _GEN_10582; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14591 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14159 : _GEN_10583; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14592 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14160 : _GEN_10584; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14593 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14161 : _GEN_10585; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14594 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14162 : _GEN_10586; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14595 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14163 : _GEN_10587; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14596 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14164 : _GEN_10588; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14597 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14165 : _GEN_10589; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14710 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14278 : _GEN_10702; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14711 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14279 : _GEN_10703; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14712 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14280 : _GEN_10704; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14713 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14281 : _GEN_10705; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14714 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14282 : _GEN_10706; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14715 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14283 : _GEN_10707; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14716 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14284 : _GEN_10708; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14717 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14285 : _GEN_10709; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14718 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14286 : _GEN_10710; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14719 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14287 : _GEN_10711; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14720 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14288 : _GEN_10712; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14721 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14289 : _GEN_10713; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14722 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14290 : _GEN_10714; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14723 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14291 : _GEN_10715; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14724 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14292 : _GEN_10716; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14725 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14293 : _GEN_10717; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14838 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_12686 : _GEN_10830; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14839 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_12687 : _GEN_10831; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14840 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_12688 : _GEN_10832; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14841 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_12689 : _GEN_10833; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14842 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_12690 : _GEN_10834; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14843 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_12691 : _GEN_10835; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14844 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_12692 : _GEN_10836; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14845 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_12693 : _GEN_10837; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14846 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_12694 : _GEN_10838; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14847 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_12695 : _GEN_10839; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14848 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_12696 : _GEN_10840; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14849 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_12697 : _GEN_10841; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14850 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_12698 : _GEN_10842; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14851 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_12699 : _GEN_10843; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14852 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_12700 : _GEN_10844; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14853 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_12701 : _GEN_10845; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14854 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_12702 : _GEN_10846; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14855 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_12703 : _GEN_10847; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14856 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_12704 : _GEN_10848; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14857 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_12705 : _GEN_10849; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14858 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_12706 : _GEN_10850; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14859 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_12707 : _GEN_10851; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14860 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_12708 : _GEN_10852; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14861 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_12709 : _GEN_10853; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14862 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_12710 : _GEN_10854; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14863 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_12711 : _GEN_10855; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14864 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_12712 : _GEN_10856; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14865 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_12713 : _GEN_10857; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14866 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_12714 : _GEN_10858; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14867 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_12715 : _GEN_10859; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14868 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_12716 : _GEN_10860; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14869 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_12717 : _GEN_10861; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14870 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_12718 : _GEN_10862; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14871 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_12719 : _GEN_10863; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14872 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_12720 : _GEN_10864; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14873 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_12721 : _GEN_10865; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14874 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_12722 : _GEN_10866; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14875 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_12723 : _GEN_10867; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14876 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_12724 : _GEN_10868; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14877 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_12725 : _GEN_10869; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14878 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_12726 : _GEN_10870; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14879 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_12727 : _GEN_10871; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14880 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_12728 : _GEN_10872; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14881 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_12729 : _GEN_10873; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14882 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_12730 : _GEN_10874; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14883 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_12731 : _GEN_10875; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14884 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_12732 : _GEN_10876; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14885 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_12733 : _GEN_10877; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14918 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_12766 : _GEN_10910; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14919 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_12767 : _GEN_10911; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14920 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_12768 : _GEN_10912; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14921 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_12769 : _GEN_10913; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14922 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_12770 : _GEN_10914; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14923 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_12771 : _GEN_10915; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14924 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_12772 : _GEN_10916; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14925 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_12773 : _GEN_10917; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14926 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_12774 : _GEN_10918; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14927 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_12775 : _GEN_10919; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14928 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_12776 : _GEN_10920; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14929 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_12777 : _GEN_10921; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14930 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_12778 : _GEN_10922; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14931 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_12779 : _GEN_10923; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14932 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_12780 : _GEN_10924; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_14933 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_12781 : _GEN_10925; // @[LoadQueueFlag.scala 204:43]
  wire [6:0] _GEN_15350 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13198 : _GEN_11342; // @[LoadQueueFlag.scala 204:43]
  wire [6:0] _GEN_15351 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13199 : _GEN_11343; // @[LoadQueueFlag.scala 204:43]
  wire [6:0] _GEN_15352 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13200 : _GEN_11344; // @[LoadQueueFlag.scala 204:43]
  wire [6:0] _GEN_15353 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13201 : _GEN_11345; // @[LoadQueueFlag.scala 204:43]
  wire [6:0] _GEN_15354 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13202 : _GEN_11346; // @[LoadQueueFlag.scala 204:43]
  wire [6:0] _GEN_15355 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13203 : _GEN_11347; // @[LoadQueueFlag.scala 204:43]
  wire [6:0] _GEN_15356 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13204 : _GEN_11348; // @[LoadQueueFlag.scala 204:43]
  wire [6:0] _GEN_15357 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13205 : _GEN_11349; // @[LoadQueueFlag.scala 204:43]
  wire [6:0] _GEN_15358 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13206 : _GEN_11350; // @[LoadQueueFlag.scala 204:43]
  wire [6:0] _GEN_15359 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13207 : _GEN_11351; // @[LoadQueueFlag.scala 204:43]
  wire [6:0] _GEN_15360 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13208 : _GEN_11352; // @[LoadQueueFlag.scala 204:43]
  wire [6:0] _GEN_15361 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13209 : _GEN_11353; // @[LoadQueueFlag.scala 204:43]
  wire [6:0] _GEN_15362 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13210 : _GEN_11354; // @[LoadQueueFlag.scala 204:43]
  wire [6:0] _GEN_15363 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13211 : _GEN_11355; // @[LoadQueueFlag.scala 204:43]
  wire [6:0] _GEN_15364 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13212 : _GEN_11356; // @[LoadQueueFlag.scala 204:43]
  wire [6:0] _GEN_15365 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13213 : _GEN_11357; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_15366 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13214 : _GEN_11358; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_15367 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13215 : _GEN_11359; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_15368 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13216 : _GEN_11360; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_15369 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13217 : _GEN_11361; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_15370 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13218 : _GEN_11362; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_15371 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13219 : _GEN_11363; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_15372 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13220 : _GEN_11364; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_15373 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13221 : _GEN_11365; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_15374 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13222 : _GEN_11366; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_15375 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13223 : _GEN_11367; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_15376 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13224 : _GEN_11368; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_15377 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13225 : _GEN_11369; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_15378 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13226 : _GEN_11370; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_15379 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13227 : _GEN_11371; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_15380 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13228 : _GEN_11372; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_15381 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13229 : _GEN_11373; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_15382 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13230 : _GEN_11374; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_15383 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13231 : _GEN_11375; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_15384 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13232 : _GEN_11376; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_15385 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13233 : _GEN_11377; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_15386 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13234 : _GEN_11378; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_15387 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13235 : _GEN_11379; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_15388 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13236 : _GEN_11380; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_15389 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13237 : _GEN_11381; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_15390 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13238 : _GEN_11382; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_15391 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13239 : _GEN_11383; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_15392 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13240 : _GEN_11384; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_15393 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13241 : _GEN_11385; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_15394 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13242 : _GEN_11386; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_15395 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13243 : _GEN_11387; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_15396 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13244 : _GEN_11388; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_15397 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13245 : _GEN_11389; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_15446 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13294 : _GEN_11438; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_15447 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13295 : _GEN_11439; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_15448 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13296 : _GEN_11440; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_15449 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13297 : _GEN_11441; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_15450 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13298 : _GEN_11442; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_15451 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13299 : _GEN_11443; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_15452 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13300 : _GEN_11444; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_15453 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13301 : _GEN_11445; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_15454 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13302 : _GEN_11446; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_15455 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13303 : _GEN_11447; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_15456 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13304 : _GEN_11448; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_15457 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13305 : _GEN_11449; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_15458 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13306 : _GEN_11450; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_15459 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13307 : _GEN_11451; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_15460 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13308 : _GEN_11452; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_15461 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13309 : _GEN_11453; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_15766 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13614 : _GEN_11758; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_15767 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13615 : _GEN_11759; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_15768 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13616 : _GEN_11760; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_15769 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13617 : _GEN_11761; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_15770 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13618 : _GEN_11762; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_15771 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13619 : _GEN_11763; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_15772 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13620 : _GEN_11764; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_15773 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13621 : _GEN_11765; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_15774 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13622 : _GEN_11766; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_15775 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13623 : _GEN_11767; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_15776 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13624 : _GEN_11768; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_15777 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13625 : _GEN_11769; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_15778 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13626 : _GEN_11770; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_15779 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13627 : _GEN_11771; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_15780 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13628 : _GEN_11772; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_15781 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13629 : _GEN_11773; // @[LoadQueueFlag.scala 204:43]
  wire [5:0] _GEN_15878 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13726 : _GEN_11870; // @[LoadQueueFlag.scala 204:43]
  wire [5:0] _GEN_15879 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13727 : _GEN_11871; // @[LoadQueueFlag.scala 204:43]
  wire [5:0] _GEN_15880 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13728 : _GEN_11872; // @[LoadQueueFlag.scala 204:43]
  wire [5:0] _GEN_15881 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13729 : _GEN_11873; // @[LoadQueueFlag.scala 204:43]
  wire [5:0] _GEN_15882 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13730 : _GEN_11874; // @[LoadQueueFlag.scala 204:43]
  wire [5:0] _GEN_15883 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13731 : _GEN_11875; // @[LoadQueueFlag.scala 204:43]
  wire [5:0] _GEN_15884 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13732 : _GEN_11876; // @[LoadQueueFlag.scala 204:43]
  wire [5:0] _GEN_15885 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13733 : _GEN_11877; // @[LoadQueueFlag.scala 204:43]
  wire [5:0] _GEN_15886 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13734 : _GEN_11878; // @[LoadQueueFlag.scala 204:43]
  wire [5:0] _GEN_15887 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13735 : _GEN_11879; // @[LoadQueueFlag.scala 204:43]
  wire [5:0] _GEN_15888 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13736 : _GEN_11880; // @[LoadQueueFlag.scala 204:43]
  wire [5:0] _GEN_15889 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13737 : _GEN_11881; // @[LoadQueueFlag.scala 204:43]
  wire [5:0] _GEN_15890 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13738 : _GEN_11882; // @[LoadQueueFlag.scala 204:43]
  wire [5:0] _GEN_15891 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13739 : _GEN_11883; // @[LoadQueueFlag.scala 204:43]
  wire [5:0] _GEN_15892 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13740 : _GEN_11884; // @[LoadQueueFlag.scala 204:43]
  wire [5:0] _GEN_15893 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_13741 : _GEN_11885; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_16182 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14326 : _GEN_12174; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_16183 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14327 : _GEN_12175; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_16184 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14328 : _GEN_12176; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_16185 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14329 : _GEN_12177; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_16186 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14330 : _GEN_12178; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_16187 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14331 : _GEN_12179; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_16188 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14332 : _GEN_12180; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_16189 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14333 : _GEN_12181; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_16190 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14334 : _GEN_12182; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_16191 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14335 : _GEN_12183; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_16192 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14336 : _GEN_12184; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_16193 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14337 : _GEN_12185; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_16194 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14338 : _GEN_12186; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_16195 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14339 : _GEN_12187; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_16196 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14340 : _GEN_12188; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_16197 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14341 : _GEN_12189; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_16198 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14342 : _GEN_12190; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_16199 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14343 : _GEN_12191; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_16200 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14344 : _GEN_12192; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_16201 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14345 : _GEN_12193; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_16202 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14346 : _GEN_12194; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_16203 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14347 : _GEN_12195; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_16204 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14348 : _GEN_12196; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_16205 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14349 : _GEN_12197; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_16206 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14350 : _GEN_12198; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_16207 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14351 : _GEN_12199; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_16208 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14352 : _GEN_12200; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_16209 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14353 : _GEN_12201; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_16210 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14354 : _GEN_12202; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_16211 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14355 : _GEN_12203; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_16212 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14356 : _GEN_12204; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_16213 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14357 : _GEN_12205; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_16214 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14358 : _GEN_12206; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_16215 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14359 : _GEN_12207; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_16216 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14360 : _GEN_12208; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_16217 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14361 : _GEN_12209; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_16218 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14362 : _GEN_12210; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_16219 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14363 : _GEN_12211; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_16220 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14364 : _GEN_12212; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_16221 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14365 : _GEN_12213; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_16222 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14366 : _GEN_12214; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_16223 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14367 : _GEN_12215; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_16224 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14368 : _GEN_12216; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_16225 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14369 : _GEN_12217; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_16226 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14370 : _GEN_12218; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_16227 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14371 : _GEN_12219; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_16228 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14372 : _GEN_12220; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_16229 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14373 : _GEN_12221; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_16230 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14374 : _GEN_12222; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_16231 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14375 : _GEN_12223; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_16232 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14376 : _GEN_12224; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_16233 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14377 : _GEN_12225; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_16234 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14378 : _GEN_12226; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_16235 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14379 : _GEN_12227; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_16236 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14380 : _GEN_12228; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_16237 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14381 : _GEN_12229; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_16238 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14382 : _GEN_12230; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_16239 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14383 : _GEN_12231; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_16240 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14384 : _GEN_12232; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_16241 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14385 : _GEN_12233; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_16242 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14386 : _GEN_12234; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_16243 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14387 : _GEN_12235; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_16244 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14388 : _GEN_12236; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_16245 = io_enq_req_3_valid & ~enqCancel_3 ? _GEN_14389 : _GEN_12237; // @[LoadQueueFlag.scala 204:43]
  wire  _GEN_16294 = 4'h0 == deqLookupVec_new_ptr_value ? 1'h0 : _GEN_14438; // @[LoadQueueFlag.scala 233:{40,40}]
  wire  _GEN_16295 = 4'h1 == deqLookupVec_new_ptr_value ? 1'h0 : _GEN_14439; // @[LoadQueueFlag.scala 233:{40,40}]
  wire  _GEN_16296 = 4'h2 == deqLookupVec_new_ptr_value ? 1'h0 : _GEN_14440; // @[LoadQueueFlag.scala 233:{40,40}]
  wire  _GEN_16297 = 4'h3 == deqLookupVec_new_ptr_value ? 1'h0 : _GEN_14441; // @[LoadQueueFlag.scala 233:{40,40}]
  wire  _GEN_16298 = 4'h4 == deqLookupVec_new_ptr_value ? 1'h0 : _GEN_14442; // @[LoadQueueFlag.scala 233:{40,40}]
  wire  _GEN_16299 = 4'h5 == deqLookupVec_new_ptr_value ? 1'h0 : _GEN_14443; // @[LoadQueueFlag.scala 233:{40,40}]
  wire  _GEN_16300 = 4'h6 == deqLookupVec_new_ptr_value ? 1'h0 : _GEN_14444; // @[LoadQueueFlag.scala 233:{40,40}]
  wire  _GEN_16301 = 4'h7 == deqLookupVec_new_ptr_value ? 1'h0 : _GEN_14445; // @[LoadQueueFlag.scala 233:{40,40}]
  wire  _GEN_16302 = 4'h8 == deqLookupVec_new_ptr_value ? 1'h0 : _GEN_14446; // @[LoadQueueFlag.scala 233:{40,40}]
  wire  _GEN_16303 = 4'h9 == deqLookupVec_new_ptr_value ? 1'h0 : _GEN_14447; // @[LoadQueueFlag.scala 233:{40,40}]
  wire  _GEN_16304 = 4'ha == deqLookupVec_new_ptr_value ? 1'h0 : _GEN_14448; // @[LoadQueueFlag.scala 233:{40,40}]
  wire  _GEN_16305 = 4'hb == deqLookupVec_new_ptr_value ? 1'h0 : _GEN_14449; // @[LoadQueueFlag.scala 233:{40,40}]
  wire  _GEN_16306 = 4'hc == deqLookupVec_new_ptr_value ? 1'h0 : _GEN_14450; // @[LoadQueueFlag.scala 233:{40,40}]
  wire  _GEN_16307 = 4'hd == deqLookupVec_new_ptr_value ? 1'h0 : _GEN_14451; // @[LoadQueueFlag.scala 233:{40,40}]
  wire  _GEN_16308 = 4'he == deqLookupVec_new_ptr_value ? 1'h0 : _GEN_14452; // @[LoadQueueFlag.scala 233:{40,40}]
  wire  _GEN_16309 = 4'hf == deqLookupVec_new_ptr_value ? 1'h0 : _GEN_14453; // @[LoadQueueFlag.scala 233:{40,40}]
  wire  _GEN_16326 = commitCount > 2'h0 ? _GEN_16294 : _GEN_14438; // @[LoadQueueFlag.scala 232:30]
  wire  _GEN_16327 = commitCount > 2'h0 ? _GEN_16295 : _GEN_14439; // @[LoadQueueFlag.scala 232:30]
  wire  _GEN_16328 = commitCount > 2'h0 ? _GEN_16296 : _GEN_14440; // @[LoadQueueFlag.scala 232:30]
  wire  _GEN_16329 = commitCount > 2'h0 ? _GEN_16297 : _GEN_14441; // @[LoadQueueFlag.scala 232:30]
  wire  _GEN_16330 = commitCount > 2'h0 ? _GEN_16298 : _GEN_14442; // @[LoadQueueFlag.scala 232:30]
  wire  _GEN_16331 = commitCount > 2'h0 ? _GEN_16299 : _GEN_14443; // @[LoadQueueFlag.scala 232:30]
  wire  _GEN_16332 = commitCount > 2'h0 ? _GEN_16300 : _GEN_14444; // @[LoadQueueFlag.scala 232:30]
  wire  _GEN_16333 = commitCount > 2'h0 ? _GEN_16301 : _GEN_14445; // @[LoadQueueFlag.scala 232:30]
  wire  _GEN_16334 = commitCount > 2'h0 ? _GEN_16302 : _GEN_14446; // @[LoadQueueFlag.scala 232:30]
  wire  _GEN_16335 = commitCount > 2'h0 ? _GEN_16303 : _GEN_14447; // @[LoadQueueFlag.scala 232:30]
  wire  _GEN_16336 = commitCount > 2'h0 ? _GEN_16304 : _GEN_14448; // @[LoadQueueFlag.scala 232:30]
  wire  _GEN_16337 = commitCount > 2'h0 ? _GEN_16305 : _GEN_14449; // @[LoadQueueFlag.scala 232:30]
  wire  _GEN_16338 = commitCount > 2'h0 ? _GEN_16306 : _GEN_14450; // @[LoadQueueFlag.scala 232:30]
  wire  _GEN_16339 = commitCount > 2'h0 ? _GEN_16307 : _GEN_14451; // @[LoadQueueFlag.scala 232:30]
  wire  _GEN_16340 = commitCount > 2'h0 ? _GEN_16308 : _GEN_14452; // @[LoadQueueFlag.scala 232:30]
  wire  _GEN_16341 = commitCount > 2'h0 ? _GEN_16309 : _GEN_14453; // @[LoadQueueFlag.scala 232:30]
  wire [15:0] _hasExceptions_T = {2'h0,io_loadIn_0_bits_uop_cf_exceptionVec_13,1'h0,4'h0,2'h0,
    io_loadIn_0_bits_uop_cf_exceptionVec_5,io_loadIn_0_bits_uop_cf_exceptionVec_4,4'h0}; // @[LoadQueueFlag.scala 287:97]
  wire  hasExceptions = |_hasExceptions_T; // @[LoadQueueFlag.scala 287:104]
  wire [7:0] _needReplay_T = {io_loadIn_0_bits_replayInfo_cause_7,io_loadIn_0_bits_replayInfo_cause_6,
    io_loadIn_0_bits_replayInfo_cause_5,io_loadIn_0_bits_replayInfo_cause_4,io_loadIn_0_bits_replayInfo_cause_3,
    io_loadIn_0_bits_replayInfo_cause_2,io_loadIn_0_bits_replayInfo_cause_1,io_loadIn_0_bits_replayInfo_cause_0}; // @[LoadUnit.scala 62:29]
  wire  needReplay = |_needReplay_T; // @[LoadUnit.scala 62:36]
  wire  _datavalidVal_T = ~io_loadIn_0_bits_mmio; // @[LoadQueueFlag.scala 295:13]
  wire  _datavalidVal_T_1 = ~io_loadIn_0_bits_miss; // @[LoadQueueFlag.scala 296:13]
  wire  datavalidVal = ~io_loadIn_0_bits_mmio & _datavalidVal_T_1; // @[LoadQueueFlag.scala 295:37]
  wire  _issued_T_1 = ~needReplay; // @[LoadQueueFlag.scala 299:29]
  wire  _issued_T_2 = ~io_loadIn_0_bits_tlbMiss; // @[LoadQueueFlag.scala 299:44]
  wire  _GEN_16502 = 4'h0 == io_loadIn_0_bits_uop_lqIdx_value ? _issued_T_2 : _GEN_16182; // @[LoadQueueFlag.scala 303:{32,32}]
  wire  _GEN_16503 = 4'h1 == io_loadIn_0_bits_uop_lqIdx_value ? _issued_T_2 : _GEN_16183; // @[LoadQueueFlag.scala 303:{32,32}]
  wire  _GEN_16504 = 4'h2 == io_loadIn_0_bits_uop_lqIdx_value ? _issued_T_2 : _GEN_16184; // @[LoadQueueFlag.scala 303:{32,32}]
  wire  _GEN_16505 = 4'h3 == io_loadIn_0_bits_uop_lqIdx_value ? _issued_T_2 : _GEN_16185; // @[LoadQueueFlag.scala 303:{32,32}]
  wire  _GEN_16506 = 4'h4 == io_loadIn_0_bits_uop_lqIdx_value ? _issued_T_2 : _GEN_16186; // @[LoadQueueFlag.scala 303:{32,32}]
  wire  _GEN_16507 = 4'h5 == io_loadIn_0_bits_uop_lqIdx_value ? _issued_T_2 : _GEN_16187; // @[LoadQueueFlag.scala 303:{32,32}]
  wire  _GEN_16508 = 4'h6 == io_loadIn_0_bits_uop_lqIdx_value ? _issued_T_2 : _GEN_16188; // @[LoadQueueFlag.scala 303:{32,32}]
  wire  _GEN_16509 = 4'h7 == io_loadIn_0_bits_uop_lqIdx_value ? _issued_T_2 : _GEN_16189; // @[LoadQueueFlag.scala 303:{32,32}]
  wire  _GEN_16510 = 4'h8 == io_loadIn_0_bits_uop_lqIdx_value ? _issued_T_2 : _GEN_16190; // @[LoadQueueFlag.scala 303:{32,32}]
  wire  _GEN_16511 = 4'h9 == io_loadIn_0_bits_uop_lqIdx_value ? _issued_T_2 : _GEN_16191; // @[LoadQueueFlag.scala 303:{32,32}]
  wire  _GEN_16512 = 4'ha == io_loadIn_0_bits_uop_lqIdx_value ? _issued_T_2 : _GEN_16192; // @[LoadQueueFlag.scala 303:{32,32}]
  wire  _GEN_16513 = 4'hb == io_loadIn_0_bits_uop_lqIdx_value ? _issued_T_2 : _GEN_16193; // @[LoadQueueFlag.scala 303:{32,32}]
  wire  _GEN_16514 = 4'hc == io_loadIn_0_bits_uop_lqIdx_value ? _issued_T_2 : _GEN_16194; // @[LoadQueueFlag.scala 303:{32,32}]
  wire  _GEN_16515 = 4'hd == io_loadIn_0_bits_uop_lqIdx_value ? _issued_T_2 : _GEN_16195; // @[LoadQueueFlag.scala 303:{32,32}]
  wire  _GEN_16516 = 4'he == io_loadIn_0_bits_uop_lqIdx_value ? _issued_T_2 : _GEN_16196; // @[LoadQueueFlag.scala 303:{32,32}]
  wire  _GEN_16517 = 4'hf == io_loadIn_0_bits_uop_lqIdx_value ? _issued_T_2 : _GEN_16197; // @[LoadQueueFlag.scala 303:{32,32}]
  wire  _GEN_16518 = 4'h0 == io_loadIn_0_bits_uop_lqIdx_value ? datavalidVal : _GEN_16198; // @[LoadQueueFlag.scala 304:{32,32}]
  wire  _GEN_16519 = 4'h1 == io_loadIn_0_bits_uop_lqIdx_value ? datavalidVal : _GEN_16199; // @[LoadQueueFlag.scala 304:{32,32}]
  wire  _GEN_16520 = 4'h2 == io_loadIn_0_bits_uop_lqIdx_value ? datavalidVal : _GEN_16200; // @[LoadQueueFlag.scala 304:{32,32}]
  wire  _GEN_16521 = 4'h3 == io_loadIn_0_bits_uop_lqIdx_value ? datavalidVal : _GEN_16201; // @[LoadQueueFlag.scala 304:{32,32}]
  wire  _GEN_16522 = 4'h4 == io_loadIn_0_bits_uop_lqIdx_value ? datavalidVal : _GEN_16202; // @[LoadQueueFlag.scala 304:{32,32}]
  wire  _GEN_16523 = 4'h5 == io_loadIn_0_bits_uop_lqIdx_value ? datavalidVal : _GEN_16203; // @[LoadQueueFlag.scala 304:{32,32}]
  wire  _GEN_16524 = 4'h6 == io_loadIn_0_bits_uop_lqIdx_value ? datavalidVal : _GEN_16204; // @[LoadQueueFlag.scala 304:{32,32}]
  wire  _GEN_16525 = 4'h7 == io_loadIn_0_bits_uop_lqIdx_value ? datavalidVal : _GEN_16205; // @[LoadQueueFlag.scala 304:{32,32}]
  wire  _GEN_16526 = 4'h8 == io_loadIn_0_bits_uop_lqIdx_value ? datavalidVal : _GEN_16206; // @[LoadQueueFlag.scala 304:{32,32}]
  wire  _GEN_16527 = 4'h9 == io_loadIn_0_bits_uop_lqIdx_value ? datavalidVal : _GEN_16207; // @[LoadQueueFlag.scala 304:{32,32}]
  wire  _GEN_16528 = 4'ha == io_loadIn_0_bits_uop_lqIdx_value ? datavalidVal : _GEN_16208; // @[LoadQueueFlag.scala 304:{32,32}]
  wire  _GEN_16529 = 4'hb == io_loadIn_0_bits_uop_lqIdx_value ? datavalidVal : _GEN_16209; // @[LoadQueueFlag.scala 304:{32,32}]
  wire  _GEN_16530 = 4'hc == io_loadIn_0_bits_uop_lqIdx_value ? datavalidVal : _GEN_16210; // @[LoadQueueFlag.scala 304:{32,32}]
  wire  _GEN_16531 = 4'hd == io_loadIn_0_bits_uop_lqIdx_value ? datavalidVal : _GEN_16211; // @[LoadQueueFlag.scala 304:{32,32}]
  wire  _GEN_16532 = 4'he == io_loadIn_0_bits_uop_lqIdx_value ? datavalidVal : _GEN_16212; // @[LoadQueueFlag.scala 304:{32,32}]
  wire  _GEN_16533 = 4'hf == io_loadIn_0_bits_uop_lqIdx_value ? datavalidVal : _GEN_16213; // @[LoadQueueFlag.scala 304:{32,32}]
  wire  _GEN_16534 = 4'h0 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_mmio : _GEN_16214; // @[LoadQueueFlag.scala 305:{30,30}]
  wire  _GEN_16535 = 4'h1 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_mmio : _GEN_16215; // @[LoadQueueFlag.scala 305:{30,30}]
  wire  _GEN_16536 = 4'h2 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_mmio : _GEN_16216; // @[LoadQueueFlag.scala 305:{30,30}]
  wire  _GEN_16537 = 4'h3 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_mmio : _GEN_16217; // @[LoadQueueFlag.scala 305:{30,30}]
  wire  _GEN_16538 = 4'h4 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_mmio : _GEN_16218; // @[LoadQueueFlag.scala 305:{30,30}]
  wire  _GEN_16539 = 4'h5 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_mmio : _GEN_16219; // @[LoadQueueFlag.scala 305:{30,30}]
  wire  _GEN_16540 = 4'h6 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_mmio : _GEN_16220; // @[LoadQueueFlag.scala 305:{30,30}]
  wire  _GEN_16541 = 4'h7 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_mmio : _GEN_16221; // @[LoadQueueFlag.scala 305:{30,30}]
  wire  _GEN_16542 = 4'h8 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_mmio : _GEN_16222; // @[LoadQueueFlag.scala 305:{30,30}]
  wire  _GEN_16543 = 4'h9 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_mmio : _GEN_16223; // @[LoadQueueFlag.scala 305:{30,30}]
  wire  _GEN_16544 = 4'ha == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_mmio : _GEN_16224; // @[LoadQueueFlag.scala 305:{30,30}]
  wire  _GEN_16545 = 4'hb == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_mmio : _GEN_16225; // @[LoadQueueFlag.scala 305:{30,30}]
  wire  _GEN_16546 = 4'hc == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_mmio : _GEN_16226; // @[LoadQueueFlag.scala 305:{30,30}]
  wire  _GEN_16547 = 4'hd == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_mmio : _GEN_16227; // @[LoadQueueFlag.scala 305:{30,30}]
  wire  _GEN_16548 = 4'he == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_mmio : _GEN_16228; // @[LoadQueueFlag.scala 305:{30,30}]
  wire  _GEN_16549 = 4'hf == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_mmio : _GEN_16229; // @[LoadQueueFlag.scala 305:{30,30}]
  wire  _GEN_16550 = 4'h0 == io_loadIn_0_bits_uop_lqIdx_value ? _datavalidVal_T & ~hasExceptions : _GEN_16230; // @[LoadQueueFlag.scala 306:{34,34}]
  wire  _GEN_16551 = 4'h1 == io_loadIn_0_bits_uop_lqIdx_value ? _datavalidVal_T & ~hasExceptions : _GEN_16231; // @[LoadQueueFlag.scala 306:{34,34}]
  wire  _GEN_16552 = 4'h2 == io_loadIn_0_bits_uop_lqIdx_value ? _datavalidVal_T & ~hasExceptions : _GEN_16232; // @[LoadQueueFlag.scala 306:{34,34}]
  wire  _GEN_16553 = 4'h3 == io_loadIn_0_bits_uop_lqIdx_value ? _datavalidVal_T & ~hasExceptions : _GEN_16233; // @[LoadQueueFlag.scala 306:{34,34}]
  wire  _GEN_16554 = 4'h4 == io_loadIn_0_bits_uop_lqIdx_value ? _datavalidVal_T & ~hasExceptions : _GEN_16234; // @[LoadQueueFlag.scala 306:{34,34}]
  wire  _GEN_16555 = 4'h5 == io_loadIn_0_bits_uop_lqIdx_value ? _datavalidVal_T & ~hasExceptions : _GEN_16235; // @[LoadQueueFlag.scala 306:{34,34}]
  wire  _GEN_16556 = 4'h6 == io_loadIn_0_bits_uop_lqIdx_value ? _datavalidVal_T & ~hasExceptions : _GEN_16236; // @[LoadQueueFlag.scala 306:{34,34}]
  wire  _GEN_16557 = 4'h7 == io_loadIn_0_bits_uop_lqIdx_value ? _datavalidVal_T & ~hasExceptions : _GEN_16237; // @[LoadQueueFlag.scala 306:{34,34}]
  wire  _GEN_16558 = 4'h8 == io_loadIn_0_bits_uop_lqIdx_value ? _datavalidVal_T & ~hasExceptions : _GEN_16238; // @[LoadQueueFlag.scala 306:{34,34}]
  wire  _GEN_16559 = 4'h9 == io_loadIn_0_bits_uop_lqIdx_value ? _datavalidVal_T & ~hasExceptions : _GEN_16239; // @[LoadQueueFlag.scala 306:{34,34}]
  wire  _GEN_16560 = 4'ha == io_loadIn_0_bits_uop_lqIdx_value ? _datavalidVal_T & ~hasExceptions : _GEN_16240; // @[LoadQueueFlag.scala 306:{34,34}]
  wire  _GEN_16561 = 4'hb == io_loadIn_0_bits_uop_lqIdx_value ? _datavalidVal_T & ~hasExceptions : _GEN_16241; // @[LoadQueueFlag.scala 306:{34,34}]
  wire  _GEN_16562 = 4'hc == io_loadIn_0_bits_uop_lqIdx_value ? _datavalidVal_T & ~hasExceptions : _GEN_16242; // @[LoadQueueFlag.scala 306:{34,34}]
  wire  _GEN_16563 = 4'hd == io_loadIn_0_bits_uop_lqIdx_value ? _datavalidVal_T & ~hasExceptions : _GEN_16243; // @[LoadQueueFlag.scala 306:{34,34}]
  wire  _GEN_16564 = 4'he == io_loadIn_0_bits_uop_lqIdx_value ? _datavalidVal_T & ~hasExceptions : _GEN_16244; // @[LoadQueueFlag.scala 306:{34,34}]
  wire  _GEN_16565 = 4'hf == io_loadIn_0_bits_uop_lqIdx_value ? _datavalidVal_T & ~hasExceptions : _GEN_16245; // @[LoadQueueFlag.scala 306:{34,34}]
  wire [5:0] _GEN_16566 = 4'h0 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_pdest : _GEN_15878; // @[LoadQueueFlag.scala 310:{34,34}]
  wire [5:0] _GEN_16567 = 4'h1 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_pdest : _GEN_15879; // @[LoadQueueFlag.scala 310:{34,34}]
  wire [5:0] _GEN_16568 = 4'h2 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_pdest : _GEN_15880; // @[LoadQueueFlag.scala 310:{34,34}]
  wire [5:0] _GEN_16569 = 4'h3 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_pdest : _GEN_15881; // @[LoadQueueFlag.scala 310:{34,34}]
  wire [5:0] _GEN_16570 = 4'h4 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_pdest : _GEN_15882; // @[LoadQueueFlag.scala 310:{34,34}]
  wire [5:0] _GEN_16571 = 4'h5 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_pdest : _GEN_15883; // @[LoadQueueFlag.scala 310:{34,34}]
  wire [5:0] _GEN_16572 = 4'h6 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_pdest : _GEN_15884; // @[LoadQueueFlag.scala 310:{34,34}]
  wire [5:0] _GEN_16573 = 4'h7 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_pdest : _GEN_15885; // @[LoadQueueFlag.scala 310:{34,34}]
  wire [5:0] _GEN_16574 = 4'h8 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_pdest : _GEN_15886; // @[LoadQueueFlag.scala 310:{34,34}]
  wire [5:0] _GEN_16575 = 4'h9 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_pdest : _GEN_15887; // @[LoadQueueFlag.scala 310:{34,34}]
  wire [5:0] _GEN_16576 = 4'ha == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_pdest : _GEN_15888; // @[LoadQueueFlag.scala 310:{34,34}]
  wire [5:0] _GEN_16577 = 4'hb == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_pdest : _GEN_15889; // @[LoadQueueFlag.scala 310:{34,34}]
  wire [5:0] _GEN_16578 = 4'hc == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_pdest : _GEN_15890; // @[LoadQueueFlag.scala 310:{34,34}]
  wire [5:0] _GEN_16579 = 4'hd == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_pdest : _GEN_15891; // @[LoadQueueFlag.scala 310:{34,34}]
  wire [5:0] _GEN_16580 = 4'he == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_pdest : _GEN_15892; // @[LoadQueueFlag.scala 310:{34,34}]
  wire [5:0] _GEN_16581 = 4'hf == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_pdest : _GEN_15893; // @[LoadQueueFlag.scala 310:{34,34}]
  wire [5:0] _GEN_16582 = io_loadIn_0_bits_lqDataWenDup_1 ? _GEN_16566 : _GEN_15878; // @[LoadQueueFlag.scala 309:50]
  wire [5:0] _GEN_16583 = io_loadIn_0_bits_lqDataWenDup_1 ? _GEN_16567 : _GEN_15879; // @[LoadQueueFlag.scala 309:50]
  wire [5:0] _GEN_16584 = io_loadIn_0_bits_lqDataWenDup_1 ? _GEN_16568 : _GEN_15880; // @[LoadQueueFlag.scala 309:50]
  wire [5:0] _GEN_16585 = io_loadIn_0_bits_lqDataWenDup_1 ? _GEN_16569 : _GEN_15881; // @[LoadQueueFlag.scala 309:50]
  wire [5:0] _GEN_16586 = io_loadIn_0_bits_lqDataWenDup_1 ? _GEN_16570 : _GEN_15882; // @[LoadQueueFlag.scala 309:50]
  wire [5:0] _GEN_16587 = io_loadIn_0_bits_lqDataWenDup_1 ? _GEN_16571 : _GEN_15883; // @[LoadQueueFlag.scala 309:50]
  wire [5:0] _GEN_16588 = io_loadIn_0_bits_lqDataWenDup_1 ? _GEN_16572 : _GEN_15884; // @[LoadQueueFlag.scala 309:50]
  wire [5:0] _GEN_16589 = io_loadIn_0_bits_lqDataWenDup_1 ? _GEN_16573 : _GEN_15885; // @[LoadQueueFlag.scala 309:50]
  wire [5:0] _GEN_16590 = io_loadIn_0_bits_lqDataWenDup_1 ? _GEN_16574 : _GEN_15886; // @[LoadQueueFlag.scala 309:50]
  wire [5:0] _GEN_16591 = io_loadIn_0_bits_lqDataWenDup_1 ? _GEN_16575 : _GEN_15887; // @[LoadQueueFlag.scala 309:50]
  wire [5:0] _GEN_16592 = io_loadIn_0_bits_lqDataWenDup_1 ? _GEN_16576 : _GEN_15888; // @[LoadQueueFlag.scala 309:50]
  wire [5:0] _GEN_16593 = io_loadIn_0_bits_lqDataWenDup_1 ? _GEN_16577 : _GEN_15889; // @[LoadQueueFlag.scala 309:50]
  wire [5:0] _GEN_16594 = io_loadIn_0_bits_lqDataWenDup_1 ? _GEN_16578 : _GEN_15890; // @[LoadQueueFlag.scala 309:50]
  wire [5:0] _GEN_16595 = io_loadIn_0_bits_lqDataWenDup_1 ? _GEN_16579 : _GEN_15891; // @[LoadQueueFlag.scala 309:50]
  wire [5:0] _GEN_16596 = io_loadIn_0_bits_lqDataWenDup_1 ? _GEN_16580 : _GEN_15892; // @[LoadQueueFlag.scala 309:50]
  wire [5:0] _GEN_16597 = io_loadIn_0_bits_lqDataWenDup_1 ? _GEN_16581 : _GEN_15893; // @[LoadQueueFlag.scala 309:50]
  wire  _GEN_16710 = 4'h0 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_exceptionVec_4 : _GEN_14566; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_16711 = 4'h1 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_exceptionVec_4 : _GEN_14567; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_16712 = 4'h2 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_exceptionVec_4 : _GEN_14568; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_16713 = 4'h3 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_exceptionVec_4 : _GEN_14569; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_16714 = 4'h4 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_exceptionVec_4 : _GEN_14570; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_16715 = 4'h5 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_exceptionVec_4 : _GEN_14571; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_16716 = 4'h6 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_exceptionVec_4 : _GEN_14572; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_16717 = 4'h7 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_exceptionVec_4 : _GEN_14573; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_16718 = 4'h8 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_exceptionVec_4 : _GEN_14574; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_16719 = 4'h9 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_exceptionVec_4 : _GEN_14575; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_16720 = 4'ha == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_exceptionVec_4 : _GEN_14576; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_16721 = 4'hb == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_exceptionVec_4 : _GEN_14577; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_16722 = 4'hc == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_exceptionVec_4 : _GEN_14578; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_16723 = 4'hd == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_exceptionVec_4 : _GEN_14579; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_16724 = 4'he == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_exceptionVec_4 : _GEN_14580; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_16725 = 4'hf == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_exceptionVec_4 : _GEN_14581; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_16726 = 4'h0 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_exceptionVec_5 : _GEN_14582; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_16727 = 4'h1 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_exceptionVec_5 : _GEN_14583; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_16728 = 4'h2 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_exceptionVec_5 : _GEN_14584; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_16729 = 4'h3 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_exceptionVec_5 : _GEN_14585; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_16730 = 4'h4 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_exceptionVec_5 : _GEN_14586; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_16731 = 4'h5 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_exceptionVec_5 : _GEN_14587; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_16732 = 4'h6 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_exceptionVec_5 : _GEN_14588; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_16733 = 4'h7 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_exceptionVec_5 : _GEN_14589; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_16734 = 4'h8 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_exceptionVec_5 : _GEN_14590; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_16735 = 4'h9 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_exceptionVec_5 : _GEN_14591; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_16736 = 4'ha == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_exceptionVec_5 : _GEN_14592; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_16737 = 4'hb == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_exceptionVec_5 : _GEN_14593; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_16738 = 4'hc == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_exceptionVec_5 : _GEN_14594; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_16739 = 4'hd == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_exceptionVec_5 : _GEN_14595; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_16740 = 4'he == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_exceptionVec_5 : _GEN_14596; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_16741 = 4'hf == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_exceptionVec_5 : _GEN_14597; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_16854 = 4'h0 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_exceptionVec_13 : _GEN_14710; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_16855 = 4'h1 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_exceptionVec_13 : _GEN_14711; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_16856 = 4'h2 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_exceptionVec_13 : _GEN_14712; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_16857 = 4'h3 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_exceptionVec_13 : _GEN_14713; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_16858 = 4'h4 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_exceptionVec_13 : _GEN_14714; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_16859 = 4'h5 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_exceptionVec_13 : _GEN_14715; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_16860 = 4'h6 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_exceptionVec_13 : _GEN_14716; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_16861 = 4'h7 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_exceptionVec_13 : _GEN_14717; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_16862 = 4'h8 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_exceptionVec_13 : _GEN_14718; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_16863 = 4'h9 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_exceptionVec_13 : _GEN_14719; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_16864 = 4'ha == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_exceptionVec_13 : _GEN_14720; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_16865 = 4'hb == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_exceptionVec_13 : _GEN_14721; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_16866 = 4'hc == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_exceptionVec_13 : _GEN_14722; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_16867 = 4'hd == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_exceptionVec_13 : _GEN_14723; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_16868 = 4'he == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_exceptionVec_13 : _GEN_14724; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_16869 = 4'hf == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_exceptionVec_13 : _GEN_14725; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_16982 = 4'h0 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_trigger_backendEn_1 : _GEN_14838
    ; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_16983 = 4'h1 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_trigger_backendEn_1 : _GEN_14839
    ; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_16984 = 4'h2 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_trigger_backendEn_1 : _GEN_14840
    ; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_16985 = 4'h3 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_trigger_backendEn_1 : _GEN_14841
    ; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_16986 = 4'h4 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_trigger_backendEn_1 : _GEN_14842
    ; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_16987 = 4'h5 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_trigger_backendEn_1 : _GEN_14843
    ; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_16988 = 4'h6 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_trigger_backendEn_1 : _GEN_14844
    ; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_16989 = 4'h7 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_trigger_backendEn_1 : _GEN_14845
    ; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_16990 = 4'h8 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_trigger_backendEn_1 : _GEN_14846
    ; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_16991 = 4'h9 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_trigger_backendEn_1 : _GEN_14847
    ; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_16992 = 4'ha == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_trigger_backendEn_1 : _GEN_14848
    ; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_16993 = 4'hb == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_trigger_backendEn_1 : _GEN_14849
    ; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_16994 = 4'hc == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_trigger_backendEn_1 : _GEN_14850
    ; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_16995 = 4'hd == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_trigger_backendEn_1 : _GEN_14851
    ; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_16996 = 4'he == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_trigger_backendEn_1 : _GEN_14852
    ; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_16997 = 4'hf == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_trigger_backendEn_1 : _GEN_14853
    ; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_16998 = 4'h0 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_trigger_backendHit_0 :
    _GEN_14854; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_16999 = 4'h1 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_trigger_backendHit_0 :
    _GEN_14855; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_17000 = 4'h2 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_trigger_backendHit_0 :
    _GEN_14856; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_17001 = 4'h3 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_trigger_backendHit_0 :
    _GEN_14857; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_17002 = 4'h4 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_trigger_backendHit_0 :
    _GEN_14858; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_17003 = 4'h5 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_trigger_backendHit_0 :
    _GEN_14859; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_17004 = 4'h6 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_trigger_backendHit_0 :
    _GEN_14860; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_17005 = 4'h7 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_trigger_backendHit_0 :
    _GEN_14861; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_17006 = 4'h8 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_trigger_backendHit_0 :
    _GEN_14862; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_17007 = 4'h9 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_trigger_backendHit_0 :
    _GEN_14863; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_17008 = 4'ha == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_trigger_backendHit_0 :
    _GEN_14864; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_17009 = 4'hb == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_trigger_backendHit_0 :
    _GEN_14865; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_17010 = 4'hc == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_trigger_backendHit_0 :
    _GEN_14866; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_17011 = 4'hd == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_trigger_backendHit_0 :
    _GEN_14867; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_17012 = 4'he == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_trigger_backendHit_0 :
    _GEN_14868; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_17013 = 4'hf == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_trigger_backendHit_0 :
    _GEN_14869; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_17014 = 4'h0 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_trigger_backendHit_1 :
    _GEN_14870; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_17015 = 4'h1 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_trigger_backendHit_1 :
    _GEN_14871; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_17016 = 4'h2 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_trigger_backendHit_1 :
    _GEN_14872; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_17017 = 4'h3 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_trigger_backendHit_1 :
    _GEN_14873; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_17018 = 4'h4 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_trigger_backendHit_1 :
    _GEN_14874; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_17019 = 4'h5 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_trigger_backendHit_1 :
    _GEN_14875; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_17020 = 4'h6 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_trigger_backendHit_1 :
    _GEN_14876; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_17021 = 4'h7 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_trigger_backendHit_1 :
    _GEN_14877; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_17022 = 4'h8 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_trigger_backendHit_1 :
    _GEN_14878; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_17023 = 4'h9 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_trigger_backendHit_1 :
    _GEN_14879; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_17024 = 4'ha == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_trigger_backendHit_1 :
    _GEN_14880; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_17025 = 4'hb == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_trigger_backendHit_1 :
    _GEN_14881; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_17026 = 4'hc == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_trigger_backendHit_1 :
    _GEN_14882; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_17027 = 4'hd == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_trigger_backendHit_1 :
    _GEN_14883; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_17028 = 4'he == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_trigger_backendHit_1 :
    _GEN_14884; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_17029 = 4'hf == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_trigger_backendHit_1 :
    _GEN_14885; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_17062 = 4'h0 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_trigger_backendHit_4 :
    _GEN_14918; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_17063 = 4'h1 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_trigger_backendHit_4 :
    _GEN_14919; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_17064 = 4'h2 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_trigger_backendHit_4 :
    _GEN_14920; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_17065 = 4'h3 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_trigger_backendHit_4 :
    _GEN_14921; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_17066 = 4'h4 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_trigger_backendHit_4 :
    _GEN_14922; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_17067 = 4'h5 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_trigger_backendHit_4 :
    _GEN_14923; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_17068 = 4'h6 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_trigger_backendHit_4 :
    _GEN_14924; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_17069 = 4'h7 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_trigger_backendHit_4 :
    _GEN_14925; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_17070 = 4'h8 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_trigger_backendHit_4 :
    _GEN_14926; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_17071 = 4'h9 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_trigger_backendHit_4 :
    _GEN_14927; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_17072 = 4'ha == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_trigger_backendHit_4 :
    _GEN_14928; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_17073 = 4'hb == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_trigger_backendHit_4 :
    _GEN_14929; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_17074 = 4'hc == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_trigger_backendHit_4 :
    _GEN_14930; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_17075 = 4'hd == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_trigger_backendHit_4 :
    _GEN_14931; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_17076 = 4'he == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_trigger_backendHit_4 :
    _GEN_14932; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_17077 = 4'hf == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_cf_trigger_backendHit_4 :
    _GEN_14933; // @[LoadQueueFlag.scala 313:{31,31}]
  wire  _GEN_17462 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_16710 : _GEN_14566; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17463 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_16711 : _GEN_14567; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17464 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_16712 : _GEN_14568; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17465 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_16713 : _GEN_14569; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17466 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_16714 : _GEN_14570; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17467 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_16715 : _GEN_14571; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17468 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_16716 : _GEN_14572; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17469 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_16717 : _GEN_14573; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17470 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_16718 : _GEN_14574; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17471 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_16719 : _GEN_14575; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17472 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_16720 : _GEN_14576; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17473 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_16721 : _GEN_14577; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17474 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_16722 : _GEN_14578; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17475 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_16723 : _GEN_14579; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17476 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_16724 : _GEN_14580; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17477 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_16725 : _GEN_14581; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17478 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_16726 : _GEN_14582; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17479 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_16727 : _GEN_14583; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17480 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_16728 : _GEN_14584; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17481 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_16729 : _GEN_14585; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17482 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_16730 : _GEN_14586; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17483 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_16731 : _GEN_14587; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17484 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_16732 : _GEN_14588; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17485 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_16733 : _GEN_14589; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17486 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_16734 : _GEN_14590; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17487 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_16735 : _GEN_14591; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17488 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_16736 : _GEN_14592; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17489 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_16737 : _GEN_14593; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17490 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_16738 : _GEN_14594; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17491 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_16739 : _GEN_14595; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17492 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_16740 : _GEN_14596; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17493 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_16741 : _GEN_14597; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17606 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_16854 : _GEN_14710; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17607 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_16855 : _GEN_14711; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17608 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_16856 : _GEN_14712; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17609 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_16857 : _GEN_14713; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17610 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_16858 : _GEN_14714; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17611 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_16859 : _GEN_14715; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17612 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_16860 : _GEN_14716; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17613 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_16861 : _GEN_14717; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17614 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_16862 : _GEN_14718; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17615 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_16863 : _GEN_14719; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17616 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_16864 : _GEN_14720; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17617 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_16865 : _GEN_14721; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17618 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_16866 : _GEN_14722; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17619 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_16867 : _GEN_14723; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17620 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_16868 : _GEN_14724; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17621 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_16869 : _GEN_14725; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17734 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_16982 : _GEN_14838; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17735 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_16983 : _GEN_14839; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17736 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_16984 : _GEN_14840; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17737 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_16985 : _GEN_14841; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17738 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_16986 : _GEN_14842; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17739 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_16987 : _GEN_14843; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17740 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_16988 : _GEN_14844; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17741 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_16989 : _GEN_14845; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17742 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_16990 : _GEN_14846; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17743 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_16991 : _GEN_14847; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17744 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_16992 : _GEN_14848; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17745 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_16993 : _GEN_14849; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17746 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_16994 : _GEN_14850; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17747 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_16995 : _GEN_14851; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17748 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_16996 : _GEN_14852; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17749 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_16997 : _GEN_14853; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17750 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_16998 : _GEN_14854; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17751 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_16999 : _GEN_14855; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17752 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_17000 : _GEN_14856; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17753 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_17001 : _GEN_14857; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17754 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_17002 : _GEN_14858; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17755 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_17003 : _GEN_14859; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17756 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_17004 : _GEN_14860; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17757 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_17005 : _GEN_14861; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17758 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_17006 : _GEN_14862; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17759 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_17007 : _GEN_14863; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17760 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_17008 : _GEN_14864; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17761 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_17009 : _GEN_14865; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17762 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_17010 : _GEN_14866; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17763 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_17011 : _GEN_14867; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17764 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_17012 : _GEN_14868; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17765 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_17013 : _GEN_14869; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17766 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_17014 : _GEN_14870; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17767 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_17015 : _GEN_14871; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17768 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_17016 : _GEN_14872; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17769 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_17017 : _GEN_14873; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17770 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_17018 : _GEN_14874; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17771 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_17019 : _GEN_14875; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17772 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_17020 : _GEN_14876; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17773 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_17021 : _GEN_14877; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17774 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_17022 : _GEN_14878; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17775 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_17023 : _GEN_14879; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17776 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_17024 : _GEN_14880; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17777 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_17025 : _GEN_14881; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17778 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_17026 : _GEN_14882; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17779 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_17027 : _GEN_14883; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17780 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_17028 : _GEN_14884; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17781 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_17029 : _GEN_14885; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17814 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_17062 : _GEN_14918; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17815 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_17063 : _GEN_14919; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17816 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_17064 : _GEN_14920; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17817 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_17065 : _GEN_14921; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17818 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_17066 : _GEN_14922; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17819 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_17067 : _GEN_14923; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17820 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_17068 : _GEN_14924; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17821 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_17069 : _GEN_14925; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17822 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_17070 : _GEN_14926; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17823 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_17071 : _GEN_14927; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17824 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_17072 : _GEN_14928; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17825 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_17073 : _GEN_14929; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17826 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_17074 : _GEN_14930; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17827 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_17075 : _GEN_14931; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17828 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_17076 : _GEN_14932; // @[LoadQueueFlag.scala 312:50]
  wire  _GEN_17829 = io_loadIn_0_bits_lqDataWenDup_2 ? _GEN_17077 : _GEN_14933; // @[LoadQueueFlag.scala 312:50]
  wire [6:0] _GEN_18246 = 4'h0 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_ctrl_fuOpType : _GEN_15350; // @[LoadQueueFlag.scala 316:{33,33}]
  wire [6:0] _GEN_18247 = 4'h1 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_ctrl_fuOpType : _GEN_15351; // @[LoadQueueFlag.scala 316:{33,33}]
  wire [6:0] _GEN_18248 = 4'h2 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_ctrl_fuOpType : _GEN_15352; // @[LoadQueueFlag.scala 316:{33,33}]
  wire [6:0] _GEN_18249 = 4'h3 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_ctrl_fuOpType : _GEN_15353; // @[LoadQueueFlag.scala 316:{33,33}]
  wire [6:0] _GEN_18250 = 4'h4 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_ctrl_fuOpType : _GEN_15354; // @[LoadQueueFlag.scala 316:{33,33}]
  wire [6:0] _GEN_18251 = 4'h5 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_ctrl_fuOpType : _GEN_15355; // @[LoadQueueFlag.scala 316:{33,33}]
  wire [6:0] _GEN_18252 = 4'h6 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_ctrl_fuOpType : _GEN_15356; // @[LoadQueueFlag.scala 316:{33,33}]
  wire [6:0] _GEN_18253 = 4'h7 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_ctrl_fuOpType : _GEN_15357; // @[LoadQueueFlag.scala 316:{33,33}]
  wire [6:0] _GEN_18254 = 4'h8 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_ctrl_fuOpType : _GEN_15358; // @[LoadQueueFlag.scala 316:{33,33}]
  wire [6:0] _GEN_18255 = 4'h9 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_ctrl_fuOpType : _GEN_15359; // @[LoadQueueFlag.scala 316:{33,33}]
  wire [6:0] _GEN_18256 = 4'ha == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_ctrl_fuOpType : _GEN_15360; // @[LoadQueueFlag.scala 316:{33,33}]
  wire [6:0] _GEN_18257 = 4'hb == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_ctrl_fuOpType : _GEN_15361; // @[LoadQueueFlag.scala 316:{33,33}]
  wire [6:0] _GEN_18258 = 4'hc == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_ctrl_fuOpType : _GEN_15362; // @[LoadQueueFlag.scala 316:{33,33}]
  wire [6:0] _GEN_18259 = 4'hd == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_ctrl_fuOpType : _GEN_15363; // @[LoadQueueFlag.scala 316:{33,33}]
  wire [6:0] _GEN_18260 = 4'he == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_ctrl_fuOpType : _GEN_15364; // @[LoadQueueFlag.scala 316:{33,33}]
  wire [6:0] _GEN_18261 = 4'hf == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_ctrl_fuOpType : _GEN_15365; // @[LoadQueueFlag.scala 316:{33,33}]
  wire  _GEN_18262 = 4'h0 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_ctrl_rfWen : _GEN_15366; // @[LoadQueueFlag.scala 316:{33,33}]
  wire  _GEN_18263 = 4'h1 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_ctrl_rfWen : _GEN_15367; // @[LoadQueueFlag.scala 316:{33,33}]
  wire  _GEN_18264 = 4'h2 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_ctrl_rfWen : _GEN_15368; // @[LoadQueueFlag.scala 316:{33,33}]
  wire  _GEN_18265 = 4'h3 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_ctrl_rfWen : _GEN_15369; // @[LoadQueueFlag.scala 316:{33,33}]
  wire  _GEN_18266 = 4'h4 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_ctrl_rfWen : _GEN_15370; // @[LoadQueueFlag.scala 316:{33,33}]
  wire  _GEN_18267 = 4'h5 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_ctrl_rfWen : _GEN_15371; // @[LoadQueueFlag.scala 316:{33,33}]
  wire  _GEN_18268 = 4'h6 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_ctrl_rfWen : _GEN_15372; // @[LoadQueueFlag.scala 316:{33,33}]
  wire  _GEN_18269 = 4'h7 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_ctrl_rfWen : _GEN_15373; // @[LoadQueueFlag.scala 316:{33,33}]
  wire  _GEN_18270 = 4'h8 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_ctrl_rfWen : _GEN_15374; // @[LoadQueueFlag.scala 316:{33,33}]
  wire  _GEN_18271 = 4'h9 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_ctrl_rfWen : _GEN_15375; // @[LoadQueueFlag.scala 316:{33,33}]
  wire  _GEN_18272 = 4'ha == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_ctrl_rfWen : _GEN_15376; // @[LoadQueueFlag.scala 316:{33,33}]
  wire  _GEN_18273 = 4'hb == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_ctrl_rfWen : _GEN_15377; // @[LoadQueueFlag.scala 316:{33,33}]
  wire  _GEN_18274 = 4'hc == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_ctrl_rfWen : _GEN_15378; // @[LoadQueueFlag.scala 316:{33,33}]
  wire  _GEN_18275 = 4'hd == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_ctrl_rfWen : _GEN_15379; // @[LoadQueueFlag.scala 316:{33,33}]
  wire  _GEN_18276 = 4'he == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_ctrl_rfWen : _GEN_15380; // @[LoadQueueFlag.scala 316:{33,33}]
  wire  _GEN_18277 = 4'hf == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_ctrl_rfWen : _GEN_15381; // @[LoadQueueFlag.scala 316:{33,33}]
  wire  _GEN_18278 = 4'h0 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_ctrl_fpWen : _GEN_15382; // @[LoadQueueFlag.scala 316:{33,33}]
  wire  _GEN_18279 = 4'h1 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_ctrl_fpWen : _GEN_15383; // @[LoadQueueFlag.scala 316:{33,33}]
  wire  _GEN_18280 = 4'h2 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_ctrl_fpWen : _GEN_15384; // @[LoadQueueFlag.scala 316:{33,33}]
  wire  _GEN_18281 = 4'h3 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_ctrl_fpWen : _GEN_15385; // @[LoadQueueFlag.scala 316:{33,33}]
  wire  _GEN_18282 = 4'h4 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_ctrl_fpWen : _GEN_15386; // @[LoadQueueFlag.scala 316:{33,33}]
  wire  _GEN_18283 = 4'h5 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_ctrl_fpWen : _GEN_15387; // @[LoadQueueFlag.scala 316:{33,33}]
  wire  _GEN_18284 = 4'h6 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_ctrl_fpWen : _GEN_15388; // @[LoadQueueFlag.scala 316:{33,33}]
  wire  _GEN_18285 = 4'h7 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_ctrl_fpWen : _GEN_15389; // @[LoadQueueFlag.scala 316:{33,33}]
  wire  _GEN_18286 = 4'h8 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_ctrl_fpWen : _GEN_15390; // @[LoadQueueFlag.scala 316:{33,33}]
  wire  _GEN_18287 = 4'h9 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_ctrl_fpWen : _GEN_15391; // @[LoadQueueFlag.scala 316:{33,33}]
  wire  _GEN_18288 = 4'ha == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_ctrl_fpWen : _GEN_15392; // @[LoadQueueFlag.scala 316:{33,33}]
  wire  _GEN_18289 = 4'hb == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_ctrl_fpWen : _GEN_15393; // @[LoadQueueFlag.scala 316:{33,33}]
  wire  _GEN_18290 = 4'hc == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_ctrl_fpWen : _GEN_15394; // @[LoadQueueFlag.scala 316:{33,33}]
  wire  _GEN_18291 = 4'hd == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_ctrl_fpWen : _GEN_15395; // @[LoadQueueFlag.scala 316:{33,33}]
  wire  _GEN_18292 = 4'he == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_ctrl_fpWen : _GEN_15396; // @[LoadQueueFlag.scala 316:{33,33}]
  wire  _GEN_18293 = 4'hf == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_ctrl_fpWen : _GEN_15397; // @[LoadQueueFlag.scala 316:{33,33}]
  wire  _GEN_18342 = 4'h0 == io_loadIn_0_bits_uop_lqIdx_value ? 1'h0 : _GEN_15446; // @[LoadQueueFlag.scala 316:{33,33}]
  wire  _GEN_18343 = 4'h1 == io_loadIn_0_bits_uop_lqIdx_value ? 1'h0 : _GEN_15447; // @[LoadQueueFlag.scala 316:{33,33}]
  wire  _GEN_18344 = 4'h2 == io_loadIn_0_bits_uop_lqIdx_value ? 1'h0 : _GEN_15448; // @[LoadQueueFlag.scala 316:{33,33}]
  wire  _GEN_18345 = 4'h3 == io_loadIn_0_bits_uop_lqIdx_value ? 1'h0 : _GEN_15449; // @[LoadQueueFlag.scala 316:{33,33}]
  wire  _GEN_18346 = 4'h4 == io_loadIn_0_bits_uop_lqIdx_value ? 1'h0 : _GEN_15450; // @[LoadQueueFlag.scala 316:{33,33}]
  wire  _GEN_18347 = 4'h5 == io_loadIn_0_bits_uop_lqIdx_value ? 1'h0 : _GEN_15451; // @[LoadQueueFlag.scala 316:{33,33}]
  wire  _GEN_18348 = 4'h6 == io_loadIn_0_bits_uop_lqIdx_value ? 1'h0 : _GEN_15452; // @[LoadQueueFlag.scala 316:{33,33}]
  wire  _GEN_18349 = 4'h7 == io_loadIn_0_bits_uop_lqIdx_value ? 1'h0 : _GEN_15453; // @[LoadQueueFlag.scala 316:{33,33}]
  wire  _GEN_18350 = 4'h8 == io_loadIn_0_bits_uop_lqIdx_value ? 1'h0 : _GEN_15454; // @[LoadQueueFlag.scala 316:{33,33}]
  wire  _GEN_18351 = 4'h9 == io_loadIn_0_bits_uop_lqIdx_value ? 1'h0 : _GEN_15455; // @[LoadQueueFlag.scala 316:{33,33}]
  wire  _GEN_18352 = 4'ha == io_loadIn_0_bits_uop_lqIdx_value ? 1'h0 : _GEN_15456; // @[LoadQueueFlag.scala 316:{33,33}]
  wire  _GEN_18353 = 4'hb == io_loadIn_0_bits_uop_lqIdx_value ? 1'h0 : _GEN_15457; // @[LoadQueueFlag.scala 316:{33,33}]
  wire  _GEN_18354 = 4'hc == io_loadIn_0_bits_uop_lqIdx_value ? 1'h0 : _GEN_15458; // @[LoadQueueFlag.scala 316:{33,33}]
  wire  _GEN_18355 = 4'hd == io_loadIn_0_bits_uop_lqIdx_value ? 1'h0 : _GEN_15459; // @[LoadQueueFlag.scala 316:{33,33}]
  wire  _GEN_18356 = 4'he == io_loadIn_0_bits_uop_lqIdx_value ? 1'h0 : _GEN_15460; // @[LoadQueueFlag.scala 316:{33,33}]
  wire  _GEN_18357 = 4'hf == io_loadIn_0_bits_uop_lqIdx_value ? 1'h0 : _GEN_15461; // @[LoadQueueFlag.scala 316:{33,33}]
  wire  _GEN_18662 = 4'h0 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_ctrl_replayInst : _GEN_15766; // @[LoadQueueFlag.scala 316:{33,33}]
  wire  _GEN_18663 = 4'h1 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_ctrl_replayInst : _GEN_15767; // @[LoadQueueFlag.scala 316:{33,33}]
  wire  _GEN_18664 = 4'h2 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_ctrl_replayInst : _GEN_15768; // @[LoadQueueFlag.scala 316:{33,33}]
  wire  _GEN_18665 = 4'h3 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_ctrl_replayInst : _GEN_15769; // @[LoadQueueFlag.scala 316:{33,33}]
  wire  _GEN_18666 = 4'h4 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_ctrl_replayInst : _GEN_15770; // @[LoadQueueFlag.scala 316:{33,33}]
  wire  _GEN_18667 = 4'h5 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_ctrl_replayInst : _GEN_15771; // @[LoadQueueFlag.scala 316:{33,33}]
  wire  _GEN_18668 = 4'h6 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_ctrl_replayInst : _GEN_15772; // @[LoadQueueFlag.scala 316:{33,33}]
  wire  _GEN_18669 = 4'h7 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_ctrl_replayInst : _GEN_15773; // @[LoadQueueFlag.scala 316:{33,33}]
  wire  _GEN_18670 = 4'h8 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_ctrl_replayInst : _GEN_15774; // @[LoadQueueFlag.scala 316:{33,33}]
  wire  _GEN_18671 = 4'h9 == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_ctrl_replayInst : _GEN_15775; // @[LoadQueueFlag.scala 316:{33,33}]
  wire  _GEN_18672 = 4'ha == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_ctrl_replayInst : _GEN_15776; // @[LoadQueueFlag.scala 316:{33,33}]
  wire  _GEN_18673 = 4'hb == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_ctrl_replayInst : _GEN_15777; // @[LoadQueueFlag.scala 316:{33,33}]
  wire  _GEN_18674 = 4'hc == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_ctrl_replayInst : _GEN_15778; // @[LoadQueueFlag.scala 316:{33,33}]
  wire  _GEN_18675 = 4'hd == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_ctrl_replayInst : _GEN_15779; // @[LoadQueueFlag.scala 316:{33,33}]
  wire  _GEN_18676 = 4'he == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_ctrl_replayInst : _GEN_15780; // @[LoadQueueFlag.scala 316:{33,33}]
  wire  _GEN_18677 = 4'hf == io_loadIn_0_bits_uop_lqIdx_value ? io_loadIn_0_bits_uop_ctrl_replayInst : _GEN_15781; // @[LoadQueueFlag.scala 316:{33,33}]
  wire [6:0] _GEN_18822 = io_loadIn_0_bits_lqDataWenDup_3 ? _GEN_18246 : _GEN_15350; // @[LoadQueueFlag.scala 315:50]
  wire [6:0] _GEN_18823 = io_loadIn_0_bits_lqDataWenDup_3 ? _GEN_18247 : _GEN_15351; // @[LoadQueueFlag.scala 315:50]
  wire [6:0] _GEN_18824 = io_loadIn_0_bits_lqDataWenDup_3 ? _GEN_18248 : _GEN_15352; // @[LoadQueueFlag.scala 315:50]
  wire [6:0] _GEN_18825 = io_loadIn_0_bits_lqDataWenDup_3 ? _GEN_18249 : _GEN_15353; // @[LoadQueueFlag.scala 315:50]
  wire [6:0] _GEN_18826 = io_loadIn_0_bits_lqDataWenDup_3 ? _GEN_18250 : _GEN_15354; // @[LoadQueueFlag.scala 315:50]
  wire [6:0] _GEN_18827 = io_loadIn_0_bits_lqDataWenDup_3 ? _GEN_18251 : _GEN_15355; // @[LoadQueueFlag.scala 315:50]
  wire [6:0] _GEN_18828 = io_loadIn_0_bits_lqDataWenDup_3 ? _GEN_18252 : _GEN_15356; // @[LoadQueueFlag.scala 315:50]
  wire [6:0] _GEN_18829 = io_loadIn_0_bits_lqDataWenDup_3 ? _GEN_18253 : _GEN_15357; // @[LoadQueueFlag.scala 315:50]
  wire [6:0] _GEN_18830 = io_loadIn_0_bits_lqDataWenDup_3 ? _GEN_18254 : _GEN_15358; // @[LoadQueueFlag.scala 315:50]
  wire [6:0] _GEN_18831 = io_loadIn_0_bits_lqDataWenDup_3 ? _GEN_18255 : _GEN_15359; // @[LoadQueueFlag.scala 315:50]
  wire [6:0] _GEN_18832 = io_loadIn_0_bits_lqDataWenDup_3 ? _GEN_18256 : _GEN_15360; // @[LoadQueueFlag.scala 315:50]
  wire [6:0] _GEN_18833 = io_loadIn_0_bits_lqDataWenDup_3 ? _GEN_18257 : _GEN_15361; // @[LoadQueueFlag.scala 315:50]
  wire [6:0] _GEN_18834 = io_loadIn_0_bits_lqDataWenDup_3 ? _GEN_18258 : _GEN_15362; // @[LoadQueueFlag.scala 315:50]
  wire [6:0] _GEN_18835 = io_loadIn_0_bits_lqDataWenDup_3 ? _GEN_18259 : _GEN_15363; // @[LoadQueueFlag.scala 315:50]
  wire [6:0] _GEN_18836 = io_loadIn_0_bits_lqDataWenDup_3 ? _GEN_18260 : _GEN_15364; // @[LoadQueueFlag.scala 315:50]
  wire [6:0] _GEN_18837 = io_loadIn_0_bits_lqDataWenDup_3 ? _GEN_18261 : _GEN_15365; // @[LoadQueueFlag.scala 315:50]
  wire  _GEN_18838 = io_loadIn_0_bits_lqDataWenDup_3 ? _GEN_18262 : _GEN_15366; // @[LoadQueueFlag.scala 315:50]
  wire  _GEN_18839 = io_loadIn_0_bits_lqDataWenDup_3 ? _GEN_18263 : _GEN_15367; // @[LoadQueueFlag.scala 315:50]
  wire  _GEN_18840 = io_loadIn_0_bits_lqDataWenDup_3 ? _GEN_18264 : _GEN_15368; // @[LoadQueueFlag.scala 315:50]
  wire  _GEN_18841 = io_loadIn_0_bits_lqDataWenDup_3 ? _GEN_18265 : _GEN_15369; // @[LoadQueueFlag.scala 315:50]
  wire  _GEN_18842 = io_loadIn_0_bits_lqDataWenDup_3 ? _GEN_18266 : _GEN_15370; // @[LoadQueueFlag.scala 315:50]
  wire  _GEN_18843 = io_loadIn_0_bits_lqDataWenDup_3 ? _GEN_18267 : _GEN_15371; // @[LoadQueueFlag.scala 315:50]
  wire  _GEN_18844 = io_loadIn_0_bits_lqDataWenDup_3 ? _GEN_18268 : _GEN_15372; // @[LoadQueueFlag.scala 315:50]
  wire  _GEN_18845 = io_loadIn_0_bits_lqDataWenDup_3 ? _GEN_18269 : _GEN_15373; // @[LoadQueueFlag.scala 315:50]
  wire  _GEN_18846 = io_loadIn_0_bits_lqDataWenDup_3 ? _GEN_18270 : _GEN_15374; // @[LoadQueueFlag.scala 315:50]
  wire  _GEN_18847 = io_loadIn_0_bits_lqDataWenDup_3 ? _GEN_18271 : _GEN_15375; // @[LoadQueueFlag.scala 315:50]
  wire  _GEN_18848 = io_loadIn_0_bits_lqDataWenDup_3 ? _GEN_18272 : _GEN_15376; // @[LoadQueueFlag.scala 315:50]
  wire  _GEN_18849 = io_loadIn_0_bits_lqDataWenDup_3 ? _GEN_18273 : _GEN_15377; // @[LoadQueueFlag.scala 315:50]
  wire  _GEN_18850 = io_loadIn_0_bits_lqDataWenDup_3 ? _GEN_18274 : _GEN_15378; // @[LoadQueueFlag.scala 315:50]
  wire  _GEN_18851 = io_loadIn_0_bits_lqDataWenDup_3 ? _GEN_18275 : _GEN_15379; // @[LoadQueueFlag.scala 315:50]
  wire  _GEN_18852 = io_loadIn_0_bits_lqDataWenDup_3 ? _GEN_18276 : _GEN_15380; // @[LoadQueueFlag.scala 315:50]
  wire  _GEN_18853 = io_loadIn_0_bits_lqDataWenDup_3 ? _GEN_18277 : _GEN_15381; // @[LoadQueueFlag.scala 315:50]
  wire  _GEN_18854 = io_loadIn_0_bits_lqDataWenDup_3 ? _GEN_18278 : _GEN_15382; // @[LoadQueueFlag.scala 315:50]
  wire  _GEN_18855 = io_loadIn_0_bits_lqDataWenDup_3 ? _GEN_18279 : _GEN_15383; // @[LoadQueueFlag.scala 315:50]
  wire  _GEN_18856 = io_loadIn_0_bits_lqDataWenDup_3 ? _GEN_18280 : _GEN_15384; // @[LoadQueueFlag.scala 315:50]
  wire  _GEN_18857 = io_loadIn_0_bits_lqDataWenDup_3 ? _GEN_18281 : _GEN_15385; // @[LoadQueueFlag.scala 315:50]
  wire  _GEN_18858 = io_loadIn_0_bits_lqDataWenDup_3 ? _GEN_18282 : _GEN_15386; // @[LoadQueueFlag.scala 315:50]
  wire  _GEN_18859 = io_loadIn_0_bits_lqDataWenDup_3 ? _GEN_18283 : _GEN_15387; // @[LoadQueueFlag.scala 315:50]
  wire  _GEN_18860 = io_loadIn_0_bits_lqDataWenDup_3 ? _GEN_18284 : _GEN_15388; // @[LoadQueueFlag.scala 315:50]
  wire  _GEN_18861 = io_loadIn_0_bits_lqDataWenDup_3 ? _GEN_18285 : _GEN_15389; // @[LoadQueueFlag.scala 315:50]
  wire  _GEN_18862 = io_loadIn_0_bits_lqDataWenDup_3 ? _GEN_18286 : _GEN_15390; // @[LoadQueueFlag.scala 315:50]
  wire  _GEN_18863 = io_loadIn_0_bits_lqDataWenDup_3 ? _GEN_18287 : _GEN_15391; // @[LoadQueueFlag.scala 315:50]
  wire  _GEN_18864 = io_loadIn_0_bits_lqDataWenDup_3 ? _GEN_18288 : _GEN_15392; // @[LoadQueueFlag.scala 315:50]
  wire  _GEN_18865 = io_loadIn_0_bits_lqDataWenDup_3 ? _GEN_18289 : _GEN_15393; // @[LoadQueueFlag.scala 315:50]
  wire  _GEN_18866 = io_loadIn_0_bits_lqDataWenDup_3 ? _GEN_18290 : _GEN_15394; // @[LoadQueueFlag.scala 315:50]
  wire  _GEN_18867 = io_loadIn_0_bits_lqDataWenDup_3 ? _GEN_18291 : _GEN_15395; // @[LoadQueueFlag.scala 315:50]
  wire  _GEN_18868 = io_loadIn_0_bits_lqDataWenDup_3 ? _GEN_18292 : _GEN_15396; // @[LoadQueueFlag.scala 315:50]
  wire  _GEN_18869 = io_loadIn_0_bits_lqDataWenDup_3 ? _GEN_18293 : _GEN_15397; // @[LoadQueueFlag.scala 315:50]
  wire  _GEN_18918 = io_loadIn_0_bits_lqDataWenDup_3 ? _GEN_18342 : _GEN_15446; // @[LoadQueueFlag.scala 315:50]
  wire  _GEN_18919 = io_loadIn_0_bits_lqDataWenDup_3 ? _GEN_18343 : _GEN_15447; // @[LoadQueueFlag.scala 315:50]
  wire  _GEN_18920 = io_loadIn_0_bits_lqDataWenDup_3 ? _GEN_18344 : _GEN_15448; // @[LoadQueueFlag.scala 315:50]
  wire  _GEN_18921 = io_loadIn_0_bits_lqDataWenDup_3 ? _GEN_18345 : _GEN_15449; // @[LoadQueueFlag.scala 315:50]
  wire  _GEN_18922 = io_loadIn_0_bits_lqDataWenDup_3 ? _GEN_18346 : _GEN_15450; // @[LoadQueueFlag.scala 315:50]
  wire  _GEN_18923 = io_loadIn_0_bits_lqDataWenDup_3 ? _GEN_18347 : _GEN_15451; // @[LoadQueueFlag.scala 315:50]
  wire  _GEN_18924 = io_loadIn_0_bits_lqDataWenDup_3 ? _GEN_18348 : _GEN_15452; // @[LoadQueueFlag.scala 315:50]
  wire  _GEN_18925 = io_loadIn_0_bits_lqDataWenDup_3 ? _GEN_18349 : _GEN_15453; // @[LoadQueueFlag.scala 315:50]
  wire  _GEN_18926 = io_loadIn_0_bits_lqDataWenDup_3 ? _GEN_18350 : _GEN_15454; // @[LoadQueueFlag.scala 315:50]
  wire  _GEN_18927 = io_loadIn_0_bits_lqDataWenDup_3 ? _GEN_18351 : _GEN_15455; // @[LoadQueueFlag.scala 315:50]
  wire  _GEN_18928 = io_loadIn_0_bits_lqDataWenDup_3 ? _GEN_18352 : _GEN_15456; // @[LoadQueueFlag.scala 315:50]
  wire  _GEN_18929 = io_loadIn_0_bits_lqDataWenDup_3 ? _GEN_18353 : _GEN_15457; // @[LoadQueueFlag.scala 315:50]
  wire  _GEN_18930 = io_loadIn_0_bits_lqDataWenDup_3 ? _GEN_18354 : _GEN_15458; // @[LoadQueueFlag.scala 315:50]
  wire  _GEN_18931 = io_loadIn_0_bits_lqDataWenDup_3 ? _GEN_18355 : _GEN_15459; // @[LoadQueueFlag.scala 315:50]
  wire  _GEN_18932 = io_loadIn_0_bits_lqDataWenDup_3 ? _GEN_18356 : _GEN_15460; // @[LoadQueueFlag.scala 315:50]
  wire  _GEN_18933 = io_loadIn_0_bits_lqDataWenDup_3 ? _GEN_18357 : _GEN_15461; // @[LoadQueueFlag.scala 315:50]
  wire  _GEN_19238 = io_loadIn_0_bits_lqDataWenDup_3 ? _GEN_18662 : _GEN_15766; // @[LoadQueueFlag.scala 315:50]
  wire  _GEN_19239 = io_loadIn_0_bits_lqDataWenDup_3 ? _GEN_18663 : _GEN_15767; // @[LoadQueueFlag.scala 315:50]
  wire  _GEN_19240 = io_loadIn_0_bits_lqDataWenDup_3 ? _GEN_18664 : _GEN_15768; // @[LoadQueueFlag.scala 315:50]
  wire  _GEN_19241 = io_loadIn_0_bits_lqDataWenDup_3 ? _GEN_18665 : _GEN_15769; // @[LoadQueueFlag.scala 315:50]
  wire  _GEN_19242 = io_loadIn_0_bits_lqDataWenDup_3 ? _GEN_18666 : _GEN_15770; // @[LoadQueueFlag.scala 315:50]
  wire  _GEN_19243 = io_loadIn_0_bits_lqDataWenDup_3 ? _GEN_18667 : _GEN_15771; // @[LoadQueueFlag.scala 315:50]
  wire  _GEN_19244 = io_loadIn_0_bits_lqDataWenDup_3 ? _GEN_18668 : _GEN_15772; // @[LoadQueueFlag.scala 315:50]
  wire  _GEN_19245 = io_loadIn_0_bits_lqDataWenDup_3 ? _GEN_18669 : _GEN_15773; // @[LoadQueueFlag.scala 315:50]
  wire  _GEN_19246 = io_loadIn_0_bits_lqDataWenDup_3 ? _GEN_18670 : _GEN_15774; // @[LoadQueueFlag.scala 315:50]
  wire  _GEN_19247 = io_loadIn_0_bits_lqDataWenDup_3 ? _GEN_18671 : _GEN_15775; // @[LoadQueueFlag.scala 315:50]
  wire  _GEN_19248 = io_loadIn_0_bits_lqDataWenDup_3 ? _GEN_18672 : _GEN_15776; // @[LoadQueueFlag.scala 315:50]
  wire  _GEN_19249 = io_loadIn_0_bits_lqDataWenDup_3 ? _GEN_18673 : _GEN_15777; // @[LoadQueueFlag.scala 315:50]
  wire  _GEN_19250 = io_loadIn_0_bits_lqDataWenDup_3 ? _GEN_18674 : _GEN_15778; // @[LoadQueueFlag.scala 315:50]
  wire  _GEN_19251 = io_loadIn_0_bits_lqDataWenDup_3 ? _GEN_18675 : _GEN_15779; // @[LoadQueueFlag.scala 315:50]
  wire  _GEN_19252 = io_loadIn_0_bits_lqDataWenDup_3 ? _GEN_18676 : _GEN_15780; // @[LoadQueueFlag.scala 315:50]
  wire  _GEN_19253 = io_loadIn_0_bits_lqDataWenDup_3 ? _GEN_18677 : _GEN_15781; // @[LoadQueueFlag.scala 315:50]
  wire  _GEN_19771 = _issued_T_1 ? _GEN_16502 : _GEN_16182; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19772 = _issued_T_1 ? _GEN_16503 : _GEN_16183; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19773 = _issued_T_1 ? _GEN_16504 : _GEN_16184; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19774 = _issued_T_1 ? _GEN_16505 : _GEN_16185; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19775 = _issued_T_1 ? _GEN_16506 : _GEN_16186; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19776 = _issued_T_1 ? _GEN_16507 : _GEN_16187; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19777 = _issued_T_1 ? _GEN_16508 : _GEN_16188; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19778 = _issued_T_1 ? _GEN_16509 : _GEN_16189; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19779 = _issued_T_1 ? _GEN_16510 : _GEN_16190; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19780 = _issued_T_1 ? _GEN_16511 : _GEN_16191; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19781 = _issued_T_1 ? _GEN_16512 : _GEN_16192; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19782 = _issued_T_1 ? _GEN_16513 : _GEN_16193; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19783 = _issued_T_1 ? _GEN_16514 : _GEN_16194; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19784 = _issued_T_1 ? _GEN_16515 : _GEN_16195; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19785 = _issued_T_1 ? _GEN_16516 : _GEN_16196; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19786 = _issued_T_1 ? _GEN_16517 : _GEN_16197; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19787 = _issued_T_1 ? _GEN_16518 : _GEN_16198; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19788 = _issued_T_1 ? _GEN_16519 : _GEN_16199; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19789 = _issued_T_1 ? _GEN_16520 : _GEN_16200; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19790 = _issued_T_1 ? _GEN_16521 : _GEN_16201; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19791 = _issued_T_1 ? _GEN_16522 : _GEN_16202; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19792 = _issued_T_1 ? _GEN_16523 : _GEN_16203; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19793 = _issued_T_1 ? _GEN_16524 : _GEN_16204; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19794 = _issued_T_1 ? _GEN_16525 : _GEN_16205; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19795 = _issued_T_1 ? _GEN_16526 : _GEN_16206; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19796 = _issued_T_1 ? _GEN_16527 : _GEN_16207; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19797 = _issued_T_1 ? _GEN_16528 : _GEN_16208; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19798 = _issued_T_1 ? _GEN_16529 : _GEN_16209; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19799 = _issued_T_1 ? _GEN_16530 : _GEN_16210; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19800 = _issued_T_1 ? _GEN_16531 : _GEN_16211; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19801 = _issued_T_1 ? _GEN_16532 : _GEN_16212; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19802 = _issued_T_1 ? _GEN_16533 : _GEN_16213; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19803 = _issued_T_1 ? _GEN_16534 : _GEN_16214; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19804 = _issued_T_1 ? _GEN_16535 : _GEN_16215; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19805 = _issued_T_1 ? _GEN_16536 : _GEN_16216; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19806 = _issued_T_1 ? _GEN_16537 : _GEN_16217; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19807 = _issued_T_1 ? _GEN_16538 : _GEN_16218; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19808 = _issued_T_1 ? _GEN_16539 : _GEN_16219; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19809 = _issued_T_1 ? _GEN_16540 : _GEN_16220; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19810 = _issued_T_1 ? _GEN_16541 : _GEN_16221; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19811 = _issued_T_1 ? _GEN_16542 : _GEN_16222; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19812 = _issued_T_1 ? _GEN_16543 : _GEN_16223; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19813 = _issued_T_1 ? _GEN_16544 : _GEN_16224; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19814 = _issued_T_1 ? _GEN_16545 : _GEN_16225; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19815 = _issued_T_1 ? _GEN_16546 : _GEN_16226; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19816 = _issued_T_1 ? _GEN_16547 : _GEN_16227; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19817 = _issued_T_1 ? _GEN_16548 : _GEN_16228; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19818 = _issued_T_1 ? _GEN_16549 : _GEN_16229; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19819 = _issued_T_1 ? _GEN_16550 : _GEN_16230; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19820 = _issued_T_1 ? _GEN_16551 : _GEN_16231; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19821 = _issued_T_1 ? _GEN_16552 : _GEN_16232; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19822 = _issued_T_1 ? _GEN_16553 : _GEN_16233; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19823 = _issued_T_1 ? _GEN_16554 : _GEN_16234; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19824 = _issued_T_1 ? _GEN_16555 : _GEN_16235; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19825 = _issued_T_1 ? _GEN_16556 : _GEN_16236; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19826 = _issued_T_1 ? _GEN_16557 : _GEN_16237; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19827 = _issued_T_1 ? _GEN_16558 : _GEN_16238; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19828 = _issued_T_1 ? _GEN_16559 : _GEN_16239; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19829 = _issued_T_1 ? _GEN_16560 : _GEN_16240; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19830 = _issued_T_1 ? _GEN_16561 : _GEN_16241; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19831 = _issued_T_1 ? _GEN_16562 : _GEN_16242; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19832 = _issued_T_1 ? _GEN_16563 : _GEN_16243; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19833 = _issued_T_1 ? _GEN_16564 : _GEN_16244; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19834 = _issued_T_1 ? _GEN_16565 : _GEN_16245; // @[LoadQueueFlag.scala 301:26]
  wire [5:0] _GEN_19835 = _issued_T_1 ? _GEN_16582 : _GEN_15878; // @[LoadQueueFlag.scala 301:26]
  wire [5:0] _GEN_19836 = _issued_T_1 ? _GEN_16583 : _GEN_15879; // @[LoadQueueFlag.scala 301:26]
  wire [5:0] _GEN_19837 = _issued_T_1 ? _GEN_16584 : _GEN_15880; // @[LoadQueueFlag.scala 301:26]
  wire [5:0] _GEN_19838 = _issued_T_1 ? _GEN_16585 : _GEN_15881; // @[LoadQueueFlag.scala 301:26]
  wire [5:0] _GEN_19839 = _issued_T_1 ? _GEN_16586 : _GEN_15882; // @[LoadQueueFlag.scala 301:26]
  wire [5:0] _GEN_19840 = _issued_T_1 ? _GEN_16587 : _GEN_15883; // @[LoadQueueFlag.scala 301:26]
  wire [5:0] _GEN_19841 = _issued_T_1 ? _GEN_16588 : _GEN_15884; // @[LoadQueueFlag.scala 301:26]
  wire [5:0] _GEN_19842 = _issued_T_1 ? _GEN_16589 : _GEN_15885; // @[LoadQueueFlag.scala 301:26]
  wire [5:0] _GEN_19843 = _issued_T_1 ? _GEN_16590 : _GEN_15886; // @[LoadQueueFlag.scala 301:26]
  wire [5:0] _GEN_19844 = _issued_T_1 ? _GEN_16591 : _GEN_15887; // @[LoadQueueFlag.scala 301:26]
  wire [5:0] _GEN_19845 = _issued_T_1 ? _GEN_16592 : _GEN_15888; // @[LoadQueueFlag.scala 301:26]
  wire [5:0] _GEN_19846 = _issued_T_1 ? _GEN_16593 : _GEN_15889; // @[LoadQueueFlag.scala 301:26]
  wire [5:0] _GEN_19847 = _issued_T_1 ? _GEN_16594 : _GEN_15890; // @[LoadQueueFlag.scala 301:26]
  wire [5:0] _GEN_19848 = _issued_T_1 ? _GEN_16595 : _GEN_15891; // @[LoadQueueFlag.scala 301:26]
  wire [5:0] _GEN_19849 = _issued_T_1 ? _GEN_16596 : _GEN_15892; // @[LoadQueueFlag.scala 301:26]
  wire [5:0] _GEN_19850 = _issued_T_1 ? _GEN_16597 : _GEN_15893; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19963 = _issued_T_1 ? _GEN_17462 : _GEN_14566; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19964 = _issued_T_1 ? _GEN_17463 : _GEN_14567; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19965 = _issued_T_1 ? _GEN_17464 : _GEN_14568; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19966 = _issued_T_1 ? _GEN_17465 : _GEN_14569; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19967 = _issued_T_1 ? _GEN_17466 : _GEN_14570; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19968 = _issued_T_1 ? _GEN_17467 : _GEN_14571; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19969 = _issued_T_1 ? _GEN_17468 : _GEN_14572; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19970 = _issued_T_1 ? _GEN_17469 : _GEN_14573; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19971 = _issued_T_1 ? _GEN_17470 : _GEN_14574; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19972 = _issued_T_1 ? _GEN_17471 : _GEN_14575; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19973 = _issued_T_1 ? _GEN_17472 : _GEN_14576; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19974 = _issued_T_1 ? _GEN_17473 : _GEN_14577; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19975 = _issued_T_1 ? _GEN_17474 : _GEN_14578; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19976 = _issued_T_1 ? _GEN_17475 : _GEN_14579; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19977 = _issued_T_1 ? _GEN_17476 : _GEN_14580; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19978 = _issued_T_1 ? _GEN_17477 : _GEN_14581; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19979 = _issued_T_1 ? _GEN_17478 : _GEN_14582; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19980 = _issued_T_1 ? _GEN_17479 : _GEN_14583; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19981 = _issued_T_1 ? _GEN_17480 : _GEN_14584; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19982 = _issued_T_1 ? _GEN_17481 : _GEN_14585; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19983 = _issued_T_1 ? _GEN_17482 : _GEN_14586; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19984 = _issued_T_1 ? _GEN_17483 : _GEN_14587; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19985 = _issued_T_1 ? _GEN_17484 : _GEN_14588; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19986 = _issued_T_1 ? _GEN_17485 : _GEN_14589; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19987 = _issued_T_1 ? _GEN_17486 : _GEN_14590; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19988 = _issued_T_1 ? _GEN_17487 : _GEN_14591; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19989 = _issued_T_1 ? _GEN_17488 : _GEN_14592; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19990 = _issued_T_1 ? _GEN_17489 : _GEN_14593; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19991 = _issued_T_1 ? _GEN_17490 : _GEN_14594; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19992 = _issued_T_1 ? _GEN_17491 : _GEN_14595; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19993 = _issued_T_1 ? _GEN_17492 : _GEN_14596; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_19994 = _issued_T_1 ? _GEN_17493 : _GEN_14597; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20107 = _issued_T_1 ? _GEN_17606 : _GEN_14710; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20108 = _issued_T_1 ? _GEN_17607 : _GEN_14711; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20109 = _issued_T_1 ? _GEN_17608 : _GEN_14712; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20110 = _issued_T_1 ? _GEN_17609 : _GEN_14713; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20111 = _issued_T_1 ? _GEN_17610 : _GEN_14714; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20112 = _issued_T_1 ? _GEN_17611 : _GEN_14715; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20113 = _issued_T_1 ? _GEN_17612 : _GEN_14716; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20114 = _issued_T_1 ? _GEN_17613 : _GEN_14717; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20115 = _issued_T_1 ? _GEN_17614 : _GEN_14718; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20116 = _issued_T_1 ? _GEN_17615 : _GEN_14719; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20117 = _issued_T_1 ? _GEN_17616 : _GEN_14720; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20118 = _issued_T_1 ? _GEN_17617 : _GEN_14721; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20119 = _issued_T_1 ? _GEN_17618 : _GEN_14722; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20120 = _issued_T_1 ? _GEN_17619 : _GEN_14723; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20121 = _issued_T_1 ? _GEN_17620 : _GEN_14724; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20122 = _issued_T_1 ? _GEN_17621 : _GEN_14725; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20235 = _issued_T_1 ? _GEN_17734 : _GEN_14838; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20236 = _issued_T_1 ? _GEN_17735 : _GEN_14839; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20237 = _issued_T_1 ? _GEN_17736 : _GEN_14840; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20238 = _issued_T_1 ? _GEN_17737 : _GEN_14841; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20239 = _issued_T_1 ? _GEN_17738 : _GEN_14842; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20240 = _issued_T_1 ? _GEN_17739 : _GEN_14843; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20241 = _issued_T_1 ? _GEN_17740 : _GEN_14844; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20242 = _issued_T_1 ? _GEN_17741 : _GEN_14845; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20243 = _issued_T_1 ? _GEN_17742 : _GEN_14846; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20244 = _issued_T_1 ? _GEN_17743 : _GEN_14847; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20245 = _issued_T_1 ? _GEN_17744 : _GEN_14848; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20246 = _issued_T_1 ? _GEN_17745 : _GEN_14849; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20247 = _issued_T_1 ? _GEN_17746 : _GEN_14850; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20248 = _issued_T_1 ? _GEN_17747 : _GEN_14851; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20249 = _issued_T_1 ? _GEN_17748 : _GEN_14852; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20250 = _issued_T_1 ? _GEN_17749 : _GEN_14853; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20251 = _issued_T_1 ? _GEN_17750 : _GEN_14854; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20252 = _issued_T_1 ? _GEN_17751 : _GEN_14855; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20253 = _issued_T_1 ? _GEN_17752 : _GEN_14856; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20254 = _issued_T_1 ? _GEN_17753 : _GEN_14857; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20255 = _issued_T_1 ? _GEN_17754 : _GEN_14858; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20256 = _issued_T_1 ? _GEN_17755 : _GEN_14859; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20257 = _issued_T_1 ? _GEN_17756 : _GEN_14860; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20258 = _issued_T_1 ? _GEN_17757 : _GEN_14861; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20259 = _issued_T_1 ? _GEN_17758 : _GEN_14862; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20260 = _issued_T_1 ? _GEN_17759 : _GEN_14863; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20261 = _issued_T_1 ? _GEN_17760 : _GEN_14864; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20262 = _issued_T_1 ? _GEN_17761 : _GEN_14865; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20263 = _issued_T_1 ? _GEN_17762 : _GEN_14866; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20264 = _issued_T_1 ? _GEN_17763 : _GEN_14867; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20265 = _issued_T_1 ? _GEN_17764 : _GEN_14868; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20266 = _issued_T_1 ? _GEN_17765 : _GEN_14869; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20267 = _issued_T_1 ? _GEN_17766 : _GEN_14870; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20268 = _issued_T_1 ? _GEN_17767 : _GEN_14871; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20269 = _issued_T_1 ? _GEN_17768 : _GEN_14872; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20270 = _issued_T_1 ? _GEN_17769 : _GEN_14873; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20271 = _issued_T_1 ? _GEN_17770 : _GEN_14874; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20272 = _issued_T_1 ? _GEN_17771 : _GEN_14875; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20273 = _issued_T_1 ? _GEN_17772 : _GEN_14876; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20274 = _issued_T_1 ? _GEN_17773 : _GEN_14877; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20275 = _issued_T_1 ? _GEN_17774 : _GEN_14878; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20276 = _issued_T_1 ? _GEN_17775 : _GEN_14879; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20277 = _issued_T_1 ? _GEN_17776 : _GEN_14880; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20278 = _issued_T_1 ? _GEN_17777 : _GEN_14881; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20279 = _issued_T_1 ? _GEN_17778 : _GEN_14882; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20280 = _issued_T_1 ? _GEN_17779 : _GEN_14883; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20281 = _issued_T_1 ? _GEN_17780 : _GEN_14884; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20282 = _issued_T_1 ? _GEN_17781 : _GEN_14885; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20315 = _issued_T_1 ? _GEN_17814 : _GEN_14918; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20316 = _issued_T_1 ? _GEN_17815 : _GEN_14919; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20317 = _issued_T_1 ? _GEN_17816 : _GEN_14920; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20318 = _issued_T_1 ? _GEN_17817 : _GEN_14921; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20319 = _issued_T_1 ? _GEN_17818 : _GEN_14922; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20320 = _issued_T_1 ? _GEN_17819 : _GEN_14923; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20321 = _issued_T_1 ? _GEN_17820 : _GEN_14924; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20322 = _issued_T_1 ? _GEN_17821 : _GEN_14925; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20323 = _issued_T_1 ? _GEN_17822 : _GEN_14926; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20324 = _issued_T_1 ? _GEN_17823 : _GEN_14927; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20325 = _issued_T_1 ? _GEN_17824 : _GEN_14928; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20326 = _issued_T_1 ? _GEN_17825 : _GEN_14929; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20327 = _issued_T_1 ? _GEN_17826 : _GEN_14930; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20328 = _issued_T_1 ? _GEN_17827 : _GEN_14931; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20329 = _issued_T_1 ? _GEN_17828 : _GEN_14932; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20330 = _issued_T_1 ? _GEN_17829 : _GEN_14933; // @[LoadQueueFlag.scala 301:26]
  wire [6:0] _GEN_20747 = _issued_T_1 ? _GEN_18822 : _GEN_15350; // @[LoadQueueFlag.scala 301:26]
  wire [6:0] _GEN_20748 = _issued_T_1 ? _GEN_18823 : _GEN_15351; // @[LoadQueueFlag.scala 301:26]
  wire [6:0] _GEN_20749 = _issued_T_1 ? _GEN_18824 : _GEN_15352; // @[LoadQueueFlag.scala 301:26]
  wire [6:0] _GEN_20750 = _issued_T_1 ? _GEN_18825 : _GEN_15353; // @[LoadQueueFlag.scala 301:26]
  wire [6:0] _GEN_20751 = _issued_T_1 ? _GEN_18826 : _GEN_15354; // @[LoadQueueFlag.scala 301:26]
  wire [6:0] _GEN_20752 = _issued_T_1 ? _GEN_18827 : _GEN_15355; // @[LoadQueueFlag.scala 301:26]
  wire [6:0] _GEN_20753 = _issued_T_1 ? _GEN_18828 : _GEN_15356; // @[LoadQueueFlag.scala 301:26]
  wire [6:0] _GEN_20754 = _issued_T_1 ? _GEN_18829 : _GEN_15357; // @[LoadQueueFlag.scala 301:26]
  wire [6:0] _GEN_20755 = _issued_T_1 ? _GEN_18830 : _GEN_15358; // @[LoadQueueFlag.scala 301:26]
  wire [6:0] _GEN_20756 = _issued_T_1 ? _GEN_18831 : _GEN_15359; // @[LoadQueueFlag.scala 301:26]
  wire [6:0] _GEN_20757 = _issued_T_1 ? _GEN_18832 : _GEN_15360; // @[LoadQueueFlag.scala 301:26]
  wire [6:0] _GEN_20758 = _issued_T_1 ? _GEN_18833 : _GEN_15361; // @[LoadQueueFlag.scala 301:26]
  wire [6:0] _GEN_20759 = _issued_T_1 ? _GEN_18834 : _GEN_15362; // @[LoadQueueFlag.scala 301:26]
  wire [6:0] _GEN_20760 = _issued_T_1 ? _GEN_18835 : _GEN_15363; // @[LoadQueueFlag.scala 301:26]
  wire [6:0] _GEN_20761 = _issued_T_1 ? _GEN_18836 : _GEN_15364; // @[LoadQueueFlag.scala 301:26]
  wire [6:0] _GEN_20762 = _issued_T_1 ? _GEN_18837 : _GEN_15365; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20763 = _issued_T_1 ? _GEN_18838 : _GEN_15366; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20764 = _issued_T_1 ? _GEN_18839 : _GEN_15367; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20765 = _issued_T_1 ? _GEN_18840 : _GEN_15368; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20766 = _issued_T_1 ? _GEN_18841 : _GEN_15369; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20767 = _issued_T_1 ? _GEN_18842 : _GEN_15370; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20768 = _issued_T_1 ? _GEN_18843 : _GEN_15371; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20769 = _issued_T_1 ? _GEN_18844 : _GEN_15372; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20770 = _issued_T_1 ? _GEN_18845 : _GEN_15373; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20771 = _issued_T_1 ? _GEN_18846 : _GEN_15374; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20772 = _issued_T_1 ? _GEN_18847 : _GEN_15375; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20773 = _issued_T_1 ? _GEN_18848 : _GEN_15376; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20774 = _issued_T_1 ? _GEN_18849 : _GEN_15377; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20775 = _issued_T_1 ? _GEN_18850 : _GEN_15378; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20776 = _issued_T_1 ? _GEN_18851 : _GEN_15379; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20777 = _issued_T_1 ? _GEN_18852 : _GEN_15380; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20778 = _issued_T_1 ? _GEN_18853 : _GEN_15381; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20779 = _issued_T_1 ? _GEN_18854 : _GEN_15382; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20780 = _issued_T_1 ? _GEN_18855 : _GEN_15383; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20781 = _issued_T_1 ? _GEN_18856 : _GEN_15384; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20782 = _issued_T_1 ? _GEN_18857 : _GEN_15385; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20783 = _issued_T_1 ? _GEN_18858 : _GEN_15386; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20784 = _issued_T_1 ? _GEN_18859 : _GEN_15387; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20785 = _issued_T_1 ? _GEN_18860 : _GEN_15388; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20786 = _issued_T_1 ? _GEN_18861 : _GEN_15389; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20787 = _issued_T_1 ? _GEN_18862 : _GEN_15390; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20788 = _issued_T_1 ? _GEN_18863 : _GEN_15391; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20789 = _issued_T_1 ? _GEN_18864 : _GEN_15392; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20790 = _issued_T_1 ? _GEN_18865 : _GEN_15393; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20791 = _issued_T_1 ? _GEN_18866 : _GEN_15394; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20792 = _issued_T_1 ? _GEN_18867 : _GEN_15395; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20793 = _issued_T_1 ? _GEN_18868 : _GEN_15396; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20794 = _issued_T_1 ? _GEN_18869 : _GEN_15397; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20843 = _issued_T_1 ? _GEN_18918 : _GEN_15446; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20844 = _issued_T_1 ? _GEN_18919 : _GEN_15447; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20845 = _issued_T_1 ? _GEN_18920 : _GEN_15448; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20846 = _issued_T_1 ? _GEN_18921 : _GEN_15449; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20847 = _issued_T_1 ? _GEN_18922 : _GEN_15450; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20848 = _issued_T_1 ? _GEN_18923 : _GEN_15451; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20849 = _issued_T_1 ? _GEN_18924 : _GEN_15452; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20850 = _issued_T_1 ? _GEN_18925 : _GEN_15453; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20851 = _issued_T_1 ? _GEN_18926 : _GEN_15454; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20852 = _issued_T_1 ? _GEN_18927 : _GEN_15455; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20853 = _issued_T_1 ? _GEN_18928 : _GEN_15456; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20854 = _issued_T_1 ? _GEN_18929 : _GEN_15457; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20855 = _issued_T_1 ? _GEN_18930 : _GEN_15458; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20856 = _issued_T_1 ? _GEN_18931 : _GEN_15459; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20857 = _issued_T_1 ? _GEN_18932 : _GEN_15460; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_20858 = _issued_T_1 ? _GEN_18933 : _GEN_15461; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_21163 = _issued_T_1 ? _GEN_19238 : _GEN_15766; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_21164 = _issued_T_1 ? _GEN_19239 : _GEN_15767; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_21165 = _issued_T_1 ? _GEN_19240 : _GEN_15768; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_21166 = _issued_T_1 ? _GEN_19241 : _GEN_15769; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_21167 = _issued_T_1 ? _GEN_19242 : _GEN_15770; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_21168 = _issued_T_1 ? _GEN_19243 : _GEN_15771; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_21169 = _issued_T_1 ? _GEN_19244 : _GEN_15772; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_21170 = _issued_T_1 ? _GEN_19245 : _GEN_15773; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_21171 = _issued_T_1 ? _GEN_19246 : _GEN_15774; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_21172 = _issued_T_1 ? _GEN_19247 : _GEN_15775; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_21173 = _issued_T_1 ? _GEN_19248 : _GEN_15776; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_21174 = _issued_T_1 ? _GEN_19249 : _GEN_15777; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_21175 = _issued_T_1 ? _GEN_19250 : _GEN_15778; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_21176 = _issued_T_1 ? _GEN_19251 : _GEN_15779; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_21177 = _issued_T_1 ? _GEN_19252 : _GEN_15780; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_21178 = _issued_T_1 ? _GEN_19253 : _GEN_15781; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_21339 = _issued_T_1 & io_loadIn_0_bits_lqDataWenDup_5; // @[LoadQueueFlag.scala 301:26 280:40]
  wire  _GEN_21397 = io_loadIn_0_valid ? _GEN_19771 : _GEN_16182; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21398 = io_loadIn_0_valid ? _GEN_19772 : _GEN_16183; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21399 = io_loadIn_0_valid ? _GEN_19773 : _GEN_16184; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21400 = io_loadIn_0_valid ? _GEN_19774 : _GEN_16185; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21401 = io_loadIn_0_valid ? _GEN_19775 : _GEN_16186; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21402 = io_loadIn_0_valid ? _GEN_19776 : _GEN_16187; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21403 = io_loadIn_0_valid ? _GEN_19777 : _GEN_16188; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21404 = io_loadIn_0_valid ? _GEN_19778 : _GEN_16189; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21405 = io_loadIn_0_valid ? _GEN_19779 : _GEN_16190; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21406 = io_loadIn_0_valid ? _GEN_19780 : _GEN_16191; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21407 = io_loadIn_0_valid ? _GEN_19781 : _GEN_16192; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21408 = io_loadIn_0_valid ? _GEN_19782 : _GEN_16193; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21409 = io_loadIn_0_valid ? _GEN_19783 : _GEN_16194; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21410 = io_loadIn_0_valid ? _GEN_19784 : _GEN_16195; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21411 = io_loadIn_0_valid ? _GEN_19785 : _GEN_16196; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21412 = io_loadIn_0_valid ? _GEN_19786 : _GEN_16197; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21413 = io_loadIn_0_valid ? _GEN_19787 : _GEN_16198; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21414 = io_loadIn_0_valid ? _GEN_19788 : _GEN_16199; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21415 = io_loadIn_0_valid ? _GEN_19789 : _GEN_16200; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21416 = io_loadIn_0_valid ? _GEN_19790 : _GEN_16201; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21417 = io_loadIn_0_valid ? _GEN_19791 : _GEN_16202; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21418 = io_loadIn_0_valid ? _GEN_19792 : _GEN_16203; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21419 = io_loadIn_0_valid ? _GEN_19793 : _GEN_16204; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21420 = io_loadIn_0_valid ? _GEN_19794 : _GEN_16205; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21421 = io_loadIn_0_valid ? _GEN_19795 : _GEN_16206; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21422 = io_loadIn_0_valid ? _GEN_19796 : _GEN_16207; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21423 = io_loadIn_0_valid ? _GEN_19797 : _GEN_16208; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21424 = io_loadIn_0_valid ? _GEN_19798 : _GEN_16209; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21425 = io_loadIn_0_valid ? _GEN_19799 : _GEN_16210; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21426 = io_loadIn_0_valid ? _GEN_19800 : _GEN_16211; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21427 = io_loadIn_0_valid ? _GEN_19801 : _GEN_16212; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21428 = io_loadIn_0_valid ? _GEN_19802 : _GEN_16213; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21429 = io_loadIn_0_valid ? _GEN_19803 : _GEN_16214; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21430 = io_loadIn_0_valid ? _GEN_19804 : _GEN_16215; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21431 = io_loadIn_0_valid ? _GEN_19805 : _GEN_16216; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21432 = io_loadIn_0_valid ? _GEN_19806 : _GEN_16217; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21433 = io_loadIn_0_valid ? _GEN_19807 : _GEN_16218; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21434 = io_loadIn_0_valid ? _GEN_19808 : _GEN_16219; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21435 = io_loadIn_0_valid ? _GEN_19809 : _GEN_16220; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21436 = io_loadIn_0_valid ? _GEN_19810 : _GEN_16221; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21437 = io_loadIn_0_valid ? _GEN_19811 : _GEN_16222; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21438 = io_loadIn_0_valid ? _GEN_19812 : _GEN_16223; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21439 = io_loadIn_0_valid ? _GEN_19813 : _GEN_16224; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21440 = io_loadIn_0_valid ? _GEN_19814 : _GEN_16225; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21441 = io_loadIn_0_valid ? _GEN_19815 : _GEN_16226; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21442 = io_loadIn_0_valid ? _GEN_19816 : _GEN_16227; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21443 = io_loadIn_0_valid ? _GEN_19817 : _GEN_16228; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21444 = io_loadIn_0_valid ? _GEN_19818 : _GEN_16229; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21445 = io_loadIn_0_valid ? _GEN_19819 : _GEN_16230; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21446 = io_loadIn_0_valid ? _GEN_19820 : _GEN_16231; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21447 = io_loadIn_0_valid ? _GEN_19821 : _GEN_16232; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21448 = io_loadIn_0_valid ? _GEN_19822 : _GEN_16233; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21449 = io_loadIn_0_valid ? _GEN_19823 : _GEN_16234; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21450 = io_loadIn_0_valid ? _GEN_19824 : _GEN_16235; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21451 = io_loadIn_0_valid ? _GEN_19825 : _GEN_16236; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21452 = io_loadIn_0_valid ? _GEN_19826 : _GEN_16237; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21453 = io_loadIn_0_valid ? _GEN_19827 : _GEN_16238; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21454 = io_loadIn_0_valid ? _GEN_19828 : _GEN_16239; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21455 = io_loadIn_0_valid ? _GEN_19829 : _GEN_16240; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21456 = io_loadIn_0_valid ? _GEN_19830 : _GEN_16241; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21457 = io_loadIn_0_valid ? _GEN_19831 : _GEN_16242; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21458 = io_loadIn_0_valid ? _GEN_19832 : _GEN_16243; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21459 = io_loadIn_0_valid ? _GEN_19833 : _GEN_16244; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21460 = io_loadIn_0_valid ? _GEN_19834 : _GEN_16245; // @[LoadQueueFlag.scala 286:31]
  wire [5:0] _GEN_21461 = io_loadIn_0_valid ? _GEN_19835 : _GEN_15878; // @[LoadQueueFlag.scala 286:31]
  wire [5:0] _GEN_21462 = io_loadIn_0_valid ? _GEN_19836 : _GEN_15879; // @[LoadQueueFlag.scala 286:31]
  wire [5:0] _GEN_21463 = io_loadIn_0_valid ? _GEN_19837 : _GEN_15880; // @[LoadQueueFlag.scala 286:31]
  wire [5:0] _GEN_21464 = io_loadIn_0_valid ? _GEN_19838 : _GEN_15881; // @[LoadQueueFlag.scala 286:31]
  wire [5:0] _GEN_21465 = io_loadIn_0_valid ? _GEN_19839 : _GEN_15882; // @[LoadQueueFlag.scala 286:31]
  wire [5:0] _GEN_21466 = io_loadIn_0_valid ? _GEN_19840 : _GEN_15883; // @[LoadQueueFlag.scala 286:31]
  wire [5:0] _GEN_21467 = io_loadIn_0_valid ? _GEN_19841 : _GEN_15884; // @[LoadQueueFlag.scala 286:31]
  wire [5:0] _GEN_21468 = io_loadIn_0_valid ? _GEN_19842 : _GEN_15885; // @[LoadQueueFlag.scala 286:31]
  wire [5:0] _GEN_21469 = io_loadIn_0_valid ? _GEN_19843 : _GEN_15886; // @[LoadQueueFlag.scala 286:31]
  wire [5:0] _GEN_21470 = io_loadIn_0_valid ? _GEN_19844 : _GEN_15887; // @[LoadQueueFlag.scala 286:31]
  wire [5:0] _GEN_21471 = io_loadIn_0_valid ? _GEN_19845 : _GEN_15888; // @[LoadQueueFlag.scala 286:31]
  wire [5:0] _GEN_21472 = io_loadIn_0_valid ? _GEN_19846 : _GEN_15889; // @[LoadQueueFlag.scala 286:31]
  wire [5:0] _GEN_21473 = io_loadIn_0_valid ? _GEN_19847 : _GEN_15890; // @[LoadQueueFlag.scala 286:31]
  wire [5:0] _GEN_21474 = io_loadIn_0_valid ? _GEN_19848 : _GEN_15891; // @[LoadQueueFlag.scala 286:31]
  wire [5:0] _GEN_21475 = io_loadIn_0_valid ? _GEN_19849 : _GEN_15892; // @[LoadQueueFlag.scala 286:31]
  wire [5:0] _GEN_21476 = io_loadIn_0_valid ? _GEN_19850 : _GEN_15893; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21589 = io_loadIn_0_valid ? _GEN_19963 : _GEN_14566; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21590 = io_loadIn_0_valid ? _GEN_19964 : _GEN_14567; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21591 = io_loadIn_0_valid ? _GEN_19965 : _GEN_14568; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21592 = io_loadIn_0_valid ? _GEN_19966 : _GEN_14569; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21593 = io_loadIn_0_valid ? _GEN_19967 : _GEN_14570; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21594 = io_loadIn_0_valid ? _GEN_19968 : _GEN_14571; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21595 = io_loadIn_0_valid ? _GEN_19969 : _GEN_14572; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21596 = io_loadIn_0_valid ? _GEN_19970 : _GEN_14573; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21597 = io_loadIn_0_valid ? _GEN_19971 : _GEN_14574; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21598 = io_loadIn_0_valid ? _GEN_19972 : _GEN_14575; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21599 = io_loadIn_0_valid ? _GEN_19973 : _GEN_14576; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21600 = io_loadIn_0_valid ? _GEN_19974 : _GEN_14577; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21601 = io_loadIn_0_valid ? _GEN_19975 : _GEN_14578; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21602 = io_loadIn_0_valid ? _GEN_19976 : _GEN_14579; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21603 = io_loadIn_0_valid ? _GEN_19977 : _GEN_14580; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21604 = io_loadIn_0_valid ? _GEN_19978 : _GEN_14581; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21605 = io_loadIn_0_valid ? _GEN_19979 : _GEN_14582; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21606 = io_loadIn_0_valid ? _GEN_19980 : _GEN_14583; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21607 = io_loadIn_0_valid ? _GEN_19981 : _GEN_14584; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21608 = io_loadIn_0_valid ? _GEN_19982 : _GEN_14585; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21609 = io_loadIn_0_valid ? _GEN_19983 : _GEN_14586; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21610 = io_loadIn_0_valid ? _GEN_19984 : _GEN_14587; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21611 = io_loadIn_0_valid ? _GEN_19985 : _GEN_14588; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21612 = io_loadIn_0_valid ? _GEN_19986 : _GEN_14589; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21613 = io_loadIn_0_valid ? _GEN_19987 : _GEN_14590; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21614 = io_loadIn_0_valid ? _GEN_19988 : _GEN_14591; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21615 = io_loadIn_0_valid ? _GEN_19989 : _GEN_14592; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21616 = io_loadIn_0_valid ? _GEN_19990 : _GEN_14593; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21617 = io_loadIn_0_valid ? _GEN_19991 : _GEN_14594; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21618 = io_loadIn_0_valid ? _GEN_19992 : _GEN_14595; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21619 = io_loadIn_0_valid ? _GEN_19993 : _GEN_14596; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21620 = io_loadIn_0_valid ? _GEN_19994 : _GEN_14597; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21733 = io_loadIn_0_valid ? _GEN_20107 : _GEN_14710; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21734 = io_loadIn_0_valid ? _GEN_20108 : _GEN_14711; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21735 = io_loadIn_0_valid ? _GEN_20109 : _GEN_14712; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21736 = io_loadIn_0_valid ? _GEN_20110 : _GEN_14713; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21737 = io_loadIn_0_valid ? _GEN_20111 : _GEN_14714; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21738 = io_loadIn_0_valid ? _GEN_20112 : _GEN_14715; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21739 = io_loadIn_0_valid ? _GEN_20113 : _GEN_14716; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21740 = io_loadIn_0_valid ? _GEN_20114 : _GEN_14717; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21741 = io_loadIn_0_valid ? _GEN_20115 : _GEN_14718; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21742 = io_loadIn_0_valid ? _GEN_20116 : _GEN_14719; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21743 = io_loadIn_0_valid ? _GEN_20117 : _GEN_14720; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21744 = io_loadIn_0_valid ? _GEN_20118 : _GEN_14721; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21745 = io_loadIn_0_valid ? _GEN_20119 : _GEN_14722; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21746 = io_loadIn_0_valid ? _GEN_20120 : _GEN_14723; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21747 = io_loadIn_0_valid ? _GEN_20121 : _GEN_14724; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21748 = io_loadIn_0_valid ? _GEN_20122 : _GEN_14725; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21861 = io_loadIn_0_valid ? _GEN_20235 : _GEN_14838; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21862 = io_loadIn_0_valid ? _GEN_20236 : _GEN_14839; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21863 = io_loadIn_0_valid ? _GEN_20237 : _GEN_14840; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21864 = io_loadIn_0_valid ? _GEN_20238 : _GEN_14841; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21865 = io_loadIn_0_valid ? _GEN_20239 : _GEN_14842; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21866 = io_loadIn_0_valid ? _GEN_20240 : _GEN_14843; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21867 = io_loadIn_0_valid ? _GEN_20241 : _GEN_14844; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21868 = io_loadIn_0_valid ? _GEN_20242 : _GEN_14845; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21869 = io_loadIn_0_valid ? _GEN_20243 : _GEN_14846; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21870 = io_loadIn_0_valid ? _GEN_20244 : _GEN_14847; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21871 = io_loadIn_0_valid ? _GEN_20245 : _GEN_14848; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21872 = io_loadIn_0_valid ? _GEN_20246 : _GEN_14849; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21873 = io_loadIn_0_valid ? _GEN_20247 : _GEN_14850; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21874 = io_loadIn_0_valid ? _GEN_20248 : _GEN_14851; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21875 = io_loadIn_0_valid ? _GEN_20249 : _GEN_14852; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21876 = io_loadIn_0_valid ? _GEN_20250 : _GEN_14853; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21877 = io_loadIn_0_valid ? _GEN_20251 : _GEN_14854; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21878 = io_loadIn_0_valid ? _GEN_20252 : _GEN_14855; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21879 = io_loadIn_0_valid ? _GEN_20253 : _GEN_14856; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21880 = io_loadIn_0_valid ? _GEN_20254 : _GEN_14857; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21881 = io_loadIn_0_valid ? _GEN_20255 : _GEN_14858; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21882 = io_loadIn_0_valid ? _GEN_20256 : _GEN_14859; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21883 = io_loadIn_0_valid ? _GEN_20257 : _GEN_14860; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21884 = io_loadIn_0_valid ? _GEN_20258 : _GEN_14861; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21885 = io_loadIn_0_valid ? _GEN_20259 : _GEN_14862; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21886 = io_loadIn_0_valid ? _GEN_20260 : _GEN_14863; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21887 = io_loadIn_0_valid ? _GEN_20261 : _GEN_14864; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21888 = io_loadIn_0_valid ? _GEN_20262 : _GEN_14865; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21889 = io_loadIn_0_valid ? _GEN_20263 : _GEN_14866; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21890 = io_loadIn_0_valid ? _GEN_20264 : _GEN_14867; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21891 = io_loadIn_0_valid ? _GEN_20265 : _GEN_14868; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21892 = io_loadIn_0_valid ? _GEN_20266 : _GEN_14869; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21893 = io_loadIn_0_valid ? _GEN_20267 : _GEN_14870; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21894 = io_loadIn_0_valid ? _GEN_20268 : _GEN_14871; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21895 = io_loadIn_0_valid ? _GEN_20269 : _GEN_14872; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21896 = io_loadIn_0_valid ? _GEN_20270 : _GEN_14873; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21897 = io_loadIn_0_valid ? _GEN_20271 : _GEN_14874; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21898 = io_loadIn_0_valid ? _GEN_20272 : _GEN_14875; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21899 = io_loadIn_0_valid ? _GEN_20273 : _GEN_14876; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21900 = io_loadIn_0_valid ? _GEN_20274 : _GEN_14877; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21901 = io_loadIn_0_valid ? _GEN_20275 : _GEN_14878; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21902 = io_loadIn_0_valid ? _GEN_20276 : _GEN_14879; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21903 = io_loadIn_0_valid ? _GEN_20277 : _GEN_14880; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21904 = io_loadIn_0_valid ? _GEN_20278 : _GEN_14881; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21905 = io_loadIn_0_valid ? _GEN_20279 : _GEN_14882; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21906 = io_loadIn_0_valid ? _GEN_20280 : _GEN_14883; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21907 = io_loadIn_0_valid ? _GEN_20281 : _GEN_14884; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21908 = io_loadIn_0_valid ? _GEN_20282 : _GEN_14885; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21941 = io_loadIn_0_valid ? _GEN_20315 : _GEN_14918; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21942 = io_loadIn_0_valid ? _GEN_20316 : _GEN_14919; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21943 = io_loadIn_0_valid ? _GEN_20317 : _GEN_14920; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21944 = io_loadIn_0_valid ? _GEN_20318 : _GEN_14921; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21945 = io_loadIn_0_valid ? _GEN_20319 : _GEN_14922; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21946 = io_loadIn_0_valid ? _GEN_20320 : _GEN_14923; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21947 = io_loadIn_0_valid ? _GEN_20321 : _GEN_14924; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21948 = io_loadIn_0_valid ? _GEN_20322 : _GEN_14925; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21949 = io_loadIn_0_valid ? _GEN_20323 : _GEN_14926; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21950 = io_loadIn_0_valid ? _GEN_20324 : _GEN_14927; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21951 = io_loadIn_0_valid ? _GEN_20325 : _GEN_14928; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21952 = io_loadIn_0_valid ? _GEN_20326 : _GEN_14929; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21953 = io_loadIn_0_valid ? _GEN_20327 : _GEN_14930; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21954 = io_loadIn_0_valid ? _GEN_20328 : _GEN_14931; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21955 = io_loadIn_0_valid ? _GEN_20329 : _GEN_14932; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_21956 = io_loadIn_0_valid ? _GEN_20330 : _GEN_14933; // @[LoadQueueFlag.scala 286:31]
  wire [6:0] _GEN_22373 = io_loadIn_0_valid ? _GEN_20747 : _GEN_15350; // @[LoadQueueFlag.scala 286:31]
  wire [6:0] _GEN_22374 = io_loadIn_0_valid ? _GEN_20748 : _GEN_15351; // @[LoadQueueFlag.scala 286:31]
  wire [6:0] _GEN_22375 = io_loadIn_0_valid ? _GEN_20749 : _GEN_15352; // @[LoadQueueFlag.scala 286:31]
  wire [6:0] _GEN_22376 = io_loadIn_0_valid ? _GEN_20750 : _GEN_15353; // @[LoadQueueFlag.scala 286:31]
  wire [6:0] _GEN_22377 = io_loadIn_0_valid ? _GEN_20751 : _GEN_15354; // @[LoadQueueFlag.scala 286:31]
  wire [6:0] _GEN_22378 = io_loadIn_0_valid ? _GEN_20752 : _GEN_15355; // @[LoadQueueFlag.scala 286:31]
  wire [6:0] _GEN_22379 = io_loadIn_0_valid ? _GEN_20753 : _GEN_15356; // @[LoadQueueFlag.scala 286:31]
  wire [6:0] _GEN_22380 = io_loadIn_0_valid ? _GEN_20754 : _GEN_15357; // @[LoadQueueFlag.scala 286:31]
  wire [6:0] _GEN_22381 = io_loadIn_0_valid ? _GEN_20755 : _GEN_15358; // @[LoadQueueFlag.scala 286:31]
  wire [6:0] _GEN_22382 = io_loadIn_0_valid ? _GEN_20756 : _GEN_15359; // @[LoadQueueFlag.scala 286:31]
  wire [6:0] _GEN_22383 = io_loadIn_0_valid ? _GEN_20757 : _GEN_15360; // @[LoadQueueFlag.scala 286:31]
  wire [6:0] _GEN_22384 = io_loadIn_0_valid ? _GEN_20758 : _GEN_15361; // @[LoadQueueFlag.scala 286:31]
  wire [6:0] _GEN_22385 = io_loadIn_0_valid ? _GEN_20759 : _GEN_15362; // @[LoadQueueFlag.scala 286:31]
  wire [6:0] _GEN_22386 = io_loadIn_0_valid ? _GEN_20760 : _GEN_15363; // @[LoadQueueFlag.scala 286:31]
  wire [6:0] _GEN_22387 = io_loadIn_0_valid ? _GEN_20761 : _GEN_15364; // @[LoadQueueFlag.scala 286:31]
  wire [6:0] _GEN_22388 = io_loadIn_0_valid ? _GEN_20762 : _GEN_15365; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_22389 = io_loadIn_0_valid ? _GEN_20763 : _GEN_15366; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_22390 = io_loadIn_0_valid ? _GEN_20764 : _GEN_15367; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_22391 = io_loadIn_0_valid ? _GEN_20765 : _GEN_15368; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_22392 = io_loadIn_0_valid ? _GEN_20766 : _GEN_15369; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_22393 = io_loadIn_0_valid ? _GEN_20767 : _GEN_15370; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_22394 = io_loadIn_0_valid ? _GEN_20768 : _GEN_15371; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_22395 = io_loadIn_0_valid ? _GEN_20769 : _GEN_15372; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_22396 = io_loadIn_0_valid ? _GEN_20770 : _GEN_15373; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_22397 = io_loadIn_0_valid ? _GEN_20771 : _GEN_15374; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_22398 = io_loadIn_0_valid ? _GEN_20772 : _GEN_15375; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_22399 = io_loadIn_0_valid ? _GEN_20773 : _GEN_15376; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_22400 = io_loadIn_0_valid ? _GEN_20774 : _GEN_15377; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_22401 = io_loadIn_0_valid ? _GEN_20775 : _GEN_15378; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_22402 = io_loadIn_0_valid ? _GEN_20776 : _GEN_15379; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_22403 = io_loadIn_0_valid ? _GEN_20777 : _GEN_15380; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_22404 = io_loadIn_0_valid ? _GEN_20778 : _GEN_15381; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_22405 = io_loadIn_0_valid ? _GEN_20779 : _GEN_15382; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_22406 = io_loadIn_0_valid ? _GEN_20780 : _GEN_15383; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_22407 = io_loadIn_0_valid ? _GEN_20781 : _GEN_15384; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_22408 = io_loadIn_0_valid ? _GEN_20782 : _GEN_15385; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_22409 = io_loadIn_0_valid ? _GEN_20783 : _GEN_15386; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_22410 = io_loadIn_0_valid ? _GEN_20784 : _GEN_15387; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_22411 = io_loadIn_0_valid ? _GEN_20785 : _GEN_15388; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_22412 = io_loadIn_0_valid ? _GEN_20786 : _GEN_15389; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_22413 = io_loadIn_0_valid ? _GEN_20787 : _GEN_15390; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_22414 = io_loadIn_0_valid ? _GEN_20788 : _GEN_15391; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_22415 = io_loadIn_0_valid ? _GEN_20789 : _GEN_15392; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_22416 = io_loadIn_0_valid ? _GEN_20790 : _GEN_15393; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_22417 = io_loadIn_0_valid ? _GEN_20791 : _GEN_15394; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_22418 = io_loadIn_0_valid ? _GEN_20792 : _GEN_15395; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_22419 = io_loadIn_0_valid ? _GEN_20793 : _GEN_15396; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_22420 = io_loadIn_0_valid ? _GEN_20794 : _GEN_15397; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_22469 = io_loadIn_0_valid ? _GEN_20843 : _GEN_15446; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_22470 = io_loadIn_0_valid ? _GEN_20844 : _GEN_15447; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_22471 = io_loadIn_0_valid ? _GEN_20845 : _GEN_15448; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_22472 = io_loadIn_0_valid ? _GEN_20846 : _GEN_15449; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_22473 = io_loadIn_0_valid ? _GEN_20847 : _GEN_15450; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_22474 = io_loadIn_0_valid ? _GEN_20848 : _GEN_15451; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_22475 = io_loadIn_0_valid ? _GEN_20849 : _GEN_15452; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_22476 = io_loadIn_0_valid ? _GEN_20850 : _GEN_15453; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_22477 = io_loadIn_0_valid ? _GEN_20851 : _GEN_15454; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_22478 = io_loadIn_0_valid ? _GEN_20852 : _GEN_15455; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_22479 = io_loadIn_0_valid ? _GEN_20853 : _GEN_15456; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_22480 = io_loadIn_0_valid ? _GEN_20854 : _GEN_15457; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_22481 = io_loadIn_0_valid ? _GEN_20855 : _GEN_15458; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_22482 = io_loadIn_0_valid ? _GEN_20856 : _GEN_15459; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_22483 = io_loadIn_0_valid ? _GEN_20857 : _GEN_15460; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_22484 = io_loadIn_0_valid ? _GEN_20858 : _GEN_15461; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_22789 = io_loadIn_0_valid ? _GEN_21163 : _GEN_15766; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_22790 = io_loadIn_0_valid ? _GEN_21164 : _GEN_15767; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_22791 = io_loadIn_0_valid ? _GEN_21165 : _GEN_15768; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_22792 = io_loadIn_0_valid ? _GEN_21166 : _GEN_15769; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_22793 = io_loadIn_0_valid ? _GEN_21167 : _GEN_15770; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_22794 = io_loadIn_0_valid ? _GEN_21168 : _GEN_15771; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_22795 = io_loadIn_0_valid ? _GEN_21169 : _GEN_15772; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_22796 = io_loadIn_0_valid ? _GEN_21170 : _GEN_15773; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_22797 = io_loadIn_0_valid ? _GEN_21171 : _GEN_15774; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_22798 = io_loadIn_0_valid ? _GEN_21172 : _GEN_15775; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_22799 = io_loadIn_0_valid ? _GEN_21173 : _GEN_15776; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_22800 = io_loadIn_0_valid ? _GEN_21174 : _GEN_15777; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_22801 = io_loadIn_0_valid ? _GEN_21175 : _GEN_15778; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_22802 = io_loadIn_0_valid ? _GEN_21176 : _GEN_15779; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_22803 = io_loadIn_0_valid ? _GEN_21177 : _GEN_15780; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_22804 = io_loadIn_0_valid ? _GEN_21178 : _GEN_15781; // @[LoadQueueFlag.scala 286:31]
  reg  io_rob_isMMIO_0_REG; // @[LoadQueueFlag.scala 358:32]
  reg [4:0] io_rob_uop_0_REG_robIdx_value; // @[LoadQueueFlag.scala 359:29]
  wire [15:0] _hasExceptions_T_1 = {2'h0,io_loadIn_1_bits_uop_cf_exceptionVec_13,1'h0,4'h0,2'h0,
    io_loadIn_1_bits_uop_cf_exceptionVec_5,io_loadIn_1_bits_uop_cf_exceptionVec_4,4'h0}; // @[LoadQueueFlag.scala 287:97]
  wire  hasExceptions_1 = |_hasExceptions_T_1; // @[LoadQueueFlag.scala 287:104]
  wire [7:0] _needReplay_T_1 = {io_loadIn_1_bits_replayInfo_cause_7,io_loadIn_1_bits_replayInfo_cause_6,
    io_loadIn_1_bits_replayInfo_cause_5,io_loadIn_1_bits_replayInfo_cause_4,io_loadIn_1_bits_replayInfo_cause_3,
    io_loadIn_1_bits_replayInfo_cause_2,io_loadIn_1_bits_replayInfo_cause_1,io_loadIn_1_bits_replayInfo_cause_0}; // @[LoadUnit.scala 62:29]
  wire  needReplay_1 = |_needReplay_T_1; // @[LoadUnit.scala 62:36]
  wire  _datavalidVal_T_2 = ~io_loadIn_1_bits_mmio; // @[LoadQueueFlag.scala 295:13]
  wire  _datavalidVal_T_3 = ~io_loadIn_1_bits_miss; // @[LoadQueueFlag.scala 296:13]
  wire  datavalidVal_1 = ~io_loadIn_1_bits_mmio & _datavalidVal_T_3; // @[LoadQueueFlag.scala 295:37]
  wire  _issued_T_7 = ~needReplay_1; // @[LoadQueueFlag.scala 299:29]
  wire  _issued_T_8 = ~io_loadIn_1_bits_tlbMiss; // @[LoadQueueFlag.scala 299:44]
  wire  _GEN_23039 = 4'h0 == io_loadIn_1_bits_uop_lqIdx_value ? datavalidVal_1 : _GEN_21413; // @[LoadQueueFlag.scala 304:{32,32}]
  wire  _GEN_23040 = 4'h1 == io_loadIn_1_bits_uop_lqIdx_value ? datavalidVal_1 : _GEN_21414; // @[LoadQueueFlag.scala 304:{32,32}]
  wire  _GEN_23041 = 4'h2 == io_loadIn_1_bits_uop_lqIdx_value ? datavalidVal_1 : _GEN_21415; // @[LoadQueueFlag.scala 304:{32,32}]
  wire  _GEN_23042 = 4'h3 == io_loadIn_1_bits_uop_lqIdx_value ? datavalidVal_1 : _GEN_21416; // @[LoadQueueFlag.scala 304:{32,32}]
  wire  _GEN_23043 = 4'h4 == io_loadIn_1_bits_uop_lqIdx_value ? datavalidVal_1 : _GEN_21417; // @[LoadQueueFlag.scala 304:{32,32}]
  wire  _GEN_23044 = 4'h5 == io_loadIn_1_bits_uop_lqIdx_value ? datavalidVal_1 : _GEN_21418; // @[LoadQueueFlag.scala 304:{32,32}]
  wire  _GEN_23045 = 4'h6 == io_loadIn_1_bits_uop_lqIdx_value ? datavalidVal_1 : _GEN_21419; // @[LoadQueueFlag.scala 304:{32,32}]
  wire  _GEN_23046 = 4'h7 == io_loadIn_1_bits_uop_lqIdx_value ? datavalidVal_1 : _GEN_21420; // @[LoadQueueFlag.scala 304:{32,32}]
  wire  _GEN_23047 = 4'h8 == io_loadIn_1_bits_uop_lqIdx_value ? datavalidVal_1 : _GEN_21421; // @[LoadQueueFlag.scala 304:{32,32}]
  wire  _GEN_23048 = 4'h9 == io_loadIn_1_bits_uop_lqIdx_value ? datavalidVal_1 : _GEN_21422; // @[LoadQueueFlag.scala 304:{32,32}]
  wire  _GEN_23049 = 4'ha == io_loadIn_1_bits_uop_lqIdx_value ? datavalidVal_1 : _GEN_21423; // @[LoadQueueFlag.scala 304:{32,32}]
  wire  _GEN_23050 = 4'hb == io_loadIn_1_bits_uop_lqIdx_value ? datavalidVal_1 : _GEN_21424; // @[LoadQueueFlag.scala 304:{32,32}]
  wire  _GEN_23051 = 4'hc == io_loadIn_1_bits_uop_lqIdx_value ? datavalidVal_1 : _GEN_21425; // @[LoadQueueFlag.scala 304:{32,32}]
  wire  _GEN_23052 = 4'hd == io_loadIn_1_bits_uop_lqIdx_value ? datavalidVal_1 : _GEN_21426; // @[LoadQueueFlag.scala 304:{32,32}]
  wire  _GEN_23053 = 4'he == io_loadIn_1_bits_uop_lqIdx_value ? datavalidVal_1 : _GEN_21427; // @[LoadQueueFlag.scala 304:{32,32}]
  wire  _GEN_23054 = 4'hf == io_loadIn_1_bits_uop_lqIdx_value ? datavalidVal_1 : _GEN_21428; // @[LoadQueueFlag.scala 304:{32,32}]
  wire  _GEN_23055 = 4'h0 == io_loadIn_1_bits_uop_lqIdx_value ? io_loadIn_1_bits_mmio : _GEN_21429; // @[LoadQueueFlag.scala 305:{30,30}]
  wire  _GEN_23056 = 4'h1 == io_loadIn_1_bits_uop_lqIdx_value ? io_loadIn_1_bits_mmio : _GEN_21430; // @[LoadQueueFlag.scala 305:{30,30}]
  wire  _GEN_23057 = 4'h2 == io_loadIn_1_bits_uop_lqIdx_value ? io_loadIn_1_bits_mmio : _GEN_21431; // @[LoadQueueFlag.scala 305:{30,30}]
  wire  _GEN_23058 = 4'h3 == io_loadIn_1_bits_uop_lqIdx_value ? io_loadIn_1_bits_mmio : _GEN_21432; // @[LoadQueueFlag.scala 305:{30,30}]
  wire  _GEN_23059 = 4'h4 == io_loadIn_1_bits_uop_lqIdx_value ? io_loadIn_1_bits_mmio : _GEN_21433; // @[LoadQueueFlag.scala 305:{30,30}]
  wire  _GEN_23060 = 4'h5 == io_loadIn_1_bits_uop_lqIdx_value ? io_loadIn_1_bits_mmio : _GEN_21434; // @[LoadQueueFlag.scala 305:{30,30}]
  wire  _GEN_23061 = 4'h6 == io_loadIn_1_bits_uop_lqIdx_value ? io_loadIn_1_bits_mmio : _GEN_21435; // @[LoadQueueFlag.scala 305:{30,30}]
  wire  _GEN_23062 = 4'h7 == io_loadIn_1_bits_uop_lqIdx_value ? io_loadIn_1_bits_mmio : _GEN_21436; // @[LoadQueueFlag.scala 305:{30,30}]
  wire  _GEN_23063 = 4'h8 == io_loadIn_1_bits_uop_lqIdx_value ? io_loadIn_1_bits_mmio : _GEN_21437; // @[LoadQueueFlag.scala 305:{30,30}]
  wire  _GEN_23064 = 4'h9 == io_loadIn_1_bits_uop_lqIdx_value ? io_loadIn_1_bits_mmio : _GEN_21438; // @[LoadQueueFlag.scala 305:{30,30}]
  wire  _GEN_23065 = 4'ha == io_loadIn_1_bits_uop_lqIdx_value ? io_loadIn_1_bits_mmio : _GEN_21439; // @[LoadQueueFlag.scala 305:{30,30}]
  wire  _GEN_23066 = 4'hb == io_loadIn_1_bits_uop_lqIdx_value ? io_loadIn_1_bits_mmio : _GEN_21440; // @[LoadQueueFlag.scala 305:{30,30}]
  wire  _GEN_23067 = 4'hc == io_loadIn_1_bits_uop_lqIdx_value ? io_loadIn_1_bits_mmio : _GEN_21441; // @[LoadQueueFlag.scala 305:{30,30}]
  wire  _GEN_23068 = 4'hd == io_loadIn_1_bits_uop_lqIdx_value ? io_loadIn_1_bits_mmio : _GEN_21442; // @[LoadQueueFlag.scala 305:{30,30}]
  wire  _GEN_23069 = 4'he == io_loadIn_1_bits_uop_lqIdx_value ? io_loadIn_1_bits_mmio : _GEN_21443; // @[LoadQueueFlag.scala 305:{30,30}]
  wire  _GEN_23070 = 4'hf == io_loadIn_1_bits_uop_lqIdx_value ? io_loadIn_1_bits_mmio : _GEN_21444; // @[LoadQueueFlag.scala 305:{30,30}]
  wire  _GEN_23071 = 4'h0 == io_loadIn_1_bits_uop_lqIdx_value ? _datavalidVal_T_2 & ~hasExceptions_1 : _GEN_21445; // @[LoadQueueFlag.scala 306:{34,34}]
  wire  _GEN_23072 = 4'h1 == io_loadIn_1_bits_uop_lqIdx_value ? _datavalidVal_T_2 & ~hasExceptions_1 : _GEN_21446; // @[LoadQueueFlag.scala 306:{34,34}]
  wire  _GEN_23073 = 4'h2 == io_loadIn_1_bits_uop_lqIdx_value ? _datavalidVal_T_2 & ~hasExceptions_1 : _GEN_21447; // @[LoadQueueFlag.scala 306:{34,34}]
  wire  _GEN_23074 = 4'h3 == io_loadIn_1_bits_uop_lqIdx_value ? _datavalidVal_T_2 & ~hasExceptions_1 : _GEN_21448; // @[LoadQueueFlag.scala 306:{34,34}]
  wire  _GEN_23075 = 4'h4 == io_loadIn_1_bits_uop_lqIdx_value ? _datavalidVal_T_2 & ~hasExceptions_1 : _GEN_21449; // @[LoadQueueFlag.scala 306:{34,34}]
  wire  _GEN_23076 = 4'h5 == io_loadIn_1_bits_uop_lqIdx_value ? _datavalidVal_T_2 & ~hasExceptions_1 : _GEN_21450; // @[LoadQueueFlag.scala 306:{34,34}]
  wire  _GEN_23077 = 4'h6 == io_loadIn_1_bits_uop_lqIdx_value ? _datavalidVal_T_2 & ~hasExceptions_1 : _GEN_21451; // @[LoadQueueFlag.scala 306:{34,34}]
  wire  _GEN_23078 = 4'h7 == io_loadIn_1_bits_uop_lqIdx_value ? _datavalidVal_T_2 & ~hasExceptions_1 : _GEN_21452; // @[LoadQueueFlag.scala 306:{34,34}]
  wire  _GEN_23079 = 4'h8 == io_loadIn_1_bits_uop_lqIdx_value ? _datavalidVal_T_2 & ~hasExceptions_1 : _GEN_21453; // @[LoadQueueFlag.scala 306:{34,34}]
  wire  _GEN_23080 = 4'h9 == io_loadIn_1_bits_uop_lqIdx_value ? _datavalidVal_T_2 & ~hasExceptions_1 : _GEN_21454; // @[LoadQueueFlag.scala 306:{34,34}]
  wire  _GEN_23081 = 4'ha == io_loadIn_1_bits_uop_lqIdx_value ? _datavalidVal_T_2 & ~hasExceptions_1 : _GEN_21455; // @[LoadQueueFlag.scala 306:{34,34}]
  wire  _GEN_23082 = 4'hb == io_loadIn_1_bits_uop_lqIdx_value ? _datavalidVal_T_2 & ~hasExceptions_1 : _GEN_21456; // @[LoadQueueFlag.scala 306:{34,34}]
  wire  _GEN_23083 = 4'hc == io_loadIn_1_bits_uop_lqIdx_value ? _datavalidVal_T_2 & ~hasExceptions_1 : _GEN_21457; // @[LoadQueueFlag.scala 306:{34,34}]
  wire  _GEN_23084 = 4'hd == io_loadIn_1_bits_uop_lqIdx_value ? _datavalidVal_T_2 & ~hasExceptions_1 : _GEN_21458; // @[LoadQueueFlag.scala 306:{34,34}]
  wire  _GEN_23085 = 4'he == io_loadIn_1_bits_uop_lqIdx_value ? _datavalidVal_T_2 & ~hasExceptions_1 : _GEN_21459; // @[LoadQueueFlag.scala 306:{34,34}]
  wire  _GEN_23086 = 4'hf == io_loadIn_1_bits_uop_lqIdx_value ? _datavalidVal_T_2 & ~hasExceptions_1 : _GEN_21460; // @[LoadQueueFlag.scala 306:{34,34}]
  wire  _GEN_26308 = _issued_T_7 ? _GEN_23039 : _GEN_21413; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_26309 = _issued_T_7 ? _GEN_23040 : _GEN_21414; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_26310 = _issued_T_7 ? _GEN_23041 : _GEN_21415; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_26311 = _issued_T_7 ? _GEN_23042 : _GEN_21416; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_26312 = _issued_T_7 ? _GEN_23043 : _GEN_21417; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_26313 = _issued_T_7 ? _GEN_23044 : _GEN_21418; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_26314 = _issued_T_7 ? _GEN_23045 : _GEN_21419; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_26315 = _issued_T_7 ? _GEN_23046 : _GEN_21420; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_26316 = _issued_T_7 ? _GEN_23047 : _GEN_21421; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_26317 = _issued_T_7 ? _GEN_23048 : _GEN_21422; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_26318 = _issued_T_7 ? _GEN_23049 : _GEN_21423; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_26319 = _issued_T_7 ? _GEN_23050 : _GEN_21424; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_26320 = _issued_T_7 ? _GEN_23051 : _GEN_21425; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_26321 = _issued_T_7 ? _GEN_23052 : _GEN_21426; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_26322 = _issued_T_7 ? _GEN_23053 : _GEN_21427; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_26323 = _issued_T_7 ? _GEN_23054 : _GEN_21428; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_26324 = _issued_T_7 ? _GEN_23055 : _GEN_21429; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_26325 = _issued_T_7 ? _GEN_23056 : _GEN_21430; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_26326 = _issued_T_7 ? _GEN_23057 : _GEN_21431; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_26327 = _issued_T_7 ? _GEN_23058 : _GEN_21432; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_26328 = _issued_T_7 ? _GEN_23059 : _GEN_21433; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_26329 = _issued_T_7 ? _GEN_23060 : _GEN_21434; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_26330 = _issued_T_7 ? _GEN_23061 : _GEN_21435; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_26331 = _issued_T_7 ? _GEN_23062 : _GEN_21436; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_26332 = _issued_T_7 ? _GEN_23063 : _GEN_21437; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_26333 = _issued_T_7 ? _GEN_23064 : _GEN_21438; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_26334 = _issued_T_7 ? _GEN_23065 : _GEN_21439; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_26335 = _issued_T_7 ? _GEN_23066 : _GEN_21440; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_26336 = _issued_T_7 ? _GEN_23067 : _GEN_21441; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_26337 = _issued_T_7 ? _GEN_23068 : _GEN_21442; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_26338 = _issued_T_7 ? _GEN_23069 : _GEN_21443; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_26339 = _issued_T_7 ? _GEN_23070 : _GEN_21444; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_26340 = _issued_T_7 ? _GEN_23071 : _GEN_21445; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_26341 = _issued_T_7 ? _GEN_23072 : _GEN_21446; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_26342 = _issued_T_7 ? _GEN_23073 : _GEN_21447; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_26343 = _issued_T_7 ? _GEN_23074 : _GEN_21448; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_26344 = _issued_T_7 ? _GEN_23075 : _GEN_21449; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_26345 = _issued_T_7 ? _GEN_23076 : _GEN_21450; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_26346 = _issued_T_7 ? _GEN_23077 : _GEN_21451; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_26347 = _issued_T_7 ? _GEN_23078 : _GEN_21452; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_26348 = _issued_T_7 ? _GEN_23079 : _GEN_21453; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_26349 = _issued_T_7 ? _GEN_23080 : _GEN_21454; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_26350 = _issued_T_7 ? _GEN_23081 : _GEN_21455; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_26351 = _issued_T_7 ? _GEN_23082 : _GEN_21456; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_26352 = _issued_T_7 ? _GEN_23083 : _GEN_21457; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_26353 = _issued_T_7 ? _GEN_23084 : _GEN_21458; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_26354 = _issued_T_7 ? _GEN_23085 : _GEN_21459; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_26355 = _issued_T_7 ? _GEN_23086 : _GEN_21460; // @[LoadQueueFlag.scala 301:26]
  wire  _GEN_27860 = _issued_T_7 & io_loadIn_1_bits_lqDataWenDup_5; // @[LoadQueueFlag.scala 301:26 280:40]
  wire  _GEN_27934 = io_loadIn_1_valid ? _GEN_26308 : _GEN_21413; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_27935 = io_loadIn_1_valid ? _GEN_26309 : _GEN_21414; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_27936 = io_loadIn_1_valid ? _GEN_26310 : _GEN_21415; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_27937 = io_loadIn_1_valid ? _GEN_26311 : _GEN_21416; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_27938 = io_loadIn_1_valid ? _GEN_26312 : _GEN_21417; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_27939 = io_loadIn_1_valid ? _GEN_26313 : _GEN_21418; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_27940 = io_loadIn_1_valid ? _GEN_26314 : _GEN_21419; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_27941 = io_loadIn_1_valid ? _GEN_26315 : _GEN_21420; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_27942 = io_loadIn_1_valid ? _GEN_26316 : _GEN_21421; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_27943 = io_loadIn_1_valid ? _GEN_26317 : _GEN_21422; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_27944 = io_loadIn_1_valid ? _GEN_26318 : _GEN_21423; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_27945 = io_loadIn_1_valid ? _GEN_26319 : _GEN_21424; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_27946 = io_loadIn_1_valid ? _GEN_26320 : _GEN_21425; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_27947 = io_loadIn_1_valid ? _GEN_26321 : _GEN_21426; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_27948 = io_loadIn_1_valid ? _GEN_26322 : _GEN_21427; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_27949 = io_loadIn_1_valid ? _GEN_26323 : _GEN_21428; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_27950 = io_loadIn_1_valid ? _GEN_26324 : _GEN_21429; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_27951 = io_loadIn_1_valid ? _GEN_26325 : _GEN_21430; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_27952 = io_loadIn_1_valid ? _GEN_26326 : _GEN_21431; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_27953 = io_loadIn_1_valid ? _GEN_26327 : _GEN_21432; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_27954 = io_loadIn_1_valid ? _GEN_26328 : _GEN_21433; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_27955 = io_loadIn_1_valid ? _GEN_26329 : _GEN_21434; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_27956 = io_loadIn_1_valid ? _GEN_26330 : _GEN_21435; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_27957 = io_loadIn_1_valid ? _GEN_26331 : _GEN_21436; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_27958 = io_loadIn_1_valid ? _GEN_26332 : _GEN_21437; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_27959 = io_loadIn_1_valid ? _GEN_26333 : _GEN_21438; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_27960 = io_loadIn_1_valid ? _GEN_26334 : _GEN_21439; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_27961 = io_loadIn_1_valid ? _GEN_26335 : _GEN_21440; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_27962 = io_loadIn_1_valid ? _GEN_26336 : _GEN_21441; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_27963 = io_loadIn_1_valid ? _GEN_26337 : _GEN_21442; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_27964 = io_loadIn_1_valid ? _GEN_26338 : _GEN_21443; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_27965 = io_loadIn_1_valid ? _GEN_26339 : _GEN_21444; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_27966 = io_loadIn_1_valid ? _GEN_26340 : _GEN_21445; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_27967 = io_loadIn_1_valid ? _GEN_26341 : _GEN_21446; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_27968 = io_loadIn_1_valid ? _GEN_26342 : _GEN_21447; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_27969 = io_loadIn_1_valid ? _GEN_26343 : _GEN_21448; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_27970 = io_loadIn_1_valid ? _GEN_26344 : _GEN_21449; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_27971 = io_loadIn_1_valid ? _GEN_26345 : _GEN_21450; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_27972 = io_loadIn_1_valid ? _GEN_26346 : _GEN_21451; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_27973 = io_loadIn_1_valid ? _GEN_26347 : _GEN_21452; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_27974 = io_loadIn_1_valid ? _GEN_26348 : _GEN_21453; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_27975 = io_loadIn_1_valid ? _GEN_26349 : _GEN_21454; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_27976 = io_loadIn_1_valid ? _GEN_26350 : _GEN_21455; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_27977 = io_loadIn_1_valid ? _GEN_26351 : _GEN_21456; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_27978 = io_loadIn_1_valid ? _GEN_26352 : _GEN_21457; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_27979 = io_loadIn_1_valid ? _GEN_26353 : _GEN_21458; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_27980 = io_loadIn_1_valid ? _GEN_26354 : _GEN_21459; // @[LoadQueueFlag.scala 286:31]
  wire  _GEN_27981 = io_loadIn_1_valid ? _GEN_26355 : _GEN_21460; // @[LoadQueueFlag.scala 286:31]
  reg  io_rob_isMMIO_1_REG; // @[LoadQueueFlag.scala 358:32]
  reg [4:0] io_rob_uop_1_REG_robIdx_value; // @[LoadQueueFlag.scala 359:29]
  wire  _GEN_29529 = 4'h1 == deqPtrExt_rvalue ? allocated_1 : allocated_0; // @[]
  wire  _GEN_29530 = 4'h2 == deqPtrExt_rvalue ? allocated_2 : _GEN_29529; // @[]
  wire  _GEN_29531 = 4'h3 == deqPtrExt_rvalue ? allocated_3 : _GEN_29530; // @[]
  wire  _GEN_29532 = 4'h4 == deqPtrExt_rvalue ? allocated_4 : _GEN_29531; // @[]
  wire  _GEN_29533 = 4'h5 == deqPtrExt_rvalue ? allocated_5 : _GEN_29532; // @[]
  wire  _GEN_29534 = 4'h6 == deqPtrExt_rvalue ? allocated_6 : _GEN_29533; // @[]
  wire  _GEN_29535 = 4'h7 == deqPtrExt_rvalue ? allocated_7 : _GEN_29534; // @[]
  wire  _GEN_29536 = 4'h8 == deqPtrExt_rvalue ? allocated_8 : _GEN_29535; // @[]
  wire  _GEN_29537 = 4'h9 == deqPtrExt_rvalue ? allocated_9 : _GEN_29536; // @[]
  wire  _GEN_29538 = 4'ha == deqPtrExt_rvalue ? allocated_10 : _GEN_29537; // @[]
  wire  _GEN_29539 = 4'hb == deqPtrExt_rvalue ? allocated_11 : _GEN_29538; // @[]
  wire  _GEN_29540 = 4'hc == deqPtrExt_rvalue ? allocated_12 : _GEN_29539; // @[]
  wire  _GEN_29541 = 4'hd == deqPtrExt_rvalue ? allocated_13 : _GEN_29540; // @[]
  wire  _GEN_29542 = 4'he == deqPtrExt_rvalue ? allocated_14 : _GEN_29541; // @[]
  wire  lqTailAllocated = 4'hf == deqPtrExt_rvalue ? allocated_15 : _GEN_29542; // @[]
  wire  _GEN_29545 = 4'h1 == deqPtrExt_rvalue ? pending_1 : pending_0; // @[]
  wire  _GEN_29546 = 4'h2 == deqPtrExt_rvalue ? pending_2 : _GEN_29545; // @[]
  wire  _GEN_29547 = 4'h3 == deqPtrExt_rvalue ? pending_3 : _GEN_29546; // @[]
  wire  _GEN_29548 = 4'h4 == deqPtrExt_rvalue ? pending_4 : _GEN_29547; // @[]
  wire  _GEN_29549 = 4'h5 == deqPtrExt_rvalue ? pending_5 : _GEN_29548; // @[]
  wire  _GEN_29550 = 4'h6 == deqPtrExt_rvalue ? pending_6 : _GEN_29549; // @[]
  wire  _GEN_29551 = 4'h7 == deqPtrExt_rvalue ? pending_7 : _GEN_29550; // @[]
  wire  _GEN_29552 = 4'h8 == deqPtrExt_rvalue ? pending_8 : _GEN_29551; // @[]
  wire  _GEN_29553 = 4'h9 == deqPtrExt_rvalue ? pending_9 : _GEN_29552; // @[]
  wire  _GEN_29554 = 4'ha == deqPtrExt_rvalue ? pending_10 : _GEN_29553; // @[]
  wire  _GEN_29555 = 4'hb == deqPtrExt_rvalue ? pending_11 : _GEN_29554; // @[]
  wire  _GEN_29556 = 4'hc == deqPtrExt_rvalue ? pending_12 : _GEN_29555; // @[]
  wire  _GEN_29557 = 4'hd == deqPtrExt_rvalue ? pending_13 : _GEN_29556; // @[]
  wire  _GEN_29558 = 4'he == deqPtrExt_rvalue ? pending_14 : _GEN_29557; // @[]
  wire  lqTailMmioPending = 4'hf == deqPtrExt_rvalue ? pending_15 : _GEN_29558; // @[]
  wire  _GEN_29561 = 4'h1 == deqPtrExt_rvalue ? writebacked_1 : writebacked_0; // @[]
  wire  _GEN_29562 = 4'h2 == deqPtrExt_rvalue ? writebacked_2 : _GEN_29561; // @[]
  wire  _GEN_29563 = 4'h3 == deqPtrExt_rvalue ? writebacked_3 : _GEN_29562; // @[]
  wire  _GEN_29564 = 4'h4 == deqPtrExt_rvalue ? writebacked_4 : _GEN_29563; // @[]
  wire  _GEN_29565 = 4'h5 == deqPtrExt_rvalue ? writebacked_5 : _GEN_29564; // @[]
  wire  _GEN_29566 = 4'h6 == deqPtrExt_rvalue ? writebacked_6 : _GEN_29565; // @[]
  wire  _GEN_29567 = 4'h7 == deqPtrExt_rvalue ? writebacked_7 : _GEN_29566; // @[]
  wire  _GEN_29568 = 4'h8 == deqPtrExt_rvalue ? writebacked_8 : _GEN_29567; // @[]
  wire  _GEN_29569 = 4'h9 == deqPtrExt_rvalue ? writebacked_9 : _GEN_29568; // @[]
  wire  _GEN_29570 = 4'ha == deqPtrExt_rvalue ? writebacked_10 : _GEN_29569; // @[]
  wire  _GEN_29571 = 4'hb == deqPtrExt_rvalue ? writebacked_11 : _GEN_29570; // @[]
  wire  _GEN_29572 = 4'hc == deqPtrExt_rvalue ? writebacked_12 : _GEN_29571; // @[]
  wire  _GEN_29573 = 4'hd == deqPtrExt_rvalue ? writebacked_13 : _GEN_29572; // @[]
  wire  _GEN_29574 = 4'he == deqPtrExt_rvalue ? writebacked_14 : _GEN_29573; // @[]
  wire  lqTailWriteback = 4'hf == deqPtrExt_rvalue ? writebacked_15 : _GEN_29574; // @[]
  reg [1:0] uncacheState; // @[LoadQueueFlag.scala 397:29]
  reg  uncacheCommitFired; // @[LoadQueueFlag.scala 398:35]
  wire  _GEN_29576 = uncacheState == 2'h1 ? 1'h0 : uncacheCommitFired; // @[LoadQueueFlag.scala 400:32 401:24 398:35]
  reg  REG; // @[LoadQueueFlag.scala 406:20]
  wire  _T_55 = io_uncache_req_ready & io_uncache_req_valid; // @[Decoupled.scala 50:35]
  wire  _T_57 = io_uncache_resp_ready & io_uncache_resp_valid; // @[Decoupled.scala 50:35]
  reg  REG_1; // @[LoadQueueFlag.scala 421:20]
  wire [1:0] _GEN_29580 = REG_1 ? 2'h0 : uncacheState; // @[LoadQueueFlag.scala 421:37 422:22 397:29]
  reg [63:0] uncacheData; // @[LoadQueueFlag.scala 455:24]
  wire  _GEN_31509 = 4'h0 == deqPtrExt_rvalue; // @[LoadQueueFlag.scala 457:{23,23}]
  wire  _GEN_29617 = 4'h0 == deqPtrExt_rvalue | _GEN_27934; // @[LoadQueueFlag.scala 457:{23,23}]
  wire  _GEN_31510 = 4'h1 == deqPtrExt_rvalue; // @[LoadQueueFlag.scala 457:{23,23}]
  wire  _GEN_29618 = 4'h1 == deqPtrExt_rvalue | _GEN_27935; // @[LoadQueueFlag.scala 457:{23,23}]
  wire  _GEN_31511 = 4'h2 == deqPtrExt_rvalue; // @[LoadQueueFlag.scala 457:{23,23}]
  wire  _GEN_29619 = 4'h2 == deqPtrExt_rvalue | _GEN_27936; // @[LoadQueueFlag.scala 457:{23,23}]
  wire  _GEN_31512 = 4'h3 == deqPtrExt_rvalue; // @[LoadQueueFlag.scala 457:{23,23}]
  wire  _GEN_29620 = 4'h3 == deqPtrExt_rvalue | _GEN_27937; // @[LoadQueueFlag.scala 457:{23,23}]
  wire  _GEN_31513 = 4'h4 == deqPtrExt_rvalue; // @[LoadQueueFlag.scala 457:{23,23}]
  wire  _GEN_29621 = 4'h4 == deqPtrExt_rvalue | _GEN_27938; // @[LoadQueueFlag.scala 457:{23,23}]
  wire  _GEN_31514 = 4'h5 == deqPtrExt_rvalue; // @[LoadQueueFlag.scala 457:{23,23}]
  wire  _GEN_29622 = 4'h5 == deqPtrExt_rvalue | _GEN_27939; // @[LoadQueueFlag.scala 457:{23,23}]
  wire  _GEN_31515 = 4'h6 == deqPtrExt_rvalue; // @[LoadQueueFlag.scala 457:{23,23}]
  wire  _GEN_29623 = 4'h6 == deqPtrExt_rvalue | _GEN_27940; // @[LoadQueueFlag.scala 457:{23,23}]
  wire  _GEN_31516 = 4'h7 == deqPtrExt_rvalue; // @[LoadQueueFlag.scala 457:{23,23}]
  wire  _GEN_29624 = 4'h7 == deqPtrExt_rvalue | _GEN_27941; // @[LoadQueueFlag.scala 457:{23,23}]
  wire  _GEN_31517 = 4'h8 == deqPtrExt_rvalue; // @[LoadQueueFlag.scala 457:{23,23}]
  wire  _GEN_29625 = 4'h8 == deqPtrExt_rvalue | _GEN_27942; // @[LoadQueueFlag.scala 457:{23,23}]
  wire  _GEN_31518 = 4'h9 == deqPtrExt_rvalue; // @[LoadQueueFlag.scala 457:{23,23}]
  wire  _GEN_29626 = 4'h9 == deqPtrExt_rvalue | _GEN_27943; // @[LoadQueueFlag.scala 457:{23,23}]
  wire  _GEN_31519 = 4'ha == deqPtrExt_rvalue; // @[LoadQueueFlag.scala 457:{23,23}]
  wire  _GEN_29627 = 4'ha == deqPtrExt_rvalue | _GEN_27944; // @[LoadQueueFlag.scala 457:{23,23}]
  wire  _GEN_31520 = 4'hb == deqPtrExt_rvalue; // @[LoadQueueFlag.scala 457:{23,23}]
  wire  _GEN_29628 = 4'hb == deqPtrExt_rvalue | _GEN_27945; // @[LoadQueueFlag.scala 457:{23,23}]
  wire  _GEN_31521 = 4'hc == deqPtrExt_rvalue; // @[LoadQueueFlag.scala 457:{23,23}]
  wire  _GEN_29629 = 4'hc == deqPtrExt_rvalue | _GEN_27946; // @[LoadQueueFlag.scala 457:{23,23}]
  wire  _GEN_31522 = 4'hd == deqPtrExt_rvalue; // @[LoadQueueFlag.scala 457:{23,23}]
  wire  _GEN_29630 = 4'hd == deqPtrExt_rvalue | _GEN_27947; // @[LoadQueueFlag.scala 457:{23,23}]
  wire  _GEN_31523 = 4'he == deqPtrExt_rvalue; // @[LoadQueueFlag.scala 457:{23,23}]
  wire  _GEN_29631 = 4'he == deqPtrExt_rvalue | _GEN_27948; // @[LoadQueueFlag.scala 457:{23,23}]
  wire  _GEN_31524 = 4'hf == deqPtrExt_rvalue; // @[LoadQueueFlag.scala 457:{23,23}]
  wire  _GEN_29632 = 4'hf == deqPtrExt_rvalue | _GEN_27949; // @[LoadQueueFlag.scala 457:{23,23}]
  wire  _GEN_29651 = 4'h1 == deqPtrExt_rvalue ? uop_1_ctrl_fpWen : uop_0_ctrl_fpWen; // @[LoadQueue.scala 59:{28,28}]
  wire  _GEN_29652 = 4'h2 == deqPtrExt_rvalue ? uop_2_ctrl_fpWen : _GEN_29651; // @[LoadQueue.scala 59:{28,28}]
  wire  _GEN_29653 = 4'h3 == deqPtrExt_rvalue ? uop_3_ctrl_fpWen : _GEN_29652; // @[LoadQueue.scala 59:{28,28}]
  wire  _GEN_29654 = 4'h4 == deqPtrExt_rvalue ? uop_4_ctrl_fpWen : _GEN_29653; // @[LoadQueue.scala 59:{28,28}]
  wire  _GEN_29655 = 4'h5 == deqPtrExt_rvalue ? uop_5_ctrl_fpWen : _GEN_29654; // @[LoadQueue.scala 59:{28,28}]
  wire  _GEN_29656 = 4'h6 == deqPtrExt_rvalue ? uop_6_ctrl_fpWen : _GEN_29655; // @[LoadQueue.scala 59:{28,28}]
  wire  _GEN_29657 = 4'h7 == deqPtrExt_rvalue ? uop_7_ctrl_fpWen : _GEN_29656; // @[LoadQueue.scala 59:{28,28}]
  wire  _GEN_29658 = 4'h8 == deqPtrExt_rvalue ? uop_8_ctrl_fpWen : _GEN_29657; // @[LoadQueue.scala 59:{28,28}]
  wire  _GEN_29659 = 4'h9 == deqPtrExt_rvalue ? uop_9_ctrl_fpWen : _GEN_29658; // @[LoadQueue.scala 59:{28,28}]
  wire  _GEN_29660 = 4'ha == deqPtrExt_rvalue ? uop_10_ctrl_fpWen : _GEN_29659; // @[LoadQueue.scala 59:{28,28}]
  wire  _GEN_29661 = 4'hb == deqPtrExt_rvalue ? uop_11_ctrl_fpWen : _GEN_29660; // @[LoadQueue.scala 59:{28,28}]
  wire  _GEN_29662 = 4'hc == deqPtrExt_rvalue ? uop_12_ctrl_fpWen : _GEN_29661; // @[LoadQueue.scala 59:{28,28}]
  wire  _GEN_29663 = 4'hd == deqPtrExt_rvalue ? uop_13_ctrl_fpWen : _GEN_29662; // @[LoadQueue.scala 59:{28,28}]
  wire  _GEN_29664 = 4'he == deqPtrExt_rvalue ? uop_14_ctrl_fpWen : _GEN_29663; // @[LoadQueue.scala 59:{28,28}]
  wire [6:0] _GEN_29667 = 4'h1 == deqPtrExt_rvalue ? uop_1_ctrl_fuOpType : uop_0_ctrl_fuOpType; // @[LookupTree.scala 24:{34,34}]
  wire [6:0] _GEN_29668 = 4'h2 == deqPtrExt_rvalue ? uop_2_ctrl_fuOpType : _GEN_29667; // @[LookupTree.scala 24:{34,34}]
  wire [6:0] _GEN_29669 = 4'h3 == deqPtrExt_rvalue ? uop_3_ctrl_fuOpType : _GEN_29668; // @[LookupTree.scala 24:{34,34}]
  wire [6:0] _GEN_29670 = 4'h4 == deqPtrExt_rvalue ? uop_4_ctrl_fuOpType : _GEN_29669; // @[LookupTree.scala 24:{34,34}]
  wire [6:0] _GEN_29671 = 4'h5 == deqPtrExt_rvalue ? uop_5_ctrl_fuOpType : _GEN_29670; // @[LookupTree.scala 24:{34,34}]
  wire [6:0] _GEN_29672 = 4'h6 == deqPtrExt_rvalue ? uop_6_ctrl_fuOpType : _GEN_29671; // @[LookupTree.scala 24:{34,34}]
  wire [6:0] _GEN_29673 = 4'h7 == deqPtrExt_rvalue ? uop_7_ctrl_fuOpType : _GEN_29672; // @[LookupTree.scala 24:{34,34}]
  wire [6:0] _GEN_29674 = 4'h8 == deqPtrExt_rvalue ? uop_8_ctrl_fuOpType : _GEN_29673; // @[LookupTree.scala 24:{34,34}]
  wire [6:0] _GEN_29675 = 4'h9 == deqPtrExt_rvalue ? uop_9_ctrl_fuOpType : _GEN_29674; // @[LookupTree.scala 24:{34,34}]
  wire [6:0] _GEN_29676 = 4'ha == deqPtrExt_rvalue ? uop_10_ctrl_fuOpType : _GEN_29675; // @[LookupTree.scala 24:{34,34}]
  wire [6:0] _GEN_29677 = 4'hb == deqPtrExt_rvalue ? uop_11_ctrl_fuOpType : _GEN_29676; // @[LookupTree.scala 24:{34,34}]
  wire [6:0] _GEN_29678 = 4'hc == deqPtrExt_rvalue ? uop_12_ctrl_fuOpType : _GEN_29677; // @[LookupTree.scala 24:{34,34}]
  wire [6:0] _GEN_29679 = 4'hd == deqPtrExt_rvalue ? uop_13_ctrl_fuOpType : _GEN_29678; // @[LookupTree.scala 24:{34,34}]
  wire [6:0] _GEN_29680 = 4'he == deqPtrExt_rvalue ? uop_14_ctrl_fuOpType : _GEN_29679; // @[LookupTree.scala 24:{34,34}]
  wire  _GEN_29795 = 4'h1 == deqPtrExt_rvalue ? uop_1_cf_exceptionVec_4 : uop_0_cf_exceptionVec_4; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_29796 = 4'h2 == deqPtrExt_rvalue ? uop_2_cf_exceptionVec_4 : _GEN_29795; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_29797 = 4'h3 == deqPtrExt_rvalue ? uop_3_cf_exceptionVec_4 : _GEN_29796; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_29798 = 4'h4 == deqPtrExt_rvalue ? uop_4_cf_exceptionVec_4 : _GEN_29797; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_29799 = 4'h5 == deqPtrExt_rvalue ? uop_5_cf_exceptionVec_4 : _GEN_29798; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_29800 = 4'h6 == deqPtrExt_rvalue ? uop_6_cf_exceptionVec_4 : _GEN_29799; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_29801 = 4'h7 == deqPtrExt_rvalue ? uop_7_cf_exceptionVec_4 : _GEN_29800; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_29802 = 4'h8 == deqPtrExt_rvalue ? uop_8_cf_exceptionVec_4 : _GEN_29801; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_29803 = 4'h9 == deqPtrExt_rvalue ? uop_9_cf_exceptionVec_4 : _GEN_29802; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_29804 = 4'ha == deqPtrExt_rvalue ? uop_10_cf_exceptionVec_4 : _GEN_29803; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_29805 = 4'hb == deqPtrExt_rvalue ? uop_11_cf_exceptionVec_4 : _GEN_29804; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_29806 = 4'hc == deqPtrExt_rvalue ? uop_12_cf_exceptionVec_4 : _GEN_29805; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_29807 = 4'hd == deqPtrExt_rvalue ? uop_13_cf_exceptionVec_4 : _GEN_29806; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_29808 = 4'he == deqPtrExt_rvalue ? uop_14_cf_exceptionVec_4 : _GEN_29807; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_29811 = 4'h1 == deqPtrExt_rvalue ? uop_1_cf_exceptionVec_5 : uop_0_cf_exceptionVec_5; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_29812 = 4'h2 == deqPtrExt_rvalue ? uop_2_cf_exceptionVec_5 : _GEN_29811; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_29813 = 4'h3 == deqPtrExt_rvalue ? uop_3_cf_exceptionVec_5 : _GEN_29812; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_29814 = 4'h4 == deqPtrExt_rvalue ? uop_4_cf_exceptionVec_5 : _GEN_29813; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_29815 = 4'h5 == deqPtrExt_rvalue ? uop_5_cf_exceptionVec_5 : _GEN_29814; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_29816 = 4'h6 == deqPtrExt_rvalue ? uop_6_cf_exceptionVec_5 : _GEN_29815; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_29817 = 4'h7 == deqPtrExt_rvalue ? uop_7_cf_exceptionVec_5 : _GEN_29816; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_29818 = 4'h8 == deqPtrExt_rvalue ? uop_8_cf_exceptionVec_5 : _GEN_29817; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_29819 = 4'h9 == deqPtrExt_rvalue ? uop_9_cf_exceptionVec_5 : _GEN_29818; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_29820 = 4'ha == deqPtrExt_rvalue ? uop_10_cf_exceptionVec_5 : _GEN_29819; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_29821 = 4'hb == deqPtrExt_rvalue ? uop_11_cf_exceptionVec_5 : _GEN_29820; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_29822 = 4'hc == deqPtrExt_rvalue ? uop_12_cf_exceptionVec_5 : _GEN_29821; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_29823 = 4'hd == deqPtrExt_rvalue ? uop_13_cf_exceptionVec_5 : _GEN_29822; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_29824 = 4'he == deqPtrExt_rvalue ? uop_14_cf_exceptionVec_5 : _GEN_29823; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_29939 = 4'h1 == deqPtrExt_rvalue ? uop_1_cf_exceptionVec_13 : uop_0_cf_exceptionVec_13; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_29940 = 4'h2 == deqPtrExt_rvalue ? uop_2_cf_exceptionVec_13 : _GEN_29939; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_29941 = 4'h3 == deqPtrExt_rvalue ? uop_3_cf_exceptionVec_13 : _GEN_29940; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_29942 = 4'h4 == deqPtrExt_rvalue ? uop_4_cf_exceptionVec_13 : _GEN_29941; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_29943 = 4'h5 == deqPtrExt_rvalue ? uop_5_cf_exceptionVec_13 : _GEN_29942; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_29944 = 4'h6 == deqPtrExt_rvalue ? uop_6_cf_exceptionVec_13 : _GEN_29943; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_29945 = 4'h7 == deqPtrExt_rvalue ? uop_7_cf_exceptionVec_13 : _GEN_29944; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_29946 = 4'h8 == deqPtrExt_rvalue ? uop_8_cf_exceptionVec_13 : _GEN_29945; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_29947 = 4'h9 == deqPtrExt_rvalue ? uop_9_cf_exceptionVec_13 : _GEN_29946; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_29948 = 4'ha == deqPtrExt_rvalue ? uop_10_cf_exceptionVec_13 : _GEN_29947; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_29949 = 4'hb == deqPtrExt_rvalue ? uop_11_cf_exceptionVec_13 : _GEN_29948; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_29950 = 4'hc == deqPtrExt_rvalue ? uop_12_cf_exceptionVec_13 : _GEN_29949; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_29951 = 4'hd == deqPtrExt_rvalue ? uop_13_cf_exceptionVec_13 : _GEN_29950; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_29952 = 4'he == deqPtrExt_rvalue ? uop_14_cf_exceptionVec_13 : _GEN_29951; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30067 = 4'h1 == deqPtrExt_rvalue ? uop_1_cf_trigger_backendEn_1 : uop_0_cf_trigger_backendEn_1; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30068 = 4'h2 == deqPtrExt_rvalue ? uop_2_cf_trigger_backendEn_1 : _GEN_30067; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30069 = 4'h3 == deqPtrExt_rvalue ? uop_3_cf_trigger_backendEn_1 : _GEN_30068; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30070 = 4'h4 == deqPtrExt_rvalue ? uop_4_cf_trigger_backendEn_1 : _GEN_30069; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30071 = 4'h5 == deqPtrExt_rvalue ? uop_5_cf_trigger_backendEn_1 : _GEN_30070; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30072 = 4'h6 == deqPtrExt_rvalue ? uop_6_cf_trigger_backendEn_1 : _GEN_30071; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30073 = 4'h7 == deqPtrExt_rvalue ? uop_7_cf_trigger_backendEn_1 : _GEN_30072; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30074 = 4'h8 == deqPtrExt_rvalue ? uop_8_cf_trigger_backendEn_1 : _GEN_30073; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30075 = 4'h9 == deqPtrExt_rvalue ? uop_9_cf_trigger_backendEn_1 : _GEN_30074; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30076 = 4'ha == deqPtrExt_rvalue ? uop_10_cf_trigger_backendEn_1 : _GEN_30075; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30077 = 4'hb == deqPtrExt_rvalue ? uop_11_cf_trigger_backendEn_1 : _GEN_30076; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30078 = 4'hc == deqPtrExt_rvalue ? uop_12_cf_trigger_backendEn_1 : _GEN_30077; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30079 = 4'hd == deqPtrExt_rvalue ? uop_13_cf_trigger_backendEn_1 : _GEN_30078; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30080 = 4'he == deqPtrExt_rvalue ? uop_14_cf_trigger_backendEn_1 : _GEN_30079; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30083 = 4'h1 == deqPtrExt_rvalue ? uop_1_cf_trigger_backendHit_0 : uop_0_cf_trigger_backendHit_0; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30084 = 4'h2 == deqPtrExt_rvalue ? uop_2_cf_trigger_backendHit_0 : _GEN_30083; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30085 = 4'h3 == deqPtrExt_rvalue ? uop_3_cf_trigger_backendHit_0 : _GEN_30084; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30086 = 4'h4 == deqPtrExt_rvalue ? uop_4_cf_trigger_backendHit_0 : _GEN_30085; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30087 = 4'h5 == deqPtrExt_rvalue ? uop_5_cf_trigger_backendHit_0 : _GEN_30086; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30088 = 4'h6 == deqPtrExt_rvalue ? uop_6_cf_trigger_backendHit_0 : _GEN_30087; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30089 = 4'h7 == deqPtrExt_rvalue ? uop_7_cf_trigger_backendHit_0 : _GEN_30088; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30090 = 4'h8 == deqPtrExt_rvalue ? uop_8_cf_trigger_backendHit_0 : _GEN_30089; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30091 = 4'h9 == deqPtrExt_rvalue ? uop_9_cf_trigger_backendHit_0 : _GEN_30090; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30092 = 4'ha == deqPtrExt_rvalue ? uop_10_cf_trigger_backendHit_0 : _GEN_30091; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30093 = 4'hb == deqPtrExt_rvalue ? uop_11_cf_trigger_backendHit_0 : _GEN_30092; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30094 = 4'hc == deqPtrExt_rvalue ? uop_12_cf_trigger_backendHit_0 : _GEN_30093; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30095 = 4'hd == deqPtrExt_rvalue ? uop_13_cf_trigger_backendHit_0 : _GEN_30094; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30096 = 4'he == deqPtrExt_rvalue ? uop_14_cf_trigger_backendHit_0 : _GEN_30095; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30099 = 4'h1 == deqPtrExt_rvalue ? uop_1_cf_trigger_backendHit_1 : uop_0_cf_trigger_backendHit_1; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30100 = 4'h2 == deqPtrExt_rvalue ? uop_2_cf_trigger_backendHit_1 : _GEN_30099; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30101 = 4'h3 == deqPtrExt_rvalue ? uop_3_cf_trigger_backendHit_1 : _GEN_30100; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30102 = 4'h4 == deqPtrExt_rvalue ? uop_4_cf_trigger_backendHit_1 : _GEN_30101; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30103 = 4'h5 == deqPtrExt_rvalue ? uop_5_cf_trigger_backendHit_1 : _GEN_30102; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30104 = 4'h6 == deqPtrExt_rvalue ? uop_6_cf_trigger_backendHit_1 : _GEN_30103; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30105 = 4'h7 == deqPtrExt_rvalue ? uop_7_cf_trigger_backendHit_1 : _GEN_30104; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30106 = 4'h8 == deqPtrExt_rvalue ? uop_8_cf_trigger_backendHit_1 : _GEN_30105; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30107 = 4'h9 == deqPtrExt_rvalue ? uop_9_cf_trigger_backendHit_1 : _GEN_30106; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30108 = 4'ha == deqPtrExt_rvalue ? uop_10_cf_trigger_backendHit_1 : _GEN_30107; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30109 = 4'hb == deqPtrExt_rvalue ? uop_11_cf_trigger_backendHit_1 : _GEN_30108; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30110 = 4'hc == deqPtrExt_rvalue ? uop_12_cf_trigger_backendHit_1 : _GEN_30109; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30111 = 4'hd == deqPtrExt_rvalue ? uop_13_cf_trigger_backendHit_1 : _GEN_30110; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30112 = 4'he == deqPtrExt_rvalue ? uop_14_cf_trigger_backendHit_1 : _GEN_30111; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30147 = 4'h1 == deqPtrExt_rvalue ? uop_1_cf_trigger_backendHit_4 : uop_0_cf_trigger_backendHit_4; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30148 = 4'h2 == deqPtrExt_rvalue ? uop_2_cf_trigger_backendHit_4 : _GEN_30147; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30149 = 4'h3 == deqPtrExt_rvalue ? uop_3_cf_trigger_backendHit_4 : _GEN_30148; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30150 = 4'h4 == deqPtrExt_rvalue ? uop_4_cf_trigger_backendHit_4 : _GEN_30149; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30151 = 4'h5 == deqPtrExt_rvalue ? uop_5_cf_trigger_backendHit_4 : _GEN_30150; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30152 = 4'h6 == deqPtrExt_rvalue ? uop_6_cf_trigger_backendHit_4 : _GEN_30151; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30153 = 4'h7 == deqPtrExt_rvalue ? uop_7_cf_trigger_backendHit_4 : _GEN_30152; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30154 = 4'h8 == deqPtrExt_rvalue ? uop_8_cf_trigger_backendHit_4 : _GEN_30153; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30155 = 4'h9 == deqPtrExt_rvalue ? uop_9_cf_trigger_backendHit_4 : _GEN_30154; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30156 = 4'ha == deqPtrExt_rvalue ? uop_10_cf_trigger_backendHit_4 : _GEN_30155; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30157 = 4'hb == deqPtrExt_rvalue ? uop_11_cf_trigger_backendHit_4 : _GEN_30156; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30158 = 4'hc == deqPtrExt_rvalue ? uop_12_cf_trigger_backendHit_4 : _GEN_30157; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30159 = 4'hd == deqPtrExt_rvalue ? uop_13_cf_trigger_backendHit_4 : _GEN_30158; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30160 = 4'he == deqPtrExt_rvalue ? uop_14_cf_trigger_backendHit_4 : _GEN_30159; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30579 = 4'h1 == deqPtrExt_rvalue ? uop_1_ctrl_rfWen : uop_0_ctrl_rfWen; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30580 = 4'h2 == deqPtrExt_rvalue ? uop_2_ctrl_rfWen : _GEN_30579; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30581 = 4'h3 == deqPtrExt_rvalue ? uop_3_ctrl_rfWen : _GEN_30580; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30582 = 4'h4 == deqPtrExt_rvalue ? uop_4_ctrl_rfWen : _GEN_30581; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30583 = 4'h5 == deqPtrExt_rvalue ? uop_5_ctrl_rfWen : _GEN_30582; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30584 = 4'h6 == deqPtrExt_rvalue ? uop_6_ctrl_rfWen : _GEN_30583; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30585 = 4'h7 == deqPtrExt_rvalue ? uop_7_ctrl_rfWen : _GEN_30584; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30586 = 4'h8 == deqPtrExt_rvalue ? uop_8_ctrl_rfWen : _GEN_30585; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30587 = 4'h9 == deqPtrExt_rvalue ? uop_9_ctrl_rfWen : _GEN_30586; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30588 = 4'ha == deqPtrExt_rvalue ? uop_10_ctrl_rfWen : _GEN_30587; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30589 = 4'hb == deqPtrExt_rvalue ? uop_11_ctrl_rfWen : _GEN_30588; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30590 = 4'hc == deqPtrExt_rvalue ? uop_12_ctrl_rfWen : _GEN_30589; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30591 = 4'hd == deqPtrExt_rvalue ? uop_13_ctrl_rfWen : _GEN_30590; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30592 = 4'he == deqPtrExt_rvalue ? uop_14_ctrl_rfWen : _GEN_30591; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30643 = 4'h1 == deqPtrExt_rvalue ? uop_1_ctrl_flushPipe : uop_0_ctrl_flushPipe; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30644 = 4'h2 == deqPtrExt_rvalue ? uop_2_ctrl_flushPipe : _GEN_30643; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30645 = 4'h3 == deqPtrExt_rvalue ? uop_3_ctrl_flushPipe : _GEN_30644; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30646 = 4'h4 == deqPtrExt_rvalue ? uop_4_ctrl_flushPipe : _GEN_30645; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30647 = 4'h5 == deqPtrExt_rvalue ? uop_5_ctrl_flushPipe : _GEN_30646; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30648 = 4'h6 == deqPtrExt_rvalue ? uop_6_ctrl_flushPipe : _GEN_30647; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30649 = 4'h7 == deqPtrExt_rvalue ? uop_7_ctrl_flushPipe : _GEN_30648; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30650 = 4'h8 == deqPtrExt_rvalue ? uop_8_ctrl_flushPipe : _GEN_30649; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30651 = 4'h9 == deqPtrExt_rvalue ? uop_9_ctrl_flushPipe : _GEN_30650; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30652 = 4'ha == deqPtrExt_rvalue ? uop_10_ctrl_flushPipe : _GEN_30651; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30653 = 4'hb == deqPtrExt_rvalue ? uop_11_ctrl_flushPipe : _GEN_30652; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30654 = 4'hc == deqPtrExt_rvalue ? uop_12_ctrl_flushPipe : _GEN_30653; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30655 = 4'hd == deqPtrExt_rvalue ? uop_13_ctrl_flushPipe : _GEN_30654; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30656 = 4'he == deqPtrExt_rvalue ? uop_14_ctrl_flushPipe : _GEN_30655; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30963 = 4'h1 == deqPtrExt_rvalue ? uop_1_ctrl_replayInst : uop_0_ctrl_replayInst; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30964 = 4'h2 == deqPtrExt_rvalue ? uop_2_ctrl_replayInst : _GEN_30963; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30965 = 4'h3 == deqPtrExt_rvalue ? uop_3_ctrl_replayInst : _GEN_30964; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30966 = 4'h4 == deqPtrExt_rvalue ? uop_4_ctrl_replayInst : _GEN_30965; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30967 = 4'h5 == deqPtrExt_rvalue ? uop_5_ctrl_replayInst : _GEN_30966; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30968 = 4'h6 == deqPtrExt_rvalue ? uop_6_ctrl_replayInst : _GEN_30967; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30969 = 4'h7 == deqPtrExt_rvalue ? uop_7_ctrl_replayInst : _GEN_30968; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30970 = 4'h8 == deqPtrExt_rvalue ? uop_8_ctrl_replayInst : _GEN_30969; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30971 = 4'h9 == deqPtrExt_rvalue ? uop_9_ctrl_replayInst : _GEN_30970; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30972 = 4'ha == deqPtrExt_rvalue ? uop_10_ctrl_replayInst : _GEN_30971; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30973 = 4'hb == deqPtrExt_rvalue ? uop_11_ctrl_replayInst : _GEN_30972; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30974 = 4'hc == deqPtrExt_rvalue ? uop_12_ctrl_replayInst : _GEN_30973; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30975 = 4'hd == deqPtrExt_rvalue ? uop_13_ctrl_replayInst : _GEN_30974; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_30976 = 4'he == deqPtrExt_rvalue ? uop_14_ctrl_replayInst : _GEN_30975; // @[LoadQueueFlag.scala 480:{26,26}]
  wire [5:0] _GEN_31075 = 4'h1 == deqPtrExt_rvalue ? uop_1_pdest : uop_0_pdest; // @[LoadQueueFlag.scala 480:{26,26}]
  wire [5:0] _GEN_31076 = 4'h2 == deqPtrExt_rvalue ? uop_2_pdest : _GEN_31075; // @[LoadQueueFlag.scala 480:{26,26}]
  wire [5:0] _GEN_31077 = 4'h3 == deqPtrExt_rvalue ? uop_3_pdest : _GEN_31076; // @[LoadQueueFlag.scala 480:{26,26}]
  wire [5:0] _GEN_31078 = 4'h4 == deqPtrExt_rvalue ? uop_4_pdest : _GEN_31077; // @[LoadQueueFlag.scala 480:{26,26}]
  wire [5:0] _GEN_31079 = 4'h5 == deqPtrExt_rvalue ? uop_5_pdest : _GEN_31078; // @[LoadQueueFlag.scala 480:{26,26}]
  wire [5:0] _GEN_31080 = 4'h6 == deqPtrExt_rvalue ? uop_6_pdest : _GEN_31079; // @[LoadQueueFlag.scala 480:{26,26}]
  wire [5:0] _GEN_31081 = 4'h7 == deqPtrExt_rvalue ? uop_7_pdest : _GEN_31080; // @[LoadQueueFlag.scala 480:{26,26}]
  wire [5:0] _GEN_31082 = 4'h8 == deqPtrExt_rvalue ? uop_8_pdest : _GEN_31081; // @[LoadQueueFlag.scala 480:{26,26}]
  wire [5:0] _GEN_31083 = 4'h9 == deqPtrExt_rvalue ? uop_9_pdest : _GEN_31082; // @[LoadQueueFlag.scala 480:{26,26}]
  wire [5:0] _GEN_31084 = 4'ha == deqPtrExt_rvalue ? uop_10_pdest : _GEN_31083; // @[LoadQueueFlag.scala 480:{26,26}]
  wire [5:0] _GEN_31085 = 4'hb == deqPtrExt_rvalue ? uop_11_pdest : _GEN_31084; // @[LoadQueueFlag.scala 480:{26,26}]
  wire [5:0] _GEN_31086 = 4'hc == deqPtrExt_rvalue ? uop_12_pdest : _GEN_31085; // @[LoadQueueFlag.scala 480:{26,26}]
  wire [5:0] _GEN_31087 = 4'hd == deqPtrExt_rvalue ? uop_13_pdest : _GEN_31086; // @[LoadQueueFlag.scala 480:{26,26}]
  wire [5:0] _GEN_31088 = 4'he == deqPtrExt_rvalue ? uop_14_pdest : _GEN_31087; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_31107 = 4'h1 == deqPtrExt_rvalue ? uop_1_robIdx_flag : uop_0_robIdx_flag; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_31108 = 4'h2 == deqPtrExt_rvalue ? uop_2_robIdx_flag : _GEN_31107; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_31109 = 4'h3 == deqPtrExt_rvalue ? uop_3_robIdx_flag : _GEN_31108; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_31110 = 4'h4 == deqPtrExt_rvalue ? uop_4_robIdx_flag : _GEN_31109; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_31111 = 4'h5 == deqPtrExt_rvalue ? uop_5_robIdx_flag : _GEN_31110; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_31112 = 4'h6 == deqPtrExt_rvalue ? uop_6_robIdx_flag : _GEN_31111; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_31113 = 4'h7 == deqPtrExt_rvalue ? uop_7_robIdx_flag : _GEN_31112; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_31114 = 4'h8 == deqPtrExt_rvalue ? uop_8_robIdx_flag : _GEN_31113; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_31115 = 4'h9 == deqPtrExt_rvalue ? uop_9_robIdx_flag : _GEN_31114; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_31116 = 4'ha == deqPtrExt_rvalue ? uop_10_robIdx_flag : _GEN_31115; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_31117 = 4'hb == deqPtrExt_rvalue ? uop_11_robIdx_flag : _GEN_31116; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_31118 = 4'hc == deqPtrExt_rvalue ? uop_12_robIdx_flag : _GEN_31117; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_31119 = 4'hd == deqPtrExt_rvalue ? uop_13_robIdx_flag : _GEN_31118; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _GEN_31120 = 4'he == deqPtrExt_rvalue ? uop_14_robIdx_flag : _GEN_31119; // @[LoadQueueFlag.scala 480:{26,26}]
  wire [4:0] _GEN_31123 = 4'h1 == deqPtrExt_rvalue ? uop_1_robIdx_value : uop_0_robIdx_value; // @[LoadQueueFlag.scala 480:{26,26}]
  wire [4:0] _GEN_31124 = 4'h2 == deqPtrExt_rvalue ? uop_2_robIdx_value : _GEN_31123; // @[LoadQueueFlag.scala 480:{26,26}]
  wire [4:0] _GEN_31125 = 4'h3 == deqPtrExt_rvalue ? uop_3_robIdx_value : _GEN_31124; // @[LoadQueueFlag.scala 480:{26,26}]
  wire [4:0] _GEN_31126 = 4'h4 == deqPtrExt_rvalue ? uop_4_robIdx_value : _GEN_31125; // @[LoadQueueFlag.scala 480:{26,26}]
  wire [4:0] _GEN_31127 = 4'h5 == deqPtrExt_rvalue ? uop_5_robIdx_value : _GEN_31126; // @[LoadQueueFlag.scala 480:{26,26}]
  wire [4:0] _GEN_31128 = 4'h6 == deqPtrExt_rvalue ? uop_6_robIdx_value : _GEN_31127; // @[LoadQueueFlag.scala 480:{26,26}]
  wire [4:0] _GEN_31129 = 4'h7 == deqPtrExt_rvalue ? uop_7_robIdx_value : _GEN_31128; // @[LoadQueueFlag.scala 480:{26,26}]
  wire [4:0] _GEN_31130 = 4'h8 == deqPtrExt_rvalue ? uop_8_robIdx_value : _GEN_31129; // @[LoadQueueFlag.scala 480:{26,26}]
  wire [4:0] _GEN_31131 = 4'h9 == deqPtrExt_rvalue ? uop_9_robIdx_value : _GEN_31130; // @[LoadQueueFlag.scala 480:{26,26}]
  wire [4:0] _GEN_31132 = 4'ha == deqPtrExt_rvalue ? uop_10_robIdx_value : _GEN_31131; // @[LoadQueueFlag.scala 480:{26,26}]
  wire [4:0] _GEN_31133 = 4'hb == deqPtrExt_rvalue ? uop_11_robIdx_value : _GEN_31132; // @[LoadQueueFlag.scala 480:{26,26}]
  wire [4:0] _GEN_31134 = 4'hc == deqPtrExt_rvalue ? uop_12_robIdx_value : _GEN_31133; // @[LoadQueueFlag.scala 480:{26,26}]
  wire [4:0] _GEN_31135 = 4'hd == deqPtrExt_rvalue ? uop_13_robIdx_value : _GEN_31134; // @[LoadQueueFlag.scala 480:{26,26}]
  wire [4:0] _GEN_31136 = 4'he == deqPtrExt_rvalue ? uop_14_robIdx_value : _GEN_31135; // @[LoadQueueFlag.scala 480:{26,26}]
  wire  _T_61 = io_loadOut_0_ready & io_loadOut_0_valid; // @[Decoupled.scala 50:35]
  wire  _GEN_31394 = _GEN_31509 | _GEN_27966; // @[LoadQueueFlag.scala 502:{25,25}]
  wire  _GEN_31395 = _GEN_31510 | _GEN_27967; // @[LoadQueueFlag.scala 502:{25,25}]
  wire  _GEN_31396 = _GEN_31511 | _GEN_27968; // @[LoadQueueFlag.scala 502:{25,25}]
  wire  _GEN_31397 = _GEN_31512 | _GEN_27969; // @[LoadQueueFlag.scala 502:{25,25}]
  wire  _GEN_31398 = _GEN_31513 | _GEN_27970; // @[LoadQueueFlag.scala 502:{25,25}]
  wire  _GEN_31399 = _GEN_31514 | _GEN_27971; // @[LoadQueueFlag.scala 502:{25,25}]
  wire  _GEN_31400 = _GEN_31515 | _GEN_27972; // @[LoadQueueFlag.scala 502:{25,25}]
  wire  _GEN_31401 = _GEN_31516 | _GEN_27973; // @[LoadQueueFlag.scala 502:{25,25}]
  wire  _GEN_31402 = _GEN_31517 | _GEN_27974; // @[LoadQueueFlag.scala 502:{25,25}]
  wire  _GEN_31403 = _GEN_31518 | _GEN_27975; // @[LoadQueueFlag.scala 502:{25,25}]
  wire  _GEN_31404 = _GEN_31519 | _GEN_27976; // @[LoadQueueFlag.scala 502:{25,25}]
  wire  _GEN_31405 = _GEN_31520 | _GEN_27977; // @[LoadQueueFlag.scala 502:{25,25}]
  wire  _GEN_31406 = _GEN_31521 | _GEN_27978; // @[LoadQueueFlag.scala 502:{25,25}]
  wire  _GEN_31407 = _GEN_31522 | _GEN_27979; // @[LoadQueueFlag.scala 502:{25,25}]
  wire  _GEN_31408 = _GEN_31523 | _GEN_27980; // @[LoadQueueFlag.scala 502:{25,25}]
  wire  _GEN_31409 = _GEN_31524 | _GEN_27981; // @[LoadQueueFlag.scala 502:{25,25}]
  wire  _T_68 = ~io_loadOut_0_ready; // @[LoadQueueFlag.scala 523:69]
  reg  io_perf_0_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg  io_perf_0_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  reg  io_perf_1_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg  io_perf_1_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  reg  io_perf_2_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg  io_perf_2_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  reg  io_perf_3_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg  io_perf_3_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  LqVAddrModule_1 vaddrModule ( // @[LoadQueueFlag.scala 63:27]
    .clock(vaddrModule_clock),
    .io_raddr_1(vaddrModule_io_raddr_1),
    .io_rdata_1(vaddrModule_io_rdata_1),
    .io_wen_0(vaddrModule_io_wen_0),
    .io_wen_1(vaddrModule_io_wen_1),
    .io_waddr_0(vaddrModule_io_waddr_0),
    .io_waddr_1(vaddrModule_io_waddr_1),
    .io_wdata_0(vaddrModule_io_wdata_0),
    .io_wdata_1(vaddrModule_io_wdata_1)
  );
  LqPAddrModule_2 paddrModule ( // @[LoadQueueFlag.scala 72:27]
    .clock(paddrModule_clock),
    .io_raddr_0(paddrModule_io_raddr_0),
    .io_rdata_0(paddrModule_io_rdata_0),
    .io_wen_0(paddrModule_io_wen_0),
    .io_wen_1(paddrModule_io_wen_1),
    .io_waddr_0(paddrModule_io_waddr_0),
    .io_waddr_1(paddrModule_io_waddr_1),
    .io_wdata_0(paddrModule_io_wdata_0),
    .io_wdata_1(paddrModule_io_wdata_1)
  );
  LqMaskModule_1 maskModule ( // @[LoadQueueFlag.scala 81:26]
    .clock(maskModule_clock),
    .io_raddr_0(maskModule_io_raddr_0),
    .io_rdata_0(maskModule_io_rdata_0),
    .io_wen_0(maskModule_io_wen_0),
    .io_wen_1(maskModule_io_wen_1),
    .io_waddr_0(maskModule_io_waddr_0),
    .io_waddr_1(maskModule_io_waddr_1),
    .io_wdata_0(maskModule_io_wdata_0),
    .io_wdata_1(maskModule_io_wdata_1)
  );
  LqTriggerResultModule vaddrTriggerResultModule ( // @[LoadQueueFlag.scala 105:40]
    .clock(vaddrTriggerResultModule_clock),
    .io_raddr_0(vaddrTriggerResultModule_io_raddr_0),
    .io_rdata_0_0(vaddrTriggerResultModule_io_rdata_0_0),
    .io_rdata_0_1(vaddrTriggerResultModule_io_rdata_0_1),
    .io_rdata_0_2(vaddrTriggerResultModule_io_rdata_0_2),
    .io_wen_0(vaddrTriggerResultModule_io_wen_0),
    .io_wen_1(vaddrTriggerResultModule_io_wen_1),
    .io_waddr_0(vaddrTriggerResultModule_io_waddr_0),
    .io_waddr_1(vaddrTriggerResultModule_io_waddr_1),
    .io_wdata_0_0(vaddrTriggerResultModule_io_wdata_0_0),
    .io_wdata_0_1(vaddrTriggerResultModule_io_wdata_0_1),
    .io_wdata_0_2(vaddrTriggerResultModule_io_wdata_0_2),
    .io_wdata_1_0(vaddrTriggerResultModule_io_wdata_1_0),
    .io_wdata_1_1(vaddrTriggerResultModule_io_wdata_1_1),
    .io_wdata_1_2(vaddrTriggerResultModule_io_wdata_1_2)
  );
  assign io_enq_canAccept = validCount <= 5'he; // @[LoadQueueFlag.scala 130:33]
  assign io_loadOut_0_valid = uncacheState == 2'h3 & ~uncacheCommitFired; // @[LoadQueueFlag.scala 478:52]
  assign io_loadOut_0_bits_uop_cf_exceptionVec_4 = 4'hf == deqPtrExt_rvalue ? uop_15_cf_exceptionVec_4 : _GEN_29808; // @[LoadQueueFlag.scala 480:{26,26}]
  assign io_loadOut_0_bits_uop_cf_exceptionVec_5 = 4'hf == deqPtrExt_rvalue ? uop_15_cf_exceptionVec_5 : _GEN_29824; // @[LoadQueueFlag.scala 480:{26,26}]
  assign io_loadOut_0_bits_uop_cf_exceptionVec_13 = 4'hf == deqPtrExt_rvalue ? uop_15_cf_exceptionVec_13 : _GEN_29952; // @[LoadQueueFlag.scala 480:{26,26}]
  assign io_loadOut_0_bits_uop_cf_trigger_backendEn_1 = 4'hf == deqPtrExt_rvalue ? uop_15_cf_trigger_backendEn_1 :
    _GEN_30080; // @[LoadQueueFlag.scala 480:{26,26}]
  assign io_loadOut_0_bits_uop_cf_trigger_backendHit_0 = 4'hf == deqPtrExt_rvalue ? uop_15_cf_trigger_backendHit_0 :
    _GEN_30096; // @[LoadQueueFlag.scala 480:{26,26}]
  assign io_loadOut_0_bits_uop_cf_trigger_backendHit_1 = 4'hf == deqPtrExt_rvalue ? uop_15_cf_trigger_backendHit_1 :
    _GEN_30112; // @[LoadQueueFlag.scala 480:{26,26}]
  assign io_loadOut_0_bits_uop_cf_trigger_backendHit_4 = 4'hf == deqPtrExt_rvalue ? uop_15_cf_trigger_backendHit_4 :
    _GEN_30160; // @[LoadQueueFlag.scala 480:{26,26}]
  assign io_loadOut_0_bits_uop_ctrl_fuOpType = 4'hf == deqPtrExt_rvalue ? uop_15_ctrl_fuOpType : _GEN_29680; // @[LookupTree.scala 24:{34,34}]
  assign io_loadOut_0_bits_uop_ctrl_rfWen = 4'hf == deqPtrExt_rvalue ? uop_15_ctrl_rfWen : _GEN_30592; // @[LoadQueueFlag.scala 480:{26,26}]
  assign io_loadOut_0_bits_uop_ctrl_fpWen = 4'hf == deqPtrExt_rvalue ? uop_15_ctrl_fpWen : _GEN_29664; // @[LoadQueue.scala 59:{28,28}]
  assign io_loadOut_0_bits_uop_ctrl_flushPipe = 4'hf == deqPtrExt_rvalue ? uop_15_ctrl_flushPipe : _GEN_30656; // @[LoadQueueFlag.scala 480:{26,26}]
  assign io_loadOut_0_bits_uop_ctrl_replayInst = 4'hf == deqPtrExt_rvalue ? uop_15_ctrl_replayInst : _GEN_30976; // @[LoadQueueFlag.scala 480:{26,26}]
  assign io_loadOut_0_bits_uop_pdest = 4'hf == deqPtrExt_rvalue ? uop_15_pdest : _GEN_31088; // @[LoadQueueFlag.scala 480:{26,26}]
  assign io_loadOut_0_bits_uop_robIdx_flag = 4'hf == deqPtrExt_rvalue ? uop_15_robIdx_flag : _GEN_31120; // @[LoadQueueFlag.scala 480:{26,26}]
  assign io_loadOut_0_bits_uop_robIdx_value = 4'hf == deqPtrExt_rvalue ? uop_15_robIdx_value : _GEN_31136; // @[LoadQueueFlag.scala 480:{26,26}]
  assign io_ldRawDataOut_0_lqData = uncacheData; // @[LoadQueueFlag.scala 495:29]
  assign io_ldRawDataOut_0_uop_ctrl_fuOpType = io_loadOut_0_bits_uop_ctrl_fuOpType; // @[LoadQueueFlag.scala 496:26]
  assign io_ldRawDataOut_0_uop_ctrl_fpWen = io_loadOut_0_bits_uop_ctrl_fpWen; // @[LoadQueueFlag.scala 496:26]
  assign io_ldRawDataOut_0_addrOffset = paddrModule_io_rdata_0[2:0]; // @[LoadQueueFlag.scala 497:33]
  assign io_rob_isMMIO_0 = io_rob_isMMIO_0_REG; // @[LoadQueueFlag.scala 358:22]
  assign io_rob_isMMIO_1 = io_rob_isMMIO_1_REG; // @[LoadQueueFlag.scala 358:22]
  assign io_rob_uop_0_robIdx_value = io_rob_uop_0_REG_robIdx_value; // @[LoadQueueFlag.scala 359:19]
  assign io_rob_uop_1_robIdx_value = io_rob_uop_1_REG_robIdx_value; // @[LoadQueueFlag.scala 359:19]
  assign io_uncache_req_valid = uncacheState == 2'h1; // @[LoadQueueFlag.scala 431:40]
  assign io_uncache_req_bits_addr = paddrModule_io_rdata_0; // @[LoadQueueFlag.scala 434:28]
  assign io_uncache_req_bits_mask = maskModule_io_rdata_0; // @[LoadQueueFlag.scala 435:28]
  assign io_uncache_resp_ready = 1'h1; // @[LoadQueueFlag.scala 441:25]
  assign io_trigger_0_lqLoadAddrTriggerHitVec_0 = io_loadOut_0_valid & vaddrTriggerResultModule_io_rdata_0_0; // @[LoadQueueFlag.scala 371:51]
  assign io_trigger_0_lqLoadAddrTriggerHitVec_1 = io_loadOut_0_valid & vaddrTriggerResultModule_io_rdata_0_1; // @[LoadQueueFlag.scala 371:51]
  assign io_trigger_0_lqLoadAddrTriggerHitVec_2 = io_loadOut_0_valid & vaddrTriggerResultModule_io_rdata_0_2; // @[LoadQueueFlag.scala 371:51]
  assign io_exceptionAddr_vaddr = vaddrModule_io_rdata_1; // @[LoadQueueFlag.scala 365:26]
  assign io_ldIssuePtr_flag = deqPtrExt_rflag; // @[LoadQueueFlag.scala 118:23 166:13]
  assign io_ldIssuePtr_value = deqPtrExt_rvalue; // @[LoadQueueFlag.scala 118:23 166:13]
  assign io_lqDeq = io_lqDeq_REG; // @[LoadQueueFlag.scala 168:12]
  assign io_lqCancelCnt = io_lqCancelCnt_REG; // @[LoadQueueFlag.scala 169:18]
  assign io_perf_0_value = {{5'd0}, io_perf_0_value_REG_1}; // @[PerfCounterUtils.scala 188:17]
  assign io_perf_1_value = {{5'd0}, io_perf_1_value_REG_1}; // @[PerfCounterUtils.scala 188:17]
  assign io_perf_2_value = {{5'd0}, io_perf_2_value_REG_1}; // @[PerfCounterUtils.scala 188:17]
  assign io_perf_3_value = {{5'd0}, io_perf_3_value_REG_1}; // @[PerfCounterUtils.scala 188:17]
  assign vaddrModule_clock = clock;
  assign vaddrModule_io_raddr_1 = _deqPtrExtNext_new_ptr_T_2[3:0]; // @[CircularQueuePtr.scala 39:59]
  assign vaddrModule_io_wen_0 = io_loadIn_0_valid & _issued_T_1; // @[LoadQueueFlag.scala 277:27 286:31]
  assign vaddrModule_io_wen_1 = io_loadIn_1_valid & _issued_T_7; // @[LoadQueueFlag.scala 277:27 286:31]
  assign vaddrModule_io_waddr_0 = io_loadIn_0_bits_uop_lqIdx_value; // @[LoadQueueFlag.scala 301:26 330:33]
  assign vaddrModule_io_waddr_1 = io_loadIn_1_bits_uop_lqIdx_value; // @[LoadQueueFlag.scala 301:26 330:33]
  assign vaddrModule_io_wdata_0 = io_loadIn_0_bits_vaddr; // @[LoadQueueFlag.scala 301:26 331:33]
  assign vaddrModule_io_wdata_1 = io_loadIn_1_bits_vaddr; // @[LoadQueueFlag.scala 301:26 331:33]
  assign paddrModule_clock = clock;
  assign paddrModule_io_raddr_0 = _deqPtrExtNext_new_ptr_T_2[3:0]; // @[CircularQueuePtr.scala 39:59]
  assign paddrModule_io_wen_0 = io_loadIn_0_valid & _issued_T_1; // @[LoadQueueFlag.scala 277:27 286:31]
  assign paddrModule_io_wen_1 = io_loadIn_1_valid & _issued_T_7; // @[LoadQueueFlag.scala 277:27 286:31]
  assign paddrModule_io_waddr_0 = io_loadIn_0_bits_uop_lqIdx_value; // @[LoadQueueFlag.scala 301:26 330:33]
  assign paddrModule_io_waddr_1 = io_loadIn_1_bits_uop_lqIdx_value; // @[LoadQueueFlag.scala 301:26 330:33]
  assign paddrModule_io_wdata_0 = io_loadIn_0_bits_paddr; // @[LoadQueueFlag.scala 301:26 335:33]
  assign paddrModule_io_wdata_1 = io_loadIn_1_bits_paddr; // @[LoadQueueFlag.scala 301:26 335:33]
  assign maskModule_clock = clock;
  assign maskModule_io_raddr_0 = _deqPtrExtNext_new_ptr_T_2[3:0]; // @[CircularQueuePtr.scala 39:59]
  assign maskModule_io_wen_0 = io_loadIn_0_valid & _issued_T_1; // @[LoadQueueFlag.scala 277:27 286:31]
  assign maskModule_io_wen_1 = io_loadIn_1_valid & _issued_T_7; // @[LoadQueueFlag.scala 277:27 286:31]
  assign maskModule_io_waddr_0 = io_loadIn_0_bits_uop_lqIdx_value; // @[LoadQueueFlag.scala 301:26 330:33]
  assign maskModule_io_waddr_1 = io_loadIn_1_bits_uop_lqIdx_value; // @[LoadQueueFlag.scala 301:26 330:33]
  assign maskModule_io_wdata_0 = io_loadIn_0_bits_mask[7:0];
  assign maskModule_io_wdata_1 = io_loadIn_1_bits_mask[7:0];
  assign vaddrTriggerResultModule_clock = clock;
  assign vaddrTriggerResultModule_io_raddr_0 = deqPtrExt_rvalue; // @[LoadQueueFlag.scala 118:23 166:13]
  assign vaddrTriggerResultModule_io_wen_0 = io_loadIn_0_valid & _GEN_21339; // @[LoadQueueFlag.scala 286:31 280:40]
  assign vaddrTriggerResultModule_io_wen_1 = io_loadIn_1_valid & _GEN_27860; // @[LoadQueueFlag.scala 286:31 280:40]
  assign vaddrTriggerResultModule_io_waddr_0 = io_loadIn_0_bits_uop_lqIdx_value; // @[LoadQueueFlag.scala 321:50 323:48]
  assign vaddrTriggerResultModule_io_waddr_1 = io_loadIn_1_bits_uop_lqIdx_value; // @[LoadQueueFlag.scala 321:50 323:48]
  assign vaddrTriggerResultModule_io_wdata_0_0 = io_trigger_0_hitLoadAddrTriggerHitVec_0; // @[LoadQueueFlag.scala 321:50 324:48]
  assign vaddrTriggerResultModule_io_wdata_0_1 = io_trigger_0_hitLoadAddrTriggerHitVec_1; // @[LoadQueueFlag.scala 321:50 324:48]
  assign vaddrTriggerResultModule_io_wdata_0_2 = io_trigger_0_hitLoadAddrTriggerHitVec_2; // @[LoadQueueFlag.scala 321:50 324:48]
  assign vaddrTriggerResultModule_io_wdata_1_0 = io_trigger_1_hitLoadAddrTriggerHitVec_0; // @[LoadQueueFlag.scala 321:50 324:48]
  assign vaddrTriggerResultModule_io_wdata_1_1 = io_trigger_1_hitLoadAddrTriggerHitVec_1; // @[LoadQueueFlag.scala 321:50 324:48]
  assign vaddrTriggerResultModule_io_wdata_1_2 = io_trigger_1_hitLoadAddrTriggerHitVec_2; // @[LoadQueueFlag.scala 321:50 324:48]
  always @(posedge clock) begin
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'h0 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_0_cf_exceptionVec_4 <= io_loadIn_1_bits_uop_cf_exceptionVec_4; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_0_cf_exceptionVec_4 <= _GEN_21589;
          end
        end else begin
          uop_0_cf_exceptionVec_4 <= _GEN_21589;
        end
      end else begin
        uop_0_cf_exceptionVec_4 <= _GEN_21589;
      end
    end else begin
      uop_0_cf_exceptionVec_4 <= _GEN_21589;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'h0 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_0_cf_exceptionVec_5 <= io_loadIn_1_bits_uop_cf_exceptionVec_5; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_0_cf_exceptionVec_5 <= _GEN_21605;
          end
        end else begin
          uop_0_cf_exceptionVec_5 <= _GEN_21605;
        end
      end else begin
        uop_0_cf_exceptionVec_5 <= _GEN_21605;
      end
    end else begin
      uop_0_cf_exceptionVec_5 <= _GEN_21605;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'h0 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_0_cf_exceptionVec_13 <= io_loadIn_1_bits_uop_cf_exceptionVec_13; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_0_cf_exceptionVec_13 <= _GEN_21733;
          end
        end else begin
          uop_0_cf_exceptionVec_13 <= _GEN_21733;
        end
      end else begin
        uop_0_cf_exceptionVec_13 <= _GEN_21733;
      end
    end else begin
      uop_0_cf_exceptionVec_13 <= _GEN_21733;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'h0 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_0_cf_trigger_backendEn_1 <= io_loadIn_1_bits_uop_cf_trigger_backendEn_1; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_0_cf_trigger_backendEn_1 <= _GEN_21861;
          end
        end else begin
          uop_0_cf_trigger_backendEn_1 <= _GEN_21861;
        end
      end else begin
        uop_0_cf_trigger_backendEn_1 <= _GEN_21861;
      end
    end else begin
      uop_0_cf_trigger_backendEn_1 <= _GEN_21861;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'h0 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_0_cf_trigger_backendHit_0 <= io_loadIn_1_bits_uop_cf_trigger_backendHit_0; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_0_cf_trigger_backendHit_0 <= _GEN_21877;
          end
        end else begin
          uop_0_cf_trigger_backendHit_0 <= _GEN_21877;
        end
      end else begin
        uop_0_cf_trigger_backendHit_0 <= _GEN_21877;
      end
    end else begin
      uop_0_cf_trigger_backendHit_0 <= _GEN_21877;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'h0 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_0_cf_trigger_backendHit_1 <= io_loadIn_1_bits_uop_cf_trigger_backendHit_1; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_0_cf_trigger_backendHit_1 <= _GEN_21893;
          end
        end else begin
          uop_0_cf_trigger_backendHit_1 <= _GEN_21893;
        end
      end else begin
        uop_0_cf_trigger_backendHit_1 <= _GEN_21893;
      end
    end else begin
      uop_0_cf_trigger_backendHit_1 <= _GEN_21893;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'h0 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_0_cf_trigger_backendHit_4 <= io_loadIn_1_bits_uop_cf_trigger_backendHit_4; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_0_cf_trigger_backendHit_4 <= _GEN_21941;
          end
        end else begin
          uop_0_cf_trigger_backendHit_4 <= _GEN_21941;
        end
      end else begin
        uop_0_cf_trigger_backendHit_4 <= _GEN_21941;
      end
    end else begin
      uop_0_cf_trigger_backendHit_4 <= _GEN_21941;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_3) begin // @[LoadQueueFlag.scala 315:50]
          if (4'h0 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 316:33]
            uop_0_ctrl_fuOpType <= io_loadIn_1_bits_uop_ctrl_fuOpType; // @[LoadQueueFlag.scala 316:33]
          end else begin
            uop_0_ctrl_fuOpType <= _GEN_22373;
          end
        end else begin
          uop_0_ctrl_fuOpType <= _GEN_22373;
        end
      end else begin
        uop_0_ctrl_fuOpType <= _GEN_22373;
      end
    end else begin
      uop_0_ctrl_fuOpType <= _GEN_22373;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_3) begin // @[LoadQueueFlag.scala 315:50]
          if (4'h0 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 316:33]
            uop_0_ctrl_rfWen <= io_loadIn_1_bits_uop_ctrl_rfWen; // @[LoadQueueFlag.scala 316:33]
          end else begin
            uop_0_ctrl_rfWen <= _GEN_22389;
          end
        end else begin
          uop_0_ctrl_rfWen <= _GEN_22389;
        end
      end else begin
        uop_0_ctrl_rfWen <= _GEN_22389;
      end
    end else begin
      uop_0_ctrl_rfWen <= _GEN_22389;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_3) begin // @[LoadQueueFlag.scala 315:50]
          if (4'h0 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 316:33]
            uop_0_ctrl_fpWen <= io_loadIn_1_bits_uop_ctrl_fpWen; // @[LoadQueueFlag.scala 316:33]
          end else begin
            uop_0_ctrl_fpWen <= _GEN_22405;
          end
        end else begin
          uop_0_ctrl_fpWen <= _GEN_22405;
        end
      end else begin
        uop_0_ctrl_fpWen <= _GEN_22405;
      end
    end else begin
      uop_0_ctrl_fpWen <= _GEN_22405;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_3) begin // @[LoadQueueFlag.scala 315:50]
          if (4'h0 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 316:33]
            uop_0_ctrl_flushPipe <= 1'h0; // @[LoadQueueFlag.scala 316:33]
          end else begin
            uop_0_ctrl_flushPipe <= _GEN_22469;
          end
        end else begin
          uop_0_ctrl_flushPipe <= _GEN_22469;
        end
      end else begin
        uop_0_ctrl_flushPipe <= _GEN_22469;
      end
    end else begin
      uop_0_ctrl_flushPipe <= _GEN_22469;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_3) begin // @[LoadQueueFlag.scala 315:50]
          if (4'h0 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 316:33]
            uop_0_ctrl_replayInst <= io_loadIn_1_bits_uop_ctrl_replayInst; // @[LoadQueueFlag.scala 316:33]
          end else begin
            uop_0_ctrl_replayInst <= _GEN_22789;
          end
        end else begin
          uop_0_ctrl_replayInst <= _GEN_22789;
        end
      end else begin
        uop_0_ctrl_replayInst <= _GEN_22789;
      end
    end else begin
      uop_0_ctrl_replayInst <= _GEN_22789;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_1) begin // @[LoadQueueFlag.scala 309:50]
          if (4'h0 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 310:34]
            uop_0_pdest <= io_loadIn_1_bits_uop_pdest; // @[LoadQueueFlag.scala 310:34]
          end else begin
            uop_0_pdest <= _GEN_21461;
          end
        end else begin
          uop_0_pdest <= _GEN_21461;
        end
      end else begin
        uop_0_pdest <= _GEN_21461;
      end
    end else begin
      uop_0_pdest <= _GEN_21461;
    end
    if (io_enq_req_3_valid & ~enqCancel_3) begin // @[LoadQueueFlag.scala 204:43]
      if (4'h0 == io_enq_req_3_bits_lqIdx_value) begin // @[LoadQueueFlag.scala 206:18]
        uop_0_robIdx_flag <= io_enq_req_3_bits_robIdx_flag; // @[LoadQueueFlag.scala 206:18]
      end else begin
        uop_0_robIdx_flag <= _GEN_11902;
      end
    end else begin
      uop_0_robIdx_flag <= _GEN_11902;
    end
    if (io_enq_req_3_valid & ~enqCancel_3) begin // @[LoadQueueFlag.scala 204:43]
      if (4'h0 == io_enq_req_3_bits_lqIdx_value) begin // @[LoadQueueFlag.scala 206:18]
        uop_0_robIdx_value <= io_enq_req_3_bits_robIdx_value; // @[LoadQueueFlag.scala 206:18]
      end else begin
        uop_0_robIdx_value <= _GEN_11918;
      end
    end else begin
      uop_0_robIdx_value <= _GEN_11918;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'h1 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_1_cf_exceptionVec_4 <= io_loadIn_1_bits_uop_cf_exceptionVec_4; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_1_cf_exceptionVec_4 <= _GEN_21590;
          end
        end else begin
          uop_1_cf_exceptionVec_4 <= _GEN_21590;
        end
      end else begin
        uop_1_cf_exceptionVec_4 <= _GEN_21590;
      end
    end else begin
      uop_1_cf_exceptionVec_4 <= _GEN_21590;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'h1 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_1_cf_exceptionVec_5 <= io_loadIn_1_bits_uop_cf_exceptionVec_5; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_1_cf_exceptionVec_5 <= _GEN_21606;
          end
        end else begin
          uop_1_cf_exceptionVec_5 <= _GEN_21606;
        end
      end else begin
        uop_1_cf_exceptionVec_5 <= _GEN_21606;
      end
    end else begin
      uop_1_cf_exceptionVec_5 <= _GEN_21606;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'h1 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_1_cf_exceptionVec_13 <= io_loadIn_1_bits_uop_cf_exceptionVec_13; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_1_cf_exceptionVec_13 <= _GEN_21734;
          end
        end else begin
          uop_1_cf_exceptionVec_13 <= _GEN_21734;
        end
      end else begin
        uop_1_cf_exceptionVec_13 <= _GEN_21734;
      end
    end else begin
      uop_1_cf_exceptionVec_13 <= _GEN_21734;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'h1 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_1_cf_trigger_backendEn_1 <= io_loadIn_1_bits_uop_cf_trigger_backendEn_1; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_1_cf_trigger_backendEn_1 <= _GEN_21862;
          end
        end else begin
          uop_1_cf_trigger_backendEn_1 <= _GEN_21862;
        end
      end else begin
        uop_1_cf_trigger_backendEn_1 <= _GEN_21862;
      end
    end else begin
      uop_1_cf_trigger_backendEn_1 <= _GEN_21862;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'h1 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_1_cf_trigger_backendHit_0 <= io_loadIn_1_bits_uop_cf_trigger_backendHit_0; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_1_cf_trigger_backendHit_0 <= _GEN_21878;
          end
        end else begin
          uop_1_cf_trigger_backendHit_0 <= _GEN_21878;
        end
      end else begin
        uop_1_cf_trigger_backendHit_0 <= _GEN_21878;
      end
    end else begin
      uop_1_cf_trigger_backendHit_0 <= _GEN_21878;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'h1 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_1_cf_trigger_backendHit_1 <= io_loadIn_1_bits_uop_cf_trigger_backendHit_1; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_1_cf_trigger_backendHit_1 <= _GEN_21894;
          end
        end else begin
          uop_1_cf_trigger_backendHit_1 <= _GEN_21894;
        end
      end else begin
        uop_1_cf_trigger_backendHit_1 <= _GEN_21894;
      end
    end else begin
      uop_1_cf_trigger_backendHit_1 <= _GEN_21894;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'h1 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_1_cf_trigger_backendHit_4 <= io_loadIn_1_bits_uop_cf_trigger_backendHit_4; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_1_cf_trigger_backendHit_4 <= _GEN_21942;
          end
        end else begin
          uop_1_cf_trigger_backendHit_4 <= _GEN_21942;
        end
      end else begin
        uop_1_cf_trigger_backendHit_4 <= _GEN_21942;
      end
    end else begin
      uop_1_cf_trigger_backendHit_4 <= _GEN_21942;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_3) begin // @[LoadQueueFlag.scala 315:50]
          if (4'h1 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 316:33]
            uop_1_ctrl_fuOpType <= io_loadIn_1_bits_uop_ctrl_fuOpType; // @[LoadQueueFlag.scala 316:33]
          end else begin
            uop_1_ctrl_fuOpType <= _GEN_22374;
          end
        end else begin
          uop_1_ctrl_fuOpType <= _GEN_22374;
        end
      end else begin
        uop_1_ctrl_fuOpType <= _GEN_22374;
      end
    end else begin
      uop_1_ctrl_fuOpType <= _GEN_22374;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_3) begin // @[LoadQueueFlag.scala 315:50]
          if (4'h1 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 316:33]
            uop_1_ctrl_rfWen <= io_loadIn_1_bits_uop_ctrl_rfWen; // @[LoadQueueFlag.scala 316:33]
          end else begin
            uop_1_ctrl_rfWen <= _GEN_22390;
          end
        end else begin
          uop_1_ctrl_rfWen <= _GEN_22390;
        end
      end else begin
        uop_1_ctrl_rfWen <= _GEN_22390;
      end
    end else begin
      uop_1_ctrl_rfWen <= _GEN_22390;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_3) begin // @[LoadQueueFlag.scala 315:50]
          if (4'h1 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 316:33]
            uop_1_ctrl_fpWen <= io_loadIn_1_bits_uop_ctrl_fpWen; // @[LoadQueueFlag.scala 316:33]
          end else begin
            uop_1_ctrl_fpWen <= _GEN_22406;
          end
        end else begin
          uop_1_ctrl_fpWen <= _GEN_22406;
        end
      end else begin
        uop_1_ctrl_fpWen <= _GEN_22406;
      end
    end else begin
      uop_1_ctrl_fpWen <= _GEN_22406;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_3) begin // @[LoadQueueFlag.scala 315:50]
          if (4'h1 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 316:33]
            uop_1_ctrl_flushPipe <= 1'h0; // @[LoadQueueFlag.scala 316:33]
          end else begin
            uop_1_ctrl_flushPipe <= _GEN_22470;
          end
        end else begin
          uop_1_ctrl_flushPipe <= _GEN_22470;
        end
      end else begin
        uop_1_ctrl_flushPipe <= _GEN_22470;
      end
    end else begin
      uop_1_ctrl_flushPipe <= _GEN_22470;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_3) begin // @[LoadQueueFlag.scala 315:50]
          if (4'h1 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 316:33]
            uop_1_ctrl_replayInst <= io_loadIn_1_bits_uop_ctrl_replayInst; // @[LoadQueueFlag.scala 316:33]
          end else begin
            uop_1_ctrl_replayInst <= _GEN_22790;
          end
        end else begin
          uop_1_ctrl_replayInst <= _GEN_22790;
        end
      end else begin
        uop_1_ctrl_replayInst <= _GEN_22790;
      end
    end else begin
      uop_1_ctrl_replayInst <= _GEN_22790;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_1) begin // @[LoadQueueFlag.scala 309:50]
          if (4'h1 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 310:34]
            uop_1_pdest <= io_loadIn_1_bits_uop_pdest; // @[LoadQueueFlag.scala 310:34]
          end else begin
            uop_1_pdest <= _GEN_21462;
          end
        end else begin
          uop_1_pdest <= _GEN_21462;
        end
      end else begin
        uop_1_pdest <= _GEN_21462;
      end
    end else begin
      uop_1_pdest <= _GEN_21462;
    end
    if (io_enq_req_3_valid & ~enqCancel_3) begin // @[LoadQueueFlag.scala 204:43]
      if (4'h1 == io_enq_req_3_bits_lqIdx_value) begin // @[LoadQueueFlag.scala 206:18]
        uop_1_robIdx_flag <= io_enq_req_3_bits_robIdx_flag; // @[LoadQueueFlag.scala 206:18]
      end else begin
        uop_1_robIdx_flag <= _GEN_11903;
      end
    end else begin
      uop_1_robIdx_flag <= _GEN_11903;
    end
    if (io_enq_req_3_valid & ~enqCancel_3) begin // @[LoadQueueFlag.scala 204:43]
      if (4'h1 == io_enq_req_3_bits_lqIdx_value) begin // @[LoadQueueFlag.scala 206:18]
        uop_1_robIdx_value <= io_enq_req_3_bits_robIdx_value; // @[LoadQueueFlag.scala 206:18]
      end else begin
        uop_1_robIdx_value <= _GEN_11919;
      end
    end else begin
      uop_1_robIdx_value <= _GEN_11919;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'h2 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_2_cf_exceptionVec_4 <= io_loadIn_1_bits_uop_cf_exceptionVec_4; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_2_cf_exceptionVec_4 <= _GEN_21591;
          end
        end else begin
          uop_2_cf_exceptionVec_4 <= _GEN_21591;
        end
      end else begin
        uop_2_cf_exceptionVec_4 <= _GEN_21591;
      end
    end else begin
      uop_2_cf_exceptionVec_4 <= _GEN_21591;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'h2 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_2_cf_exceptionVec_5 <= io_loadIn_1_bits_uop_cf_exceptionVec_5; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_2_cf_exceptionVec_5 <= _GEN_21607;
          end
        end else begin
          uop_2_cf_exceptionVec_5 <= _GEN_21607;
        end
      end else begin
        uop_2_cf_exceptionVec_5 <= _GEN_21607;
      end
    end else begin
      uop_2_cf_exceptionVec_5 <= _GEN_21607;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'h2 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_2_cf_exceptionVec_13 <= io_loadIn_1_bits_uop_cf_exceptionVec_13; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_2_cf_exceptionVec_13 <= _GEN_21735;
          end
        end else begin
          uop_2_cf_exceptionVec_13 <= _GEN_21735;
        end
      end else begin
        uop_2_cf_exceptionVec_13 <= _GEN_21735;
      end
    end else begin
      uop_2_cf_exceptionVec_13 <= _GEN_21735;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'h2 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_2_cf_trigger_backendEn_1 <= io_loadIn_1_bits_uop_cf_trigger_backendEn_1; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_2_cf_trigger_backendEn_1 <= _GEN_21863;
          end
        end else begin
          uop_2_cf_trigger_backendEn_1 <= _GEN_21863;
        end
      end else begin
        uop_2_cf_trigger_backendEn_1 <= _GEN_21863;
      end
    end else begin
      uop_2_cf_trigger_backendEn_1 <= _GEN_21863;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'h2 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_2_cf_trigger_backendHit_0 <= io_loadIn_1_bits_uop_cf_trigger_backendHit_0; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_2_cf_trigger_backendHit_0 <= _GEN_21879;
          end
        end else begin
          uop_2_cf_trigger_backendHit_0 <= _GEN_21879;
        end
      end else begin
        uop_2_cf_trigger_backendHit_0 <= _GEN_21879;
      end
    end else begin
      uop_2_cf_trigger_backendHit_0 <= _GEN_21879;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'h2 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_2_cf_trigger_backendHit_1 <= io_loadIn_1_bits_uop_cf_trigger_backendHit_1; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_2_cf_trigger_backendHit_1 <= _GEN_21895;
          end
        end else begin
          uop_2_cf_trigger_backendHit_1 <= _GEN_21895;
        end
      end else begin
        uop_2_cf_trigger_backendHit_1 <= _GEN_21895;
      end
    end else begin
      uop_2_cf_trigger_backendHit_1 <= _GEN_21895;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'h2 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_2_cf_trigger_backendHit_4 <= io_loadIn_1_bits_uop_cf_trigger_backendHit_4; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_2_cf_trigger_backendHit_4 <= _GEN_21943;
          end
        end else begin
          uop_2_cf_trigger_backendHit_4 <= _GEN_21943;
        end
      end else begin
        uop_2_cf_trigger_backendHit_4 <= _GEN_21943;
      end
    end else begin
      uop_2_cf_trigger_backendHit_4 <= _GEN_21943;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_3) begin // @[LoadQueueFlag.scala 315:50]
          if (4'h2 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 316:33]
            uop_2_ctrl_fuOpType <= io_loadIn_1_bits_uop_ctrl_fuOpType; // @[LoadQueueFlag.scala 316:33]
          end else begin
            uop_2_ctrl_fuOpType <= _GEN_22375;
          end
        end else begin
          uop_2_ctrl_fuOpType <= _GEN_22375;
        end
      end else begin
        uop_2_ctrl_fuOpType <= _GEN_22375;
      end
    end else begin
      uop_2_ctrl_fuOpType <= _GEN_22375;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_3) begin // @[LoadQueueFlag.scala 315:50]
          if (4'h2 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 316:33]
            uop_2_ctrl_rfWen <= io_loadIn_1_bits_uop_ctrl_rfWen; // @[LoadQueueFlag.scala 316:33]
          end else begin
            uop_2_ctrl_rfWen <= _GEN_22391;
          end
        end else begin
          uop_2_ctrl_rfWen <= _GEN_22391;
        end
      end else begin
        uop_2_ctrl_rfWen <= _GEN_22391;
      end
    end else begin
      uop_2_ctrl_rfWen <= _GEN_22391;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_3) begin // @[LoadQueueFlag.scala 315:50]
          if (4'h2 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 316:33]
            uop_2_ctrl_fpWen <= io_loadIn_1_bits_uop_ctrl_fpWen; // @[LoadQueueFlag.scala 316:33]
          end else begin
            uop_2_ctrl_fpWen <= _GEN_22407;
          end
        end else begin
          uop_2_ctrl_fpWen <= _GEN_22407;
        end
      end else begin
        uop_2_ctrl_fpWen <= _GEN_22407;
      end
    end else begin
      uop_2_ctrl_fpWen <= _GEN_22407;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_3) begin // @[LoadQueueFlag.scala 315:50]
          if (4'h2 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 316:33]
            uop_2_ctrl_flushPipe <= 1'h0; // @[LoadQueueFlag.scala 316:33]
          end else begin
            uop_2_ctrl_flushPipe <= _GEN_22471;
          end
        end else begin
          uop_2_ctrl_flushPipe <= _GEN_22471;
        end
      end else begin
        uop_2_ctrl_flushPipe <= _GEN_22471;
      end
    end else begin
      uop_2_ctrl_flushPipe <= _GEN_22471;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_3) begin // @[LoadQueueFlag.scala 315:50]
          if (4'h2 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 316:33]
            uop_2_ctrl_replayInst <= io_loadIn_1_bits_uop_ctrl_replayInst; // @[LoadQueueFlag.scala 316:33]
          end else begin
            uop_2_ctrl_replayInst <= _GEN_22791;
          end
        end else begin
          uop_2_ctrl_replayInst <= _GEN_22791;
        end
      end else begin
        uop_2_ctrl_replayInst <= _GEN_22791;
      end
    end else begin
      uop_2_ctrl_replayInst <= _GEN_22791;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_1) begin // @[LoadQueueFlag.scala 309:50]
          if (4'h2 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 310:34]
            uop_2_pdest <= io_loadIn_1_bits_uop_pdest; // @[LoadQueueFlag.scala 310:34]
          end else begin
            uop_2_pdest <= _GEN_21463;
          end
        end else begin
          uop_2_pdest <= _GEN_21463;
        end
      end else begin
        uop_2_pdest <= _GEN_21463;
      end
    end else begin
      uop_2_pdest <= _GEN_21463;
    end
    if (io_enq_req_3_valid & ~enqCancel_3) begin // @[LoadQueueFlag.scala 204:43]
      if (4'h2 == io_enq_req_3_bits_lqIdx_value) begin // @[LoadQueueFlag.scala 206:18]
        uop_2_robIdx_flag <= io_enq_req_3_bits_robIdx_flag; // @[LoadQueueFlag.scala 206:18]
      end else begin
        uop_2_robIdx_flag <= _GEN_11904;
      end
    end else begin
      uop_2_robIdx_flag <= _GEN_11904;
    end
    if (io_enq_req_3_valid & ~enqCancel_3) begin // @[LoadQueueFlag.scala 204:43]
      if (4'h2 == io_enq_req_3_bits_lqIdx_value) begin // @[LoadQueueFlag.scala 206:18]
        uop_2_robIdx_value <= io_enq_req_3_bits_robIdx_value; // @[LoadQueueFlag.scala 206:18]
      end else begin
        uop_2_robIdx_value <= _GEN_11920;
      end
    end else begin
      uop_2_robIdx_value <= _GEN_11920;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'h3 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_3_cf_exceptionVec_4 <= io_loadIn_1_bits_uop_cf_exceptionVec_4; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_3_cf_exceptionVec_4 <= _GEN_21592;
          end
        end else begin
          uop_3_cf_exceptionVec_4 <= _GEN_21592;
        end
      end else begin
        uop_3_cf_exceptionVec_4 <= _GEN_21592;
      end
    end else begin
      uop_3_cf_exceptionVec_4 <= _GEN_21592;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'h3 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_3_cf_exceptionVec_5 <= io_loadIn_1_bits_uop_cf_exceptionVec_5; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_3_cf_exceptionVec_5 <= _GEN_21608;
          end
        end else begin
          uop_3_cf_exceptionVec_5 <= _GEN_21608;
        end
      end else begin
        uop_3_cf_exceptionVec_5 <= _GEN_21608;
      end
    end else begin
      uop_3_cf_exceptionVec_5 <= _GEN_21608;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'h3 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_3_cf_exceptionVec_13 <= io_loadIn_1_bits_uop_cf_exceptionVec_13; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_3_cf_exceptionVec_13 <= _GEN_21736;
          end
        end else begin
          uop_3_cf_exceptionVec_13 <= _GEN_21736;
        end
      end else begin
        uop_3_cf_exceptionVec_13 <= _GEN_21736;
      end
    end else begin
      uop_3_cf_exceptionVec_13 <= _GEN_21736;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'h3 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_3_cf_trigger_backendEn_1 <= io_loadIn_1_bits_uop_cf_trigger_backendEn_1; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_3_cf_trigger_backendEn_1 <= _GEN_21864;
          end
        end else begin
          uop_3_cf_trigger_backendEn_1 <= _GEN_21864;
        end
      end else begin
        uop_3_cf_trigger_backendEn_1 <= _GEN_21864;
      end
    end else begin
      uop_3_cf_trigger_backendEn_1 <= _GEN_21864;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'h3 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_3_cf_trigger_backendHit_0 <= io_loadIn_1_bits_uop_cf_trigger_backendHit_0; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_3_cf_trigger_backendHit_0 <= _GEN_21880;
          end
        end else begin
          uop_3_cf_trigger_backendHit_0 <= _GEN_21880;
        end
      end else begin
        uop_3_cf_trigger_backendHit_0 <= _GEN_21880;
      end
    end else begin
      uop_3_cf_trigger_backendHit_0 <= _GEN_21880;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'h3 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_3_cf_trigger_backendHit_1 <= io_loadIn_1_bits_uop_cf_trigger_backendHit_1; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_3_cf_trigger_backendHit_1 <= _GEN_21896;
          end
        end else begin
          uop_3_cf_trigger_backendHit_1 <= _GEN_21896;
        end
      end else begin
        uop_3_cf_trigger_backendHit_1 <= _GEN_21896;
      end
    end else begin
      uop_3_cf_trigger_backendHit_1 <= _GEN_21896;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'h3 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_3_cf_trigger_backendHit_4 <= io_loadIn_1_bits_uop_cf_trigger_backendHit_4; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_3_cf_trigger_backendHit_4 <= _GEN_21944;
          end
        end else begin
          uop_3_cf_trigger_backendHit_4 <= _GEN_21944;
        end
      end else begin
        uop_3_cf_trigger_backendHit_4 <= _GEN_21944;
      end
    end else begin
      uop_3_cf_trigger_backendHit_4 <= _GEN_21944;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_3) begin // @[LoadQueueFlag.scala 315:50]
          if (4'h3 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 316:33]
            uop_3_ctrl_fuOpType <= io_loadIn_1_bits_uop_ctrl_fuOpType; // @[LoadQueueFlag.scala 316:33]
          end else begin
            uop_3_ctrl_fuOpType <= _GEN_22376;
          end
        end else begin
          uop_3_ctrl_fuOpType <= _GEN_22376;
        end
      end else begin
        uop_3_ctrl_fuOpType <= _GEN_22376;
      end
    end else begin
      uop_3_ctrl_fuOpType <= _GEN_22376;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_3) begin // @[LoadQueueFlag.scala 315:50]
          if (4'h3 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 316:33]
            uop_3_ctrl_rfWen <= io_loadIn_1_bits_uop_ctrl_rfWen; // @[LoadQueueFlag.scala 316:33]
          end else begin
            uop_3_ctrl_rfWen <= _GEN_22392;
          end
        end else begin
          uop_3_ctrl_rfWen <= _GEN_22392;
        end
      end else begin
        uop_3_ctrl_rfWen <= _GEN_22392;
      end
    end else begin
      uop_3_ctrl_rfWen <= _GEN_22392;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_3) begin // @[LoadQueueFlag.scala 315:50]
          if (4'h3 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 316:33]
            uop_3_ctrl_fpWen <= io_loadIn_1_bits_uop_ctrl_fpWen; // @[LoadQueueFlag.scala 316:33]
          end else begin
            uop_3_ctrl_fpWen <= _GEN_22408;
          end
        end else begin
          uop_3_ctrl_fpWen <= _GEN_22408;
        end
      end else begin
        uop_3_ctrl_fpWen <= _GEN_22408;
      end
    end else begin
      uop_3_ctrl_fpWen <= _GEN_22408;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_3) begin // @[LoadQueueFlag.scala 315:50]
          if (4'h3 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 316:33]
            uop_3_ctrl_flushPipe <= 1'h0; // @[LoadQueueFlag.scala 316:33]
          end else begin
            uop_3_ctrl_flushPipe <= _GEN_22472;
          end
        end else begin
          uop_3_ctrl_flushPipe <= _GEN_22472;
        end
      end else begin
        uop_3_ctrl_flushPipe <= _GEN_22472;
      end
    end else begin
      uop_3_ctrl_flushPipe <= _GEN_22472;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_3) begin // @[LoadQueueFlag.scala 315:50]
          if (4'h3 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 316:33]
            uop_3_ctrl_replayInst <= io_loadIn_1_bits_uop_ctrl_replayInst; // @[LoadQueueFlag.scala 316:33]
          end else begin
            uop_3_ctrl_replayInst <= _GEN_22792;
          end
        end else begin
          uop_3_ctrl_replayInst <= _GEN_22792;
        end
      end else begin
        uop_3_ctrl_replayInst <= _GEN_22792;
      end
    end else begin
      uop_3_ctrl_replayInst <= _GEN_22792;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_1) begin // @[LoadQueueFlag.scala 309:50]
          if (4'h3 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 310:34]
            uop_3_pdest <= io_loadIn_1_bits_uop_pdest; // @[LoadQueueFlag.scala 310:34]
          end else begin
            uop_3_pdest <= _GEN_21464;
          end
        end else begin
          uop_3_pdest <= _GEN_21464;
        end
      end else begin
        uop_3_pdest <= _GEN_21464;
      end
    end else begin
      uop_3_pdest <= _GEN_21464;
    end
    if (io_enq_req_3_valid & ~enqCancel_3) begin // @[LoadQueueFlag.scala 204:43]
      if (4'h3 == io_enq_req_3_bits_lqIdx_value) begin // @[LoadQueueFlag.scala 206:18]
        uop_3_robIdx_flag <= io_enq_req_3_bits_robIdx_flag; // @[LoadQueueFlag.scala 206:18]
      end else begin
        uop_3_robIdx_flag <= _GEN_11905;
      end
    end else begin
      uop_3_robIdx_flag <= _GEN_11905;
    end
    if (io_enq_req_3_valid & ~enqCancel_3) begin // @[LoadQueueFlag.scala 204:43]
      if (4'h3 == io_enq_req_3_bits_lqIdx_value) begin // @[LoadQueueFlag.scala 206:18]
        uop_3_robIdx_value <= io_enq_req_3_bits_robIdx_value; // @[LoadQueueFlag.scala 206:18]
      end else begin
        uop_3_robIdx_value <= _GEN_11921;
      end
    end else begin
      uop_3_robIdx_value <= _GEN_11921;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'h4 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_4_cf_exceptionVec_4 <= io_loadIn_1_bits_uop_cf_exceptionVec_4; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_4_cf_exceptionVec_4 <= _GEN_21593;
          end
        end else begin
          uop_4_cf_exceptionVec_4 <= _GEN_21593;
        end
      end else begin
        uop_4_cf_exceptionVec_4 <= _GEN_21593;
      end
    end else begin
      uop_4_cf_exceptionVec_4 <= _GEN_21593;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'h4 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_4_cf_exceptionVec_5 <= io_loadIn_1_bits_uop_cf_exceptionVec_5; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_4_cf_exceptionVec_5 <= _GEN_21609;
          end
        end else begin
          uop_4_cf_exceptionVec_5 <= _GEN_21609;
        end
      end else begin
        uop_4_cf_exceptionVec_5 <= _GEN_21609;
      end
    end else begin
      uop_4_cf_exceptionVec_5 <= _GEN_21609;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'h4 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_4_cf_exceptionVec_13 <= io_loadIn_1_bits_uop_cf_exceptionVec_13; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_4_cf_exceptionVec_13 <= _GEN_21737;
          end
        end else begin
          uop_4_cf_exceptionVec_13 <= _GEN_21737;
        end
      end else begin
        uop_4_cf_exceptionVec_13 <= _GEN_21737;
      end
    end else begin
      uop_4_cf_exceptionVec_13 <= _GEN_21737;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'h4 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_4_cf_trigger_backendEn_1 <= io_loadIn_1_bits_uop_cf_trigger_backendEn_1; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_4_cf_trigger_backendEn_1 <= _GEN_21865;
          end
        end else begin
          uop_4_cf_trigger_backendEn_1 <= _GEN_21865;
        end
      end else begin
        uop_4_cf_trigger_backendEn_1 <= _GEN_21865;
      end
    end else begin
      uop_4_cf_trigger_backendEn_1 <= _GEN_21865;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'h4 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_4_cf_trigger_backendHit_0 <= io_loadIn_1_bits_uop_cf_trigger_backendHit_0; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_4_cf_trigger_backendHit_0 <= _GEN_21881;
          end
        end else begin
          uop_4_cf_trigger_backendHit_0 <= _GEN_21881;
        end
      end else begin
        uop_4_cf_trigger_backendHit_0 <= _GEN_21881;
      end
    end else begin
      uop_4_cf_trigger_backendHit_0 <= _GEN_21881;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'h4 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_4_cf_trigger_backendHit_1 <= io_loadIn_1_bits_uop_cf_trigger_backendHit_1; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_4_cf_trigger_backendHit_1 <= _GEN_21897;
          end
        end else begin
          uop_4_cf_trigger_backendHit_1 <= _GEN_21897;
        end
      end else begin
        uop_4_cf_trigger_backendHit_1 <= _GEN_21897;
      end
    end else begin
      uop_4_cf_trigger_backendHit_1 <= _GEN_21897;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'h4 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_4_cf_trigger_backendHit_4 <= io_loadIn_1_bits_uop_cf_trigger_backendHit_4; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_4_cf_trigger_backendHit_4 <= _GEN_21945;
          end
        end else begin
          uop_4_cf_trigger_backendHit_4 <= _GEN_21945;
        end
      end else begin
        uop_4_cf_trigger_backendHit_4 <= _GEN_21945;
      end
    end else begin
      uop_4_cf_trigger_backendHit_4 <= _GEN_21945;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_3) begin // @[LoadQueueFlag.scala 315:50]
          if (4'h4 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 316:33]
            uop_4_ctrl_fuOpType <= io_loadIn_1_bits_uop_ctrl_fuOpType; // @[LoadQueueFlag.scala 316:33]
          end else begin
            uop_4_ctrl_fuOpType <= _GEN_22377;
          end
        end else begin
          uop_4_ctrl_fuOpType <= _GEN_22377;
        end
      end else begin
        uop_4_ctrl_fuOpType <= _GEN_22377;
      end
    end else begin
      uop_4_ctrl_fuOpType <= _GEN_22377;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_3) begin // @[LoadQueueFlag.scala 315:50]
          if (4'h4 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 316:33]
            uop_4_ctrl_rfWen <= io_loadIn_1_bits_uop_ctrl_rfWen; // @[LoadQueueFlag.scala 316:33]
          end else begin
            uop_4_ctrl_rfWen <= _GEN_22393;
          end
        end else begin
          uop_4_ctrl_rfWen <= _GEN_22393;
        end
      end else begin
        uop_4_ctrl_rfWen <= _GEN_22393;
      end
    end else begin
      uop_4_ctrl_rfWen <= _GEN_22393;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_3) begin // @[LoadQueueFlag.scala 315:50]
          if (4'h4 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 316:33]
            uop_4_ctrl_fpWen <= io_loadIn_1_bits_uop_ctrl_fpWen; // @[LoadQueueFlag.scala 316:33]
          end else begin
            uop_4_ctrl_fpWen <= _GEN_22409;
          end
        end else begin
          uop_4_ctrl_fpWen <= _GEN_22409;
        end
      end else begin
        uop_4_ctrl_fpWen <= _GEN_22409;
      end
    end else begin
      uop_4_ctrl_fpWen <= _GEN_22409;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_3) begin // @[LoadQueueFlag.scala 315:50]
          if (4'h4 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 316:33]
            uop_4_ctrl_flushPipe <= 1'h0; // @[LoadQueueFlag.scala 316:33]
          end else begin
            uop_4_ctrl_flushPipe <= _GEN_22473;
          end
        end else begin
          uop_4_ctrl_flushPipe <= _GEN_22473;
        end
      end else begin
        uop_4_ctrl_flushPipe <= _GEN_22473;
      end
    end else begin
      uop_4_ctrl_flushPipe <= _GEN_22473;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_3) begin // @[LoadQueueFlag.scala 315:50]
          if (4'h4 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 316:33]
            uop_4_ctrl_replayInst <= io_loadIn_1_bits_uop_ctrl_replayInst; // @[LoadQueueFlag.scala 316:33]
          end else begin
            uop_4_ctrl_replayInst <= _GEN_22793;
          end
        end else begin
          uop_4_ctrl_replayInst <= _GEN_22793;
        end
      end else begin
        uop_4_ctrl_replayInst <= _GEN_22793;
      end
    end else begin
      uop_4_ctrl_replayInst <= _GEN_22793;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_1) begin // @[LoadQueueFlag.scala 309:50]
          if (4'h4 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 310:34]
            uop_4_pdest <= io_loadIn_1_bits_uop_pdest; // @[LoadQueueFlag.scala 310:34]
          end else begin
            uop_4_pdest <= _GEN_21465;
          end
        end else begin
          uop_4_pdest <= _GEN_21465;
        end
      end else begin
        uop_4_pdest <= _GEN_21465;
      end
    end else begin
      uop_4_pdest <= _GEN_21465;
    end
    if (io_enq_req_3_valid & ~enqCancel_3) begin // @[LoadQueueFlag.scala 204:43]
      if (4'h4 == io_enq_req_3_bits_lqIdx_value) begin // @[LoadQueueFlag.scala 206:18]
        uop_4_robIdx_flag <= io_enq_req_3_bits_robIdx_flag; // @[LoadQueueFlag.scala 206:18]
      end else begin
        uop_4_robIdx_flag <= _GEN_11906;
      end
    end else begin
      uop_4_robIdx_flag <= _GEN_11906;
    end
    if (io_enq_req_3_valid & ~enqCancel_3) begin // @[LoadQueueFlag.scala 204:43]
      if (4'h4 == io_enq_req_3_bits_lqIdx_value) begin // @[LoadQueueFlag.scala 206:18]
        uop_4_robIdx_value <= io_enq_req_3_bits_robIdx_value; // @[LoadQueueFlag.scala 206:18]
      end else begin
        uop_4_robIdx_value <= _GEN_11922;
      end
    end else begin
      uop_4_robIdx_value <= _GEN_11922;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'h5 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_5_cf_exceptionVec_4 <= io_loadIn_1_bits_uop_cf_exceptionVec_4; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_5_cf_exceptionVec_4 <= _GEN_21594;
          end
        end else begin
          uop_5_cf_exceptionVec_4 <= _GEN_21594;
        end
      end else begin
        uop_5_cf_exceptionVec_4 <= _GEN_21594;
      end
    end else begin
      uop_5_cf_exceptionVec_4 <= _GEN_21594;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'h5 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_5_cf_exceptionVec_5 <= io_loadIn_1_bits_uop_cf_exceptionVec_5; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_5_cf_exceptionVec_5 <= _GEN_21610;
          end
        end else begin
          uop_5_cf_exceptionVec_5 <= _GEN_21610;
        end
      end else begin
        uop_5_cf_exceptionVec_5 <= _GEN_21610;
      end
    end else begin
      uop_5_cf_exceptionVec_5 <= _GEN_21610;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'h5 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_5_cf_exceptionVec_13 <= io_loadIn_1_bits_uop_cf_exceptionVec_13; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_5_cf_exceptionVec_13 <= _GEN_21738;
          end
        end else begin
          uop_5_cf_exceptionVec_13 <= _GEN_21738;
        end
      end else begin
        uop_5_cf_exceptionVec_13 <= _GEN_21738;
      end
    end else begin
      uop_5_cf_exceptionVec_13 <= _GEN_21738;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'h5 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_5_cf_trigger_backendEn_1 <= io_loadIn_1_bits_uop_cf_trigger_backendEn_1; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_5_cf_trigger_backendEn_1 <= _GEN_21866;
          end
        end else begin
          uop_5_cf_trigger_backendEn_1 <= _GEN_21866;
        end
      end else begin
        uop_5_cf_trigger_backendEn_1 <= _GEN_21866;
      end
    end else begin
      uop_5_cf_trigger_backendEn_1 <= _GEN_21866;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'h5 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_5_cf_trigger_backendHit_0 <= io_loadIn_1_bits_uop_cf_trigger_backendHit_0; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_5_cf_trigger_backendHit_0 <= _GEN_21882;
          end
        end else begin
          uop_5_cf_trigger_backendHit_0 <= _GEN_21882;
        end
      end else begin
        uop_5_cf_trigger_backendHit_0 <= _GEN_21882;
      end
    end else begin
      uop_5_cf_trigger_backendHit_0 <= _GEN_21882;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'h5 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_5_cf_trigger_backendHit_1 <= io_loadIn_1_bits_uop_cf_trigger_backendHit_1; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_5_cf_trigger_backendHit_1 <= _GEN_21898;
          end
        end else begin
          uop_5_cf_trigger_backendHit_1 <= _GEN_21898;
        end
      end else begin
        uop_5_cf_trigger_backendHit_1 <= _GEN_21898;
      end
    end else begin
      uop_5_cf_trigger_backendHit_1 <= _GEN_21898;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'h5 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_5_cf_trigger_backendHit_4 <= io_loadIn_1_bits_uop_cf_trigger_backendHit_4; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_5_cf_trigger_backendHit_4 <= _GEN_21946;
          end
        end else begin
          uop_5_cf_trigger_backendHit_4 <= _GEN_21946;
        end
      end else begin
        uop_5_cf_trigger_backendHit_4 <= _GEN_21946;
      end
    end else begin
      uop_5_cf_trigger_backendHit_4 <= _GEN_21946;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_3) begin // @[LoadQueueFlag.scala 315:50]
          if (4'h5 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 316:33]
            uop_5_ctrl_fuOpType <= io_loadIn_1_bits_uop_ctrl_fuOpType; // @[LoadQueueFlag.scala 316:33]
          end else begin
            uop_5_ctrl_fuOpType <= _GEN_22378;
          end
        end else begin
          uop_5_ctrl_fuOpType <= _GEN_22378;
        end
      end else begin
        uop_5_ctrl_fuOpType <= _GEN_22378;
      end
    end else begin
      uop_5_ctrl_fuOpType <= _GEN_22378;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_3) begin // @[LoadQueueFlag.scala 315:50]
          if (4'h5 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 316:33]
            uop_5_ctrl_rfWen <= io_loadIn_1_bits_uop_ctrl_rfWen; // @[LoadQueueFlag.scala 316:33]
          end else begin
            uop_5_ctrl_rfWen <= _GEN_22394;
          end
        end else begin
          uop_5_ctrl_rfWen <= _GEN_22394;
        end
      end else begin
        uop_5_ctrl_rfWen <= _GEN_22394;
      end
    end else begin
      uop_5_ctrl_rfWen <= _GEN_22394;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_3) begin // @[LoadQueueFlag.scala 315:50]
          if (4'h5 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 316:33]
            uop_5_ctrl_fpWen <= io_loadIn_1_bits_uop_ctrl_fpWen; // @[LoadQueueFlag.scala 316:33]
          end else begin
            uop_5_ctrl_fpWen <= _GEN_22410;
          end
        end else begin
          uop_5_ctrl_fpWen <= _GEN_22410;
        end
      end else begin
        uop_5_ctrl_fpWen <= _GEN_22410;
      end
    end else begin
      uop_5_ctrl_fpWen <= _GEN_22410;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_3) begin // @[LoadQueueFlag.scala 315:50]
          if (4'h5 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 316:33]
            uop_5_ctrl_flushPipe <= 1'h0; // @[LoadQueueFlag.scala 316:33]
          end else begin
            uop_5_ctrl_flushPipe <= _GEN_22474;
          end
        end else begin
          uop_5_ctrl_flushPipe <= _GEN_22474;
        end
      end else begin
        uop_5_ctrl_flushPipe <= _GEN_22474;
      end
    end else begin
      uop_5_ctrl_flushPipe <= _GEN_22474;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_3) begin // @[LoadQueueFlag.scala 315:50]
          if (4'h5 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 316:33]
            uop_5_ctrl_replayInst <= io_loadIn_1_bits_uop_ctrl_replayInst; // @[LoadQueueFlag.scala 316:33]
          end else begin
            uop_5_ctrl_replayInst <= _GEN_22794;
          end
        end else begin
          uop_5_ctrl_replayInst <= _GEN_22794;
        end
      end else begin
        uop_5_ctrl_replayInst <= _GEN_22794;
      end
    end else begin
      uop_5_ctrl_replayInst <= _GEN_22794;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_1) begin // @[LoadQueueFlag.scala 309:50]
          if (4'h5 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 310:34]
            uop_5_pdest <= io_loadIn_1_bits_uop_pdest; // @[LoadQueueFlag.scala 310:34]
          end else begin
            uop_5_pdest <= _GEN_21466;
          end
        end else begin
          uop_5_pdest <= _GEN_21466;
        end
      end else begin
        uop_5_pdest <= _GEN_21466;
      end
    end else begin
      uop_5_pdest <= _GEN_21466;
    end
    if (io_enq_req_3_valid & ~enqCancel_3) begin // @[LoadQueueFlag.scala 204:43]
      if (4'h5 == io_enq_req_3_bits_lqIdx_value) begin // @[LoadQueueFlag.scala 206:18]
        uop_5_robIdx_flag <= io_enq_req_3_bits_robIdx_flag; // @[LoadQueueFlag.scala 206:18]
      end else begin
        uop_5_robIdx_flag <= _GEN_11907;
      end
    end else begin
      uop_5_robIdx_flag <= _GEN_11907;
    end
    if (io_enq_req_3_valid & ~enqCancel_3) begin // @[LoadQueueFlag.scala 204:43]
      if (4'h5 == io_enq_req_3_bits_lqIdx_value) begin // @[LoadQueueFlag.scala 206:18]
        uop_5_robIdx_value <= io_enq_req_3_bits_robIdx_value; // @[LoadQueueFlag.scala 206:18]
      end else begin
        uop_5_robIdx_value <= _GEN_11923;
      end
    end else begin
      uop_5_robIdx_value <= _GEN_11923;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'h6 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_6_cf_exceptionVec_4 <= io_loadIn_1_bits_uop_cf_exceptionVec_4; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_6_cf_exceptionVec_4 <= _GEN_21595;
          end
        end else begin
          uop_6_cf_exceptionVec_4 <= _GEN_21595;
        end
      end else begin
        uop_6_cf_exceptionVec_4 <= _GEN_21595;
      end
    end else begin
      uop_6_cf_exceptionVec_4 <= _GEN_21595;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'h6 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_6_cf_exceptionVec_5 <= io_loadIn_1_bits_uop_cf_exceptionVec_5; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_6_cf_exceptionVec_5 <= _GEN_21611;
          end
        end else begin
          uop_6_cf_exceptionVec_5 <= _GEN_21611;
        end
      end else begin
        uop_6_cf_exceptionVec_5 <= _GEN_21611;
      end
    end else begin
      uop_6_cf_exceptionVec_5 <= _GEN_21611;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'h6 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_6_cf_exceptionVec_13 <= io_loadIn_1_bits_uop_cf_exceptionVec_13; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_6_cf_exceptionVec_13 <= _GEN_21739;
          end
        end else begin
          uop_6_cf_exceptionVec_13 <= _GEN_21739;
        end
      end else begin
        uop_6_cf_exceptionVec_13 <= _GEN_21739;
      end
    end else begin
      uop_6_cf_exceptionVec_13 <= _GEN_21739;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'h6 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_6_cf_trigger_backendEn_1 <= io_loadIn_1_bits_uop_cf_trigger_backendEn_1; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_6_cf_trigger_backendEn_1 <= _GEN_21867;
          end
        end else begin
          uop_6_cf_trigger_backendEn_1 <= _GEN_21867;
        end
      end else begin
        uop_6_cf_trigger_backendEn_1 <= _GEN_21867;
      end
    end else begin
      uop_6_cf_trigger_backendEn_1 <= _GEN_21867;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'h6 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_6_cf_trigger_backendHit_0 <= io_loadIn_1_bits_uop_cf_trigger_backendHit_0; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_6_cf_trigger_backendHit_0 <= _GEN_21883;
          end
        end else begin
          uop_6_cf_trigger_backendHit_0 <= _GEN_21883;
        end
      end else begin
        uop_6_cf_trigger_backendHit_0 <= _GEN_21883;
      end
    end else begin
      uop_6_cf_trigger_backendHit_0 <= _GEN_21883;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'h6 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_6_cf_trigger_backendHit_1 <= io_loadIn_1_bits_uop_cf_trigger_backendHit_1; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_6_cf_trigger_backendHit_1 <= _GEN_21899;
          end
        end else begin
          uop_6_cf_trigger_backendHit_1 <= _GEN_21899;
        end
      end else begin
        uop_6_cf_trigger_backendHit_1 <= _GEN_21899;
      end
    end else begin
      uop_6_cf_trigger_backendHit_1 <= _GEN_21899;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'h6 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_6_cf_trigger_backendHit_4 <= io_loadIn_1_bits_uop_cf_trigger_backendHit_4; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_6_cf_trigger_backendHit_4 <= _GEN_21947;
          end
        end else begin
          uop_6_cf_trigger_backendHit_4 <= _GEN_21947;
        end
      end else begin
        uop_6_cf_trigger_backendHit_4 <= _GEN_21947;
      end
    end else begin
      uop_6_cf_trigger_backendHit_4 <= _GEN_21947;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_3) begin // @[LoadQueueFlag.scala 315:50]
          if (4'h6 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 316:33]
            uop_6_ctrl_fuOpType <= io_loadIn_1_bits_uop_ctrl_fuOpType; // @[LoadQueueFlag.scala 316:33]
          end else begin
            uop_6_ctrl_fuOpType <= _GEN_22379;
          end
        end else begin
          uop_6_ctrl_fuOpType <= _GEN_22379;
        end
      end else begin
        uop_6_ctrl_fuOpType <= _GEN_22379;
      end
    end else begin
      uop_6_ctrl_fuOpType <= _GEN_22379;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_3) begin // @[LoadQueueFlag.scala 315:50]
          if (4'h6 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 316:33]
            uop_6_ctrl_rfWen <= io_loadIn_1_bits_uop_ctrl_rfWen; // @[LoadQueueFlag.scala 316:33]
          end else begin
            uop_6_ctrl_rfWen <= _GEN_22395;
          end
        end else begin
          uop_6_ctrl_rfWen <= _GEN_22395;
        end
      end else begin
        uop_6_ctrl_rfWen <= _GEN_22395;
      end
    end else begin
      uop_6_ctrl_rfWen <= _GEN_22395;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_3) begin // @[LoadQueueFlag.scala 315:50]
          if (4'h6 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 316:33]
            uop_6_ctrl_fpWen <= io_loadIn_1_bits_uop_ctrl_fpWen; // @[LoadQueueFlag.scala 316:33]
          end else begin
            uop_6_ctrl_fpWen <= _GEN_22411;
          end
        end else begin
          uop_6_ctrl_fpWen <= _GEN_22411;
        end
      end else begin
        uop_6_ctrl_fpWen <= _GEN_22411;
      end
    end else begin
      uop_6_ctrl_fpWen <= _GEN_22411;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_3) begin // @[LoadQueueFlag.scala 315:50]
          if (4'h6 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 316:33]
            uop_6_ctrl_flushPipe <= 1'h0; // @[LoadQueueFlag.scala 316:33]
          end else begin
            uop_6_ctrl_flushPipe <= _GEN_22475;
          end
        end else begin
          uop_6_ctrl_flushPipe <= _GEN_22475;
        end
      end else begin
        uop_6_ctrl_flushPipe <= _GEN_22475;
      end
    end else begin
      uop_6_ctrl_flushPipe <= _GEN_22475;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_3) begin // @[LoadQueueFlag.scala 315:50]
          if (4'h6 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 316:33]
            uop_6_ctrl_replayInst <= io_loadIn_1_bits_uop_ctrl_replayInst; // @[LoadQueueFlag.scala 316:33]
          end else begin
            uop_6_ctrl_replayInst <= _GEN_22795;
          end
        end else begin
          uop_6_ctrl_replayInst <= _GEN_22795;
        end
      end else begin
        uop_6_ctrl_replayInst <= _GEN_22795;
      end
    end else begin
      uop_6_ctrl_replayInst <= _GEN_22795;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_1) begin // @[LoadQueueFlag.scala 309:50]
          if (4'h6 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 310:34]
            uop_6_pdest <= io_loadIn_1_bits_uop_pdest; // @[LoadQueueFlag.scala 310:34]
          end else begin
            uop_6_pdest <= _GEN_21467;
          end
        end else begin
          uop_6_pdest <= _GEN_21467;
        end
      end else begin
        uop_6_pdest <= _GEN_21467;
      end
    end else begin
      uop_6_pdest <= _GEN_21467;
    end
    if (io_enq_req_3_valid & ~enqCancel_3) begin // @[LoadQueueFlag.scala 204:43]
      if (4'h6 == io_enq_req_3_bits_lqIdx_value) begin // @[LoadQueueFlag.scala 206:18]
        uop_6_robIdx_flag <= io_enq_req_3_bits_robIdx_flag; // @[LoadQueueFlag.scala 206:18]
      end else begin
        uop_6_robIdx_flag <= _GEN_11908;
      end
    end else begin
      uop_6_robIdx_flag <= _GEN_11908;
    end
    if (io_enq_req_3_valid & ~enqCancel_3) begin // @[LoadQueueFlag.scala 204:43]
      if (4'h6 == io_enq_req_3_bits_lqIdx_value) begin // @[LoadQueueFlag.scala 206:18]
        uop_6_robIdx_value <= io_enq_req_3_bits_robIdx_value; // @[LoadQueueFlag.scala 206:18]
      end else begin
        uop_6_robIdx_value <= _GEN_11924;
      end
    end else begin
      uop_6_robIdx_value <= _GEN_11924;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'h7 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_7_cf_exceptionVec_4 <= io_loadIn_1_bits_uop_cf_exceptionVec_4; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_7_cf_exceptionVec_4 <= _GEN_21596;
          end
        end else begin
          uop_7_cf_exceptionVec_4 <= _GEN_21596;
        end
      end else begin
        uop_7_cf_exceptionVec_4 <= _GEN_21596;
      end
    end else begin
      uop_7_cf_exceptionVec_4 <= _GEN_21596;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'h7 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_7_cf_exceptionVec_5 <= io_loadIn_1_bits_uop_cf_exceptionVec_5; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_7_cf_exceptionVec_5 <= _GEN_21612;
          end
        end else begin
          uop_7_cf_exceptionVec_5 <= _GEN_21612;
        end
      end else begin
        uop_7_cf_exceptionVec_5 <= _GEN_21612;
      end
    end else begin
      uop_7_cf_exceptionVec_5 <= _GEN_21612;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'h7 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_7_cf_exceptionVec_13 <= io_loadIn_1_bits_uop_cf_exceptionVec_13; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_7_cf_exceptionVec_13 <= _GEN_21740;
          end
        end else begin
          uop_7_cf_exceptionVec_13 <= _GEN_21740;
        end
      end else begin
        uop_7_cf_exceptionVec_13 <= _GEN_21740;
      end
    end else begin
      uop_7_cf_exceptionVec_13 <= _GEN_21740;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'h7 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_7_cf_trigger_backendEn_1 <= io_loadIn_1_bits_uop_cf_trigger_backendEn_1; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_7_cf_trigger_backendEn_1 <= _GEN_21868;
          end
        end else begin
          uop_7_cf_trigger_backendEn_1 <= _GEN_21868;
        end
      end else begin
        uop_7_cf_trigger_backendEn_1 <= _GEN_21868;
      end
    end else begin
      uop_7_cf_trigger_backendEn_1 <= _GEN_21868;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'h7 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_7_cf_trigger_backendHit_0 <= io_loadIn_1_bits_uop_cf_trigger_backendHit_0; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_7_cf_trigger_backendHit_0 <= _GEN_21884;
          end
        end else begin
          uop_7_cf_trigger_backendHit_0 <= _GEN_21884;
        end
      end else begin
        uop_7_cf_trigger_backendHit_0 <= _GEN_21884;
      end
    end else begin
      uop_7_cf_trigger_backendHit_0 <= _GEN_21884;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'h7 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_7_cf_trigger_backendHit_1 <= io_loadIn_1_bits_uop_cf_trigger_backendHit_1; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_7_cf_trigger_backendHit_1 <= _GEN_21900;
          end
        end else begin
          uop_7_cf_trigger_backendHit_1 <= _GEN_21900;
        end
      end else begin
        uop_7_cf_trigger_backendHit_1 <= _GEN_21900;
      end
    end else begin
      uop_7_cf_trigger_backendHit_1 <= _GEN_21900;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'h7 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_7_cf_trigger_backendHit_4 <= io_loadIn_1_bits_uop_cf_trigger_backendHit_4; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_7_cf_trigger_backendHit_4 <= _GEN_21948;
          end
        end else begin
          uop_7_cf_trigger_backendHit_4 <= _GEN_21948;
        end
      end else begin
        uop_7_cf_trigger_backendHit_4 <= _GEN_21948;
      end
    end else begin
      uop_7_cf_trigger_backendHit_4 <= _GEN_21948;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_3) begin // @[LoadQueueFlag.scala 315:50]
          if (4'h7 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 316:33]
            uop_7_ctrl_fuOpType <= io_loadIn_1_bits_uop_ctrl_fuOpType; // @[LoadQueueFlag.scala 316:33]
          end else begin
            uop_7_ctrl_fuOpType <= _GEN_22380;
          end
        end else begin
          uop_7_ctrl_fuOpType <= _GEN_22380;
        end
      end else begin
        uop_7_ctrl_fuOpType <= _GEN_22380;
      end
    end else begin
      uop_7_ctrl_fuOpType <= _GEN_22380;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_3) begin // @[LoadQueueFlag.scala 315:50]
          if (4'h7 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 316:33]
            uop_7_ctrl_rfWen <= io_loadIn_1_bits_uop_ctrl_rfWen; // @[LoadQueueFlag.scala 316:33]
          end else begin
            uop_7_ctrl_rfWen <= _GEN_22396;
          end
        end else begin
          uop_7_ctrl_rfWen <= _GEN_22396;
        end
      end else begin
        uop_7_ctrl_rfWen <= _GEN_22396;
      end
    end else begin
      uop_7_ctrl_rfWen <= _GEN_22396;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_3) begin // @[LoadQueueFlag.scala 315:50]
          if (4'h7 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 316:33]
            uop_7_ctrl_fpWen <= io_loadIn_1_bits_uop_ctrl_fpWen; // @[LoadQueueFlag.scala 316:33]
          end else begin
            uop_7_ctrl_fpWen <= _GEN_22412;
          end
        end else begin
          uop_7_ctrl_fpWen <= _GEN_22412;
        end
      end else begin
        uop_7_ctrl_fpWen <= _GEN_22412;
      end
    end else begin
      uop_7_ctrl_fpWen <= _GEN_22412;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_3) begin // @[LoadQueueFlag.scala 315:50]
          if (4'h7 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 316:33]
            uop_7_ctrl_flushPipe <= 1'h0; // @[LoadQueueFlag.scala 316:33]
          end else begin
            uop_7_ctrl_flushPipe <= _GEN_22476;
          end
        end else begin
          uop_7_ctrl_flushPipe <= _GEN_22476;
        end
      end else begin
        uop_7_ctrl_flushPipe <= _GEN_22476;
      end
    end else begin
      uop_7_ctrl_flushPipe <= _GEN_22476;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_3) begin // @[LoadQueueFlag.scala 315:50]
          if (4'h7 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 316:33]
            uop_7_ctrl_replayInst <= io_loadIn_1_bits_uop_ctrl_replayInst; // @[LoadQueueFlag.scala 316:33]
          end else begin
            uop_7_ctrl_replayInst <= _GEN_22796;
          end
        end else begin
          uop_7_ctrl_replayInst <= _GEN_22796;
        end
      end else begin
        uop_7_ctrl_replayInst <= _GEN_22796;
      end
    end else begin
      uop_7_ctrl_replayInst <= _GEN_22796;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_1) begin // @[LoadQueueFlag.scala 309:50]
          if (4'h7 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 310:34]
            uop_7_pdest <= io_loadIn_1_bits_uop_pdest; // @[LoadQueueFlag.scala 310:34]
          end else begin
            uop_7_pdest <= _GEN_21468;
          end
        end else begin
          uop_7_pdest <= _GEN_21468;
        end
      end else begin
        uop_7_pdest <= _GEN_21468;
      end
    end else begin
      uop_7_pdest <= _GEN_21468;
    end
    if (io_enq_req_3_valid & ~enqCancel_3) begin // @[LoadQueueFlag.scala 204:43]
      if (4'h7 == io_enq_req_3_bits_lqIdx_value) begin // @[LoadQueueFlag.scala 206:18]
        uop_7_robIdx_flag <= io_enq_req_3_bits_robIdx_flag; // @[LoadQueueFlag.scala 206:18]
      end else begin
        uop_7_robIdx_flag <= _GEN_11909;
      end
    end else begin
      uop_7_robIdx_flag <= _GEN_11909;
    end
    if (io_enq_req_3_valid & ~enqCancel_3) begin // @[LoadQueueFlag.scala 204:43]
      if (4'h7 == io_enq_req_3_bits_lqIdx_value) begin // @[LoadQueueFlag.scala 206:18]
        uop_7_robIdx_value <= io_enq_req_3_bits_robIdx_value; // @[LoadQueueFlag.scala 206:18]
      end else begin
        uop_7_robIdx_value <= _GEN_11925;
      end
    end else begin
      uop_7_robIdx_value <= _GEN_11925;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'h8 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_8_cf_exceptionVec_4 <= io_loadIn_1_bits_uop_cf_exceptionVec_4; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_8_cf_exceptionVec_4 <= _GEN_21597;
          end
        end else begin
          uop_8_cf_exceptionVec_4 <= _GEN_21597;
        end
      end else begin
        uop_8_cf_exceptionVec_4 <= _GEN_21597;
      end
    end else begin
      uop_8_cf_exceptionVec_4 <= _GEN_21597;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'h8 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_8_cf_exceptionVec_5 <= io_loadIn_1_bits_uop_cf_exceptionVec_5; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_8_cf_exceptionVec_5 <= _GEN_21613;
          end
        end else begin
          uop_8_cf_exceptionVec_5 <= _GEN_21613;
        end
      end else begin
        uop_8_cf_exceptionVec_5 <= _GEN_21613;
      end
    end else begin
      uop_8_cf_exceptionVec_5 <= _GEN_21613;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'h8 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_8_cf_exceptionVec_13 <= io_loadIn_1_bits_uop_cf_exceptionVec_13; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_8_cf_exceptionVec_13 <= _GEN_21741;
          end
        end else begin
          uop_8_cf_exceptionVec_13 <= _GEN_21741;
        end
      end else begin
        uop_8_cf_exceptionVec_13 <= _GEN_21741;
      end
    end else begin
      uop_8_cf_exceptionVec_13 <= _GEN_21741;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'h8 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_8_cf_trigger_backendEn_1 <= io_loadIn_1_bits_uop_cf_trigger_backendEn_1; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_8_cf_trigger_backendEn_1 <= _GEN_21869;
          end
        end else begin
          uop_8_cf_trigger_backendEn_1 <= _GEN_21869;
        end
      end else begin
        uop_8_cf_trigger_backendEn_1 <= _GEN_21869;
      end
    end else begin
      uop_8_cf_trigger_backendEn_1 <= _GEN_21869;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'h8 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_8_cf_trigger_backendHit_0 <= io_loadIn_1_bits_uop_cf_trigger_backendHit_0; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_8_cf_trigger_backendHit_0 <= _GEN_21885;
          end
        end else begin
          uop_8_cf_trigger_backendHit_0 <= _GEN_21885;
        end
      end else begin
        uop_8_cf_trigger_backendHit_0 <= _GEN_21885;
      end
    end else begin
      uop_8_cf_trigger_backendHit_0 <= _GEN_21885;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'h8 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_8_cf_trigger_backendHit_1 <= io_loadIn_1_bits_uop_cf_trigger_backendHit_1; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_8_cf_trigger_backendHit_1 <= _GEN_21901;
          end
        end else begin
          uop_8_cf_trigger_backendHit_1 <= _GEN_21901;
        end
      end else begin
        uop_8_cf_trigger_backendHit_1 <= _GEN_21901;
      end
    end else begin
      uop_8_cf_trigger_backendHit_1 <= _GEN_21901;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'h8 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_8_cf_trigger_backendHit_4 <= io_loadIn_1_bits_uop_cf_trigger_backendHit_4; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_8_cf_trigger_backendHit_4 <= _GEN_21949;
          end
        end else begin
          uop_8_cf_trigger_backendHit_4 <= _GEN_21949;
        end
      end else begin
        uop_8_cf_trigger_backendHit_4 <= _GEN_21949;
      end
    end else begin
      uop_8_cf_trigger_backendHit_4 <= _GEN_21949;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_3) begin // @[LoadQueueFlag.scala 315:50]
          if (4'h8 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 316:33]
            uop_8_ctrl_fuOpType <= io_loadIn_1_bits_uop_ctrl_fuOpType; // @[LoadQueueFlag.scala 316:33]
          end else begin
            uop_8_ctrl_fuOpType <= _GEN_22381;
          end
        end else begin
          uop_8_ctrl_fuOpType <= _GEN_22381;
        end
      end else begin
        uop_8_ctrl_fuOpType <= _GEN_22381;
      end
    end else begin
      uop_8_ctrl_fuOpType <= _GEN_22381;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_3) begin // @[LoadQueueFlag.scala 315:50]
          if (4'h8 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 316:33]
            uop_8_ctrl_rfWen <= io_loadIn_1_bits_uop_ctrl_rfWen; // @[LoadQueueFlag.scala 316:33]
          end else begin
            uop_8_ctrl_rfWen <= _GEN_22397;
          end
        end else begin
          uop_8_ctrl_rfWen <= _GEN_22397;
        end
      end else begin
        uop_8_ctrl_rfWen <= _GEN_22397;
      end
    end else begin
      uop_8_ctrl_rfWen <= _GEN_22397;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_3) begin // @[LoadQueueFlag.scala 315:50]
          if (4'h8 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 316:33]
            uop_8_ctrl_fpWen <= io_loadIn_1_bits_uop_ctrl_fpWen; // @[LoadQueueFlag.scala 316:33]
          end else begin
            uop_8_ctrl_fpWen <= _GEN_22413;
          end
        end else begin
          uop_8_ctrl_fpWen <= _GEN_22413;
        end
      end else begin
        uop_8_ctrl_fpWen <= _GEN_22413;
      end
    end else begin
      uop_8_ctrl_fpWen <= _GEN_22413;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_3) begin // @[LoadQueueFlag.scala 315:50]
          if (4'h8 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 316:33]
            uop_8_ctrl_flushPipe <= 1'h0; // @[LoadQueueFlag.scala 316:33]
          end else begin
            uop_8_ctrl_flushPipe <= _GEN_22477;
          end
        end else begin
          uop_8_ctrl_flushPipe <= _GEN_22477;
        end
      end else begin
        uop_8_ctrl_flushPipe <= _GEN_22477;
      end
    end else begin
      uop_8_ctrl_flushPipe <= _GEN_22477;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_3) begin // @[LoadQueueFlag.scala 315:50]
          if (4'h8 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 316:33]
            uop_8_ctrl_replayInst <= io_loadIn_1_bits_uop_ctrl_replayInst; // @[LoadQueueFlag.scala 316:33]
          end else begin
            uop_8_ctrl_replayInst <= _GEN_22797;
          end
        end else begin
          uop_8_ctrl_replayInst <= _GEN_22797;
        end
      end else begin
        uop_8_ctrl_replayInst <= _GEN_22797;
      end
    end else begin
      uop_8_ctrl_replayInst <= _GEN_22797;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_1) begin // @[LoadQueueFlag.scala 309:50]
          if (4'h8 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 310:34]
            uop_8_pdest <= io_loadIn_1_bits_uop_pdest; // @[LoadQueueFlag.scala 310:34]
          end else begin
            uop_8_pdest <= _GEN_21469;
          end
        end else begin
          uop_8_pdest <= _GEN_21469;
        end
      end else begin
        uop_8_pdest <= _GEN_21469;
      end
    end else begin
      uop_8_pdest <= _GEN_21469;
    end
    if (io_enq_req_3_valid & ~enqCancel_3) begin // @[LoadQueueFlag.scala 204:43]
      if (4'h8 == io_enq_req_3_bits_lqIdx_value) begin // @[LoadQueueFlag.scala 206:18]
        uop_8_robIdx_flag <= io_enq_req_3_bits_robIdx_flag; // @[LoadQueueFlag.scala 206:18]
      end else begin
        uop_8_robIdx_flag <= _GEN_11910;
      end
    end else begin
      uop_8_robIdx_flag <= _GEN_11910;
    end
    if (io_enq_req_3_valid & ~enqCancel_3) begin // @[LoadQueueFlag.scala 204:43]
      if (4'h8 == io_enq_req_3_bits_lqIdx_value) begin // @[LoadQueueFlag.scala 206:18]
        uop_8_robIdx_value <= io_enq_req_3_bits_robIdx_value; // @[LoadQueueFlag.scala 206:18]
      end else begin
        uop_8_robIdx_value <= _GEN_11926;
      end
    end else begin
      uop_8_robIdx_value <= _GEN_11926;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'h9 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_9_cf_exceptionVec_4 <= io_loadIn_1_bits_uop_cf_exceptionVec_4; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_9_cf_exceptionVec_4 <= _GEN_21598;
          end
        end else begin
          uop_9_cf_exceptionVec_4 <= _GEN_21598;
        end
      end else begin
        uop_9_cf_exceptionVec_4 <= _GEN_21598;
      end
    end else begin
      uop_9_cf_exceptionVec_4 <= _GEN_21598;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'h9 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_9_cf_exceptionVec_5 <= io_loadIn_1_bits_uop_cf_exceptionVec_5; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_9_cf_exceptionVec_5 <= _GEN_21614;
          end
        end else begin
          uop_9_cf_exceptionVec_5 <= _GEN_21614;
        end
      end else begin
        uop_9_cf_exceptionVec_5 <= _GEN_21614;
      end
    end else begin
      uop_9_cf_exceptionVec_5 <= _GEN_21614;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'h9 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_9_cf_exceptionVec_13 <= io_loadIn_1_bits_uop_cf_exceptionVec_13; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_9_cf_exceptionVec_13 <= _GEN_21742;
          end
        end else begin
          uop_9_cf_exceptionVec_13 <= _GEN_21742;
        end
      end else begin
        uop_9_cf_exceptionVec_13 <= _GEN_21742;
      end
    end else begin
      uop_9_cf_exceptionVec_13 <= _GEN_21742;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'h9 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_9_cf_trigger_backendEn_1 <= io_loadIn_1_bits_uop_cf_trigger_backendEn_1; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_9_cf_trigger_backendEn_1 <= _GEN_21870;
          end
        end else begin
          uop_9_cf_trigger_backendEn_1 <= _GEN_21870;
        end
      end else begin
        uop_9_cf_trigger_backendEn_1 <= _GEN_21870;
      end
    end else begin
      uop_9_cf_trigger_backendEn_1 <= _GEN_21870;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'h9 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_9_cf_trigger_backendHit_0 <= io_loadIn_1_bits_uop_cf_trigger_backendHit_0; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_9_cf_trigger_backendHit_0 <= _GEN_21886;
          end
        end else begin
          uop_9_cf_trigger_backendHit_0 <= _GEN_21886;
        end
      end else begin
        uop_9_cf_trigger_backendHit_0 <= _GEN_21886;
      end
    end else begin
      uop_9_cf_trigger_backendHit_0 <= _GEN_21886;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'h9 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_9_cf_trigger_backendHit_1 <= io_loadIn_1_bits_uop_cf_trigger_backendHit_1; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_9_cf_trigger_backendHit_1 <= _GEN_21902;
          end
        end else begin
          uop_9_cf_trigger_backendHit_1 <= _GEN_21902;
        end
      end else begin
        uop_9_cf_trigger_backendHit_1 <= _GEN_21902;
      end
    end else begin
      uop_9_cf_trigger_backendHit_1 <= _GEN_21902;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'h9 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_9_cf_trigger_backendHit_4 <= io_loadIn_1_bits_uop_cf_trigger_backendHit_4; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_9_cf_trigger_backendHit_4 <= _GEN_21950;
          end
        end else begin
          uop_9_cf_trigger_backendHit_4 <= _GEN_21950;
        end
      end else begin
        uop_9_cf_trigger_backendHit_4 <= _GEN_21950;
      end
    end else begin
      uop_9_cf_trigger_backendHit_4 <= _GEN_21950;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_3) begin // @[LoadQueueFlag.scala 315:50]
          if (4'h9 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 316:33]
            uop_9_ctrl_fuOpType <= io_loadIn_1_bits_uop_ctrl_fuOpType; // @[LoadQueueFlag.scala 316:33]
          end else begin
            uop_9_ctrl_fuOpType <= _GEN_22382;
          end
        end else begin
          uop_9_ctrl_fuOpType <= _GEN_22382;
        end
      end else begin
        uop_9_ctrl_fuOpType <= _GEN_22382;
      end
    end else begin
      uop_9_ctrl_fuOpType <= _GEN_22382;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_3) begin // @[LoadQueueFlag.scala 315:50]
          if (4'h9 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 316:33]
            uop_9_ctrl_rfWen <= io_loadIn_1_bits_uop_ctrl_rfWen; // @[LoadQueueFlag.scala 316:33]
          end else begin
            uop_9_ctrl_rfWen <= _GEN_22398;
          end
        end else begin
          uop_9_ctrl_rfWen <= _GEN_22398;
        end
      end else begin
        uop_9_ctrl_rfWen <= _GEN_22398;
      end
    end else begin
      uop_9_ctrl_rfWen <= _GEN_22398;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_3) begin // @[LoadQueueFlag.scala 315:50]
          if (4'h9 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 316:33]
            uop_9_ctrl_fpWen <= io_loadIn_1_bits_uop_ctrl_fpWen; // @[LoadQueueFlag.scala 316:33]
          end else begin
            uop_9_ctrl_fpWen <= _GEN_22414;
          end
        end else begin
          uop_9_ctrl_fpWen <= _GEN_22414;
        end
      end else begin
        uop_9_ctrl_fpWen <= _GEN_22414;
      end
    end else begin
      uop_9_ctrl_fpWen <= _GEN_22414;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_3) begin // @[LoadQueueFlag.scala 315:50]
          if (4'h9 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 316:33]
            uop_9_ctrl_flushPipe <= 1'h0; // @[LoadQueueFlag.scala 316:33]
          end else begin
            uop_9_ctrl_flushPipe <= _GEN_22478;
          end
        end else begin
          uop_9_ctrl_flushPipe <= _GEN_22478;
        end
      end else begin
        uop_9_ctrl_flushPipe <= _GEN_22478;
      end
    end else begin
      uop_9_ctrl_flushPipe <= _GEN_22478;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_3) begin // @[LoadQueueFlag.scala 315:50]
          if (4'h9 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 316:33]
            uop_9_ctrl_replayInst <= io_loadIn_1_bits_uop_ctrl_replayInst; // @[LoadQueueFlag.scala 316:33]
          end else begin
            uop_9_ctrl_replayInst <= _GEN_22798;
          end
        end else begin
          uop_9_ctrl_replayInst <= _GEN_22798;
        end
      end else begin
        uop_9_ctrl_replayInst <= _GEN_22798;
      end
    end else begin
      uop_9_ctrl_replayInst <= _GEN_22798;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_1) begin // @[LoadQueueFlag.scala 309:50]
          if (4'h9 == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 310:34]
            uop_9_pdest <= io_loadIn_1_bits_uop_pdest; // @[LoadQueueFlag.scala 310:34]
          end else begin
            uop_9_pdest <= _GEN_21470;
          end
        end else begin
          uop_9_pdest <= _GEN_21470;
        end
      end else begin
        uop_9_pdest <= _GEN_21470;
      end
    end else begin
      uop_9_pdest <= _GEN_21470;
    end
    if (io_enq_req_3_valid & ~enqCancel_3) begin // @[LoadQueueFlag.scala 204:43]
      if (4'h9 == io_enq_req_3_bits_lqIdx_value) begin // @[LoadQueueFlag.scala 206:18]
        uop_9_robIdx_flag <= io_enq_req_3_bits_robIdx_flag; // @[LoadQueueFlag.scala 206:18]
      end else begin
        uop_9_robIdx_flag <= _GEN_11911;
      end
    end else begin
      uop_9_robIdx_flag <= _GEN_11911;
    end
    if (io_enq_req_3_valid & ~enqCancel_3) begin // @[LoadQueueFlag.scala 204:43]
      if (4'h9 == io_enq_req_3_bits_lqIdx_value) begin // @[LoadQueueFlag.scala 206:18]
        uop_9_robIdx_value <= io_enq_req_3_bits_robIdx_value; // @[LoadQueueFlag.scala 206:18]
      end else begin
        uop_9_robIdx_value <= _GEN_11927;
      end
    end else begin
      uop_9_robIdx_value <= _GEN_11927;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'ha == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_10_cf_exceptionVec_4 <= io_loadIn_1_bits_uop_cf_exceptionVec_4; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_10_cf_exceptionVec_4 <= _GEN_21599;
          end
        end else begin
          uop_10_cf_exceptionVec_4 <= _GEN_21599;
        end
      end else begin
        uop_10_cf_exceptionVec_4 <= _GEN_21599;
      end
    end else begin
      uop_10_cf_exceptionVec_4 <= _GEN_21599;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'ha == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_10_cf_exceptionVec_5 <= io_loadIn_1_bits_uop_cf_exceptionVec_5; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_10_cf_exceptionVec_5 <= _GEN_21615;
          end
        end else begin
          uop_10_cf_exceptionVec_5 <= _GEN_21615;
        end
      end else begin
        uop_10_cf_exceptionVec_5 <= _GEN_21615;
      end
    end else begin
      uop_10_cf_exceptionVec_5 <= _GEN_21615;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'ha == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_10_cf_exceptionVec_13 <= io_loadIn_1_bits_uop_cf_exceptionVec_13; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_10_cf_exceptionVec_13 <= _GEN_21743;
          end
        end else begin
          uop_10_cf_exceptionVec_13 <= _GEN_21743;
        end
      end else begin
        uop_10_cf_exceptionVec_13 <= _GEN_21743;
      end
    end else begin
      uop_10_cf_exceptionVec_13 <= _GEN_21743;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'ha == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_10_cf_trigger_backendEn_1 <= io_loadIn_1_bits_uop_cf_trigger_backendEn_1; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_10_cf_trigger_backendEn_1 <= _GEN_21871;
          end
        end else begin
          uop_10_cf_trigger_backendEn_1 <= _GEN_21871;
        end
      end else begin
        uop_10_cf_trigger_backendEn_1 <= _GEN_21871;
      end
    end else begin
      uop_10_cf_trigger_backendEn_1 <= _GEN_21871;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'ha == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_10_cf_trigger_backendHit_0 <= io_loadIn_1_bits_uop_cf_trigger_backendHit_0; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_10_cf_trigger_backendHit_0 <= _GEN_21887;
          end
        end else begin
          uop_10_cf_trigger_backendHit_0 <= _GEN_21887;
        end
      end else begin
        uop_10_cf_trigger_backendHit_0 <= _GEN_21887;
      end
    end else begin
      uop_10_cf_trigger_backendHit_0 <= _GEN_21887;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'ha == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_10_cf_trigger_backendHit_1 <= io_loadIn_1_bits_uop_cf_trigger_backendHit_1; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_10_cf_trigger_backendHit_1 <= _GEN_21903;
          end
        end else begin
          uop_10_cf_trigger_backendHit_1 <= _GEN_21903;
        end
      end else begin
        uop_10_cf_trigger_backendHit_1 <= _GEN_21903;
      end
    end else begin
      uop_10_cf_trigger_backendHit_1 <= _GEN_21903;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'ha == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_10_cf_trigger_backendHit_4 <= io_loadIn_1_bits_uop_cf_trigger_backendHit_4; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_10_cf_trigger_backendHit_4 <= _GEN_21951;
          end
        end else begin
          uop_10_cf_trigger_backendHit_4 <= _GEN_21951;
        end
      end else begin
        uop_10_cf_trigger_backendHit_4 <= _GEN_21951;
      end
    end else begin
      uop_10_cf_trigger_backendHit_4 <= _GEN_21951;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_3) begin // @[LoadQueueFlag.scala 315:50]
          if (4'ha == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 316:33]
            uop_10_ctrl_fuOpType <= io_loadIn_1_bits_uop_ctrl_fuOpType; // @[LoadQueueFlag.scala 316:33]
          end else begin
            uop_10_ctrl_fuOpType <= _GEN_22383;
          end
        end else begin
          uop_10_ctrl_fuOpType <= _GEN_22383;
        end
      end else begin
        uop_10_ctrl_fuOpType <= _GEN_22383;
      end
    end else begin
      uop_10_ctrl_fuOpType <= _GEN_22383;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_3) begin // @[LoadQueueFlag.scala 315:50]
          if (4'ha == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 316:33]
            uop_10_ctrl_rfWen <= io_loadIn_1_bits_uop_ctrl_rfWen; // @[LoadQueueFlag.scala 316:33]
          end else begin
            uop_10_ctrl_rfWen <= _GEN_22399;
          end
        end else begin
          uop_10_ctrl_rfWen <= _GEN_22399;
        end
      end else begin
        uop_10_ctrl_rfWen <= _GEN_22399;
      end
    end else begin
      uop_10_ctrl_rfWen <= _GEN_22399;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_3) begin // @[LoadQueueFlag.scala 315:50]
          if (4'ha == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 316:33]
            uop_10_ctrl_fpWen <= io_loadIn_1_bits_uop_ctrl_fpWen; // @[LoadQueueFlag.scala 316:33]
          end else begin
            uop_10_ctrl_fpWen <= _GEN_22415;
          end
        end else begin
          uop_10_ctrl_fpWen <= _GEN_22415;
        end
      end else begin
        uop_10_ctrl_fpWen <= _GEN_22415;
      end
    end else begin
      uop_10_ctrl_fpWen <= _GEN_22415;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_3) begin // @[LoadQueueFlag.scala 315:50]
          if (4'ha == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 316:33]
            uop_10_ctrl_flushPipe <= 1'h0; // @[LoadQueueFlag.scala 316:33]
          end else begin
            uop_10_ctrl_flushPipe <= _GEN_22479;
          end
        end else begin
          uop_10_ctrl_flushPipe <= _GEN_22479;
        end
      end else begin
        uop_10_ctrl_flushPipe <= _GEN_22479;
      end
    end else begin
      uop_10_ctrl_flushPipe <= _GEN_22479;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_3) begin // @[LoadQueueFlag.scala 315:50]
          if (4'ha == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 316:33]
            uop_10_ctrl_replayInst <= io_loadIn_1_bits_uop_ctrl_replayInst; // @[LoadQueueFlag.scala 316:33]
          end else begin
            uop_10_ctrl_replayInst <= _GEN_22799;
          end
        end else begin
          uop_10_ctrl_replayInst <= _GEN_22799;
        end
      end else begin
        uop_10_ctrl_replayInst <= _GEN_22799;
      end
    end else begin
      uop_10_ctrl_replayInst <= _GEN_22799;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_1) begin // @[LoadQueueFlag.scala 309:50]
          if (4'ha == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 310:34]
            uop_10_pdest <= io_loadIn_1_bits_uop_pdest; // @[LoadQueueFlag.scala 310:34]
          end else begin
            uop_10_pdest <= _GEN_21471;
          end
        end else begin
          uop_10_pdest <= _GEN_21471;
        end
      end else begin
        uop_10_pdest <= _GEN_21471;
      end
    end else begin
      uop_10_pdest <= _GEN_21471;
    end
    if (io_enq_req_3_valid & ~enqCancel_3) begin // @[LoadQueueFlag.scala 204:43]
      if (4'ha == io_enq_req_3_bits_lqIdx_value) begin // @[LoadQueueFlag.scala 206:18]
        uop_10_robIdx_flag <= io_enq_req_3_bits_robIdx_flag; // @[LoadQueueFlag.scala 206:18]
      end else begin
        uop_10_robIdx_flag <= _GEN_11912;
      end
    end else begin
      uop_10_robIdx_flag <= _GEN_11912;
    end
    if (io_enq_req_3_valid & ~enqCancel_3) begin // @[LoadQueueFlag.scala 204:43]
      if (4'ha == io_enq_req_3_bits_lqIdx_value) begin // @[LoadQueueFlag.scala 206:18]
        uop_10_robIdx_value <= io_enq_req_3_bits_robIdx_value; // @[LoadQueueFlag.scala 206:18]
      end else begin
        uop_10_robIdx_value <= _GEN_11928;
      end
    end else begin
      uop_10_robIdx_value <= _GEN_11928;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'hb == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_11_cf_exceptionVec_4 <= io_loadIn_1_bits_uop_cf_exceptionVec_4; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_11_cf_exceptionVec_4 <= _GEN_21600;
          end
        end else begin
          uop_11_cf_exceptionVec_4 <= _GEN_21600;
        end
      end else begin
        uop_11_cf_exceptionVec_4 <= _GEN_21600;
      end
    end else begin
      uop_11_cf_exceptionVec_4 <= _GEN_21600;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'hb == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_11_cf_exceptionVec_5 <= io_loadIn_1_bits_uop_cf_exceptionVec_5; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_11_cf_exceptionVec_5 <= _GEN_21616;
          end
        end else begin
          uop_11_cf_exceptionVec_5 <= _GEN_21616;
        end
      end else begin
        uop_11_cf_exceptionVec_5 <= _GEN_21616;
      end
    end else begin
      uop_11_cf_exceptionVec_5 <= _GEN_21616;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'hb == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_11_cf_exceptionVec_13 <= io_loadIn_1_bits_uop_cf_exceptionVec_13; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_11_cf_exceptionVec_13 <= _GEN_21744;
          end
        end else begin
          uop_11_cf_exceptionVec_13 <= _GEN_21744;
        end
      end else begin
        uop_11_cf_exceptionVec_13 <= _GEN_21744;
      end
    end else begin
      uop_11_cf_exceptionVec_13 <= _GEN_21744;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'hb == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_11_cf_trigger_backendEn_1 <= io_loadIn_1_bits_uop_cf_trigger_backendEn_1; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_11_cf_trigger_backendEn_1 <= _GEN_21872;
          end
        end else begin
          uop_11_cf_trigger_backendEn_1 <= _GEN_21872;
        end
      end else begin
        uop_11_cf_trigger_backendEn_1 <= _GEN_21872;
      end
    end else begin
      uop_11_cf_trigger_backendEn_1 <= _GEN_21872;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'hb == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_11_cf_trigger_backendHit_0 <= io_loadIn_1_bits_uop_cf_trigger_backendHit_0; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_11_cf_trigger_backendHit_0 <= _GEN_21888;
          end
        end else begin
          uop_11_cf_trigger_backendHit_0 <= _GEN_21888;
        end
      end else begin
        uop_11_cf_trigger_backendHit_0 <= _GEN_21888;
      end
    end else begin
      uop_11_cf_trigger_backendHit_0 <= _GEN_21888;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'hb == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_11_cf_trigger_backendHit_1 <= io_loadIn_1_bits_uop_cf_trigger_backendHit_1; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_11_cf_trigger_backendHit_1 <= _GEN_21904;
          end
        end else begin
          uop_11_cf_trigger_backendHit_1 <= _GEN_21904;
        end
      end else begin
        uop_11_cf_trigger_backendHit_1 <= _GEN_21904;
      end
    end else begin
      uop_11_cf_trigger_backendHit_1 <= _GEN_21904;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'hb == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_11_cf_trigger_backendHit_4 <= io_loadIn_1_bits_uop_cf_trigger_backendHit_4; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_11_cf_trigger_backendHit_4 <= _GEN_21952;
          end
        end else begin
          uop_11_cf_trigger_backendHit_4 <= _GEN_21952;
        end
      end else begin
        uop_11_cf_trigger_backendHit_4 <= _GEN_21952;
      end
    end else begin
      uop_11_cf_trigger_backendHit_4 <= _GEN_21952;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_3) begin // @[LoadQueueFlag.scala 315:50]
          if (4'hb == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 316:33]
            uop_11_ctrl_fuOpType <= io_loadIn_1_bits_uop_ctrl_fuOpType; // @[LoadQueueFlag.scala 316:33]
          end else begin
            uop_11_ctrl_fuOpType <= _GEN_22384;
          end
        end else begin
          uop_11_ctrl_fuOpType <= _GEN_22384;
        end
      end else begin
        uop_11_ctrl_fuOpType <= _GEN_22384;
      end
    end else begin
      uop_11_ctrl_fuOpType <= _GEN_22384;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_3) begin // @[LoadQueueFlag.scala 315:50]
          if (4'hb == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 316:33]
            uop_11_ctrl_rfWen <= io_loadIn_1_bits_uop_ctrl_rfWen; // @[LoadQueueFlag.scala 316:33]
          end else begin
            uop_11_ctrl_rfWen <= _GEN_22400;
          end
        end else begin
          uop_11_ctrl_rfWen <= _GEN_22400;
        end
      end else begin
        uop_11_ctrl_rfWen <= _GEN_22400;
      end
    end else begin
      uop_11_ctrl_rfWen <= _GEN_22400;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_3) begin // @[LoadQueueFlag.scala 315:50]
          if (4'hb == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 316:33]
            uop_11_ctrl_fpWen <= io_loadIn_1_bits_uop_ctrl_fpWen; // @[LoadQueueFlag.scala 316:33]
          end else begin
            uop_11_ctrl_fpWen <= _GEN_22416;
          end
        end else begin
          uop_11_ctrl_fpWen <= _GEN_22416;
        end
      end else begin
        uop_11_ctrl_fpWen <= _GEN_22416;
      end
    end else begin
      uop_11_ctrl_fpWen <= _GEN_22416;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_3) begin // @[LoadQueueFlag.scala 315:50]
          if (4'hb == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 316:33]
            uop_11_ctrl_flushPipe <= 1'h0; // @[LoadQueueFlag.scala 316:33]
          end else begin
            uop_11_ctrl_flushPipe <= _GEN_22480;
          end
        end else begin
          uop_11_ctrl_flushPipe <= _GEN_22480;
        end
      end else begin
        uop_11_ctrl_flushPipe <= _GEN_22480;
      end
    end else begin
      uop_11_ctrl_flushPipe <= _GEN_22480;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_3) begin // @[LoadQueueFlag.scala 315:50]
          if (4'hb == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 316:33]
            uop_11_ctrl_replayInst <= io_loadIn_1_bits_uop_ctrl_replayInst; // @[LoadQueueFlag.scala 316:33]
          end else begin
            uop_11_ctrl_replayInst <= _GEN_22800;
          end
        end else begin
          uop_11_ctrl_replayInst <= _GEN_22800;
        end
      end else begin
        uop_11_ctrl_replayInst <= _GEN_22800;
      end
    end else begin
      uop_11_ctrl_replayInst <= _GEN_22800;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_1) begin // @[LoadQueueFlag.scala 309:50]
          if (4'hb == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 310:34]
            uop_11_pdest <= io_loadIn_1_bits_uop_pdest; // @[LoadQueueFlag.scala 310:34]
          end else begin
            uop_11_pdest <= _GEN_21472;
          end
        end else begin
          uop_11_pdest <= _GEN_21472;
        end
      end else begin
        uop_11_pdest <= _GEN_21472;
      end
    end else begin
      uop_11_pdest <= _GEN_21472;
    end
    if (io_enq_req_3_valid & ~enqCancel_3) begin // @[LoadQueueFlag.scala 204:43]
      if (4'hb == io_enq_req_3_bits_lqIdx_value) begin // @[LoadQueueFlag.scala 206:18]
        uop_11_robIdx_flag <= io_enq_req_3_bits_robIdx_flag; // @[LoadQueueFlag.scala 206:18]
      end else begin
        uop_11_robIdx_flag <= _GEN_11913;
      end
    end else begin
      uop_11_robIdx_flag <= _GEN_11913;
    end
    if (io_enq_req_3_valid & ~enqCancel_3) begin // @[LoadQueueFlag.scala 204:43]
      if (4'hb == io_enq_req_3_bits_lqIdx_value) begin // @[LoadQueueFlag.scala 206:18]
        uop_11_robIdx_value <= io_enq_req_3_bits_robIdx_value; // @[LoadQueueFlag.scala 206:18]
      end else begin
        uop_11_robIdx_value <= _GEN_11929;
      end
    end else begin
      uop_11_robIdx_value <= _GEN_11929;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'hc == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_12_cf_exceptionVec_4 <= io_loadIn_1_bits_uop_cf_exceptionVec_4; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_12_cf_exceptionVec_4 <= _GEN_21601;
          end
        end else begin
          uop_12_cf_exceptionVec_4 <= _GEN_21601;
        end
      end else begin
        uop_12_cf_exceptionVec_4 <= _GEN_21601;
      end
    end else begin
      uop_12_cf_exceptionVec_4 <= _GEN_21601;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'hc == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_12_cf_exceptionVec_5 <= io_loadIn_1_bits_uop_cf_exceptionVec_5; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_12_cf_exceptionVec_5 <= _GEN_21617;
          end
        end else begin
          uop_12_cf_exceptionVec_5 <= _GEN_21617;
        end
      end else begin
        uop_12_cf_exceptionVec_5 <= _GEN_21617;
      end
    end else begin
      uop_12_cf_exceptionVec_5 <= _GEN_21617;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'hc == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_12_cf_exceptionVec_13 <= io_loadIn_1_bits_uop_cf_exceptionVec_13; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_12_cf_exceptionVec_13 <= _GEN_21745;
          end
        end else begin
          uop_12_cf_exceptionVec_13 <= _GEN_21745;
        end
      end else begin
        uop_12_cf_exceptionVec_13 <= _GEN_21745;
      end
    end else begin
      uop_12_cf_exceptionVec_13 <= _GEN_21745;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'hc == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_12_cf_trigger_backendEn_1 <= io_loadIn_1_bits_uop_cf_trigger_backendEn_1; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_12_cf_trigger_backendEn_1 <= _GEN_21873;
          end
        end else begin
          uop_12_cf_trigger_backendEn_1 <= _GEN_21873;
        end
      end else begin
        uop_12_cf_trigger_backendEn_1 <= _GEN_21873;
      end
    end else begin
      uop_12_cf_trigger_backendEn_1 <= _GEN_21873;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'hc == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_12_cf_trigger_backendHit_0 <= io_loadIn_1_bits_uop_cf_trigger_backendHit_0; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_12_cf_trigger_backendHit_0 <= _GEN_21889;
          end
        end else begin
          uop_12_cf_trigger_backendHit_0 <= _GEN_21889;
        end
      end else begin
        uop_12_cf_trigger_backendHit_0 <= _GEN_21889;
      end
    end else begin
      uop_12_cf_trigger_backendHit_0 <= _GEN_21889;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'hc == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_12_cf_trigger_backendHit_1 <= io_loadIn_1_bits_uop_cf_trigger_backendHit_1; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_12_cf_trigger_backendHit_1 <= _GEN_21905;
          end
        end else begin
          uop_12_cf_trigger_backendHit_1 <= _GEN_21905;
        end
      end else begin
        uop_12_cf_trigger_backendHit_1 <= _GEN_21905;
      end
    end else begin
      uop_12_cf_trigger_backendHit_1 <= _GEN_21905;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'hc == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_12_cf_trigger_backendHit_4 <= io_loadIn_1_bits_uop_cf_trigger_backendHit_4; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_12_cf_trigger_backendHit_4 <= _GEN_21953;
          end
        end else begin
          uop_12_cf_trigger_backendHit_4 <= _GEN_21953;
        end
      end else begin
        uop_12_cf_trigger_backendHit_4 <= _GEN_21953;
      end
    end else begin
      uop_12_cf_trigger_backendHit_4 <= _GEN_21953;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_3) begin // @[LoadQueueFlag.scala 315:50]
          if (4'hc == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 316:33]
            uop_12_ctrl_fuOpType <= io_loadIn_1_bits_uop_ctrl_fuOpType; // @[LoadQueueFlag.scala 316:33]
          end else begin
            uop_12_ctrl_fuOpType <= _GEN_22385;
          end
        end else begin
          uop_12_ctrl_fuOpType <= _GEN_22385;
        end
      end else begin
        uop_12_ctrl_fuOpType <= _GEN_22385;
      end
    end else begin
      uop_12_ctrl_fuOpType <= _GEN_22385;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_3) begin // @[LoadQueueFlag.scala 315:50]
          if (4'hc == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 316:33]
            uop_12_ctrl_rfWen <= io_loadIn_1_bits_uop_ctrl_rfWen; // @[LoadQueueFlag.scala 316:33]
          end else begin
            uop_12_ctrl_rfWen <= _GEN_22401;
          end
        end else begin
          uop_12_ctrl_rfWen <= _GEN_22401;
        end
      end else begin
        uop_12_ctrl_rfWen <= _GEN_22401;
      end
    end else begin
      uop_12_ctrl_rfWen <= _GEN_22401;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_3) begin // @[LoadQueueFlag.scala 315:50]
          if (4'hc == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 316:33]
            uop_12_ctrl_fpWen <= io_loadIn_1_bits_uop_ctrl_fpWen; // @[LoadQueueFlag.scala 316:33]
          end else begin
            uop_12_ctrl_fpWen <= _GEN_22417;
          end
        end else begin
          uop_12_ctrl_fpWen <= _GEN_22417;
        end
      end else begin
        uop_12_ctrl_fpWen <= _GEN_22417;
      end
    end else begin
      uop_12_ctrl_fpWen <= _GEN_22417;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_3) begin // @[LoadQueueFlag.scala 315:50]
          if (4'hc == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 316:33]
            uop_12_ctrl_flushPipe <= 1'h0; // @[LoadQueueFlag.scala 316:33]
          end else begin
            uop_12_ctrl_flushPipe <= _GEN_22481;
          end
        end else begin
          uop_12_ctrl_flushPipe <= _GEN_22481;
        end
      end else begin
        uop_12_ctrl_flushPipe <= _GEN_22481;
      end
    end else begin
      uop_12_ctrl_flushPipe <= _GEN_22481;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_3) begin // @[LoadQueueFlag.scala 315:50]
          if (4'hc == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 316:33]
            uop_12_ctrl_replayInst <= io_loadIn_1_bits_uop_ctrl_replayInst; // @[LoadQueueFlag.scala 316:33]
          end else begin
            uop_12_ctrl_replayInst <= _GEN_22801;
          end
        end else begin
          uop_12_ctrl_replayInst <= _GEN_22801;
        end
      end else begin
        uop_12_ctrl_replayInst <= _GEN_22801;
      end
    end else begin
      uop_12_ctrl_replayInst <= _GEN_22801;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_1) begin // @[LoadQueueFlag.scala 309:50]
          if (4'hc == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 310:34]
            uop_12_pdest <= io_loadIn_1_bits_uop_pdest; // @[LoadQueueFlag.scala 310:34]
          end else begin
            uop_12_pdest <= _GEN_21473;
          end
        end else begin
          uop_12_pdest <= _GEN_21473;
        end
      end else begin
        uop_12_pdest <= _GEN_21473;
      end
    end else begin
      uop_12_pdest <= _GEN_21473;
    end
    if (io_enq_req_3_valid & ~enqCancel_3) begin // @[LoadQueueFlag.scala 204:43]
      if (4'hc == io_enq_req_3_bits_lqIdx_value) begin // @[LoadQueueFlag.scala 206:18]
        uop_12_robIdx_flag <= io_enq_req_3_bits_robIdx_flag; // @[LoadQueueFlag.scala 206:18]
      end else begin
        uop_12_robIdx_flag <= _GEN_11914;
      end
    end else begin
      uop_12_robIdx_flag <= _GEN_11914;
    end
    if (io_enq_req_3_valid & ~enqCancel_3) begin // @[LoadQueueFlag.scala 204:43]
      if (4'hc == io_enq_req_3_bits_lqIdx_value) begin // @[LoadQueueFlag.scala 206:18]
        uop_12_robIdx_value <= io_enq_req_3_bits_robIdx_value; // @[LoadQueueFlag.scala 206:18]
      end else begin
        uop_12_robIdx_value <= _GEN_11930;
      end
    end else begin
      uop_12_robIdx_value <= _GEN_11930;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'hd == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_13_cf_exceptionVec_4 <= io_loadIn_1_bits_uop_cf_exceptionVec_4; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_13_cf_exceptionVec_4 <= _GEN_21602;
          end
        end else begin
          uop_13_cf_exceptionVec_4 <= _GEN_21602;
        end
      end else begin
        uop_13_cf_exceptionVec_4 <= _GEN_21602;
      end
    end else begin
      uop_13_cf_exceptionVec_4 <= _GEN_21602;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'hd == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_13_cf_exceptionVec_5 <= io_loadIn_1_bits_uop_cf_exceptionVec_5; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_13_cf_exceptionVec_5 <= _GEN_21618;
          end
        end else begin
          uop_13_cf_exceptionVec_5 <= _GEN_21618;
        end
      end else begin
        uop_13_cf_exceptionVec_5 <= _GEN_21618;
      end
    end else begin
      uop_13_cf_exceptionVec_5 <= _GEN_21618;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'hd == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_13_cf_exceptionVec_13 <= io_loadIn_1_bits_uop_cf_exceptionVec_13; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_13_cf_exceptionVec_13 <= _GEN_21746;
          end
        end else begin
          uop_13_cf_exceptionVec_13 <= _GEN_21746;
        end
      end else begin
        uop_13_cf_exceptionVec_13 <= _GEN_21746;
      end
    end else begin
      uop_13_cf_exceptionVec_13 <= _GEN_21746;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'hd == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_13_cf_trigger_backendEn_1 <= io_loadIn_1_bits_uop_cf_trigger_backendEn_1; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_13_cf_trigger_backendEn_1 <= _GEN_21874;
          end
        end else begin
          uop_13_cf_trigger_backendEn_1 <= _GEN_21874;
        end
      end else begin
        uop_13_cf_trigger_backendEn_1 <= _GEN_21874;
      end
    end else begin
      uop_13_cf_trigger_backendEn_1 <= _GEN_21874;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'hd == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_13_cf_trigger_backendHit_0 <= io_loadIn_1_bits_uop_cf_trigger_backendHit_0; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_13_cf_trigger_backendHit_0 <= _GEN_21890;
          end
        end else begin
          uop_13_cf_trigger_backendHit_0 <= _GEN_21890;
        end
      end else begin
        uop_13_cf_trigger_backendHit_0 <= _GEN_21890;
      end
    end else begin
      uop_13_cf_trigger_backendHit_0 <= _GEN_21890;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'hd == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_13_cf_trigger_backendHit_1 <= io_loadIn_1_bits_uop_cf_trigger_backendHit_1; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_13_cf_trigger_backendHit_1 <= _GEN_21906;
          end
        end else begin
          uop_13_cf_trigger_backendHit_1 <= _GEN_21906;
        end
      end else begin
        uop_13_cf_trigger_backendHit_1 <= _GEN_21906;
      end
    end else begin
      uop_13_cf_trigger_backendHit_1 <= _GEN_21906;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'hd == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_13_cf_trigger_backendHit_4 <= io_loadIn_1_bits_uop_cf_trigger_backendHit_4; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_13_cf_trigger_backendHit_4 <= _GEN_21954;
          end
        end else begin
          uop_13_cf_trigger_backendHit_4 <= _GEN_21954;
        end
      end else begin
        uop_13_cf_trigger_backendHit_4 <= _GEN_21954;
      end
    end else begin
      uop_13_cf_trigger_backendHit_4 <= _GEN_21954;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_3) begin // @[LoadQueueFlag.scala 315:50]
          if (4'hd == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 316:33]
            uop_13_ctrl_fuOpType <= io_loadIn_1_bits_uop_ctrl_fuOpType; // @[LoadQueueFlag.scala 316:33]
          end else begin
            uop_13_ctrl_fuOpType <= _GEN_22386;
          end
        end else begin
          uop_13_ctrl_fuOpType <= _GEN_22386;
        end
      end else begin
        uop_13_ctrl_fuOpType <= _GEN_22386;
      end
    end else begin
      uop_13_ctrl_fuOpType <= _GEN_22386;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_3) begin // @[LoadQueueFlag.scala 315:50]
          if (4'hd == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 316:33]
            uop_13_ctrl_rfWen <= io_loadIn_1_bits_uop_ctrl_rfWen; // @[LoadQueueFlag.scala 316:33]
          end else begin
            uop_13_ctrl_rfWen <= _GEN_22402;
          end
        end else begin
          uop_13_ctrl_rfWen <= _GEN_22402;
        end
      end else begin
        uop_13_ctrl_rfWen <= _GEN_22402;
      end
    end else begin
      uop_13_ctrl_rfWen <= _GEN_22402;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_3) begin // @[LoadQueueFlag.scala 315:50]
          if (4'hd == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 316:33]
            uop_13_ctrl_fpWen <= io_loadIn_1_bits_uop_ctrl_fpWen; // @[LoadQueueFlag.scala 316:33]
          end else begin
            uop_13_ctrl_fpWen <= _GEN_22418;
          end
        end else begin
          uop_13_ctrl_fpWen <= _GEN_22418;
        end
      end else begin
        uop_13_ctrl_fpWen <= _GEN_22418;
      end
    end else begin
      uop_13_ctrl_fpWen <= _GEN_22418;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_3) begin // @[LoadQueueFlag.scala 315:50]
          if (4'hd == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 316:33]
            uop_13_ctrl_flushPipe <= 1'h0; // @[LoadQueueFlag.scala 316:33]
          end else begin
            uop_13_ctrl_flushPipe <= _GEN_22482;
          end
        end else begin
          uop_13_ctrl_flushPipe <= _GEN_22482;
        end
      end else begin
        uop_13_ctrl_flushPipe <= _GEN_22482;
      end
    end else begin
      uop_13_ctrl_flushPipe <= _GEN_22482;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_3) begin // @[LoadQueueFlag.scala 315:50]
          if (4'hd == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 316:33]
            uop_13_ctrl_replayInst <= io_loadIn_1_bits_uop_ctrl_replayInst; // @[LoadQueueFlag.scala 316:33]
          end else begin
            uop_13_ctrl_replayInst <= _GEN_22802;
          end
        end else begin
          uop_13_ctrl_replayInst <= _GEN_22802;
        end
      end else begin
        uop_13_ctrl_replayInst <= _GEN_22802;
      end
    end else begin
      uop_13_ctrl_replayInst <= _GEN_22802;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_1) begin // @[LoadQueueFlag.scala 309:50]
          if (4'hd == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 310:34]
            uop_13_pdest <= io_loadIn_1_bits_uop_pdest; // @[LoadQueueFlag.scala 310:34]
          end else begin
            uop_13_pdest <= _GEN_21474;
          end
        end else begin
          uop_13_pdest <= _GEN_21474;
        end
      end else begin
        uop_13_pdest <= _GEN_21474;
      end
    end else begin
      uop_13_pdest <= _GEN_21474;
    end
    if (io_enq_req_3_valid & ~enqCancel_3) begin // @[LoadQueueFlag.scala 204:43]
      if (4'hd == io_enq_req_3_bits_lqIdx_value) begin // @[LoadQueueFlag.scala 206:18]
        uop_13_robIdx_flag <= io_enq_req_3_bits_robIdx_flag; // @[LoadQueueFlag.scala 206:18]
      end else begin
        uop_13_robIdx_flag <= _GEN_11915;
      end
    end else begin
      uop_13_robIdx_flag <= _GEN_11915;
    end
    if (io_enq_req_3_valid & ~enqCancel_3) begin // @[LoadQueueFlag.scala 204:43]
      if (4'hd == io_enq_req_3_bits_lqIdx_value) begin // @[LoadQueueFlag.scala 206:18]
        uop_13_robIdx_value <= io_enq_req_3_bits_robIdx_value; // @[LoadQueueFlag.scala 206:18]
      end else begin
        uop_13_robIdx_value <= _GEN_11931;
      end
    end else begin
      uop_13_robIdx_value <= _GEN_11931;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'he == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_14_cf_exceptionVec_4 <= io_loadIn_1_bits_uop_cf_exceptionVec_4; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_14_cf_exceptionVec_4 <= _GEN_21603;
          end
        end else begin
          uop_14_cf_exceptionVec_4 <= _GEN_21603;
        end
      end else begin
        uop_14_cf_exceptionVec_4 <= _GEN_21603;
      end
    end else begin
      uop_14_cf_exceptionVec_4 <= _GEN_21603;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'he == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_14_cf_exceptionVec_5 <= io_loadIn_1_bits_uop_cf_exceptionVec_5; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_14_cf_exceptionVec_5 <= _GEN_21619;
          end
        end else begin
          uop_14_cf_exceptionVec_5 <= _GEN_21619;
        end
      end else begin
        uop_14_cf_exceptionVec_5 <= _GEN_21619;
      end
    end else begin
      uop_14_cf_exceptionVec_5 <= _GEN_21619;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'he == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_14_cf_exceptionVec_13 <= io_loadIn_1_bits_uop_cf_exceptionVec_13; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_14_cf_exceptionVec_13 <= _GEN_21747;
          end
        end else begin
          uop_14_cf_exceptionVec_13 <= _GEN_21747;
        end
      end else begin
        uop_14_cf_exceptionVec_13 <= _GEN_21747;
      end
    end else begin
      uop_14_cf_exceptionVec_13 <= _GEN_21747;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'he == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_14_cf_trigger_backendEn_1 <= io_loadIn_1_bits_uop_cf_trigger_backendEn_1; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_14_cf_trigger_backendEn_1 <= _GEN_21875;
          end
        end else begin
          uop_14_cf_trigger_backendEn_1 <= _GEN_21875;
        end
      end else begin
        uop_14_cf_trigger_backendEn_1 <= _GEN_21875;
      end
    end else begin
      uop_14_cf_trigger_backendEn_1 <= _GEN_21875;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'he == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_14_cf_trigger_backendHit_0 <= io_loadIn_1_bits_uop_cf_trigger_backendHit_0; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_14_cf_trigger_backendHit_0 <= _GEN_21891;
          end
        end else begin
          uop_14_cf_trigger_backendHit_0 <= _GEN_21891;
        end
      end else begin
        uop_14_cf_trigger_backendHit_0 <= _GEN_21891;
      end
    end else begin
      uop_14_cf_trigger_backendHit_0 <= _GEN_21891;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'he == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_14_cf_trigger_backendHit_1 <= io_loadIn_1_bits_uop_cf_trigger_backendHit_1; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_14_cf_trigger_backendHit_1 <= _GEN_21907;
          end
        end else begin
          uop_14_cf_trigger_backendHit_1 <= _GEN_21907;
        end
      end else begin
        uop_14_cf_trigger_backendHit_1 <= _GEN_21907;
      end
    end else begin
      uop_14_cf_trigger_backendHit_1 <= _GEN_21907;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'he == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_14_cf_trigger_backendHit_4 <= io_loadIn_1_bits_uop_cf_trigger_backendHit_4; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_14_cf_trigger_backendHit_4 <= _GEN_21955;
          end
        end else begin
          uop_14_cf_trigger_backendHit_4 <= _GEN_21955;
        end
      end else begin
        uop_14_cf_trigger_backendHit_4 <= _GEN_21955;
      end
    end else begin
      uop_14_cf_trigger_backendHit_4 <= _GEN_21955;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_3) begin // @[LoadQueueFlag.scala 315:50]
          if (4'he == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 316:33]
            uop_14_ctrl_fuOpType <= io_loadIn_1_bits_uop_ctrl_fuOpType; // @[LoadQueueFlag.scala 316:33]
          end else begin
            uop_14_ctrl_fuOpType <= _GEN_22387;
          end
        end else begin
          uop_14_ctrl_fuOpType <= _GEN_22387;
        end
      end else begin
        uop_14_ctrl_fuOpType <= _GEN_22387;
      end
    end else begin
      uop_14_ctrl_fuOpType <= _GEN_22387;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_3) begin // @[LoadQueueFlag.scala 315:50]
          if (4'he == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 316:33]
            uop_14_ctrl_rfWen <= io_loadIn_1_bits_uop_ctrl_rfWen; // @[LoadQueueFlag.scala 316:33]
          end else begin
            uop_14_ctrl_rfWen <= _GEN_22403;
          end
        end else begin
          uop_14_ctrl_rfWen <= _GEN_22403;
        end
      end else begin
        uop_14_ctrl_rfWen <= _GEN_22403;
      end
    end else begin
      uop_14_ctrl_rfWen <= _GEN_22403;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_3) begin // @[LoadQueueFlag.scala 315:50]
          if (4'he == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 316:33]
            uop_14_ctrl_fpWen <= io_loadIn_1_bits_uop_ctrl_fpWen; // @[LoadQueueFlag.scala 316:33]
          end else begin
            uop_14_ctrl_fpWen <= _GEN_22419;
          end
        end else begin
          uop_14_ctrl_fpWen <= _GEN_22419;
        end
      end else begin
        uop_14_ctrl_fpWen <= _GEN_22419;
      end
    end else begin
      uop_14_ctrl_fpWen <= _GEN_22419;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_3) begin // @[LoadQueueFlag.scala 315:50]
          if (4'he == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 316:33]
            uop_14_ctrl_flushPipe <= 1'h0; // @[LoadQueueFlag.scala 316:33]
          end else begin
            uop_14_ctrl_flushPipe <= _GEN_22483;
          end
        end else begin
          uop_14_ctrl_flushPipe <= _GEN_22483;
        end
      end else begin
        uop_14_ctrl_flushPipe <= _GEN_22483;
      end
    end else begin
      uop_14_ctrl_flushPipe <= _GEN_22483;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_3) begin // @[LoadQueueFlag.scala 315:50]
          if (4'he == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 316:33]
            uop_14_ctrl_replayInst <= io_loadIn_1_bits_uop_ctrl_replayInst; // @[LoadQueueFlag.scala 316:33]
          end else begin
            uop_14_ctrl_replayInst <= _GEN_22803;
          end
        end else begin
          uop_14_ctrl_replayInst <= _GEN_22803;
        end
      end else begin
        uop_14_ctrl_replayInst <= _GEN_22803;
      end
    end else begin
      uop_14_ctrl_replayInst <= _GEN_22803;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_1) begin // @[LoadQueueFlag.scala 309:50]
          if (4'he == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 310:34]
            uop_14_pdest <= io_loadIn_1_bits_uop_pdest; // @[LoadQueueFlag.scala 310:34]
          end else begin
            uop_14_pdest <= _GEN_21475;
          end
        end else begin
          uop_14_pdest <= _GEN_21475;
        end
      end else begin
        uop_14_pdest <= _GEN_21475;
      end
    end else begin
      uop_14_pdest <= _GEN_21475;
    end
    if (io_enq_req_3_valid & ~enqCancel_3) begin // @[LoadQueueFlag.scala 204:43]
      if (4'he == io_enq_req_3_bits_lqIdx_value) begin // @[LoadQueueFlag.scala 206:18]
        uop_14_robIdx_flag <= io_enq_req_3_bits_robIdx_flag; // @[LoadQueueFlag.scala 206:18]
      end else begin
        uop_14_robIdx_flag <= _GEN_11916;
      end
    end else begin
      uop_14_robIdx_flag <= _GEN_11916;
    end
    if (io_enq_req_3_valid & ~enqCancel_3) begin // @[LoadQueueFlag.scala 204:43]
      if (4'he == io_enq_req_3_bits_lqIdx_value) begin // @[LoadQueueFlag.scala 206:18]
        uop_14_robIdx_value <= io_enq_req_3_bits_robIdx_value; // @[LoadQueueFlag.scala 206:18]
      end else begin
        uop_14_robIdx_value <= _GEN_11932;
      end
    end else begin
      uop_14_robIdx_value <= _GEN_11932;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'hf == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_15_cf_exceptionVec_4 <= io_loadIn_1_bits_uop_cf_exceptionVec_4; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_15_cf_exceptionVec_4 <= _GEN_21604;
          end
        end else begin
          uop_15_cf_exceptionVec_4 <= _GEN_21604;
        end
      end else begin
        uop_15_cf_exceptionVec_4 <= _GEN_21604;
      end
    end else begin
      uop_15_cf_exceptionVec_4 <= _GEN_21604;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'hf == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_15_cf_exceptionVec_5 <= io_loadIn_1_bits_uop_cf_exceptionVec_5; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_15_cf_exceptionVec_5 <= _GEN_21620;
          end
        end else begin
          uop_15_cf_exceptionVec_5 <= _GEN_21620;
        end
      end else begin
        uop_15_cf_exceptionVec_5 <= _GEN_21620;
      end
    end else begin
      uop_15_cf_exceptionVec_5 <= _GEN_21620;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'hf == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_15_cf_exceptionVec_13 <= io_loadIn_1_bits_uop_cf_exceptionVec_13; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_15_cf_exceptionVec_13 <= _GEN_21748;
          end
        end else begin
          uop_15_cf_exceptionVec_13 <= _GEN_21748;
        end
      end else begin
        uop_15_cf_exceptionVec_13 <= _GEN_21748;
      end
    end else begin
      uop_15_cf_exceptionVec_13 <= _GEN_21748;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'hf == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_15_cf_trigger_backendEn_1 <= io_loadIn_1_bits_uop_cf_trigger_backendEn_1; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_15_cf_trigger_backendEn_1 <= _GEN_21876;
          end
        end else begin
          uop_15_cf_trigger_backendEn_1 <= _GEN_21876;
        end
      end else begin
        uop_15_cf_trigger_backendEn_1 <= _GEN_21876;
      end
    end else begin
      uop_15_cf_trigger_backendEn_1 <= _GEN_21876;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'hf == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_15_cf_trigger_backendHit_0 <= io_loadIn_1_bits_uop_cf_trigger_backendHit_0; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_15_cf_trigger_backendHit_0 <= _GEN_21892;
          end
        end else begin
          uop_15_cf_trigger_backendHit_0 <= _GEN_21892;
        end
      end else begin
        uop_15_cf_trigger_backendHit_0 <= _GEN_21892;
      end
    end else begin
      uop_15_cf_trigger_backendHit_0 <= _GEN_21892;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'hf == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_15_cf_trigger_backendHit_1 <= io_loadIn_1_bits_uop_cf_trigger_backendHit_1; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_15_cf_trigger_backendHit_1 <= _GEN_21908;
          end
        end else begin
          uop_15_cf_trigger_backendHit_1 <= _GEN_21908;
        end
      end else begin
        uop_15_cf_trigger_backendHit_1 <= _GEN_21908;
      end
    end else begin
      uop_15_cf_trigger_backendHit_1 <= _GEN_21908;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_2) begin // @[LoadQueueFlag.scala 312:50]
          if (4'hf == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 313:31]
            uop_15_cf_trigger_backendHit_4 <= io_loadIn_1_bits_uop_cf_trigger_backendHit_4; // @[LoadQueueFlag.scala 313:31]
          end else begin
            uop_15_cf_trigger_backendHit_4 <= _GEN_21956;
          end
        end else begin
          uop_15_cf_trigger_backendHit_4 <= _GEN_21956;
        end
      end else begin
        uop_15_cf_trigger_backendHit_4 <= _GEN_21956;
      end
    end else begin
      uop_15_cf_trigger_backendHit_4 <= _GEN_21956;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_3) begin // @[LoadQueueFlag.scala 315:50]
          if (4'hf == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 316:33]
            uop_15_ctrl_fuOpType <= io_loadIn_1_bits_uop_ctrl_fuOpType; // @[LoadQueueFlag.scala 316:33]
          end else begin
            uop_15_ctrl_fuOpType <= _GEN_22388;
          end
        end else begin
          uop_15_ctrl_fuOpType <= _GEN_22388;
        end
      end else begin
        uop_15_ctrl_fuOpType <= _GEN_22388;
      end
    end else begin
      uop_15_ctrl_fuOpType <= _GEN_22388;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_3) begin // @[LoadQueueFlag.scala 315:50]
          if (4'hf == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 316:33]
            uop_15_ctrl_rfWen <= io_loadIn_1_bits_uop_ctrl_rfWen; // @[LoadQueueFlag.scala 316:33]
          end else begin
            uop_15_ctrl_rfWen <= _GEN_22404;
          end
        end else begin
          uop_15_ctrl_rfWen <= _GEN_22404;
        end
      end else begin
        uop_15_ctrl_rfWen <= _GEN_22404;
      end
    end else begin
      uop_15_ctrl_rfWen <= _GEN_22404;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_3) begin // @[LoadQueueFlag.scala 315:50]
          if (4'hf == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 316:33]
            uop_15_ctrl_fpWen <= io_loadIn_1_bits_uop_ctrl_fpWen; // @[LoadQueueFlag.scala 316:33]
          end else begin
            uop_15_ctrl_fpWen <= _GEN_22420;
          end
        end else begin
          uop_15_ctrl_fpWen <= _GEN_22420;
        end
      end else begin
        uop_15_ctrl_fpWen <= _GEN_22420;
      end
    end else begin
      uop_15_ctrl_fpWen <= _GEN_22420;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_3) begin // @[LoadQueueFlag.scala 315:50]
          if (4'hf == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 316:33]
            uop_15_ctrl_flushPipe <= 1'h0; // @[LoadQueueFlag.scala 316:33]
          end else begin
            uop_15_ctrl_flushPipe <= _GEN_22484;
          end
        end else begin
          uop_15_ctrl_flushPipe <= _GEN_22484;
        end
      end else begin
        uop_15_ctrl_flushPipe <= _GEN_22484;
      end
    end else begin
      uop_15_ctrl_flushPipe <= _GEN_22484;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_3) begin // @[LoadQueueFlag.scala 315:50]
          if (4'hf == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 316:33]
            uop_15_ctrl_replayInst <= io_loadIn_1_bits_uop_ctrl_replayInst; // @[LoadQueueFlag.scala 316:33]
          end else begin
            uop_15_ctrl_replayInst <= _GEN_22804;
          end
        end else begin
          uop_15_ctrl_replayInst <= _GEN_22804;
        end
      end else begin
        uop_15_ctrl_replayInst <= _GEN_22804;
      end
    end else begin
      uop_15_ctrl_replayInst <= _GEN_22804;
    end
    if (io_loadIn_1_valid) begin // @[LoadQueueFlag.scala 286:31]
      if (_issued_T_7) begin // @[LoadQueueFlag.scala 301:26]
        if (io_loadIn_1_bits_lqDataWenDup_1) begin // @[LoadQueueFlag.scala 309:50]
          if (4'hf == io_loadIn_1_bits_uop_lqIdx_value) begin // @[LoadQueueFlag.scala 310:34]
            uop_15_pdest <= io_loadIn_1_bits_uop_pdest; // @[LoadQueueFlag.scala 310:34]
          end else begin
            uop_15_pdest <= _GEN_21476;
          end
        end else begin
          uop_15_pdest <= _GEN_21476;
        end
      end else begin
        uop_15_pdest <= _GEN_21476;
      end
    end else begin
      uop_15_pdest <= _GEN_21476;
    end
    if (io_enq_req_3_valid & ~enqCancel_3) begin // @[LoadQueueFlag.scala 204:43]
      if (4'hf == io_enq_req_3_bits_lqIdx_value) begin // @[LoadQueueFlag.scala 206:18]
        uop_15_robIdx_flag <= io_enq_req_3_bits_robIdx_flag; // @[LoadQueueFlag.scala 206:18]
      end else begin
        uop_15_robIdx_flag <= _GEN_11917;
      end
    end else begin
      uop_15_robIdx_flag <= _GEN_11917;
    end
    if (io_enq_req_3_valid & ~enqCancel_3) begin // @[LoadQueueFlag.scala 204:43]
      if (4'hf == io_enq_req_3_bits_lqIdx_value) begin // @[LoadQueueFlag.scala 206:18]
        uop_15_robIdx_value <= io_enq_req_3_bits_robIdx_value; // @[LoadQueueFlag.scala 206:18]
      end else begin
        uop_15_robIdx_value <= _GEN_11933;
      end
    end else begin
      uop_15_robIdx_value <= _GEN_11933;
    end
    lastCycleRedirect_valid <= io_redirect_valid; // @[LoadQueueFlag.scala 126:34]
    lastNeedCancel_0 <= _needCancel_T_2 & allocated_0; // @[LoadQueueFlag.scala 133:42]
    lastNeedCancel_1 <= _needCancel_T_6 & allocated_1; // @[LoadQueueFlag.scala 133:42]
    lastNeedCancel_2 <= _needCancel_T_10 & allocated_2; // @[LoadQueueFlag.scala 133:42]
    lastNeedCancel_3 <= _needCancel_T_14 & allocated_3; // @[LoadQueueFlag.scala 133:42]
    lastNeedCancel_4 <= _needCancel_T_18 & allocated_4; // @[LoadQueueFlag.scala 133:42]
    lastNeedCancel_5 <= _needCancel_T_22 & allocated_5; // @[LoadQueueFlag.scala 133:42]
    lastNeedCancel_6 <= _needCancel_T_26 & allocated_6; // @[LoadQueueFlag.scala 133:42]
    lastNeedCancel_7 <= _needCancel_T_30 & allocated_7; // @[LoadQueueFlag.scala 133:42]
    lastNeedCancel_8 <= _needCancel_T_34 & allocated_8; // @[LoadQueueFlag.scala 133:42]
    lastNeedCancel_9 <= _needCancel_T_38 & allocated_9; // @[LoadQueueFlag.scala 133:42]
    lastNeedCancel_10 <= _needCancel_T_42 & allocated_10; // @[LoadQueueFlag.scala 133:42]
    lastNeedCancel_11 <= _needCancel_T_46 & allocated_11; // @[LoadQueueFlag.scala 133:42]
    lastNeedCancel_12 <= _needCancel_T_50 & allocated_12; // @[LoadQueueFlag.scala 133:42]
    lastNeedCancel_13 <= _needCancel_T_54 & allocated_13; // @[LoadQueueFlag.scala 133:42]
    lastNeedCancel_14 <= _needCancel_T_58 & allocated_14; // @[LoadQueueFlag.scala 133:42]
    lastNeedCancel_15 <= _needCancel_T_62 & allocated_15; // @[LoadQueueFlag.scala 133:42]
    lastEnqCancel_REG_0 <= io_enq_req_0_valid & enqCancel_0; // @[LoadQueueFlag.scala 137:88]
    lastEnqCancel_REG_1 <= io_enq_req_1_valid & enqCancel_1; // @[LoadQueueFlag.scala 137:88]
    lastEnqCancel_REG_2 <= io_enq_req_2_valid & enqCancel_2; // @[LoadQueueFlag.scala 137:88]
    lastEnqCancel_REG_3 <= io_enq_req_3_valid & enqCancel_3; // @[LoadQueueFlag.scala 137:88]
    lastCommitCount <= _commitCount_T_6[0] + _commitCount_T_6[1]; // @[Bitwise.scala 48:55]
    io_lqDeq_REG <= lastCommitCount; // @[LoadQueueFlag.scala 168:22]
    io_lqCancelCnt_REG <= lastCycleCancelCount + _GEN_31429; // @[LoadQueueFlag.scala 169:50]
    io_rob_isMMIO_0_REG <= io_loadIn_0_valid & io_loadIn_0_bits_mmio; // @[LoadQueueFlag.scala 358:52]
    io_rob_uop_0_REG_robIdx_value <= io_loadIn_0_bits_uop_robIdx_value; // @[LoadQueueFlag.scala 359:29]
    io_rob_isMMIO_1_REG <= io_loadIn_1_valid & io_loadIn_1_bits_mmio; // @[LoadQueueFlag.scala 358:52]
    io_rob_uop_1_REG_robIdx_value <= io_loadIn_1_bits_uop_robIdx_value; // @[LoadQueueFlag.scala 359:29]
    REG <= io_rob_pendingld & lqTailMmioPending & lqTailAllocated & ~lqTailWriteback; // @[LoadQueueFlag.scala 406:78]
    REG_1 <= io_rob_commit; // @[LoadQueueFlag.scala 421:20]
    if (_T_57) begin // @[LoadQueueFlag.scala 456:31]
      uncacheData <= io_uncache_resp_bits_data; // @[LoadQueueFlag.scala 458:17]
    end
    io_perf_0_value_REG <= uncacheState != 2'h0; // @[LoadQueueFlag.scala 526:32]
    io_perf_0_value_REG_1 <= io_perf_0_value_REG; // @[PerfCounterUtils.scala 188:27]
    io_perf_1_value_REG <= io_uncache_req_ready & io_uncache_req_valid; // @[Decoupled.scala 50:35]
    io_perf_1_value_REG_1 <= io_perf_1_value_REG; // @[PerfCounterUtils.scala 188:27]
    io_perf_2_value_REG <= io_loadOut_0_ready & io_loadOut_0_valid; // @[Decoupled.scala 50:35]
    io_perf_2_value_REG_1 <= io_perf_2_value_REG; // @[PerfCounterUtils.scala 188:27]
    io_perf_3_value_REG <= io_loadOut_0_valid & _T_68; // @[LoadQueueFlag.scala 529:52]
    io_perf_3_value_REG_1 <= io_perf_3_value_REG; // @[PerfCounterUtils.scala 188:27]
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[LoadQueueFlag.scala 250:26]
      allocated_0 <= 1'h0; // @[LoadQueueFlag.scala 251:20]
    end else if (needCancel_0) begin // @[LoadQueueFlag.scala 232:30]
      allocated_0 <= 1'h0; // @[LoadQueueFlag.scala 233:{40,40}]
    end else if (commitCount > 2'h1) begin
      if (4'h0 == deqLookupVec_new_ptr_1_value) begin
        allocated_0 <= 1'h0;
      end else begin
        allocated_0 <= _GEN_16326;
      end
    end else begin
      allocated_0 <= _GEN_16326;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[LoadQueueFlag.scala 250:26]
      allocated_1 <= 1'h0; // @[LoadQueueFlag.scala 251:20]
    end else if (needCancel_1) begin // @[LoadQueueFlag.scala 232:30]
      allocated_1 <= 1'h0; // @[LoadQueueFlag.scala 233:{40,40}]
    end else if (commitCount > 2'h1) begin
      if (4'h1 == deqLookupVec_new_ptr_1_value) begin
        allocated_1 <= 1'h0;
      end else begin
        allocated_1 <= _GEN_16327;
      end
    end else begin
      allocated_1 <= _GEN_16327;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[LoadQueueFlag.scala 250:26]
      allocated_2 <= 1'h0; // @[LoadQueueFlag.scala 251:20]
    end else if (needCancel_2) begin // @[LoadQueueFlag.scala 232:30]
      allocated_2 <= 1'h0; // @[LoadQueueFlag.scala 233:{40,40}]
    end else if (commitCount > 2'h1) begin
      if (4'h2 == deqLookupVec_new_ptr_1_value) begin
        allocated_2 <= 1'h0;
      end else begin
        allocated_2 <= _GEN_16328;
      end
    end else begin
      allocated_2 <= _GEN_16328;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[LoadQueueFlag.scala 250:26]
      allocated_3 <= 1'h0; // @[LoadQueueFlag.scala 251:20]
    end else if (needCancel_3) begin // @[LoadQueueFlag.scala 232:30]
      allocated_3 <= 1'h0; // @[LoadQueueFlag.scala 233:{40,40}]
    end else if (commitCount > 2'h1) begin
      if (4'h3 == deqLookupVec_new_ptr_1_value) begin
        allocated_3 <= 1'h0;
      end else begin
        allocated_3 <= _GEN_16329;
      end
    end else begin
      allocated_3 <= _GEN_16329;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[LoadQueueFlag.scala 250:26]
      allocated_4 <= 1'h0; // @[LoadQueueFlag.scala 251:20]
    end else if (needCancel_4) begin // @[LoadQueueFlag.scala 232:30]
      allocated_4 <= 1'h0; // @[LoadQueueFlag.scala 233:{40,40}]
    end else if (commitCount > 2'h1) begin
      if (4'h4 == deqLookupVec_new_ptr_1_value) begin
        allocated_4 <= 1'h0;
      end else begin
        allocated_4 <= _GEN_16330;
      end
    end else begin
      allocated_4 <= _GEN_16330;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[LoadQueueFlag.scala 250:26]
      allocated_5 <= 1'h0; // @[LoadQueueFlag.scala 251:20]
    end else if (needCancel_5) begin // @[LoadQueueFlag.scala 232:30]
      allocated_5 <= 1'h0; // @[LoadQueueFlag.scala 233:{40,40}]
    end else if (commitCount > 2'h1) begin
      if (4'h5 == deqLookupVec_new_ptr_1_value) begin
        allocated_5 <= 1'h0;
      end else begin
        allocated_5 <= _GEN_16331;
      end
    end else begin
      allocated_5 <= _GEN_16331;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[LoadQueueFlag.scala 250:26]
      allocated_6 <= 1'h0; // @[LoadQueueFlag.scala 251:20]
    end else if (needCancel_6) begin // @[LoadQueueFlag.scala 232:30]
      allocated_6 <= 1'h0; // @[LoadQueueFlag.scala 233:{40,40}]
    end else if (commitCount > 2'h1) begin
      if (4'h6 == deqLookupVec_new_ptr_1_value) begin
        allocated_6 <= 1'h0;
      end else begin
        allocated_6 <= _GEN_16332;
      end
    end else begin
      allocated_6 <= _GEN_16332;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[LoadQueueFlag.scala 250:26]
      allocated_7 <= 1'h0; // @[LoadQueueFlag.scala 251:20]
    end else if (needCancel_7) begin // @[LoadQueueFlag.scala 232:30]
      allocated_7 <= 1'h0; // @[LoadQueueFlag.scala 233:{40,40}]
    end else if (commitCount > 2'h1) begin
      if (4'h7 == deqLookupVec_new_ptr_1_value) begin
        allocated_7 <= 1'h0;
      end else begin
        allocated_7 <= _GEN_16333;
      end
    end else begin
      allocated_7 <= _GEN_16333;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[LoadQueueFlag.scala 250:26]
      allocated_8 <= 1'h0; // @[LoadQueueFlag.scala 251:20]
    end else if (needCancel_8) begin // @[LoadQueueFlag.scala 232:30]
      allocated_8 <= 1'h0; // @[LoadQueueFlag.scala 233:{40,40}]
    end else if (commitCount > 2'h1) begin
      if (4'h8 == deqLookupVec_new_ptr_1_value) begin
        allocated_8 <= 1'h0;
      end else begin
        allocated_8 <= _GEN_16334;
      end
    end else begin
      allocated_8 <= _GEN_16334;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[LoadQueueFlag.scala 250:26]
      allocated_9 <= 1'h0; // @[LoadQueueFlag.scala 251:20]
    end else if (needCancel_9) begin // @[LoadQueueFlag.scala 232:30]
      allocated_9 <= 1'h0; // @[LoadQueueFlag.scala 233:{40,40}]
    end else if (commitCount > 2'h1) begin
      if (4'h9 == deqLookupVec_new_ptr_1_value) begin
        allocated_9 <= 1'h0;
      end else begin
        allocated_9 <= _GEN_16335;
      end
    end else begin
      allocated_9 <= _GEN_16335;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[LoadQueueFlag.scala 250:26]
      allocated_10 <= 1'h0; // @[LoadQueueFlag.scala 251:20]
    end else if (needCancel_10) begin // @[LoadQueueFlag.scala 232:30]
      allocated_10 <= 1'h0; // @[LoadQueueFlag.scala 233:{40,40}]
    end else if (commitCount > 2'h1) begin
      if (4'ha == deqLookupVec_new_ptr_1_value) begin
        allocated_10 <= 1'h0;
      end else begin
        allocated_10 <= _GEN_16336;
      end
    end else begin
      allocated_10 <= _GEN_16336;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[LoadQueueFlag.scala 250:26]
      allocated_11 <= 1'h0; // @[LoadQueueFlag.scala 251:20]
    end else if (needCancel_11) begin // @[LoadQueueFlag.scala 232:30]
      allocated_11 <= 1'h0; // @[LoadQueueFlag.scala 233:{40,40}]
    end else if (commitCount > 2'h1) begin
      if (4'hb == deqLookupVec_new_ptr_1_value) begin
        allocated_11 <= 1'h0;
      end else begin
        allocated_11 <= _GEN_16337;
      end
    end else begin
      allocated_11 <= _GEN_16337;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[LoadQueueFlag.scala 250:26]
      allocated_12 <= 1'h0; // @[LoadQueueFlag.scala 251:20]
    end else if (needCancel_12) begin // @[LoadQueueFlag.scala 232:30]
      allocated_12 <= 1'h0; // @[LoadQueueFlag.scala 233:{40,40}]
    end else if (commitCount > 2'h1) begin
      if (4'hc == deqLookupVec_new_ptr_1_value) begin
        allocated_12 <= 1'h0;
      end else begin
        allocated_12 <= _GEN_16338;
      end
    end else begin
      allocated_12 <= _GEN_16338;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[LoadQueueFlag.scala 250:26]
      allocated_13 <= 1'h0; // @[LoadQueueFlag.scala 251:20]
    end else if (needCancel_13) begin // @[LoadQueueFlag.scala 232:30]
      allocated_13 <= 1'h0; // @[LoadQueueFlag.scala 233:{40,40}]
    end else if (commitCount > 2'h1) begin
      if (4'hd == deqLookupVec_new_ptr_1_value) begin
        allocated_13 <= 1'h0;
      end else begin
        allocated_13 <= _GEN_16339;
      end
    end else begin
      allocated_13 <= _GEN_16339;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[LoadQueueFlag.scala 250:26]
      allocated_14 <= 1'h0; // @[LoadQueueFlag.scala 251:20]
    end else if (needCancel_14) begin // @[LoadQueueFlag.scala 232:30]
      allocated_14 <= 1'h0; // @[LoadQueueFlag.scala 233:{40,40}]
    end else if (commitCount > 2'h1) begin
      if (4'he == deqLookupVec_new_ptr_1_value) begin
        allocated_14 <= 1'h0;
      end else begin
        allocated_14 <= _GEN_16340;
      end
    end else begin
      allocated_14 <= _GEN_16340;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[LoadQueueFlag.scala 250:26]
      allocated_15 <= 1'h0; // @[LoadQueueFlag.scala 251:20]
    end else if (needCancel_15) begin // @[LoadQueueFlag.scala 232:30]
      allocated_15 <= 1'h0; // @[LoadQueueFlag.scala 233:{40,40}]
    end else if (commitCount > 2'h1) begin
      if (4'hf == deqLookupVec_new_ptr_1_value) begin
        allocated_15 <= 1'h0;
      end else begin
        allocated_15 <= _GEN_16341;
      end
    end else begin
      allocated_15 <= _GEN_16341;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[LoadQueueFlag.scala 286:31]
      addrvalid_0 <= 1'h0; // @[LoadQueueFlag.scala 301:26 303:{32,32}]
    end else if (io_loadIn_1_valid) begin
      if (_issued_T_7) begin
        if (4'h0 == io_loadIn_1_bits_uop_lqIdx_value) begin
          addrvalid_0 <= _issued_T_8;
        end else begin
          addrvalid_0 <= _GEN_21397;
        end
      end else begin
        addrvalid_0 <= _GEN_21397;
      end
    end else begin
      addrvalid_0 <= _GEN_21397;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[LoadQueueFlag.scala 286:31]
      addrvalid_1 <= 1'h0; // @[LoadQueueFlag.scala 301:26 303:{32,32}]
    end else if (io_loadIn_1_valid) begin
      if (_issued_T_7) begin
        if (4'h1 == io_loadIn_1_bits_uop_lqIdx_value) begin
          addrvalid_1 <= _issued_T_8;
        end else begin
          addrvalid_1 <= _GEN_21398;
        end
      end else begin
        addrvalid_1 <= _GEN_21398;
      end
    end else begin
      addrvalid_1 <= _GEN_21398;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[LoadQueueFlag.scala 286:31]
      addrvalid_2 <= 1'h0; // @[LoadQueueFlag.scala 301:26 303:{32,32}]
    end else if (io_loadIn_1_valid) begin
      if (_issued_T_7) begin
        if (4'h2 == io_loadIn_1_bits_uop_lqIdx_value) begin
          addrvalid_2 <= _issued_T_8;
        end else begin
          addrvalid_2 <= _GEN_21399;
        end
      end else begin
        addrvalid_2 <= _GEN_21399;
      end
    end else begin
      addrvalid_2 <= _GEN_21399;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[LoadQueueFlag.scala 286:31]
      addrvalid_3 <= 1'h0; // @[LoadQueueFlag.scala 301:26 303:{32,32}]
    end else if (io_loadIn_1_valid) begin
      if (_issued_T_7) begin
        if (4'h3 == io_loadIn_1_bits_uop_lqIdx_value) begin
          addrvalid_3 <= _issued_T_8;
        end else begin
          addrvalid_3 <= _GEN_21400;
        end
      end else begin
        addrvalid_3 <= _GEN_21400;
      end
    end else begin
      addrvalid_3 <= _GEN_21400;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[LoadQueueFlag.scala 286:31]
      addrvalid_4 <= 1'h0; // @[LoadQueueFlag.scala 301:26 303:{32,32}]
    end else if (io_loadIn_1_valid) begin
      if (_issued_T_7) begin
        if (4'h4 == io_loadIn_1_bits_uop_lqIdx_value) begin
          addrvalid_4 <= _issued_T_8;
        end else begin
          addrvalid_4 <= _GEN_21401;
        end
      end else begin
        addrvalid_4 <= _GEN_21401;
      end
    end else begin
      addrvalid_4 <= _GEN_21401;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[LoadQueueFlag.scala 286:31]
      addrvalid_5 <= 1'h0; // @[LoadQueueFlag.scala 301:26 303:{32,32}]
    end else if (io_loadIn_1_valid) begin
      if (_issued_T_7) begin
        if (4'h5 == io_loadIn_1_bits_uop_lqIdx_value) begin
          addrvalid_5 <= _issued_T_8;
        end else begin
          addrvalid_5 <= _GEN_21402;
        end
      end else begin
        addrvalid_5 <= _GEN_21402;
      end
    end else begin
      addrvalid_5 <= _GEN_21402;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[LoadQueueFlag.scala 286:31]
      addrvalid_6 <= 1'h0; // @[LoadQueueFlag.scala 301:26 303:{32,32}]
    end else if (io_loadIn_1_valid) begin
      if (_issued_T_7) begin
        if (4'h6 == io_loadIn_1_bits_uop_lqIdx_value) begin
          addrvalid_6 <= _issued_T_8;
        end else begin
          addrvalid_6 <= _GEN_21403;
        end
      end else begin
        addrvalid_6 <= _GEN_21403;
      end
    end else begin
      addrvalid_6 <= _GEN_21403;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[LoadQueueFlag.scala 286:31]
      addrvalid_7 <= 1'h0; // @[LoadQueueFlag.scala 301:26 303:{32,32}]
    end else if (io_loadIn_1_valid) begin
      if (_issued_T_7) begin
        if (4'h7 == io_loadIn_1_bits_uop_lqIdx_value) begin
          addrvalid_7 <= _issued_T_8;
        end else begin
          addrvalid_7 <= _GEN_21404;
        end
      end else begin
        addrvalid_7 <= _GEN_21404;
      end
    end else begin
      addrvalid_7 <= _GEN_21404;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[LoadQueueFlag.scala 286:31]
      addrvalid_8 <= 1'h0; // @[LoadQueueFlag.scala 301:26 303:{32,32}]
    end else if (io_loadIn_1_valid) begin
      if (_issued_T_7) begin
        if (4'h8 == io_loadIn_1_bits_uop_lqIdx_value) begin
          addrvalid_8 <= _issued_T_8;
        end else begin
          addrvalid_8 <= _GEN_21405;
        end
      end else begin
        addrvalid_8 <= _GEN_21405;
      end
    end else begin
      addrvalid_8 <= _GEN_21405;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[LoadQueueFlag.scala 286:31]
      addrvalid_9 <= 1'h0; // @[LoadQueueFlag.scala 301:26 303:{32,32}]
    end else if (io_loadIn_1_valid) begin
      if (_issued_T_7) begin
        if (4'h9 == io_loadIn_1_bits_uop_lqIdx_value) begin
          addrvalid_9 <= _issued_T_8;
        end else begin
          addrvalid_9 <= _GEN_21406;
        end
      end else begin
        addrvalid_9 <= _GEN_21406;
      end
    end else begin
      addrvalid_9 <= _GEN_21406;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[LoadQueueFlag.scala 286:31]
      addrvalid_10 <= 1'h0; // @[LoadQueueFlag.scala 301:26 303:{32,32}]
    end else if (io_loadIn_1_valid) begin
      if (_issued_T_7) begin
        if (4'ha == io_loadIn_1_bits_uop_lqIdx_value) begin
          addrvalid_10 <= _issued_T_8;
        end else begin
          addrvalid_10 <= _GEN_21407;
        end
      end else begin
        addrvalid_10 <= _GEN_21407;
      end
    end else begin
      addrvalid_10 <= _GEN_21407;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[LoadQueueFlag.scala 286:31]
      addrvalid_11 <= 1'h0; // @[LoadQueueFlag.scala 301:26 303:{32,32}]
    end else if (io_loadIn_1_valid) begin
      if (_issued_T_7) begin
        if (4'hb == io_loadIn_1_bits_uop_lqIdx_value) begin
          addrvalid_11 <= _issued_T_8;
        end else begin
          addrvalid_11 <= _GEN_21408;
        end
      end else begin
        addrvalid_11 <= _GEN_21408;
      end
    end else begin
      addrvalid_11 <= _GEN_21408;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[LoadQueueFlag.scala 286:31]
      addrvalid_12 <= 1'h0; // @[LoadQueueFlag.scala 301:26 303:{32,32}]
    end else if (io_loadIn_1_valid) begin
      if (_issued_T_7) begin
        if (4'hc == io_loadIn_1_bits_uop_lqIdx_value) begin
          addrvalid_12 <= _issued_T_8;
        end else begin
          addrvalid_12 <= _GEN_21409;
        end
      end else begin
        addrvalid_12 <= _GEN_21409;
      end
    end else begin
      addrvalid_12 <= _GEN_21409;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[LoadQueueFlag.scala 286:31]
      addrvalid_13 <= 1'h0; // @[LoadQueueFlag.scala 301:26 303:{32,32}]
    end else if (io_loadIn_1_valid) begin
      if (_issued_T_7) begin
        if (4'hd == io_loadIn_1_bits_uop_lqIdx_value) begin
          addrvalid_13 <= _issued_T_8;
        end else begin
          addrvalid_13 <= _GEN_21410;
        end
      end else begin
        addrvalid_13 <= _GEN_21410;
      end
    end else begin
      addrvalid_13 <= _GEN_21410;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[LoadQueueFlag.scala 286:31]
      addrvalid_14 <= 1'h0; // @[LoadQueueFlag.scala 301:26 303:{32,32}]
    end else if (io_loadIn_1_valid) begin
      if (_issued_T_7) begin
        if (4'he == io_loadIn_1_bits_uop_lqIdx_value) begin
          addrvalid_14 <= _issued_T_8;
        end else begin
          addrvalid_14 <= _GEN_21411;
        end
      end else begin
        addrvalid_14 <= _GEN_21411;
      end
    end else begin
      addrvalid_14 <= _GEN_21411;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[LoadQueueFlag.scala 286:31]
      addrvalid_15 <= 1'h0; // @[LoadQueueFlag.scala 301:26 303:{32,32}]
    end else if (io_loadIn_1_valid) begin
      if (_issued_T_7) begin
        if (4'hf == io_loadIn_1_bits_uop_lqIdx_value) begin
          addrvalid_15 <= _issued_T_8;
        end else begin
          addrvalid_15 <= _GEN_21412;
        end
      end else begin
        addrvalid_15 <= _GEN_21412;
      end
    end else begin
      addrvalid_15 <= _GEN_21412;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[LoadQueueFlag.scala 456:31]
      datavalid_0 <= 1'h0;
    end else if (_T_57) begin // @[LoadQueueFlag.scala 286:31]
      datavalid_0 <= _GEN_29617; // @[LoadQueueFlag.scala 301:26 304:{32,32}]
    end else if (io_loadIn_1_valid) begin
      if (_issued_T_7) begin
        if (4'h0 == io_loadIn_1_bits_uop_lqIdx_value) begin
          datavalid_0 <= datavalidVal_1;
        end else begin
          datavalid_0 <= _GEN_21413;
        end
      end else begin
        datavalid_0 <= _GEN_21413;
      end
    end else begin
      datavalid_0 <= _GEN_21413;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[LoadQueueFlag.scala 456:31]
      datavalid_1 <= 1'h0;
    end else if (_T_57) begin // @[LoadQueueFlag.scala 286:31]
      datavalid_1 <= _GEN_29618; // @[LoadQueueFlag.scala 301:26 304:{32,32}]
    end else if (io_loadIn_1_valid) begin
      if (_issued_T_7) begin
        if (4'h1 == io_loadIn_1_bits_uop_lqIdx_value) begin
          datavalid_1 <= datavalidVal_1;
        end else begin
          datavalid_1 <= _GEN_21414;
        end
      end else begin
        datavalid_1 <= _GEN_21414;
      end
    end else begin
      datavalid_1 <= _GEN_21414;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[LoadQueueFlag.scala 456:31]
      datavalid_2 <= 1'h0;
    end else if (_T_57) begin // @[LoadQueueFlag.scala 286:31]
      datavalid_2 <= _GEN_29619; // @[LoadQueueFlag.scala 301:26 304:{32,32}]
    end else if (io_loadIn_1_valid) begin
      if (_issued_T_7) begin
        if (4'h2 == io_loadIn_1_bits_uop_lqIdx_value) begin
          datavalid_2 <= datavalidVal_1;
        end else begin
          datavalid_2 <= _GEN_21415;
        end
      end else begin
        datavalid_2 <= _GEN_21415;
      end
    end else begin
      datavalid_2 <= _GEN_21415;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[LoadQueueFlag.scala 456:31]
      datavalid_3 <= 1'h0;
    end else if (_T_57) begin // @[LoadQueueFlag.scala 286:31]
      datavalid_3 <= _GEN_29620; // @[LoadQueueFlag.scala 301:26 304:{32,32}]
    end else if (io_loadIn_1_valid) begin
      if (_issued_T_7) begin
        if (4'h3 == io_loadIn_1_bits_uop_lqIdx_value) begin
          datavalid_3 <= datavalidVal_1;
        end else begin
          datavalid_3 <= _GEN_21416;
        end
      end else begin
        datavalid_3 <= _GEN_21416;
      end
    end else begin
      datavalid_3 <= _GEN_21416;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[LoadQueueFlag.scala 456:31]
      datavalid_4 <= 1'h0;
    end else if (_T_57) begin // @[LoadQueueFlag.scala 286:31]
      datavalid_4 <= _GEN_29621; // @[LoadQueueFlag.scala 301:26 304:{32,32}]
    end else if (io_loadIn_1_valid) begin
      if (_issued_T_7) begin
        if (4'h4 == io_loadIn_1_bits_uop_lqIdx_value) begin
          datavalid_4 <= datavalidVal_1;
        end else begin
          datavalid_4 <= _GEN_21417;
        end
      end else begin
        datavalid_4 <= _GEN_21417;
      end
    end else begin
      datavalid_4 <= _GEN_21417;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[LoadQueueFlag.scala 456:31]
      datavalid_5 <= 1'h0;
    end else if (_T_57) begin // @[LoadQueueFlag.scala 286:31]
      datavalid_5 <= _GEN_29622; // @[LoadQueueFlag.scala 301:26 304:{32,32}]
    end else if (io_loadIn_1_valid) begin
      if (_issued_T_7) begin
        if (4'h5 == io_loadIn_1_bits_uop_lqIdx_value) begin
          datavalid_5 <= datavalidVal_1;
        end else begin
          datavalid_5 <= _GEN_21418;
        end
      end else begin
        datavalid_5 <= _GEN_21418;
      end
    end else begin
      datavalid_5 <= _GEN_21418;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[LoadQueueFlag.scala 456:31]
      datavalid_6 <= 1'h0;
    end else if (_T_57) begin // @[LoadQueueFlag.scala 286:31]
      datavalid_6 <= _GEN_29623; // @[LoadQueueFlag.scala 301:26 304:{32,32}]
    end else if (io_loadIn_1_valid) begin
      if (_issued_T_7) begin
        if (4'h6 == io_loadIn_1_bits_uop_lqIdx_value) begin
          datavalid_6 <= datavalidVal_1;
        end else begin
          datavalid_6 <= _GEN_21419;
        end
      end else begin
        datavalid_6 <= _GEN_21419;
      end
    end else begin
      datavalid_6 <= _GEN_21419;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[LoadQueueFlag.scala 456:31]
      datavalid_7 <= 1'h0;
    end else if (_T_57) begin // @[LoadQueueFlag.scala 286:31]
      datavalid_7 <= _GEN_29624; // @[LoadQueueFlag.scala 301:26 304:{32,32}]
    end else if (io_loadIn_1_valid) begin
      if (_issued_T_7) begin
        if (4'h7 == io_loadIn_1_bits_uop_lqIdx_value) begin
          datavalid_7 <= datavalidVal_1;
        end else begin
          datavalid_7 <= _GEN_21420;
        end
      end else begin
        datavalid_7 <= _GEN_21420;
      end
    end else begin
      datavalid_7 <= _GEN_21420;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[LoadQueueFlag.scala 456:31]
      datavalid_8 <= 1'h0;
    end else if (_T_57) begin // @[LoadQueueFlag.scala 286:31]
      datavalid_8 <= _GEN_29625; // @[LoadQueueFlag.scala 301:26 304:{32,32}]
    end else if (io_loadIn_1_valid) begin
      if (_issued_T_7) begin
        if (4'h8 == io_loadIn_1_bits_uop_lqIdx_value) begin
          datavalid_8 <= datavalidVal_1;
        end else begin
          datavalid_8 <= _GEN_21421;
        end
      end else begin
        datavalid_8 <= _GEN_21421;
      end
    end else begin
      datavalid_8 <= _GEN_21421;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[LoadQueueFlag.scala 456:31]
      datavalid_9 <= 1'h0;
    end else if (_T_57) begin // @[LoadQueueFlag.scala 286:31]
      datavalid_9 <= _GEN_29626; // @[LoadQueueFlag.scala 301:26 304:{32,32}]
    end else if (io_loadIn_1_valid) begin
      if (_issued_T_7) begin
        if (4'h9 == io_loadIn_1_bits_uop_lqIdx_value) begin
          datavalid_9 <= datavalidVal_1;
        end else begin
          datavalid_9 <= _GEN_21422;
        end
      end else begin
        datavalid_9 <= _GEN_21422;
      end
    end else begin
      datavalid_9 <= _GEN_21422;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[LoadQueueFlag.scala 456:31]
      datavalid_10 <= 1'h0;
    end else if (_T_57) begin // @[LoadQueueFlag.scala 286:31]
      datavalid_10 <= _GEN_29627; // @[LoadQueueFlag.scala 301:26 304:{32,32}]
    end else if (io_loadIn_1_valid) begin
      if (_issued_T_7) begin
        if (4'ha == io_loadIn_1_bits_uop_lqIdx_value) begin
          datavalid_10 <= datavalidVal_1;
        end else begin
          datavalid_10 <= _GEN_21423;
        end
      end else begin
        datavalid_10 <= _GEN_21423;
      end
    end else begin
      datavalid_10 <= _GEN_21423;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[LoadQueueFlag.scala 456:31]
      datavalid_11 <= 1'h0;
    end else if (_T_57) begin // @[LoadQueueFlag.scala 286:31]
      datavalid_11 <= _GEN_29628; // @[LoadQueueFlag.scala 301:26 304:{32,32}]
    end else if (io_loadIn_1_valid) begin
      if (_issued_T_7) begin
        if (4'hb == io_loadIn_1_bits_uop_lqIdx_value) begin
          datavalid_11 <= datavalidVal_1;
        end else begin
          datavalid_11 <= _GEN_21424;
        end
      end else begin
        datavalid_11 <= _GEN_21424;
      end
    end else begin
      datavalid_11 <= _GEN_21424;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[LoadQueueFlag.scala 456:31]
      datavalid_12 <= 1'h0;
    end else if (_T_57) begin // @[LoadQueueFlag.scala 286:31]
      datavalid_12 <= _GEN_29629; // @[LoadQueueFlag.scala 301:26 304:{32,32}]
    end else if (io_loadIn_1_valid) begin
      if (_issued_T_7) begin
        if (4'hc == io_loadIn_1_bits_uop_lqIdx_value) begin
          datavalid_12 <= datavalidVal_1;
        end else begin
          datavalid_12 <= _GEN_21425;
        end
      end else begin
        datavalid_12 <= _GEN_21425;
      end
    end else begin
      datavalid_12 <= _GEN_21425;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[LoadQueueFlag.scala 456:31]
      datavalid_13 <= 1'h0;
    end else if (_T_57) begin // @[LoadQueueFlag.scala 286:31]
      datavalid_13 <= _GEN_29630; // @[LoadQueueFlag.scala 301:26 304:{32,32}]
    end else if (io_loadIn_1_valid) begin
      if (_issued_T_7) begin
        if (4'hd == io_loadIn_1_bits_uop_lqIdx_value) begin
          datavalid_13 <= datavalidVal_1;
        end else begin
          datavalid_13 <= _GEN_21426;
        end
      end else begin
        datavalid_13 <= _GEN_21426;
      end
    end else begin
      datavalid_13 <= _GEN_21426;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[LoadQueueFlag.scala 456:31]
      datavalid_14 <= 1'h0;
    end else if (_T_57) begin // @[LoadQueueFlag.scala 286:31]
      datavalid_14 <= _GEN_29631; // @[LoadQueueFlag.scala 301:26 304:{32,32}]
    end else if (io_loadIn_1_valid) begin
      if (_issued_T_7) begin
        if (4'he == io_loadIn_1_bits_uop_lqIdx_value) begin
          datavalid_14 <= datavalidVal_1;
        end else begin
          datavalid_14 <= _GEN_21427;
        end
      end else begin
        datavalid_14 <= _GEN_21427;
      end
    end else begin
      datavalid_14 <= _GEN_21427;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[LoadQueueFlag.scala 456:31]
      datavalid_15 <= 1'h0;
    end else if (_T_57) begin // @[LoadQueueFlag.scala 286:31]
      datavalid_15 <= _GEN_29632; // @[LoadQueueFlag.scala 301:26 304:{32,32}]
    end else if (io_loadIn_1_valid) begin
      if (_issued_T_7) begin
        if (4'hf == io_loadIn_1_bits_uop_lqIdx_value) begin
          datavalid_15 <= datavalidVal_1;
        end else begin
          datavalid_15 <= _GEN_21428;
        end
      end else begin
        datavalid_15 <= _GEN_21428;
      end
    end else begin
      datavalid_15 <= _GEN_21428;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[LoadQueueFlag.scala 443:30]
      pending_0 <= 1'h0; // @[LoadQueueFlag.scala 444:{21,21}]
    end else if (_T_55) begin
      if (4'h0 == deqPtrExt_rvalue) begin
        pending_0 <= 1'h0;
      end else begin
        pending_0 <= _GEN_27950;
      end
    end else begin
      pending_0 <= _GEN_27950;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[LoadQueueFlag.scala 443:30]
      pending_1 <= 1'h0; // @[LoadQueueFlag.scala 444:{21,21}]
    end else if (_T_55) begin
      if (4'h1 == deqPtrExt_rvalue) begin
        pending_1 <= 1'h0;
      end else begin
        pending_1 <= _GEN_27951;
      end
    end else begin
      pending_1 <= _GEN_27951;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[LoadQueueFlag.scala 443:30]
      pending_2 <= 1'h0; // @[LoadQueueFlag.scala 444:{21,21}]
    end else if (_T_55) begin
      if (4'h2 == deqPtrExt_rvalue) begin
        pending_2 <= 1'h0;
      end else begin
        pending_2 <= _GEN_27952;
      end
    end else begin
      pending_2 <= _GEN_27952;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[LoadQueueFlag.scala 443:30]
      pending_3 <= 1'h0; // @[LoadQueueFlag.scala 444:{21,21}]
    end else if (_T_55) begin
      if (4'h3 == deqPtrExt_rvalue) begin
        pending_3 <= 1'h0;
      end else begin
        pending_3 <= _GEN_27953;
      end
    end else begin
      pending_3 <= _GEN_27953;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[LoadQueueFlag.scala 443:30]
      pending_4 <= 1'h0; // @[LoadQueueFlag.scala 444:{21,21}]
    end else if (_T_55) begin
      if (4'h4 == deqPtrExt_rvalue) begin
        pending_4 <= 1'h0;
      end else begin
        pending_4 <= _GEN_27954;
      end
    end else begin
      pending_4 <= _GEN_27954;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[LoadQueueFlag.scala 443:30]
      pending_5 <= 1'h0; // @[LoadQueueFlag.scala 444:{21,21}]
    end else if (_T_55) begin
      if (4'h5 == deqPtrExt_rvalue) begin
        pending_5 <= 1'h0;
      end else begin
        pending_5 <= _GEN_27955;
      end
    end else begin
      pending_5 <= _GEN_27955;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[LoadQueueFlag.scala 443:30]
      pending_6 <= 1'h0; // @[LoadQueueFlag.scala 444:{21,21}]
    end else if (_T_55) begin
      if (4'h6 == deqPtrExt_rvalue) begin
        pending_6 <= 1'h0;
      end else begin
        pending_6 <= _GEN_27956;
      end
    end else begin
      pending_6 <= _GEN_27956;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[LoadQueueFlag.scala 443:30]
      pending_7 <= 1'h0; // @[LoadQueueFlag.scala 444:{21,21}]
    end else if (_T_55) begin
      if (4'h7 == deqPtrExt_rvalue) begin
        pending_7 <= 1'h0;
      end else begin
        pending_7 <= _GEN_27957;
      end
    end else begin
      pending_7 <= _GEN_27957;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[LoadQueueFlag.scala 443:30]
      pending_8 <= 1'h0; // @[LoadQueueFlag.scala 444:{21,21}]
    end else if (_T_55) begin
      if (4'h8 == deqPtrExt_rvalue) begin
        pending_8 <= 1'h0;
      end else begin
        pending_8 <= _GEN_27958;
      end
    end else begin
      pending_8 <= _GEN_27958;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[LoadQueueFlag.scala 443:30]
      pending_9 <= 1'h0; // @[LoadQueueFlag.scala 444:{21,21}]
    end else if (_T_55) begin
      if (4'h9 == deqPtrExt_rvalue) begin
        pending_9 <= 1'h0;
      end else begin
        pending_9 <= _GEN_27959;
      end
    end else begin
      pending_9 <= _GEN_27959;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[LoadQueueFlag.scala 443:30]
      pending_10 <= 1'h0; // @[LoadQueueFlag.scala 444:{21,21}]
    end else if (_T_55) begin
      if (4'ha == deqPtrExt_rvalue) begin
        pending_10 <= 1'h0;
      end else begin
        pending_10 <= _GEN_27960;
      end
    end else begin
      pending_10 <= _GEN_27960;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[LoadQueueFlag.scala 443:30]
      pending_11 <= 1'h0; // @[LoadQueueFlag.scala 444:{21,21}]
    end else if (_T_55) begin
      if (4'hb == deqPtrExt_rvalue) begin
        pending_11 <= 1'h0;
      end else begin
        pending_11 <= _GEN_27961;
      end
    end else begin
      pending_11 <= _GEN_27961;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[LoadQueueFlag.scala 443:30]
      pending_12 <= 1'h0; // @[LoadQueueFlag.scala 444:{21,21}]
    end else if (_T_55) begin
      if (4'hc == deqPtrExt_rvalue) begin
        pending_12 <= 1'h0;
      end else begin
        pending_12 <= _GEN_27962;
      end
    end else begin
      pending_12 <= _GEN_27962;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[LoadQueueFlag.scala 443:30]
      pending_13 <= 1'h0; // @[LoadQueueFlag.scala 444:{21,21}]
    end else if (_T_55) begin
      if (4'hd == deqPtrExt_rvalue) begin
        pending_13 <= 1'h0;
      end else begin
        pending_13 <= _GEN_27963;
      end
    end else begin
      pending_13 <= _GEN_27963;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[LoadQueueFlag.scala 443:30]
      pending_14 <= 1'h0; // @[LoadQueueFlag.scala 444:{21,21}]
    end else if (_T_55) begin
      if (4'he == deqPtrExt_rvalue) begin
        pending_14 <= 1'h0;
      end else begin
        pending_14 <= _GEN_27964;
      end
    end else begin
      pending_14 <= _GEN_27964;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[LoadQueueFlag.scala 443:30]
      pending_15 <= 1'h0; // @[LoadQueueFlag.scala 444:{21,21}]
    end else if (_T_55) begin
      if (4'hf == deqPtrExt_rvalue) begin
        pending_15 <= 1'h0;
      end else begin
        pending_15 <= _GEN_27965;
      end
    end else begin
      pending_15 <= _GEN_27965;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[LoadQueueFlag.scala 501:29]
      writebacked_0 <= 1'h0;
    end else if (_T_61) begin // @[LoadQueueFlag.scala 286:31]
      writebacked_0 <= _GEN_31394; // @[LoadQueueFlag.scala 301:26 306:{34,34}]
    end else if (io_loadIn_1_valid) begin
      if (_issued_T_7) begin
        if (4'h0 == io_loadIn_1_bits_uop_lqIdx_value) begin
          writebacked_0 <= _datavalidVal_T_2 & ~hasExceptions_1;
        end else begin
          writebacked_0 <= _GEN_21445;
        end
      end else begin
        writebacked_0 <= _GEN_21445;
      end
    end else begin
      writebacked_0 <= _GEN_21445;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[LoadQueueFlag.scala 501:29]
      writebacked_1 <= 1'h0;
    end else if (_T_61) begin // @[LoadQueueFlag.scala 286:31]
      writebacked_1 <= _GEN_31395; // @[LoadQueueFlag.scala 301:26 306:{34,34}]
    end else if (io_loadIn_1_valid) begin
      if (_issued_T_7) begin
        if (4'h1 == io_loadIn_1_bits_uop_lqIdx_value) begin
          writebacked_1 <= _datavalidVal_T_2 & ~hasExceptions_1;
        end else begin
          writebacked_1 <= _GEN_21446;
        end
      end else begin
        writebacked_1 <= _GEN_21446;
      end
    end else begin
      writebacked_1 <= _GEN_21446;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[LoadQueueFlag.scala 501:29]
      writebacked_2 <= 1'h0;
    end else if (_T_61) begin // @[LoadQueueFlag.scala 286:31]
      writebacked_2 <= _GEN_31396; // @[LoadQueueFlag.scala 301:26 306:{34,34}]
    end else if (io_loadIn_1_valid) begin
      if (_issued_T_7) begin
        if (4'h2 == io_loadIn_1_bits_uop_lqIdx_value) begin
          writebacked_2 <= _datavalidVal_T_2 & ~hasExceptions_1;
        end else begin
          writebacked_2 <= _GEN_21447;
        end
      end else begin
        writebacked_2 <= _GEN_21447;
      end
    end else begin
      writebacked_2 <= _GEN_21447;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[LoadQueueFlag.scala 501:29]
      writebacked_3 <= 1'h0;
    end else if (_T_61) begin // @[LoadQueueFlag.scala 286:31]
      writebacked_3 <= _GEN_31397; // @[LoadQueueFlag.scala 301:26 306:{34,34}]
    end else if (io_loadIn_1_valid) begin
      if (_issued_T_7) begin
        if (4'h3 == io_loadIn_1_bits_uop_lqIdx_value) begin
          writebacked_3 <= _datavalidVal_T_2 & ~hasExceptions_1;
        end else begin
          writebacked_3 <= _GEN_21448;
        end
      end else begin
        writebacked_3 <= _GEN_21448;
      end
    end else begin
      writebacked_3 <= _GEN_21448;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[LoadQueueFlag.scala 501:29]
      writebacked_4 <= 1'h0;
    end else if (_T_61) begin // @[LoadQueueFlag.scala 286:31]
      writebacked_4 <= _GEN_31398; // @[LoadQueueFlag.scala 301:26 306:{34,34}]
    end else if (io_loadIn_1_valid) begin
      if (_issued_T_7) begin
        if (4'h4 == io_loadIn_1_bits_uop_lqIdx_value) begin
          writebacked_4 <= _datavalidVal_T_2 & ~hasExceptions_1;
        end else begin
          writebacked_4 <= _GEN_21449;
        end
      end else begin
        writebacked_4 <= _GEN_21449;
      end
    end else begin
      writebacked_4 <= _GEN_21449;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[LoadQueueFlag.scala 501:29]
      writebacked_5 <= 1'h0;
    end else if (_T_61) begin // @[LoadQueueFlag.scala 286:31]
      writebacked_5 <= _GEN_31399; // @[LoadQueueFlag.scala 301:26 306:{34,34}]
    end else if (io_loadIn_1_valid) begin
      if (_issued_T_7) begin
        if (4'h5 == io_loadIn_1_bits_uop_lqIdx_value) begin
          writebacked_5 <= _datavalidVal_T_2 & ~hasExceptions_1;
        end else begin
          writebacked_5 <= _GEN_21450;
        end
      end else begin
        writebacked_5 <= _GEN_21450;
      end
    end else begin
      writebacked_5 <= _GEN_21450;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[LoadQueueFlag.scala 501:29]
      writebacked_6 <= 1'h0;
    end else if (_T_61) begin // @[LoadQueueFlag.scala 286:31]
      writebacked_6 <= _GEN_31400; // @[LoadQueueFlag.scala 301:26 306:{34,34}]
    end else if (io_loadIn_1_valid) begin
      if (_issued_T_7) begin
        if (4'h6 == io_loadIn_1_bits_uop_lqIdx_value) begin
          writebacked_6 <= _datavalidVal_T_2 & ~hasExceptions_1;
        end else begin
          writebacked_6 <= _GEN_21451;
        end
      end else begin
        writebacked_6 <= _GEN_21451;
      end
    end else begin
      writebacked_6 <= _GEN_21451;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[LoadQueueFlag.scala 501:29]
      writebacked_7 <= 1'h0;
    end else if (_T_61) begin // @[LoadQueueFlag.scala 286:31]
      writebacked_7 <= _GEN_31401; // @[LoadQueueFlag.scala 301:26 306:{34,34}]
    end else if (io_loadIn_1_valid) begin
      if (_issued_T_7) begin
        if (4'h7 == io_loadIn_1_bits_uop_lqIdx_value) begin
          writebacked_7 <= _datavalidVal_T_2 & ~hasExceptions_1;
        end else begin
          writebacked_7 <= _GEN_21452;
        end
      end else begin
        writebacked_7 <= _GEN_21452;
      end
    end else begin
      writebacked_7 <= _GEN_21452;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[LoadQueueFlag.scala 501:29]
      writebacked_8 <= 1'h0;
    end else if (_T_61) begin // @[LoadQueueFlag.scala 286:31]
      writebacked_8 <= _GEN_31402; // @[LoadQueueFlag.scala 301:26 306:{34,34}]
    end else if (io_loadIn_1_valid) begin
      if (_issued_T_7) begin
        if (4'h8 == io_loadIn_1_bits_uop_lqIdx_value) begin
          writebacked_8 <= _datavalidVal_T_2 & ~hasExceptions_1;
        end else begin
          writebacked_8 <= _GEN_21453;
        end
      end else begin
        writebacked_8 <= _GEN_21453;
      end
    end else begin
      writebacked_8 <= _GEN_21453;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[LoadQueueFlag.scala 501:29]
      writebacked_9 <= 1'h0;
    end else if (_T_61) begin // @[LoadQueueFlag.scala 286:31]
      writebacked_9 <= _GEN_31403; // @[LoadQueueFlag.scala 301:26 306:{34,34}]
    end else if (io_loadIn_1_valid) begin
      if (_issued_T_7) begin
        if (4'h9 == io_loadIn_1_bits_uop_lqIdx_value) begin
          writebacked_9 <= _datavalidVal_T_2 & ~hasExceptions_1;
        end else begin
          writebacked_9 <= _GEN_21454;
        end
      end else begin
        writebacked_9 <= _GEN_21454;
      end
    end else begin
      writebacked_9 <= _GEN_21454;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[LoadQueueFlag.scala 501:29]
      writebacked_10 <= 1'h0;
    end else if (_T_61) begin // @[LoadQueueFlag.scala 286:31]
      writebacked_10 <= _GEN_31404; // @[LoadQueueFlag.scala 301:26 306:{34,34}]
    end else if (io_loadIn_1_valid) begin
      if (_issued_T_7) begin
        if (4'ha == io_loadIn_1_bits_uop_lqIdx_value) begin
          writebacked_10 <= _datavalidVal_T_2 & ~hasExceptions_1;
        end else begin
          writebacked_10 <= _GEN_21455;
        end
      end else begin
        writebacked_10 <= _GEN_21455;
      end
    end else begin
      writebacked_10 <= _GEN_21455;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[LoadQueueFlag.scala 501:29]
      writebacked_11 <= 1'h0;
    end else if (_T_61) begin // @[LoadQueueFlag.scala 286:31]
      writebacked_11 <= _GEN_31405; // @[LoadQueueFlag.scala 301:26 306:{34,34}]
    end else if (io_loadIn_1_valid) begin
      if (_issued_T_7) begin
        if (4'hb == io_loadIn_1_bits_uop_lqIdx_value) begin
          writebacked_11 <= _datavalidVal_T_2 & ~hasExceptions_1;
        end else begin
          writebacked_11 <= _GEN_21456;
        end
      end else begin
        writebacked_11 <= _GEN_21456;
      end
    end else begin
      writebacked_11 <= _GEN_21456;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[LoadQueueFlag.scala 501:29]
      writebacked_12 <= 1'h0;
    end else if (_T_61) begin // @[LoadQueueFlag.scala 286:31]
      writebacked_12 <= _GEN_31406; // @[LoadQueueFlag.scala 301:26 306:{34,34}]
    end else if (io_loadIn_1_valid) begin
      if (_issued_T_7) begin
        if (4'hc == io_loadIn_1_bits_uop_lqIdx_value) begin
          writebacked_12 <= _datavalidVal_T_2 & ~hasExceptions_1;
        end else begin
          writebacked_12 <= _GEN_21457;
        end
      end else begin
        writebacked_12 <= _GEN_21457;
      end
    end else begin
      writebacked_12 <= _GEN_21457;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[LoadQueueFlag.scala 501:29]
      writebacked_13 <= 1'h0;
    end else if (_T_61) begin // @[LoadQueueFlag.scala 286:31]
      writebacked_13 <= _GEN_31407; // @[LoadQueueFlag.scala 301:26 306:{34,34}]
    end else if (io_loadIn_1_valid) begin
      if (_issued_T_7) begin
        if (4'hd == io_loadIn_1_bits_uop_lqIdx_value) begin
          writebacked_13 <= _datavalidVal_T_2 & ~hasExceptions_1;
        end else begin
          writebacked_13 <= _GEN_21458;
        end
      end else begin
        writebacked_13 <= _GEN_21458;
      end
    end else begin
      writebacked_13 <= _GEN_21458;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[LoadQueueFlag.scala 501:29]
      writebacked_14 <= 1'h0;
    end else if (_T_61) begin // @[LoadQueueFlag.scala 286:31]
      writebacked_14 <= _GEN_31408; // @[LoadQueueFlag.scala 301:26 306:{34,34}]
    end else if (io_loadIn_1_valid) begin
      if (_issued_T_7) begin
        if (4'he == io_loadIn_1_bits_uop_lqIdx_value) begin
          writebacked_14 <= _datavalidVal_T_2 & ~hasExceptions_1;
        end else begin
          writebacked_14 <= _GEN_21459;
        end
      end else begin
        writebacked_14 <= _GEN_21459;
      end
    end else begin
      writebacked_14 <= _GEN_21459;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[LoadQueueFlag.scala 501:29]
      writebacked_15 <= 1'h0;
    end else if (_T_61) begin // @[LoadQueueFlag.scala 286:31]
      writebacked_15 <= _GEN_31409; // @[LoadQueueFlag.scala 301:26 306:{34,34}]
    end else if (io_loadIn_1_valid) begin
      if (_issued_T_7) begin
        if (4'hf == io_loadIn_1_bits_uop_lqIdx_value) begin
          writebacked_15 <= _datavalidVal_T_2 & ~hasExceptions_1;
        end else begin
          writebacked_15 <= _GEN_21460;
        end
      end else begin
        writebacked_15 <= _GEN_21460;
      end
    end else begin
      writebacked_15 <= _GEN_21460;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[LoadQueueFlag.scala 141:34]
      enqPtrExt_0_flag <= 1'h0; // @[LoadQueueFlag.scala 143:19]
    end else if (lastCycleRedirect_valid) begin // @[LoadQueueFlag.scala 145:19]
      enqPtrExt_0_flag <= new_ptr_flag;
    end else begin
      enqPtrExt_0_flag <= new_ptr_4_flag;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[LoadQueueFlag.scala 141:34]
      enqPtrExt_0_value <= 4'h0; // @[LoadQueueFlag.scala 143:19]
    end else if (lastCycleRedirect_valid) begin // @[LoadQueueFlag.scala 145:19]
      enqPtrExt_0_value <= flipped_new_ptr_value;
    end else begin
      enqPtrExt_0_value <= new_ptr_4_value;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      deqPtrExt_rflag <= 1'h0; // @[Reg.scala 29:22]
    end else if (deqPtrUpdateEna) begin // @[Reg.scala 28:20]
      deqPtrExt_rflag <= deqPtrExtNext_new_ptr_flag;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      deqPtrExt_rvalue <= 4'h0; // @[Reg.scala 29:22]
    end else if (deqPtrUpdateEna) begin // @[Reg.scala 28:20]
      deqPtrExt_rvalue <= deqPtrExtNext_new_ptr_value;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[LoadQueueFlag.scala 404:25]
      uncacheState <= 2'h0; // @[LoadQueueFlag.scala 406:100 407:22 397:29]
    end else if (2'h0 == uncacheState) begin // @[LoadQueueFlag.scala 404:25]
      if (REG) begin // @[LoadQueueFlag.scala 411:34]
        uncacheState <= 2'h1; // @[LoadQueueFlag.scala 412:22]
      end
    end else if (2'h1 == uncacheState) begin // @[LoadQueueFlag.scala 404:25]
      if (_T_55) begin // @[LoadQueueFlag.scala 416:35]
        uncacheState <= 2'h2; // @[LoadQueueFlag.scala 417:22]
      end
    end else if (2'h2 == uncacheState) begin // @[LoadQueueFlag.scala 404:25]
      if (_T_57) begin
        uncacheState <= 2'h3;
      end
    end else if (2'h3 == uncacheState) begin // @[LoadQueueFlag.scala 397:29]
      uncacheState <= _GEN_29580;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[LoadQueueFlag.scala 501:29]
      uncacheCommitFired <= 1'h0; // @[LoadQueueFlag.scala 503:24]
    end else begin
      uncacheCommitFired <= _T_61 | _GEN_29576;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  allocated_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  allocated_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  allocated_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  allocated_3 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  allocated_4 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  allocated_5 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  allocated_6 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  allocated_7 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  allocated_8 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  allocated_9 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  allocated_10 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  allocated_11 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  allocated_12 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  allocated_13 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  allocated_14 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  allocated_15 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  uop_0_cf_exceptionVec_4 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  uop_0_cf_exceptionVec_5 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  uop_0_cf_exceptionVec_13 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  uop_0_cf_trigger_backendEn_1 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  uop_0_cf_trigger_backendHit_0 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  uop_0_cf_trigger_backendHit_1 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  uop_0_cf_trigger_backendHit_4 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  uop_0_ctrl_fuOpType = _RAND_23[6:0];
  _RAND_24 = {1{`RANDOM}};
  uop_0_ctrl_rfWen = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  uop_0_ctrl_fpWen = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  uop_0_ctrl_flushPipe = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  uop_0_ctrl_replayInst = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  uop_0_pdest = _RAND_28[5:0];
  _RAND_29 = {1{`RANDOM}};
  uop_0_robIdx_flag = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  uop_0_robIdx_value = _RAND_30[4:0];
  _RAND_31 = {1{`RANDOM}};
  uop_1_cf_exceptionVec_4 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  uop_1_cf_exceptionVec_5 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  uop_1_cf_exceptionVec_13 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  uop_1_cf_trigger_backendEn_1 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  uop_1_cf_trigger_backendHit_0 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  uop_1_cf_trigger_backendHit_1 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  uop_1_cf_trigger_backendHit_4 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  uop_1_ctrl_fuOpType = _RAND_38[6:0];
  _RAND_39 = {1{`RANDOM}};
  uop_1_ctrl_rfWen = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  uop_1_ctrl_fpWen = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  uop_1_ctrl_flushPipe = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  uop_1_ctrl_replayInst = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  uop_1_pdest = _RAND_43[5:0];
  _RAND_44 = {1{`RANDOM}};
  uop_1_robIdx_flag = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  uop_1_robIdx_value = _RAND_45[4:0];
  _RAND_46 = {1{`RANDOM}};
  uop_2_cf_exceptionVec_4 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  uop_2_cf_exceptionVec_5 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  uop_2_cf_exceptionVec_13 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  uop_2_cf_trigger_backendEn_1 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  uop_2_cf_trigger_backendHit_0 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  uop_2_cf_trigger_backendHit_1 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  uop_2_cf_trigger_backendHit_4 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  uop_2_ctrl_fuOpType = _RAND_53[6:0];
  _RAND_54 = {1{`RANDOM}};
  uop_2_ctrl_rfWen = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  uop_2_ctrl_fpWen = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  uop_2_ctrl_flushPipe = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  uop_2_ctrl_replayInst = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  uop_2_pdest = _RAND_58[5:0];
  _RAND_59 = {1{`RANDOM}};
  uop_2_robIdx_flag = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  uop_2_robIdx_value = _RAND_60[4:0];
  _RAND_61 = {1{`RANDOM}};
  uop_3_cf_exceptionVec_4 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  uop_3_cf_exceptionVec_5 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  uop_3_cf_exceptionVec_13 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  uop_3_cf_trigger_backendEn_1 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  uop_3_cf_trigger_backendHit_0 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  uop_3_cf_trigger_backendHit_1 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  uop_3_cf_trigger_backendHit_4 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  uop_3_ctrl_fuOpType = _RAND_68[6:0];
  _RAND_69 = {1{`RANDOM}};
  uop_3_ctrl_rfWen = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  uop_3_ctrl_fpWen = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  uop_3_ctrl_flushPipe = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  uop_3_ctrl_replayInst = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  uop_3_pdest = _RAND_73[5:0];
  _RAND_74 = {1{`RANDOM}};
  uop_3_robIdx_flag = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  uop_3_robIdx_value = _RAND_75[4:0];
  _RAND_76 = {1{`RANDOM}};
  uop_4_cf_exceptionVec_4 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  uop_4_cf_exceptionVec_5 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  uop_4_cf_exceptionVec_13 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  uop_4_cf_trigger_backendEn_1 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  uop_4_cf_trigger_backendHit_0 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  uop_4_cf_trigger_backendHit_1 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  uop_4_cf_trigger_backendHit_4 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  uop_4_ctrl_fuOpType = _RAND_83[6:0];
  _RAND_84 = {1{`RANDOM}};
  uop_4_ctrl_rfWen = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  uop_4_ctrl_fpWen = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  uop_4_ctrl_flushPipe = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  uop_4_ctrl_replayInst = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  uop_4_pdest = _RAND_88[5:0];
  _RAND_89 = {1{`RANDOM}};
  uop_4_robIdx_flag = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  uop_4_robIdx_value = _RAND_90[4:0];
  _RAND_91 = {1{`RANDOM}};
  uop_5_cf_exceptionVec_4 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  uop_5_cf_exceptionVec_5 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  uop_5_cf_exceptionVec_13 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  uop_5_cf_trigger_backendEn_1 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  uop_5_cf_trigger_backendHit_0 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  uop_5_cf_trigger_backendHit_1 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  uop_5_cf_trigger_backendHit_4 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  uop_5_ctrl_fuOpType = _RAND_98[6:0];
  _RAND_99 = {1{`RANDOM}};
  uop_5_ctrl_rfWen = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  uop_5_ctrl_fpWen = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  uop_5_ctrl_flushPipe = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  uop_5_ctrl_replayInst = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  uop_5_pdest = _RAND_103[5:0];
  _RAND_104 = {1{`RANDOM}};
  uop_5_robIdx_flag = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  uop_5_robIdx_value = _RAND_105[4:0];
  _RAND_106 = {1{`RANDOM}};
  uop_6_cf_exceptionVec_4 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  uop_6_cf_exceptionVec_5 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  uop_6_cf_exceptionVec_13 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  uop_6_cf_trigger_backendEn_1 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  uop_6_cf_trigger_backendHit_0 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  uop_6_cf_trigger_backendHit_1 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  uop_6_cf_trigger_backendHit_4 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  uop_6_ctrl_fuOpType = _RAND_113[6:0];
  _RAND_114 = {1{`RANDOM}};
  uop_6_ctrl_rfWen = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  uop_6_ctrl_fpWen = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  uop_6_ctrl_flushPipe = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  uop_6_ctrl_replayInst = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  uop_6_pdest = _RAND_118[5:0];
  _RAND_119 = {1{`RANDOM}};
  uop_6_robIdx_flag = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  uop_6_robIdx_value = _RAND_120[4:0];
  _RAND_121 = {1{`RANDOM}};
  uop_7_cf_exceptionVec_4 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  uop_7_cf_exceptionVec_5 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  uop_7_cf_exceptionVec_13 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  uop_7_cf_trigger_backendEn_1 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  uop_7_cf_trigger_backendHit_0 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  uop_7_cf_trigger_backendHit_1 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  uop_7_cf_trigger_backendHit_4 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  uop_7_ctrl_fuOpType = _RAND_128[6:0];
  _RAND_129 = {1{`RANDOM}};
  uop_7_ctrl_rfWen = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  uop_7_ctrl_fpWen = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  uop_7_ctrl_flushPipe = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  uop_7_ctrl_replayInst = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  uop_7_pdest = _RAND_133[5:0];
  _RAND_134 = {1{`RANDOM}};
  uop_7_robIdx_flag = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  uop_7_robIdx_value = _RAND_135[4:0];
  _RAND_136 = {1{`RANDOM}};
  uop_8_cf_exceptionVec_4 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  uop_8_cf_exceptionVec_5 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  uop_8_cf_exceptionVec_13 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  uop_8_cf_trigger_backendEn_1 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  uop_8_cf_trigger_backendHit_0 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  uop_8_cf_trigger_backendHit_1 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  uop_8_cf_trigger_backendHit_4 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  uop_8_ctrl_fuOpType = _RAND_143[6:0];
  _RAND_144 = {1{`RANDOM}};
  uop_8_ctrl_rfWen = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  uop_8_ctrl_fpWen = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  uop_8_ctrl_flushPipe = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  uop_8_ctrl_replayInst = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  uop_8_pdest = _RAND_148[5:0];
  _RAND_149 = {1{`RANDOM}};
  uop_8_robIdx_flag = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  uop_8_robIdx_value = _RAND_150[4:0];
  _RAND_151 = {1{`RANDOM}};
  uop_9_cf_exceptionVec_4 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  uop_9_cf_exceptionVec_5 = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  uop_9_cf_exceptionVec_13 = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  uop_9_cf_trigger_backendEn_1 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  uop_9_cf_trigger_backendHit_0 = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  uop_9_cf_trigger_backendHit_1 = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  uop_9_cf_trigger_backendHit_4 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  uop_9_ctrl_fuOpType = _RAND_158[6:0];
  _RAND_159 = {1{`RANDOM}};
  uop_9_ctrl_rfWen = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  uop_9_ctrl_fpWen = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  uop_9_ctrl_flushPipe = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  uop_9_ctrl_replayInst = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  uop_9_pdest = _RAND_163[5:0];
  _RAND_164 = {1{`RANDOM}};
  uop_9_robIdx_flag = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  uop_9_robIdx_value = _RAND_165[4:0];
  _RAND_166 = {1{`RANDOM}};
  uop_10_cf_exceptionVec_4 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  uop_10_cf_exceptionVec_5 = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  uop_10_cf_exceptionVec_13 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  uop_10_cf_trigger_backendEn_1 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  uop_10_cf_trigger_backendHit_0 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  uop_10_cf_trigger_backendHit_1 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  uop_10_cf_trigger_backendHit_4 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  uop_10_ctrl_fuOpType = _RAND_173[6:0];
  _RAND_174 = {1{`RANDOM}};
  uop_10_ctrl_rfWen = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  uop_10_ctrl_fpWen = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  uop_10_ctrl_flushPipe = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  uop_10_ctrl_replayInst = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  uop_10_pdest = _RAND_178[5:0];
  _RAND_179 = {1{`RANDOM}};
  uop_10_robIdx_flag = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  uop_10_robIdx_value = _RAND_180[4:0];
  _RAND_181 = {1{`RANDOM}};
  uop_11_cf_exceptionVec_4 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  uop_11_cf_exceptionVec_5 = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  uop_11_cf_exceptionVec_13 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  uop_11_cf_trigger_backendEn_1 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  uop_11_cf_trigger_backendHit_0 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  uop_11_cf_trigger_backendHit_1 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  uop_11_cf_trigger_backendHit_4 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  uop_11_ctrl_fuOpType = _RAND_188[6:0];
  _RAND_189 = {1{`RANDOM}};
  uop_11_ctrl_rfWen = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  uop_11_ctrl_fpWen = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  uop_11_ctrl_flushPipe = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  uop_11_ctrl_replayInst = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  uop_11_pdest = _RAND_193[5:0];
  _RAND_194 = {1{`RANDOM}};
  uop_11_robIdx_flag = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  uop_11_robIdx_value = _RAND_195[4:0];
  _RAND_196 = {1{`RANDOM}};
  uop_12_cf_exceptionVec_4 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  uop_12_cf_exceptionVec_5 = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  uop_12_cf_exceptionVec_13 = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  uop_12_cf_trigger_backendEn_1 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  uop_12_cf_trigger_backendHit_0 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  uop_12_cf_trigger_backendHit_1 = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  uop_12_cf_trigger_backendHit_4 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  uop_12_ctrl_fuOpType = _RAND_203[6:0];
  _RAND_204 = {1{`RANDOM}};
  uop_12_ctrl_rfWen = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  uop_12_ctrl_fpWen = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  uop_12_ctrl_flushPipe = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  uop_12_ctrl_replayInst = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  uop_12_pdest = _RAND_208[5:0];
  _RAND_209 = {1{`RANDOM}};
  uop_12_robIdx_flag = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  uop_12_robIdx_value = _RAND_210[4:0];
  _RAND_211 = {1{`RANDOM}};
  uop_13_cf_exceptionVec_4 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  uop_13_cf_exceptionVec_5 = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  uop_13_cf_exceptionVec_13 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  uop_13_cf_trigger_backendEn_1 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  uop_13_cf_trigger_backendHit_0 = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  uop_13_cf_trigger_backendHit_1 = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  uop_13_cf_trigger_backendHit_4 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  uop_13_ctrl_fuOpType = _RAND_218[6:0];
  _RAND_219 = {1{`RANDOM}};
  uop_13_ctrl_rfWen = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  uop_13_ctrl_fpWen = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  uop_13_ctrl_flushPipe = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  uop_13_ctrl_replayInst = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  uop_13_pdest = _RAND_223[5:0];
  _RAND_224 = {1{`RANDOM}};
  uop_13_robIdx_flag = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  uop_13_robIdx_value = _RAND_225[4:0];
  _RAND_226 = {1{`RANDOM}};
  uop_14_cf_exceptionVec_4 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  uop_14_cf_exceptionVec_5 = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  uop_14_cf_exceptionVec_13 = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  uop_14_cf_trigger_backendEn_1 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  uop_14_cf_trigger_backendHit_0 = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  uop_14_cf_trigger_backendHit_1 = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  uop_14_cf_trigger_backendHit_4 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  uop_14_ctrl_fuOpType = _RAND_233[6:0];
  _RAND_234 = {1{`RANDOM}};
  uop_14_ctrl_rfWen = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  uop_14_ctrl_fpWen = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  uop_14_ctrl_flushPipe = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  uop_14_ctrl_replayInst = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  uop_14_pdest = _RAND_238[5:0];
  _RAND_239 = {1{`RANDOM}};
  uop_14_robIdx_flag = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  uop_14_robIdx_value = _RAND_240[4:0];
  _RAND_241 = {1{`RANDOM}};
  uop_15_cf_exceptionVec_4 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  uop_15_cf_exceptionVec_5 = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  uop_15_cf_exceptionVec_13 = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  uop_15_cf_trigger_backendEn_1 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  uop_15_cf_trigger_backendHit_0 = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  uop_15_cf_trigger_backendHit_1 = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  uop_15_cf_trigger_backendHit_4 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  uop_15_ctrl_fuOpType = _RAND_248[6:0];
  _RAND_249 = {1{`RANDOM}};
  uop_15_ctrl_rfWen = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  uop_15_ctrl_fpWen = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  uop_15_ctrl_flushPipe = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  uop_15_ctrl_replayInst = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  uop_15_pdest = _RAND_253[5:0];
  _RAND_254 = {1{`RANDOM}};
  uop_15_robIdx_flag = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  uop_15_robIdx_value = _RAND_255[4:0];
  _RAND_256 = {1{`RANDOM}};
  addrvalid_0 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  addrvalid_1 = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  addrvalid_2 = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  addrvalid_3 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  addrvalid_4 = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  addrvalid_5 = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  addrvalid_6 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  addrvalid_7 = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  addrvalid_8 = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  addrvalid_9 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  addrvalid_10 = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  addrvalid_11 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  addrvalid_12 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  addrvalid_13 = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  addrvalid_14 = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  addrvalid_15 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  datavalid_0 = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  datavalid_1 = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  datavalid_2 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  datavalid_3 = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  datavalid_4 = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  datavalid_5 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  datavalid_6 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  datavalid_7 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  datavalid_8 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  datavalid_9 = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  datavalid_10 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  datavalid_11 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  datavalid_12 = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  datavalid_13 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  datavalid_14 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  datavalid_15 = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  pending_0 = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  pending_1 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  pending_2 = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  pending_3 = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  pending_4 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  pending_5 = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  pending_6 = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  pending_7 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  pending_8 = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  pending_9 = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  pending_10 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  pending_11 = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  pending_12 = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  pending_13 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  pending_14 = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  pending_15 = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  writebacked_0 = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  writebacked_1 = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  writebacked_2 = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  writebacked_3 = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  writebacked_4 = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  writebacked_5 = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  writebacked_6 = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  writebacked_7 = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  writebacked_8 = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  writebacked_9 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  writebacked_10 = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  writebacked_11 = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  writebacked_12 = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  writebacked_13 = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  writebacked_14 = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  writebacked_15 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  enqPtrExt_0_flag = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  enqPtrExt_0_value = _RAND_321[3:0];
  _RAND_322 = {1{`RANDOM}};
  lastCycleRedirect_valid = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  deqPtrExt_rflag = _RAND_323[0:0];
  _RAND_324 = {1{`RANDOM}};
  deqPtrExt_rvalue = _RAND_324[3:0];
  _RAND_325 = {1{`RANDOM}};
  lastNeedCancel_0 = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  lastNeedCancel_1 = _RAND_326[0:0];
  _RAND_327 = {1{`RANDOM}};
  lastNeedCancel_2 = _RAND_327[0:0];
  _RAND_328 = {1{`RANDOM}};
  lastNeedCancel_3 = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  lastNeedCancel_4 = _RAND_329[0:0];
  _RAND_330 = {1{`RANDOM}};
  lastNeedCancel_5 = _RAND_330[0:0];
  _RAND_331 = {1{`RANDOM}};
  lastNeedCancel_6 = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  lastNeedCancel_7 = _RAND_332[0:0];
  _RAND_333 = {1{`RANDOM}};
  lastNeedCancel_8 = _RAND_333[0:0];
  _RAND_334 = {1{`RANDOM}};
  lastNeedCancel_9 = _RAND_334[0:0];
  _RAND_335 = {1{`RANDOM}};
  lastNeedCancel_10 = _RAND_335[0:0];
  _RAND_336 = {1{`RANDOM}};
  lastNeedCancel_11 = _RAND_336[0:0];
  _RAND_337 = {1{`RANDOM}};
  lastNeedCancel_12 = _RAND_337[0:0];
  _RAND_338 = {1{`RANDOM}};
  lastNeedCancel_13 = _RAND_338[0:0];
  _RAND_339 = {1{`RANDOM}};
  lastNeedCancel_14 = _RAND_339[0:0];
  _RAND_340 = {1{`RANDOM}};
  lastNeedCancel_15 = _RAND_340[0:0];
  _RAND_341 = {1{`RANDOM}};
  lastEnqCancel_REG_0 = _RAND_341[0:0];
  _RAND_342 = {1{`RANDOM}};
  lastEnqCancel_REG_1 = _RAND_342[0:0];
  _RAND_343 = {1{`RANDOM}};
  lastEnqCancel_REG_2 = _RAND_343[0:0];
  _RAND_344 = {1{`RANDOM}};
  lastEnqCancel_REG_3 = _RAND_344[0:0];
  _RAND_345 = {1{`RANDOM}};
  lastCommitCount = _RAND_345[1:0];
  _RAND_346 = {1{`RANDOM}};
  io_lqDeq_REG = _RAND_346[1:0];
  _RAND_347 = {1{`RANDOM}};
  io_lqCancelCnt_REG = _RAND_347[4:0];
  _RAND_348 = {1{`RANDOM}};
  io_rob_isMMIO_0_REG = _RAND_348[0:0];
  _RAND_349 = {1{`RANDOM}};
  io_rob_uop_0_REG_robIdx_value = _RAND_349[4:0];
  _RAND_350 = {1{`RANDOM}};
  io_rob_isMMIO_1_REG = _RAND_350[0:0];
  _RAND_351 = {1{`RANDOM}};
  io_rob_uop_1_REG_robIdx_value = _RAND_351[4:0];
  _RAND_352 = {1{`RANDOM}};
  uncacheState = _RAND_352[1:0];
  _RAND_353 = {1{`RANDOM}};
  uncacheCommitFired = _RAND_353[0:0];
  _RAND_354 = {1{`RANDOM}};
  REG = _RAND_354[0:0];
  _RAND_355 = {1{`RANDOM}};
  REG_1 = _RAND_355[0:0];
  _RAND_356 = {2{`RANDOM}};
  uncacheData = _RAND_356[63:0];
  _RAND_357 = {1{`RANDOM}};
  io_perf_0_value_REG = _RAND_357[0:0];
  _RAND_358 = {1{`RANDOM}};
  io_perf_0_value_REG_1 = _RAND_358[0:0];
  _RAND_359 = {1{`RANDOM}};
  io_perf_1_value_REG = _RAND_359[0:0];
  _RAND_360 = {1{`RANDOM}};
  io_perf_1_value_REG_1 = _RAND_360[0:0];
  _RAND_361 = {1{`RANDOM}};
  io_perf_2_value_REG = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  io_perf_2_value_REG_1 = _RAND_362[0:0];
  _RAND_363 = {1{`RANDOM}};
  io_perf_3_value_REG = _RAND_363[0:0];
  _RAND_364 = {1{`RANDOM}};
  io_perf_3_value_REG_1 = _RAND_364[0:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    allocated_0 = 1'h0;
  end
  if (reset) begin
    allocated_1 = 1'h0;
  end
  if (reset) begin
    allocated_2 = 1'h0;
  end
  if (reset) begin
    allocated_3 = 1'h0;
  end
  if (reset) begin
    allocated_4 = 1'h0;
  end
  if (reset) begin
    allocated_5 = 1'h0;
  end
  if (reset) begin
    allocated_6 = 1'h0;
  end
  if (reset) begin
    allocated_7 = 1'h0;
  end
  if (reset) begin
    allocated_8 = 1'h0;
  end
  if (reset) begin
    allocated_9 = 1'h0;
  end
  if (reset) begin
    allocated_10 = 1'h0;
  end
  if (reset) begin
    allocated_11 = 1'h0;
  end
  if (reset) begin
    allocated_12 = 1'h0;
  end
  if (reset) begin
    allocated_13 = 1'h0;
  end
  if (reset) begin
    allocated_14 = 1'h0;
  end
  if (reset) begin
    allocated_15 = 1'h0;
  end
  if (reset) begin
    addrvalid_0 = 1'h0;
  end
  if (reset) begin
    addrvalid_1 = 1'h0;
  end
  if (reset) begin
    addrvalid_2 = 1'h0;
  end
  if (reset) begin
    addrvalid_3 = 1'h0;
  end
  if (reset) begin
    addrvalid_4 = 1'h0;
  end
  if (reset) begin
    addrvalid_5 = 1'h0;
  end
  if (reset) begin
    addrvalid_6 = 1'h0;
  end
  if (reset) begin
    addrvalid_7 = 1'h0;
  end
  if (reset) begin
    addrvalid_8 = 1'h0;
  end
  if (reset) begin
    addrvalid_9 = 1'h0;
  end
  if (reset) begin
    addrvalid_10 = 1'h0;
  end
  if (reset) begin
    addrvalid_11 = 1'h0;
  end
  if (reset) begin
    addrvalid_12 = 1'h0;
  end
  if (reset) begin
    addrvalid_13 = 1'h0;
  end
  if (reset) begin
    addrvalid_14 = 1'h0;
  end
  if (reset) begin
    addrvalid_15 = 1'h0;
  end
  if (reset) begin
    datavalid_0 = 1'h0;
  end
  if (reset) begin
    datavalid_1 = 1'h0;
  end
  if (reset) begin
    datavalid_2 = 1'h0;
  end
  if (reset) begin
    datavalid_3 = 1'h0;
  end
  if (reset) begin
    datavalid_4 = 1'h0;
  end
  if (reset) begin
    datavalid_5 = 1'h0;
  end
  if (reset) begin
    datavalid_6 = 1'h0;
  end
  if (reset) begin
    datavalid_7 = 1'h0;
  end
  if (reset) begin
    datavalid_8 = 1'h0;
  end
  if (reset) begin
    datavalid_9 = 1'h0;
  end
  if (reset) begin
    datavalid_10 = 1'h0;
  end
  if (reset) begin
    datavalid_11 = 1'h0;
  end
  if (reset) begin
    datavalid_12 = 1'h0;
  end
  if (reset) begin
    datavalid_13 = 1'h0;
  end
  if (reset) begin
    datavalid_14 = 1'h0;
  end
  if (reset) begin
    datavalid_15 = 1'h0;
  end
  if (reset) begin
    pending_0 = 1'h0;
  end
  if (reset) begin
    pending_1 = 1'h0;
  end
  if (reset) begin
    pending_2 = 1'h0;
  end
  if (reset) begin
    pending_3 = 1'h0;
  end
  if (reset) begin
    pending_4 = 1'h0;
  end
  if (reset) begin
    pending_5 = 1'h0;
  end
  if (reset) begin
    pending_6 = 1'h0;
  end
  if (reset) begin
    pending_7 = 1'h0;
  end
  if (reset) begin
    pending_8 = 1'h0;
  end
  if (reset) begin
    pending_9 = 1'h0;
  end
  if (reset) begin
    pending_10 = 1'h0;
  end
  if (reset) begin
    pending_11 = 1'h0;
  end
  if (reset) begin
    pending_12 = 1'h0;
  end
  if (reset) begin
    pending_13 = 1'h0;
  end
  if (reset) begin
    pending_14 = 1'h0;
  end
  if (reset) begin
    pending_15 = 1'h0;
  end
  if (reset) begin
    writebacked_0 = 1'h0;
  end
  if (reset) begin
    writebacked_1 = 1'h0;
  end
  if (reset) begin
    writebacked_2 = 1'h0;
  end
  if (reset) begin
    writebacked_3 = 1'h0;
  end
  if (reset) begin
    writebacked_4 = 1'h0;
  end
  if (reset) begin
    writebacked_5 = 1'h0;
  end
  if (reset) begin
    writebacked_6 = 1'h0;
  end
  if (reset) begin
    writebacked_7 = 1'h0;
  end
  if (reset) begin
    writebacked_8 = 1'h0;
  end
  if (reset) begin
    writebacked_9 = 1'h0;
  end
  if (reset) begin
    writebacked_10 = 1'h0;
  end
  if (reset) begin
    writebacked_11 = 1'h0;
  end
  if (reset) begin
    writebacked_12 = 1'h0;
  end
  if (reset) begin
    writebacked_13 = 1'h0;
  end
  if (reset) begin
    writebacked_14 = 1'h0;
  end
  if (reset) begin
    writebacked_15 = 1'h0;
  end
  if (reset) begin
    enqPtrExt_0_flag = 1'h0;
  end
  if (reset) begin
    enqPtrExt_0_value = 4'h0;
  end
  if (reset) begin
    deqPtrExt_rflag = 1'h0;
  end
  if (reset) begin
    deqPtrExt_rvalue = 4'h0;
  end
  if (reset) begin
    uncacheState = 2'h0;
  end
  if (reset) begin
    uncacheCommitFired = 1'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule

