module FTBBank(
  input         clock,
  input         reset,
  input         io_s1_fire,
  output        io_req_pc_ready,
  input         io_req_pc_valid,
  input  [38:0] io_req_pc_bits,
  output        io_read_resp_valid,
  output [2:0]  io_read_resp_brSlots_0_offset,
  output [11:0] io_read_resp_brSlots_0_lower,
  output [1:0]  io_read_resp_brSlots_0_tarStat,
  output        io_read_resp_brSlots_0_sharing,
  output        io_read_resp_brSlots_0_valid,
  output [2:0]  io_read_resp_tailSlot_offset,
  output [19:0] io_read_resp_tailSlot_lower,
  output [1:0]  io_read_resp_tailSlot_tarStat,
  output        io_read_resp_tailSlot_sharing,
  output        io_read_resp_tailSlot_valid,
  output [2:0]  io_read_resp_pftAddr,
  output        io_read_resp_carry,
  output        io_read_resp_isCall,
  output        io_read_resp_isRet,
  output        io_read_resp_isJalr,
  output        io_read_resp_last_may_be_rvi_call,
  output        io_read_resp_always_taken_0,
  output        io_read_resp_always_taken_1,
  output        io_read_hits_valid,
  output [1:0]  io_read_hits_bits,
  input         io_u_req_pc_valid,
  input  [38:0] io_u_req_pc_bits,
  output        io_update_hits_valid,
  output [1:0]  io_update_hits_bits,
  input         io_update_access,
  input  [38:0] io_update_pc,
  input         io_update_write_data_valid,
  input         io_update_write_data_bits_entry_valid,
  input  [2:0]  io_update_write_data_bits_entry_brSlots_0_offset,
  input  [11:0] io_update_write_data_bits_entry_brSlots_0_lower,
  input  [1:0]  io_update_write_data_bits_entry_brSlots_0_tarStat,
  input         io_update_write_data_bits_entry_brSlots_0_sharing,
  input         io_update_write_data_bits_entry_brSlots_0_valid,
  input  [2:0]  io_update_write_data_bits_entry_tailSlot_offset,
  input  [19:0] io_update_write_data_bits_entry_tailSlot_lower,
  input  [1:0]  io_update_write_data_bits_entry_tailSlot_tarStat,
  input         io_update_write_data_bits_entry_tailSlot_sharing,
  input         io_update_write_data_bits_entry_tailSlot_valid,
  input  [2:0]  io_update_write_data_bits_entry_pftAddr,
  input         io_update_write_data_bits_entry_carry,
  input         io_update_write_data_bits_entry_isCall,
  input         io_update_write_data_bits_entry_isRet,
  input         io_update_write_data_bits_entry_isJalr,
  input         io_update_write_data_bits_entry_last_may_be_rvi_call,
  input         io_update_write_data_bits_entry_always_taken_0,
  input         io_update_write_data_bits_entry_always_taken_1,
  input  [19:0] io_update_write_data_bits_tag,
  input  [1:0]  io_update_write_way,
  input         io_update_write_alloc
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
`endif // RANDOMIZE_REG_INIT
  wire  ftb_clock; // @[FTB.scala 302:21]
  wire  ftb_reset; // @[FTB.scala 302:21]
  wire  ftb_io_rreq_ready; // @[FTB.scala 302:21]
  wire  ftb_io_rreq_valid; // @[FTB.scala 302:21]
  wire [8:0] ftb_io_rreq_bits_setIdx; // @[FTB.scala 302:21]
  wire  ftb_io_rresp_data_0_entry_valid; // @[FTB.scala 302:21]
  wire [2:0] ftb_io_rresp_data_0_entry_brSlots_0_offset; // @[FTB.scala 302:21]
  wire [11:0] ftb_io_rresp_data_0_entry_brSlots_0_lower; // @[FTB.scala 302:21]
  wire [1:0] ftb_io_rresp_data_0_entry_brSlots_0_tarStat; // @[FTB.scala 302:21]
  wire  ftb_io_rresp_data_0_entry_brSlots_0_sharing; // @[FTB.scala 302:21]
  wire  ftb_io_rresp_data_0_entry_brSlots_0_valid; // @[FTB.scala 302:21]
  wire [2:0] ftb_io_rresp_data_0_entry_tailSlot_offset; // @[FTB.scala 302:21]
  wire [19:0] ftb_io_rresp_data_0_entry_tailSlot_lower; // @[FTB.scala 302:21]
  wire [1:0] ftb_io_rresp_data_0_entry_tailSlot_tarStat; // @[FTB.scala 302:21]
  wire  ftb_io_rresp_data_0_entry_tailSlot_sharing; // @[FTB.scala 302:21]
  wire  ftb_io_rresp_data_0_entry_tailSlot_valid; // @[FTB.scala 302:21]
  wire [2:0] ftb_io_rresp_data_0_entry_pftAddr; // @[FTB.scala 302:21]
  wire  ftb_io_rresp_data_0_entry_carry; // @[FTB.scala 302:21]
  wire  ftb_io_rresp_data_0_entry_isCall; // @[FTB.scala 302:21]
  wire  ftb_io_rresp_data_0_entry_isRet; // @[FTB.scala 302:21]
  wire  ftb_io_rresp_data_0_entry_isJalr; // @[FTB.scala 302:21]
  wire  ftb_io_rresp_data_0_entry_last_may_be_rvi_call; // @[FTB.scala 302:21]
  wire  ftb_io_rresp_data_0_entry_always_taken_0; // @[FTB.scala 302:21]
  wire  ftb_io_rresp_data_0_entry_always_taken_1; // @[FTB.scala 302:21]
  wire [19:0] ftb_io_rresp_data_0_tag; // @[FTB.scala 302:21]
  wire  ftb_io_rresp_data_1_entry_valid; // @[FTB.scala 302:21]
  wire [2:0] ftb_io_rresp_data_1_entry_brSlots_0_offset; // @[FTB.scala 302:21]
  wire [11:0] ftb_io_rresp_data_1_entry_brSlots_0_lower; // @[FTB.scala 302:21]
  wire [1:0] ftb_io_rresp_data_1_entry_brSlots_0_tarStat; // @[FTB.scala 302:21]
  wire  ftb_io_rresp_data_1_entry_brSlots_0_sharing; // @[FTB.scala 302:21]
  wire  ftb_io_rresp_data_1_entry_brSlots_0_valid; // @[FTB.scala 302:21]
  wire [2:0] ftb_io_rresp_data_1_entry_tailSlot_offset; // @[FTB.scala 302:21]
  wire [19:0] ftb_io_rresp_data_1_entry_tailSlot_lower; // @[FTB.scala 302:21]
  wire [1:0] ftb_io_rresp_data_1_entry_tailSlot_tarStat; // @[FTB.scala 302:21]
  wire  ftb_io_rresp_data_1_entry_tailSlot_sharing; // @[FTB.scala 302:21]
  wire  ftb_io_rresp_data_1_entry_tailSlot_valid; // @[FTB.scala 302:21]
  wire [2:0] ftb_io_rresp_data_1_entry_pftAddr; // @[FTB.scala 302:21]
  wire  ftb_io_rresp_data_1_entry_carry; // @[FTB.scala 302:21]
  wire  ftb_io_rresp_data_1_entry_isCall; // @[FTB.scala 302:21]
  wire  ftb_io_rresp_data_1_entry_isRet; // @[FTB.scala 302:21]
  wire  ftb_io_rresp_data_1_entry_isJalr; // @[FTB.scala 302:21]
  wire  ftb_io_rresp_data_1_entry_last_may_be_rvi_call; // @[FTB.scala 302:21]
  wire  ftb_io_rresp_data_1_entry_always_taken_0; // @[FTB.scala 302:21]
  wire  ftb_io_rresp_data_1_entry_always_taken_1; // @[FTB.scala 302:21]
  wire [19:0] ftb_io_rresp_data_1_tag; // @[FTB.scala 302:21]
  wire  ftb_io_rresp_data_2_entry_valid; // @[FTB.scala 302:21]
  wire [2:0] ftb_io_rresp_data_2_entry_brSlots_0_offset; // @[FTB.scala 302:21]
  wire [11:0] ftb_io_rresp_data_2_entry_brSlots_0_lower; // @[FTB.scala 302:21]
  wire [1:0] ftb_io_rresp_data_2_entry_brSlots_0_tarStat; // @[FTB.scala 302:21]
  wire  ftb_io_rresp_data_2_entry_brSlots_0_sharing; // @[FTB.scala 302:21]
  wire  ftb_io_rresp_data_2_entry_brSlots_0_valid; // @[FTB.scala 302:21]
  wire [2:0] ftb_io_rresp_data_2_entry_tailSlot_offset; // @[FTB.scala 302:21]
  wire [19:0] ftb_io_rresp_data_2_entry_tailSlot_lower; // @[FTB.scala 302:21]
  wire [1:0] ftb_io_rresp_data_2_entry_tailSlot_tarStat; // @[FTB.scala 302:21]
  wire  ftb_io_rresp_data_2_entry_tailSlot_sharing; // @[FTB.scala 302:21]
  wire  ftb_io_rresp_data_2_entry_tailSlot_valid; // @[FTB.scala 302:21]
  wire [2:0] ftb_io_rresp_data_2_entry_pftAddr; // @[FTB.scala 302:21]
  wire  ftb_io_rresp_data_2_entry_carry; // @[FTB.scala 302:21]
  wire  ftb_io_rresp_data_2_entry_isCall; // @[FTB.scala 302:21]
  wire  ftb_io_rresp_data_2_entry_isRet; // @[FTB.scala 302:21]
  wire  ftb_io_rresp_data_2_entry_isJalr; // @[FTB.scala 302:21]
  wire  ftb_io_rresp_data_2_entry_last_may_be_rvi_call; // @[FTB.scala 302:21]
  wire  ftb_io_rresp_data_2_entry_always_taken_0; // @[FTB.scala 302:21]
  wire  ftb_io_rresp_data_2_entry_always_taken_1; // @[FTB.scala 302:21]
  wire [19:0] ftb_io_rresp_data_2_tag; // @[FTB.scala 302:21]
  wire  ftb_io_rresp_data_3_entry_valid; // @[FTB.scala 302:21]
  wire [2:0] ftb_io_rresp_data_3_entry_brSlots_0_offset; // @[FTB.scala 302:21]
  wire [11:0] ftb_io_rresp_data_3_entry_brSlots_0_lower; // @[FTB.scala 302:21]
  wire [1:0] ftb_io_rresp_data_3_entry_brSlots_0_tarStat; // @[FTB.scala 302:21]
  wire  ftb_io_rresp_data_3_entry_brSlots_0_sharing; // @[FTB.scala 302:21]
  wire  ftb_io_rresp_data_3_entry_brSlots_0_valid; // @[FTB.scala 302:21]
  wire [2:0] ftb_io_rresp_data_3_entry_tailSlot_offset; // @[FTB.scala 302:21]
  wire [19:0] ftb_io_rresp_data_3_entry_tailSlot_lower; // @[FTB.scala 302:21]
  wire [1:0] ftb_io_rresp_data_3_entry_tailSlot_tarStat; // @[FTB.scala 302:21]
  wire  ftb_io_rresp_data_3_entry_tailSlot_sharing; // @[FTB.scala 302:21]
  wire  ftb_io_rresp_data_3_entry_tailSlot_valid; // @[FTB.scala 302:21]
  wire [2:0] ftb_io_rresp_data_3_entry_pftAddr; // @[FTB.scala 302:21]
  wire  ftb_io_rresp_data_3_entry_carry; // @[FTB.scala 302:21]
  wire  ftb_io_rresp_data_3_entry_isCall; // @[FTB.scala 302:21]
  wire  ftb_io_rresp_data_3_entry_isRet; // @[FTB.scala 302:21]
  wire  ftb_io_rresp_data_3_entry_isJalr; // @[FTB.scala 302:21]
  wire  ftb_io_rresp_data_3_entry_last_may_be_rvi_call; // @[FTB.scala 302:21]
  wire  ftb_io_rresp_data_3_entry_always_taken_0; // @[FTB.scala 302:21]
  wire  ftb_io_rresp_data_3_entry_always_taken_1; // @[FTB.scala 302:21]
  wire [19:0] ftb_io_rresp_data_3_tag; // @[FTB.scala 302:21]
  wire  ftb_io_wreq_valid; // @[FTB.scala 302:21]
  wire [8:0] ftb_io_wreq_bits_setIdx; // @[FTB.scala 302:21]
  wire  ftb_io_wreq_bits_data_0_entry_valid; // @[FTB.scala 302:21]
  wire [2:0] ftb_io_wreq_bits_data_0_entry_brSlots_0_offset; // @[FTB.scala 302:21]
  wire [11:0] ftb_io_wreq_bits_data_0_entry_brSlots_0_lower; // @[FTB.scala 302:21]
  wire [1:0] ftb_io_wreq_bits_data_0_entry_brSlots_0_tarStat; // @[FTB.scala 302:21]
  wire  ftb_io_wreq_bits_data_0_entry_brSlots_0_sharing; // @[FTB.scala 302:21]
  wire  ftb_io_wreq_bits_data_0_entry_brSlots_0_valid; // @[FTB.scala 302:21]
  wire [2:0] ftb_io_wreq_bits_data_0_entry_tailSlot_offset; // @[FTB.scala 302:21]
  wire [19:0] ftb_io_wreq_bits_data_0_entry_tailSlot_lower; // @[FTB.scala 302:21]
  wire [1:0] ftb_io_wreq_bits_data_0_entry_tailSlot_tarStat; // @[FTB.scala 302:21]
  wire  ftb_io_wreq_bits_data_0_entry_tailSlot_sharing; // @[FTB.scala 302:21]
  wire  ftb_io_wreq_bits_data_0_entry_tailSlot_valid; // @[FTB.scala 302:21]
  wire [2:0] ftb_io_wreq_bits_data_0_entry_pftAddr; // @[FTB.scala 302:21]
  wire  ftb_io_wreq_bits_data_0_entry_carry; // @[FTB.scala 302:21]
  wire  ftb_io_wreq_bits_data_0_entry_isCall; // @[FTB.scala 302:21]
  wire  ftb_io_wreq_bits_data_0_entry_isRet; // @[FTB.scala 302:21]
  wire  ftb_io_wreq_bits_data_0_entry_isJalr; // @[FTB.scala 302:21]
  wire  ftb_io_wreq_bits_data_0_entry_last_may_be_rvi_call; // @[FTB.scala 302:21]
  wire  ftb_io_wreq_bits_data_0_entry_always_taken_0; // @[FTB.scala 302:21]
  wire  ftb_io_wreq_bits_data_0_entry_always_taken_1; // @[FTB.scala 302:21]
  wire [19:0] ftb_io_wreq_bits_data_0_tag; // @[FTB.scala 302:21]
  wire  ftb_io_wreq_bits_data_1_entry_valid; // @[FTB.scala 302:21]
  wire [2:0] ftb_io_wreq_bits_data_1_entry_brSlots_0_offset; // @[FTB.scala 302:21]
  wire [11:0] ftb_io_wreq_bits_data_1_entry_brSlots_0_lower; // @[FTB.scala 302:21]
  wire [1:0] ftb_io_wreq_bits_data_1_entry_brSlots_0_tarStat; // @[FTB.scala 302:21]
  wire  ftb_io_wreq_bits_data_1_entry_brSlots_0_sharing; // @[FTB.scala 302:21]
  wire  ftb_io_wreq_bits_data_1_entry_brSlots_0_valid; // @[FTB.scala 302:21]
  wire [2:0] ftb_io_wreq_bits_data_1_entry_tailSlot_offset; // @[FTB.scala 302:21]
  wire [19:0] ftb_io_wreq_bits_data_1_entry_tailSlot_lower; // @[FTB.scala 302:21]
  wire [1:0] ftb_io_wreq_bits_data_1_entry_tailSlot_tarStat; // @[FTB.scala 302:21]
  wire  ftb_io_wreq_bits_data_1_entry_tailSlot_sharing; // @[FTB.scala 302:21]
  wire  ftb_io_wreq_bits_data_1_entry_tailSlot_valid; // @[FTB.scala 302:21]
  wire [2:0] ftb_io_wreq_bits_data_1_entry_pftAddr; // @[FTB.scala 302:21]
  wire  ftb_io_wreq_bits_data_1_entry_carry; // @[FTB.scala 302:21]
  wire  ftb_io_wreq_bits_data_1_entry_isCall; // @[FTB.scala 302:21]
  wire  ftb_io_wreq_bits_data_1_entry_isRet; // @[FTB.scala 302:21]
  wire  ftb_io_wreq_bits_data_1_entry_isJalr; // @[FTB.scala 302:21]
  wire  ftb_io_wreq_bits_data_1_entry_last_may_be_rvi_call; // @[FTB.scala 302:21]
  wire  ftb_io_wreq_bits_data_1_entry_always_taken_0; // @[FTB.scala 302:21]
  wire  ftb_io_wreq_bits_data_1_entry_always_taken_1; // @[FTB.scala 302:21]
  wire [19:0] ftb_io_wreq_bits_data_1_tag; // @[FTB.scala 302:21]
  wire  ftb_io_wreq_bits_data_2_entry_valid; // @[FTB.scala 302:21]
  wire [2:0] ftb_io_wreq_bits_data_2_entry_brSlots_0_offset; // @[FTB.scala 302:21]
  wire [11:0] ftb_io_wreq_bits_data_2_entry_brSlots_0_lower; // @[FTB.scala 302:21]
  wire [1:0] ftb_io_wreq_bits_data_2_entry_brSlots_0_tarStat; // @[FTB.scala 302:21]
  wire  ftb_io_wreq_bits_data_2_entry_brSlots_0_sharing; // @[FTB.scala 302:21]
  wire  ftb_io_wreq_bits_data_2_entry_brSlots_0_valid; // @[FTB.scala 302:21]
  wire [2:0] ftb_io_wreq_bits_data_2_entry_tailSlot_offset; // @[FTB.scala 302:21]
  wire [19:0] ftb_io_wreq_bits_data_2_entry_tailSlot_lower; // @[FTB.scala 302:21]
  wire [1:0] ftb_io_wreq_bits_data_2_entry_tailSlot_tarStat; // @[FTB.scala 302:21]
  wire  ftb_io_wreq_bits_data_2_entry_tailSlot_sharing; // @[FTB.scala 302:21]
  wire  ftb_io_wreq_bits_data_2_entry_tailSlot_valid; // @[FTB.scala 302:21]
  wire [2:0] ftb_io_wreq_bits_data_2_entry_pftAddr; // @[FTB.scala 302:21]
  wire  ftb_io_wreq_bits_data_2_entry_carry; // @[FTB.scala 302:21]
  wire  ftb_io_wreq_bits_data_2_entry_isCall; // @[FTB.scala 302:21]
  wire  ftb_io_wreq_bits_data_2_entry_isRet; // @[FTB.scala 302:21]
  wire  ftb_io_wreq_bits_data_2_entry_isJalr; // @[FTB.scala 302:21]
  wire  ftb_io_wreq_bits_data_2_entry_last_may_be_rvi_call; // @[FTB.scala 302:21]
  wire  ftb_io_wreq_bits_data_2_entry_always_taken_0; // @[FTB.scala 302:21]
  wire  ftb_io_wreq_bits_data_2_entry_always_taken_1; // @[FTB.scala 302:21]
  wire [19:0] ftb_io_wreq_bits_data_2_tag; // @[FTB.scala 302:21]
  wire  ftb_io_wreq_bits_data_3_entry_valid; // @[FTB.scala 302:21]
  wire [2:0] ftb_io_wreq_bits_data_3_entry_brSlots_0_offset; // @[FTB.scala 302:21]
  wire [11:0] ftb_io_wreq_bits_data_3_entry_brSlots_0_lower; // @[FTB.scala 302:21]
  wire [1:0] ftb_io_wreq_bits_data_3_entry_brSlots_0_tarStat; // @[FTB.scala 302:21]
  wire  ftb_io_wreq_bits_data_3_entry_brSlots_0_sharing; // @[FTB.scala 302:21]
  wire  ftb_io_wreq_bits_data_3_entry_brSlots_0_valid; // @[FTB.scala 302:21]
  wire [2:0] ftb_io_wreq_bits_data_3_entry_tailSlot_offset; // @[FTB.scala 302:21]
  wire [19:0] ftb_io_wreq_bits_data_3_entry_tailSlot_lower; // @[FTB.scala 302:21]
  wire [1:0] ftb_io_wreq_bits_data_3_entry_tailSlot_tarStat; // @[FTB.scala 302:21]
  wire  ftb_io_wreq_bits_data_3_entry_tailSlot_sharing; // @[FTB.scala 302:21]
  wire  ftb_io_wreq_bits_data_3_entry_tailSlot_valid; // @[FTB.scala 302:21]
  wire [2:0] ftb_io_wreq_bits_data_3_entry_pftAddr; // @[FTB.scala 302:21]
  wire  ftb_io_wreq_bits_data_3_entry_carry; // @[FTB.scala 302:21]
  wire  ftb_io_wreq_bits_data_3_entry_isCall; // @[FTB.scala 302:21]
  wire  ftb_io_wreq_bits_data_3_entry_isRet; // @[FTB.scala 302:21]
  wire  ftb_io_wreq_bits_data_3_entry_isJalr; // @[FTB.scala 302:21]
  wire  ftb_io_wreq_bits_data_3_entry_last_may_be_rvi_call; // @[FTB.scala 302:21]
  wire  ftb_io_wreq_bits_data_3_entry_always_taken_0; // @[FTB.scala 302:21]
  wire  ftb_io_wreq_bits_data_3_entry_always_taken_1; // @[FTB.scala 302:21]
  wire [19:0] ftb_io_wreq_bits_data_3_tag; // @[FTB.scala 302:21]
  wire [3:0] ftb_io_wreq_bits_waymask; // @[FTB.scala 302:21]
  reg  pred_rdata_REG; // @[FTB.scala 305:62]
  reg  pred_rdata_hold_data_0_entry_valid; // @[Reg.scala 16:16]
  reg [2:0] pred_rdata_hold_data_0_entry_brSlots_0_offset; // @[Reg.scala 16:16]
  reg [11:0] pred_rdata_hold_data_0_entry_brSlots_0_lower; // @[Reg.scala 16:16]
  reg [1:0] pred_rdata_hold_data_0_entry_brSlots_0_tarStat; // @[Reg.scala 16:16]
  reg  pred_rdata_hold_data_0_entry_brSlots_0_sharing; // @[Reg.scala 16:16]
  reg  pred_rdata_hold_data_0_entry_brSlots_0_valid; // @[Reg.scala 16:16]
  reg [2:0] pred_rdata_hold_data_0_entry_tailSlot_offset; // @[Reg.scala 16:16]
  reg [19:0] pred_rdata_hold_data_0_entry_tailSlot_lower; // @[Reg.scala 16:16]
  reg [1:0] pred_rdata_hold_data_0_entry_tailSlot_tarStat; // @[Reg.scala 16:16]
  reg  pred_rdata_hold_data_0_entry_tailSlot_sharing; // @[Reg.scala 16:16]
  reg  pred_rdata_hold_data_0_entry_tailSlot_valid; // @[Reg.scala 16:16]
  reg [2:0] pred_rdata_hold_data_0_entry_pftAddr; // @[Reg.scala 16:16]
  reg  pred_rdata_hold_data_0_entry_carry; // @[Reg.scala 16:16]
  reg  pred_rdata_hold_data_0_entry_isCall; // @[Reg.scala 16:16]
  reg  pred_rdata_hold_data_0_entry_isRet; // @[Reg.scala 16:16]
  reg  pred_rdata_hold_data_0_entry_isJalr; // @[Reg.scala 16:16]
  reg  pred_rdata_hold_data_0_entry_last_may_be_rvi_call; // @[Reg.scala 16:16]
  reg  pred_rdata_hold_data_0_entry_always_taken_0; // @[Reg.scala 16:16]
  reg  pred_rdata_hold_data_0_entry_always_taken_1; // @[Reg.scala 16:16]
  reg [19:0] pred_rdata_hold_data_0_tag; // @[Reg.scala 16:16]
  reg  pred_rdata_hold_data_1_entry_valid; // @[Reg.scala 16:16]
  reg [2:0] pred_rdata_hold_data_1_entry_brSlots_0_offset; // @[Reg.scala 16:16]
  reg [11:0] pred_rdata_hold_data_1_entry_brSlots_0_lower; // @[Reg.scala 16:16]
  reg [1:0] pred_rdata_hold_data_1_entry_brSlots_0_tarStat; // @[Reg.scala 16:16]
  reg  pred_rdata_hold_data_1_entry_brSlots_0_sharing; // @[Reg.scala 16:16]
  reg  pred_rdata_hold_data_1_entry_brSlots_0_valid; // @[Reg.scala 16:16]
  reg [2:0] pred_rdata_hold_data_1_entry_tailSlot_offset; // @[Reg.scala 16:16]
  reg [19:0] pred_rdata_hold_data_1_entry_tailSlot_lower; // @[Reg.scala 16:16]
  reg [1:0] pred_rdata_hold_data_1_entry_tailSlot_tarStat; // @[Reg.scala 16:16]
  reg  pred_rdata_hold_data_1_entry_tailSlot_sharing; // @[Reg.scala 16:16]
  reg  pred_rdata_hold_data_1_entry_tailSlot_valid; // @[Reg.scala 16:16]
  reg [2:0] pred_rdata_hold_data_1_entry_pftAddr; // @[Reg.scala 16:16]
  reg  pred_rdata_hold_data_1_entry_carry; // @[Reg.scala 16:16]
  reg  pred_rdata_hold_data_1_entry_isCall; // @[Reg.scala 16:16]
  reg  pred_rdata_hold_data_1_entry_isRet; // @[Reg.scala 16:16]
  reg  pred_rdata_hold_data_1_entry_isJalr; // @[Reg.scala 16:16]
  reg  pred_rdata_hold_data_1_entry_last_may_be_rvi_call; // @[Reg.scala 16:16]
  reg  pred_rdata_hold_data_1_entry_always_taken_0; // @[Reg.scala 16:16]
  reg  pred_rdata_hold_data_1_entry_always_taken_1; // @[Reg.scala 16:16]
  reg [19:0] pred_rdata_hold_data_1_tag; // @[Reg.scala 16:16]
  reg  pred_rdata_hold_data_2_entry_valid; // @[Reg.scala 16:16]
  reg [2:0] pred_rdata_hold_data_2_entry_brSlots_0_offset; // @[Reg.scala 16:16]
  reg [11:0] pred_rdata_hold_data_2_entry_brSlots_0_lower; // @[Reg.scala 16:16]
  reg [1:0] pred_rdata_hold_data_2_entry_brSlots_0_tarStat; // @[Reg.scala 16:16]
  reg  pred_rdata_hold_data_2_entry_brSlots_0_sharing; // @[Reg.scala 16:16]
  reg  pred_rdata_hold_data_2_entry_brSlots_0_valid; // @[Reg.scala 16:16]
  reg [2:0] pred_rdata_hold_data_2_entry_tailSlot_offset; // @[Reg.scala 16:16]
  reg [19:0] pred_rdata_hold_data_2_entry_tailSlot_lower; // @[Reg.scala 16:16]
  reg [1:0] pred_rdata_hold_data_2_entry_tailSlot_tarStat; // @[Reg.scala 16:16]
  reg  pred_rdata_hold_data_2_entry_tailSlot_sharing; // @[Reg.scala 16:16]
  reg  pred_rdata_hold_data_2_entry_tailSlot_valid; // @[Reg.scala 16:16]
  reg [2:0] pred_rdata_hold_data_2_entry_pftAddr; // @[Reg.scala 16:16]
  reg  pred_rdata_hold_data_2_entry_carry; // @[Reg.scala 16:16]
  reg  pred_rdata_hold_data_2_entry_isCall; // @[Reg.scala 16:16]
  reg  pred_rdata_hold_data_2_entry_isRet; // @[Reg.scala 16:16]
  reg  pred_rdata_hold_data_2_entry_isJalr; // @[Reg.scala 16:16]
  reg  pred_rdata_hold_data_2_entry_last_may_be_rvi_call; // @[Reg.scala 16:16]
  reg  pred_rdata_hold_data_2_entry_always_taken_0; // @[Reg.scala 16:16]
  reg  pred_rdata_hold_data_2_entry_always_taken_1; // @[Reg.scala 16:16]
  reg [19:0] pred_rdata_hold_data_2_tag; // @[Reg.scala 16:16]
  reg  pred_rdata_hold_data_3_entry_valid; // @[Reg.scala 16:16]
  reg [2:0] pred_rdata_hold_data_3_entry_brSlots_0_offset; // @[Reg.scala 16:16]
  reg [11:0] pred_rdata_hold_data_3_entry_brSlots_0_lower; // @[Reg.scala 16:16]
  reg [1:0] pred_rdata_hold_data_3_entry_brSlots_0_tarStat; // @[Reg.scala 16:16]
  reg  pred_rdata_hold_data_3_entry_brSlots_0_sharing; // @[Reg.scala 16:16]
  reg  pred_rdata_hold_data_3_entry_brSlots_0_valid; // @[Reg.scala 16:16]
  reg [2:0] pred_rdata_hold_data_3_entry_tailSlot_offset; // @[Reg.scala 16:16]
  reg [19:0] pred_rdata_hold_data_3_entry_tailSlot_lower; // @[Reg.scala 16:16]
  reg [1:0] pred_rdata_hold_data_3_entry_tailSlot_tarStat; // @[Reg.scala 16:16]
  reg  pred_rdata_hold_data_3_entry_tailSlot_sharing; // @[Reg.scala 16:16]
  reg  pred_rdata_hold_data_3_entry_tailSlot_valid; // @[Reg.scala 16:16]
  reg [2:0] pred_rdata_hold_data_3_entry_pftAddr; // @[Reg.scala 16:16]
  reg  pred_rdata_hold_data_3_entry_carry; // @[Reg.scala 16:16]
  reg  pred_rdata_hold_data_3_entry_isCall; // @[Reg.scala 16:16]
  reg  pred_rdata_hold_data_3_entry_isRet; // @[Reg.scala 16:16]
  reg  pred_rdata_hold_data_3_entry_isJalr; // @[Reg.scala 16:16]
  reg  pred_rdata_hold_data_3_entry_last_may_be_rvi_call; // @[Reg.scala 16:16]
  reg  pred_rdata_hold_data_3_entry_always_taken_0; // @[Reg.scala 16:16]
  reg  pred_rdata_hold_data_3_entry_always_taken_1; // @[Reg.scala 16:16]
  reg [19:0] pred_rdata_hold_data_3_tag; // @[Reg.scala 16:16]
  wire  _GEN_0 = pred_rdata_REG ? ftb_io_rresp_data_0_entry_valid : pred_rdata_hold_data_0_entry_valid; // @[Reg.scala 16:16 17:{18,22}]
  wire [2:0] _GEN_1 = pred_rdata_REG ? ftb_io_rresp_data_0_entry_brSlots_0_offset :
    pred_rdata_hold_data_0_entry_brSlots_0_offset; // @[Reg.scala 16:16 17:{18,22}]
  wire [11:0] _GEN_2 = pred_rdata_REG ? ftb_io_rresp_data_0_entry_brSlots_0_lower :
    pred_rdata_hold_data_0_entry_brSlots_0_lower; // @[Reg.scala 16:16 17:{18,22}]
  wire [1:0] _GEN_3 = pred_rdata_REG ? ftb_io_rresp_data_0_entry_brSlots_0_tarStat :
    pred_rdata_hold_data_0_entry_brSlots_0_tarStat; // @[Reg.scala 16:16 17:{18,22}]
  wire  _GEN_4 = pred_rdata_REG ? ftb_io_rresp_data_0_entry_brSlots_0_sharing :
    pred_rdata_hold_data_0_entry_brSlots_0_sharing; // @[Reg.scala 16:16 17:{18,22}]
  wire  _GEN_5 = pred_rdata_REG ? ftb_io_rresp_data_0_entry_brSlots_0_valid :
    pred_rdata_hold_data_0_entry_brSlots_0_valid; // @[Reg.scala 16:16 17:{18,22}]
  wire [2:0] _GEN_6 = pred_rdata_REG ? ftb_io_rresp_data_0_entry_tailSlot_offset :
    pred_rdata_hold_data_0_entry_tailSlot_offset; // @[Reg.scala 16:16 17:{18,22}]
  wire [19:0] _GEN_7 = pred_rdata_REG ? ftb_io_rresp_data_0_entry_tailSlot_lower :
    pred_rdata_hold_data_0_entry_tailSlot_lower; // @[Reg.scala 16:16 17:{18,22}]
  wire [1:0] _GEN_8 = pred_rdata_REG ? ftb_io_rresp_data_0_entry_tailSlot_tarStat :
    pred_rdata_hold_data_0_entry_tailSlot_tarStat; // @[Reg.scala 16:16 17:{18,22}]
  wire  _GEN_9 = pred_rdata_REG ? ftb_io_rresp_data_0_entry_tailSlot_sharing :
    pred_rdata_hold_data_0_entry_tailSlot_sharing; // @[Reg.scala 16:16 17:{18,22}]
  wire  _GEN_10 = pred_rdata_REG ? ftb_io_rresp_data_0_entry_tailSlot_valid :
    pred_rdata_hold_data_0_entry_tailSlot_valid; // @[Reg.scala 16:16 17:{18,22}]
  wire [2:0] _GEN_11 = pred_rdata_REG ? ftb_io_rresp_data_0_entry_pftAddr : pred_rdata_hold_data_0_entry_pftAddr; // @[Reg.scala 16:16 17:{18,22}]
  wire  _GEN_12 = pred_rdata_REG ? ftb_io_rresp_data_0_entry_carry : pred_rdata_hold_data_0_entry_carry; // @[Reg.scala 16:16 17:{18,22}]
  wire  _GEN_13 = pred_rdata_REG ? ftb_io_rresp_data_0_entry_isCall : pred_rdata_hold_data_0_entry_isCall; // @[Reg.scala 16:16 17:{18,22}]
  wire  _GEN_14 = pred_rdata_REG ? ftb_io_rresp_data_0_entry_isRet : pred_rdata_hold_data_0_entry_isRet; // @[Reg.scala 16:16 17:{18,22}]
  wire  _GEN_15 = pred_rdata_REG ? ftb_io_rresp_data_0_entry_isJalr : pred_rdata_hold_data_0_entry_isJalr; // @[Reg.scala 16:16 17:{18,22}]
  wire  _GEN_16 = pred_rdata_REG ? ftb_io_rresp_data_0_entry_last_may_be_rvi_call :
    pred_rdata_hold_data_0_entry_last_may_be_rvi_call; // @[Reg.scala 16:16 17:{18,22}]
  wire  _GEN_17 = pred_rdata_REG ? ftb_io_rresp_data_0_entry_always_taken_0 :
    pred_rdata_hold_data_0_entry_always_taken_0; // @[Reg.scala 16:16 17:{18,22}]
  wire  _GEN_18 = pred_rdata_REG ? ftb_io_rresp_data_0_entry_always_taken_1 :
    pred_rdata_hold_data_0_entry_always_taken_1; // @[Reg.scala 16:16 17:{18,22}]
  wire [19:0] _GEN_19 = pred_rdata_REG ? ftb_io_rresp_data_0_tag : pred_rdata_hold_data_0_tag; // @[Reg.scala 16:16 17:{18,22}]
  wire  _GEN_20 = pred_rdata_REG ? ftb_io_rresp_data_1_entry_valid : pred_rdata_hold_data_1_entry_valid; // @[Reg.scala 16:16 17:{18,22}]
  wire [2:0] _GEN_21 = pred_rdata_REG ? ftb_io_rresp_data_1_entry_brSlots_0_offset :
    pred_rdata_hold_data_1_entry_brSlots_0_offset; // @[Reg.scala 16:16 17:{18,22}]
  wire [11:0] _GEN_22 = pred_rdata_REG ? ftb_io_rresp_data_1_entry_brSlots_0_lower :
    pred_rdata_hold_data_1_entry_brSlots_0_lower; // @[Reg.scala 16:16 17:{18,22}]
  wire [1:0] _GEN_23 = pred_rdata_REG ? ftb_io_rresp_data_1_entry_brSlots_0_tarStat :
    pred_rdata_hold_data_1_entry_brSlots_0_tarStat; // @[Reg.scala 16:16 17:{18,22}]
  wire  _GEN_24 = pred_rdata_REG ? ftb_io_rresp_data_1_entry_brSlots_0_sharing :
    pred_rdata_hold_data_1_entry_brSlots_0_sharing; // @[Reg.scala 16:16 17:{18,22}]
  wire  _GEN_25 = pred_rdata_REG ? ftb_io_rresp_data_1_entry_brSlots_0_valid :
    pred_rdata_hold_data_1_entry_brSlots_0_valid; // @[Reg.scala 16:16 17:{18,22}]
  wire [2:0] _GEN_26 = pred_rdata_REG ? ftb_io_rresp_data_1_entry_tailSlot_offset :
    pred_rdata_hold_data_1_entry_tailSlot_offset; // @[Reg.scala 16:16 17:{18,22}]
  wire [19:0] _GEN_27 = pred_rdata_REG ? ftb_io_rresp_data_1_entry_tailSlot_lower :
    pred_rdata_hold_data_1_entry_tailSlot_lower; // @[Reg.scala 16:16 17:{18,22}]
  wire [1:0] _GEN_28 = pred_rdata_REG ? ftb_io_rresp_data_1_entry_tailSlot_tarStat :
    pred_rdata_hold_data_1_entry_tailSlot_tarStat; // @[Reg.scala 16:16 17:{18,22}]
  wire  _GEN_29 = pred_rdata_REG ? ftb_io_rresp_data_1_entry_tailSlot_sharing :
    pred_rdata_hold_data_1_entry_tailSlot_sharing; // @[Reg.scala 16:16 17:{18,22}]
  wire  _GEN_30 = pred_rdata_REG ? ftb_io_rresp_data_1_entry_tailSlot_valid :
    pred_rdata_hold_data_1_entry_tailSlot_valid; // @[Reg.scala 16:16 17:{18,22}]
  wire [2:0] _GEN_31 = pred_rdata_REG ? ftb_io_rresp_data_1_entry_pftAddr : pred_rdata_hold_data_1_entry_pftAddr; // @[Reg.scala 16:16 17:{18,22}]
  wire  _GEN_32 = pred_rdata_REG ? ftb_io_rresp_data_1_entry_carry : pred_rdata_hold_data_1_entry_carry; // @[Reg.scala 16:16 17:{18,22}]
  wire  _GEN_33 = pred_rdata_REG ? ftb_io_rresp_data_1_entry_isCall : pred_rdata_hold_data_1_entry_isCall; // @[Reg.scala 16:16 17:{18,22}]
  wire  _GEN_34 = pred_rdata_REG ? ftb_io_rresp_data_1_entry_isRet : pred_rdata_hold_data_1_entry_isRet; // @[Reg.scala 16:16 17:{18,22}]
  wire  _GEN_35 = pred_rdata_REG ? ftb_io_rresp_data_1_entry_isJalr : pred_rdata_hold_data_1_entry_isJalr; // @[Reg.scala 16:16 17:{18,22}]
  wire  _GEN_36 = pred_rdata_REG ? ftb_io_rresp_data_1_entry_last_may_be_rvi_call :
    pred_rdata_hold_data_1_entry_last_may_be_rvi_call; // @[Reg.scala 16:16 17:{18,22}]
  wire  _GEN_37 = pred_rdata_REG ? ftb_io_rresp_data_1_entry_always_taken_0 :
    pred_rdata_hold_data_1_entry_always_taken_0; // @[Reg.scala 16:16 17:{18,22}]
  wire  _GEN_38 = pred_rdata_REG ? ftb_io_rresp_data_1_entry_always_taken_1 :
    pred_rdata_hold_data_1_entry_always_taken_1; // @[Reg.scala 16:16 17:{18,22}]
  wire [19:0] _GEN_39 = pred_rdata_REG ? ftb_io_rresp_data_1_tag : pred_rdata_hold_data_1_tag; // @[Reg.scala 16:16 17:{18,22}]
  wire  _GEN_40 = pred_rdata_REG ? ftb_io_rresp_data_2_entry_valid : pred_rdata_hold_data_2_entry_valid; // @[Reg.scala 16:16 17:{18,22}]
  wire [2:0] _GEN_41 = pred_rdata_REG ? ftb_io_rresp_data_2_entry_brSlots_0_offset :
    pred_rdata_hold_data_2_entry_brSlots_0_offset; // @[Reg.scala 16:16 17:{18,22}]
  wire [11:0] _GEN_42 = pred_rdata_REG ? ftb_io_rresp_data_2_entry_brSlots_0_lower :
    pred_rdata_hold_data_2_entry_brSlots_0_lower; // @[Reg.scala 16:16 17:{18,22}]
  wire [1:0] _GEN_43 = pred_rdata_REG ? ftb_io_rresp_data_2_entry_brSlots_0_tarStat :
    pred_rdata_hold_data_2_entry_brSlots_0_tarStat; // @[Reg.scala 16:16 17:{18,22}]
  wire  _GEN_44 = pred_rdata_REG ? ftb_io_rresp_data_2_entry_brSlots_0_sharing :
    pred_rdata_hold_data_2_entry_brSlots_0_sharing; // @[Reg.scala 16:16 17:{18,22}]
  wire  _GEN_45 = pred_rdata_REG ? ftb_io_rresp_data_2_entry_brSlots_0_valid :
    pred_rdata_hold_data_2_entry_brSlots_0_valid; // @[Reg.scala 16:16 17:{18,22}]
  wire [2:0] _GEN_46 = pred_rdata_REG ? ftb_io_rresp_data_2_entry_tailSlot_offset :
    pred_rdata_hold_data_2_entry_tailSlot_offset; // @[Reg.scala 16:16 17:{18,22}]
  wire [19:0] _GEN_47 = pred_rdata_REG ? ftb_io_rresp_data_2_entry_tailSlot_lower :
    pred_rdata_hold_data_2_entry_tailSlot_lower; // @[Reg.scala 16:16 17:{18,22}]
  wire [1:0] _GEN_48 = pred_rdata_REG ? ftb_io_rresp_data_2_entry_tailSlot_tarStat :
    pred_rdata_hold_data_2_entry_tailSlot_tarStat; // @[Reg.scala 16:16 17:{18,22}]
  wire  _GEN_49 = pred_rdata_REG ? ftb_io_rresp_data_2_entry_tailSlot_sharing :
    pred_rdata_hold_data_2_entry_tailSlot_sharing; // @[Reg.scala 16:16 17:{18,22}]
  wire  _GEN_50 = pred_rdata_REG ? ftb_io_rresp_data_2_entry_tailSlot_valid :
    pred_rdata_hold_data_2_entry_tailSlot_valid; // @[Reg.scala 16:16 17:{18,22}]
  wire [2:0] _GEN_51 = pred_rdata_REG ? ftb_io_rresp_data_2_entry_pftAddr : pred_rdata_hold_data_2_entry_pftAddr; // @[Reg.scala 16:16 17:{18,22}]
  wire  _GEN_52 = pred_rdata_REG ? ftb_io_rresp_data_2_entry_carry : pred_rdata_hold_data_2_entry_carry; // @[Reg.scala 16:16 17:{18,22}]
  wire  _GEN_53 = pred_rdata_REG ? ftb_io_rresp_data_2_entry_isCall : pred_rdata_hold_data_2_entry_isCall; // @[Reg.scala 16:16 17:{18,22}]
  wire  _GEN_54 = pred_rdata_REG ? ftb_io_rresp_data_2_entry_isRet : pred_rdata_hold_data_2_entry_isRet; // @[Reg.scala 16:16 17:{18,22}]
  wire  _GEN_55 = pred_rdata_REG ? ftb_io_rresp_data_2_entry_isJalr : pred_rdata_hold_data_2_entry_isJalr; // @[Reg.scala 16:16 17:{18,22}]
  wire  _GEN_56 = pred_rdata_REG ? ftb_io_rresp_data_2_entry_last_may_be_rvi_call :
    pred_rdata_hold_data_2_entry_last_may_be_rvi_call; // @[Reg.scala 16:16 17:{18,22}]
  wire  _GEN_57 = pred_rdata_REG ? ftb_io_rresp_data_2_entry_always_taken_0 :
    pred_rdata_hold_data_2_entry_always_taken_0; // @[Reg.scala 16:16 17:{18,22}]
  wire  _GEN_58 = pred_rdata_REG ? ftb_io_rresp_data_2_entry_always_taken_1 :
    pred_rdata_hold_data_2_entry_always_taken_1; // @[Reg.scala 16:16 17:{18,22}]
  wire [19:0] _GEN_59 = pred_rdata_REG ? ftb_io_rresp_data_2_tag : pred_rdata_hold_data_2_tag; // @[Reg.scala 16:16 17:{18,22}]
  wire  _GEN_60 = pred_rdata_REG ? ftb_io_rresp_data_3_entry_valid : pred_rdata_hold_data_3_entry_valid; // @[Reg.scala 16:16 17:{18,22}]
  wire [2:0] _GEN_61 = pred_rdata_REG ? ftb_io_rresp_data_3_entry_brSlots_0_offset :
    pred_rdata_hold_data_3_entry_brSlots_0_offset; // @[Reg.scala 16:16 17:{18,22}]
  wire [11:0] _GEN_62 = pred_rdata_REG ? ftb_io_rresp_data_3_entry_brSlots_0_lower :
    pred_rdata_hold_data_3_entry_brSlots_0_lower; // @[Reg.scala 16:16 17:{18,22}]
  wire [1:0] _GEN_63 = pred_rdata_REG ? ftb_io_rresp_data_3_entry_brSlots_0_tarStat :
    pred_rdata_hold_data_3_entry_brSlots_0_tarStat; // @[Reg.scala 16:16 17:{18,22}]
  wire  _GEN_64 = pred_rdata_REG ? ftb_io_rresp_data_3_entry_brSlots_0_sharing :
    pred_rdata_hold_data_3_entry_brSlots_0_sharing; // @[Reg.scala 16:16 17:{18,22}]
  wire  _GEN_65 = pred_rdata_REG ? ftb_io_rresp_data_3_entry_brSlots_0_valid :
    pred_rdata_hold_data_3_entry_brSlots_0_valid; // @[Reg.scala 16:16 17:{18,22}]
  wire [2:0] _GEN_66 = pred_rdata_REG ? ftb_io_rresp_data_3_entry_tailSlot_offset :
    pred_rdata_hold_data_3_entry_tailSlot_offset; // @[Reg.scala 16:16 17:{18,22}]
  wire [19:0] _GEN_67 = pred_rdata_REG ? ftb_io_rresp_data_3_entry_tailSlot_lower :
    pred_rdata_hold_data_3_entry_tailSlot_lower; // @[Reg.scala 16:16 17:{18,22}]
  wire [1:0] _GEN_68 = pred_rdata_REG ? ftb_io_rresp_data_3_entry_tailSlot_tarStat :
    pred_rdata_hold_data_3_entry_tailSlot_tarStat; // @[Reg.scala 16:16 17:{18,22}]
  wire  _GEN_69 = pred_rdata_REG ? ftb_io_rresp_data_3_entry_tailSlot_sharing :
    pred_rdata_hold_data_3_entry_tailSlot_sharing; // @[Reg.scala 16:16 17:{18,22}]
  wire  _GEN_70 = pred_rdata_REG ? ftb_io_rresp_data_3_entry_tailSlot_valid :
    pred_rdata_hold_data_3_entry_tailSlot_valid; // @[Reg.scala 16:16 17:{18,22}]
  wire [2:0] _GEN_71 = pred_rdata_REG ? ftb_io_rresp_data_3_entry_pftAddr : pred_rdata_hold_data_3_entry_pftAddr; // @[Reg.scala 16:16 17:{18,22}]
  wire  _GEN_72 = pred_rdata_REG ? ftb_io_rresp_data_3_entry_carry : pred_rdata_hold_data_3_entry_carry; // @[Reg.scala 16:16 17:{18,22}]
  wire  _GEN_73 = pred_rdata_REG ? ftb_io_rresp_data_3_entry_isCall : pred_rdata_hold_data_3_entry_isCall; // @[Reg.scala 16:16 17:{18,22}]
  wire  _GEN_74 = pred_rdata_REG ? ftb_io_rresp_data_3_entry_isRet : pred_rdata_hold_data_3_entry_isRet; // @[Reg.scala 16:16 17:{18,22}]
  wire  _GEN_75 = pred_rdata_REG ? ftb_io_rresp_data_3_entry_isJalr : pred_rdata_hold_data_3_entry_isJalr; // @[Reg.scala 16:16 17:{18,22}]
  wire  _GEN_76 = pred_rdata_REG ? ftb_io_rresp_data_3_entry_last_may_be_rvi_call :
    pred_rdata_hold_data_3_entry_last_may_be_rvi_call; // @[Reg.scala 16:16 17:{18,22}]
  wire  _GEN_77 = pred_rdata_REG ? ftb_io_rresp_data_3_entry_always_taken_0 :
    pred_rdata_hold_data_3_entry_always_taken_0; // @[Reg.scala 16:16 17:{18,22}]
  wire  _GEN_78 = pred_rdata_REG ? ftb_io_rresp_data_3_entry_always_taken_1 :
    pred_rdata_hold_data_3_entry_always_taken_1; // @[Reg.scala 16:16 17:{18,22}]
  wire [19:0] _GEN_79 = pred_rdata_REG ? ftb_io_rresp_data_3_tag : pred_rdata_hold_data_3_tag; // @[Reg.scala 16:16 17:{18,22}]
  reg [19:0] req_tag; // @[Reg.scala 16:16]
  reg [8:0] req_idx; // @[Reg.scala 16:16]
  reg [19:0] u_req_tag; // @[Reg.scala 16:16]
  wire  total_hits_0 = _GEN_19 == req_tag & _GEN_0 & io_s1_fire; // @[FTB.scala 322:107]
  wire  total_hits_1 = _GEN_39 == req_tag & _GEN_20 & io_s1_fire; // @[FTB.scala 322:107]
  wire  total_hits_2 = _GEN_59 == req_tag & _GEN_40 & io_s1_fire; // @[FTB.scala 322:107]
  wire  total_hits_3 = _GEN_79 == req_tag & _GEN_60 & io_s1_fire; // @[FTB.scala 322:107]
  wire  hit = total_hits_0 | total_hits_1 | total_hits_2 | total_hits_3; // @[FTB.scala 323:34]
  wire [3:0] _hit_way_T = {total_hits_3,total_hits_2,total_hits_1,total_hits_0}; // @[OneHot.scala 22:45]
  wire [1:0] hit_way_hi_1 = _hit_way_T[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] hit_way_lo_1 = _hit_way_T[1:0]; // @[OneHot.scala 31:18]
  wire  _hit_way_T_1 = |hit_way_hi_1; // @[OneHot.scala 32:14]
  wire [1:0] _hit_way_T_2 = hit_way_hi_1 | hit_way_lo_1; // @[OneHot.scala 32:28]
  wire [1:0] hit_way = {_hit_way_T_1,_hit_way_T_2[1]}; // @[Cat.scala 31:58]
  reg  u_total_hits_REG; // @[FTB.scala 328:96]
  wire  u_total_hits_0 = ftb_io_rresp_data_0_tag == u_req_tag & ftb_io_rresp_data_0_entry_valid & u_total_hits_REG; // @[FTB.scala 328:86]
  reg  u_total_hits_REG_1; // @[FTB.scala 328:96]
  wire  u_total_hits_1 = ftb_io_rresp_data_1_tag == u_req_tag & ftb_io_rresp_data_1_entry_valid & u_total_hits_REG_1; // @[FTB.scala 328:86]
  reg  u_total_hits_REG_2; // @[FTB.scala 328:96]
  wire  u_total_hits_2 = ftb_io_rresp_data_2_tag == u_req_tag & ftb_io_rresp_data_2_entry_valid & u_total_hits_REG_2; // @[FTB.scala 328:86]
  reg  u_total_hits_REG_3; // @[FTB.scala 328:96]
  wire  u_total_hits_3 = ftb_io_rresp_data_3_tag == u_req_tag & ftb_io_rresp_data_3_entry_valid & u_total_hits_REG_3; // @[FTB.scala 328:86]
  wire [3:0] _u_hit_way_T = {u_total_hits_3,u_total_hits_2,u_total_hits_1,u_total_hits_0}; // @[OneHot.scala 22:45]
  wire [1:0] u_hit_way_hi_1 = _u_hit_way_T[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] u_hit_way_lo_1 = _u_hit_way_T[1:0]; // @[OneHot.scala 31:18]
  wire  _u_hit_way_T_1 = |u_hit_way_hi_1; // @[OneHot.scala 32:14]
  wire [1:0] _u_hit_way_T_2 = u_hit_way_hi_1 | u_hit_way_lo_1; // @[OneHot.scala 32:28]
  reg [2:0] state_vec_0; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_1; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_2; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_3; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_4; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_5; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_6; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_7; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_8; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_9; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_10; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_11; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_12; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_13; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_14; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_15; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_16; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_17; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_18; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_19; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_20; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_21; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_22; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_23; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_24; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_25; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_26; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_27; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_28; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_29; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_30; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_31; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_32; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_33; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_34; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_35; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_36; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_37; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_38; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_39; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_40; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_41; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_42; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_43; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_44; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_45; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_46; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_47; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_48; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_49; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_50; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_51; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_52; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_53; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_54; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_55; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_56; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_57; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_58; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_59; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_60; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_61; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_62; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_63; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_64; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_65; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_66; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_67; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_68; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_69; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_70; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_71; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_72; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_73; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_74; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_75; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_76; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_77; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_78; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_79; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_80; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_81; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_82; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_83; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_84; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_85; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_86; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_87; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_88; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_89; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_90; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_91; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_92; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_93; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_94; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_95; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_96; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_97; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_98; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_99; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_100; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_101; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_102; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_103; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_104; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_105; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_106; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_107; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_108; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_109; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_110; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_111; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_112; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_113; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_114; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_115; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_116; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_117; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_118; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_119; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_120; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_121; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_122; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_123; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_124; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_125; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_126; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_127; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_128; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_129; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_130; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_131; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_132; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_133; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_134; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_135; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_136; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_137; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_138; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_139; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_140; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_141; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_142; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_143; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_144; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_145; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_146; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_147; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_148; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_149; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_150; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_151; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_152; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_153; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_154; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_155; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_156; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_157; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_158; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_159; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_160; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_161; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_162; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_163; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_164; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_165; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_166; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_167; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_168; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_169; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_170; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_171; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_172; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_173; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_174; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_175; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_176; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_177; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_178; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_179; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_180; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_181; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_182; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_183; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_184; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_185; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_186; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_187; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_188; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_189; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_190; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_191; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_192; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_193; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_194; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_195; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_196; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_197; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_198; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_199; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_200; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_201; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_202; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_203; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_204; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_205; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_206; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_207; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_208; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_209; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_210; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_211; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_212; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_213; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_214; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_215; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_216; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_217; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_218; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_219; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_220; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_221; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_222; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_223; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_224; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_225; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_226; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_227; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_228; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_229; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_230; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_231; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_232; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_233; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_234; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_235; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_236; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_237; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_238; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_239; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_240; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_241; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_242; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_243; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_244; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_245; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_246; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_247; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_248; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_249; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_250; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_251; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_252; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_253; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_254; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_255; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_256; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_257; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_258; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_259; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_260; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_261; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_262; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_263; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_264; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_265; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_266; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_267; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_268; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_269; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_270; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_271; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_272; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_273; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_274; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_275; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_276; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_277; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_278; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_279; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_280; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_281; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_282; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_283; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_284; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_285; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_286; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_287; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_288; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_289; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_290; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_291; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_292; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_293; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_294; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_295; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_296; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_297; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_298; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_299; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_300; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_301; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_302; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_303; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_304; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_305; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_306; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_307; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_308; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_309; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_310; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_311; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_312; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_313; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_314; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_315; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_316; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_317; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_318; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_319; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_320; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_321; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_322; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_323; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_324; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_325; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_326; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_327; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_328; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_329; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_330; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_331; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_332; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_333; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_334; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_335; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_336; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_337; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_338; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_339; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_340; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_341; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_342; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_343; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_344; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_345; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_346; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_347; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_348; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_349; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_350; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_351; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_352; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_353; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_354; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_355; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_356; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_357; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_358; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_359; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_360; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_361; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_362; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_363; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_364; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_365; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_366; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_367; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_368; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_369; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_370; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_371; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_372; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_373; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_374; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_375; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_376; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_377; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_378; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_379; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_380; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_381; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_382; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_383; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_384; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_385; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_386; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_387; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_388; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_389; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_390; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_391; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_392; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_393; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_394; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_395; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_396; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_397; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_398; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_399; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_400; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_401; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_402; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_403; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_404; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_405; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_406; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_407; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_408; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_409; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_410; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_411; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_412; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_413; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_414; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_415; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_416; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_417; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_418; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_419; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_420; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_421; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_422; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_423; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_424; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_425; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_426; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_427; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_428; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_429; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_430; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_431; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_432; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_433; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_434; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_435; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_436; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_437; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_438; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_439; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_440; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_441; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_442; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_443; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_444; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_445; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_446; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_447; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_448; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_449; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_450; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_451; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_452; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_453; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_454; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_455; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_456; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_457; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_458; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_459; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_460; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_461; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_462; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_463; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_464; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_465; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_466; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_467; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_468; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_469; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_470; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_471; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_472; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_473; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_474; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_475; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_476; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_477; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_478; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_479; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_480; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_481; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_482; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_483; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_484; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_485; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_486; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_487; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_488; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_489; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_490; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_491; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_492; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_493; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_494; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_495; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_496; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_497; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_498; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_499; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_500; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_501; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_502; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_503; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_504; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_505; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_506; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_507; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_508; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_509; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_510; // @[Replacement.scala 305:17]
  reg [2:0] state_vec_511; // @[Replacement.scala 305:17]
  wire [8:0] write_set = io_update_pc[9:1]; // @[FrontendBundle.scala 389:65]
  wire [8:0] touch_set_0 = io_update_write_data_valid ? write_set : req_idx; // @[FTB.scala 356:24]
  wire  touch_way_0_valid = io_update_write_data_valid | hit; // @[FTB.scala 358:43]
  reg  allocWriteWay_REG_3; // @[FTB.scala 386:41]
  reg  allocWriteWay_REG_2; // @[FTB.scala 386:41]
  reg  allocWriteWay_REG_1; // @[FTB.scala 386:41]
  reg  allocWriteWay_REG_0; // @[FTB.scala 386:41]
  wire [3:0] _allocWriteWay_T = {allocWriteWay_REG_3,allocWriteWay_REG_2,allocWriteWay_REG_1,allocWriteWay_REG_0}; // @[FTB.scala 386:79]
  wire  allocWriteWay_valid = &_allocWriteWay_T; // @[FTB.scala 366:37]
  wire [2:0] _GEN_596 = 9'h1 == write_set ? state_vec_1 : state_vec_0; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_597 = 9'h2 == write_set ? state_vec_2 : _GEN_596; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_598 = 9'h3 == write_set ? state_vec_3 : _GEN_597; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_599 = 9'h4 == write_set ? state_vec_4 : _GEN_598; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_600 = 9'h5 == write_set ? state_vec_5 : _GEN_599; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_601 = 9'h6 == write_set ? state_vec_6 : _GEN_600; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_602 = 9'h7 == write_set ? state_vec_7 : _GEN_601; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_603 = 9'h8 == write_set ? state_vec_8 : _GEN_602; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_604 = 9'h9 == write_set ? state_vec_9 : _GEN_603; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_605 = 9'ha == write_set ? state_vec_10 : _GEN_604; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_606 = 9'hb == write_set ? state_vec_11 : _GEN_605; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_607 = 9'hc == write_set ? state_vec_12 : _GEN_606; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_608 = 9'hd == write_set ? state_vec_13 : _GEN_607; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_609 = 9'he == write_set ? state_vec_14 : _GEN_608; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_610 = 9'hf == write_set ? state_vec_15 : _GEN_609; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_611 = 9'h10 == write_set ? state_vec_16 : _GEN_610; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_612 = 9'h11 == write_set ? state_vec_17 : _GEN_611; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_613 = 9'h12 == write_set ? state_vec_18 : _GEN_612; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_614 = 9'h13 == write_set ? state_vec_19 : _GEN_613; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_615 = 9'h14 == write_set ? state_vec_20 : _GEN_614; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_616 = 9'h15 == write_set ? state_vec_21 : _GEN_615; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_617 = 9'h16 == write_set ? state_vec_22 : _GEN_616; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_618 = 9'h17 == write_set ? state_vec_23 : _GEN_617; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_619 = 9'h18 == write_set ? state_vec_24 : _GEN_618; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_620 = 9'h19 == write_set ? state_vec_25 : _GEN_619; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_621 = 9'h1a == write_set ? state_vec_26 : _GEN_620; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_622 = 9'h1b == write_set ? state_vec_27 : _GEN_621; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_623 = 9'h1c == write_set ? state_vec_28 : _GEN_622; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_624 = 9'h1d == write_set ? state_vec_29 : _GEN_623; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_625 = 9'h1e == write_set ? state_vec_30 : _GEN_624; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_626 = 9'h1f == write_set ? state_vec_31 : _GEN_625; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_627 = 9'h20 == write_set ? state_vec_32 : _GEN_626; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_628 = 9'h21 == write_set ? state_vec_33 : _GEN_627; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_629 = 9'h22 == write_set ? state_vec_34 : _GEN_628; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_630 = 9'h23 == write_set ? state_vec_35 : _GEN_629; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_631 = 9'h24 == write_set ? state_vec_36 : _GEN_630; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_632 = 9'h25 == write_set ? state_vec_37 : _GEN_631; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_633 = 9'h26 == write_set ? state_vec_38 : _GEN_632; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_634 = 9'h27 == write_set ? state_vec_39 : _GEN_633; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_635 = 9'h28 == write_set ? state_vec_40 : _GEN_634; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_636 = 9'h29 == write_set ? state_vec_41 : _GEN_635; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_637 = 9'h2a == write_set ? state_vec_42 : _GEN_636; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_638 = 9'h2b == write_set ? state_vec_43 : _GEN_637; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_639 = 9'h2c == write_set ? state_vec_44 : _GEN_638; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_640 = 9'h2d == write_set ? state_vec_45 : _GEN_639; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_641 = 9'h2e == write_set ? state_vec_46 : _GEN_640; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_642 = 9'h2f == write_set ? state_vec_47 : _GEN_641; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_643 = 9'h30 == write_set ? state_vec_48 : _GEN_642; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_644 = 9'h31 == write_set ? state_vec_49 : _GEN_643; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_645 = 9'h32 == write_set ? state_vec_50 : _GEN_644; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_646 = 9'h33 == write_set ? state_vec_51 : _GEN_645; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_647 = 9'h34 == write_set ? state_vec_52 : _GEN_646; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_648 = 9'h35 == write_set ? state_vec_53 : _GEN_647; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_649 = 9'h36 == write_set ? state_vec_54 : _GEN_648; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_650 = 9'h37 == write_set ? state_vec_55 : _GEN_649; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_651 = 9'h38 == write_set ? state_vec_56 : _GEN_650; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_652 = 9'h39 == write_set ? state_vec_57 : _GEN_651; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_653 = 9'h3a == write_set ? state_vec_58 : _GEN_652; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_654 = 9'h3b == write_set ? state_vec_59 : _GEN_653; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_655 = 9'h3c == write_set ? state_vec_60 : _GEN_654; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_656 = 9'h3d == write_set ? state_vec_61 : _GEN_655; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_657 = 9'h3e == write_set ? state_vec_62 : _GEN_656; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_658 = 9'h3f == write_set ? state_vec_63 : _GEN_657; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_659 = 9'h40 == write_set ? state_vec_64 : _GEN_658; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_660 = 9'h41 == write_set ? state_vec_65 : _GEN_659; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_661 = 9'h42 == write_set ? state_vec_66 : _GEN_660; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_662 = 9'h43 == write_set ? state_vec_67 : _GEN_661; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_663 = 9'h44 == write_set ? state_vec_68 : _GEN_662; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_664 = 9'h45 == write_set ? state_vec_69 : _GEN_663; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_665 = 9'h46 == write_set ? state_vec_70 : _GEN_664; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_666 = 9'h47 == write_set ? state_vec_71 : _GEN_665; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_667 = 9'h48 == write_set ? state_vec_72 : _GEN_666; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_668 = 9'h49 == write_set ? state_vec_73 : _GEN_667; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_669 = 9'h4a == write_set ? state_vec_74 : _GEN_668; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_670 = 9'h4b == write_set ? state_vec_75 : _GEN_669; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_671 = 9'h4c == write_set ? state_vec_76 : _GEN_670; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_672 = 9'h4d == write_set ? state_vec_77 : _GEN_671; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_673 = 9'h4e == write_set ? state_vec_78 : _GEN_672; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_674 = 9'h4f == write_set ? state_vec_79 : _GEN_673; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_675 = 9'h50 == write_set ? state_vec_80 : _GEN_674; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_676 = 9'h51 == write_set ? state_vec_81 : _GEN_675; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_677 = 9'h52 == write_set ? state_vec_82 : _GEN_676; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_678 = 9'h53 == write_set ? state_vec_83 : _GEN_677; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_679 = 9'h54 == write_set ? state_vec_84 : _GEN_678; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_680 = 9'h55 == write_set ? state_vec_85 : _GEN_679; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_681 = 9'h56 == write_set ? state_vec_86 : _GEN_680; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_682 = 9'h57 == write_set ? state_vec_87 : _GEN_681; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_683 = 9'h58 == write_set ? state_vec_88 : _GEN_682; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_684 = 9'h59 == write_set ? state_vec_89 : _GEN_683; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_685 = 9'h5a == write_set ? state_vec_90 : _GEN_684; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_686 = 9'h5b == write_set ? state_vec_91 : _GEN_685; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_687 = 9'h5c == write_set ? state_vec_92 : _GEN_686; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_688 = 9'h5d == write_set ? state_vec_93 : _GEN_687; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_689 = 9'h5e == write_set ? state_vec_94 : _GEN_688; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_690 = 9'h5f == write_set ? state_vec_95 : _GEN_689; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_691 = 9'h60 == write_set ? state_vec_96 : _GEN_690; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_692 = 9'h61 == write_set ? state_vec_97 : _GEN_691; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_693 = 9'h62 == write_set ? state_vec_98 : _GEN_692; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_694 = 9'h63 == write_set ? state_vec_99 : _GEN_693; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_695 = 9'h64 == write_set ? state_vec_100 : _GEN_694; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_696 = 9'h65 == write_set ? state_vec_101 : _GEN_695; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_697 = 9'h66 == write_set ? state_vec_102 : _GEN_696; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_698 = 9'h67 == write_set ? state_vec_103 : _GEN_697; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_699 = 9'h68 == write_set ? state_vec_104 : _GEN_698; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_700 = 9'h69 == write_set ? state_vec_105 : _GEN_699; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_701 = 9'h6a == write_set ? state_vec_106 : _GEN_700; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_702 = 9'h6b == write_set ? state_vec_107 : _GEN_701; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_703 = 9'h6c == write_set ? state_vec_108 : _GEN_702; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_704 = 9'h6d == write_set ? state_vec_109 : _GEN_703; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_705 = 9'h6e == write_set ? state_vec_110 : _GEN_704; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_706 = 9'h6f == write_set ? state_vec_111 : _GEN_705; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_707 = 9'h70 == write_set ? state_vec_112 : _GEN_706; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_708 = 9'h71 == write_set ? state_vec_113 : _GEN_707; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_709 = 9'h72 == write_set ? state_vec_114 : _GEN_708; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_710 = 9'h73 == write_set ? state_vec_115 : _GEN_709; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_711 = 9'h74 == write_set ? state_vec_116 : _GEN_710; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_712 = 9'h75 == write_set ? state_vec_117 : _GEN_711; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_713 = 9'h76 == write_set ? state_vec_118 : _GEN_712; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_714 = 9'h77 == write_set ? state_vec_119 : _GEN_713; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_715 = 9'h78 == write_set ? state_vec_120 : _GEN_714; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_716 = 9'h79 == write_set ? state_vec_121 : _GEN_715; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_717 = 9'h7a == write_set ? state_vec_122 : _GEN_716; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_718 = 9'h7b == write_set ? state_vec_123 : _GEN_717; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_719 = 9'h7c == write_set ? state_vec_124 : _GEN_718; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_720 = 9'h7d == write_set ? state_vec_125 : _GEN_719; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_721 = 9'h7e == write_set ? state_vec_126 : _GEN_720; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_722 = 9'h7f == write_set ? state_vec_127 : _GEN_721; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_723 = 9'h80 == write_set ? state_vec_128 : _GEN_722; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_724 = 9'h81 == write_set ? state_vec_129 : _GEN_723; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_725 = 9'h82 == write_set ? state_vec_130 : _GEN_724; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_726 = 9'h83 == write_set ? state_vec_131 : _GEN_725; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_727 = 9'h84 == write_set ? state_vec_132 : _GEN_726; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_728 = 9'h85 == write_set ? state_vec_133 : _GEN_727; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_729 = 9'h86 == write_set ? state_vec_134 : _GEN_728; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_730 = 9'h87 == write_set ? state_vec_135 : _GEN_729; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_731 = 9'h88 == write_set ? state_vec_136 : _GEN_730; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_732 = 9'h89 == write_set ? state_vec_137 : _GEN_731; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_733 = 9'h8a == write_set ? state_vec_138 : _GEN_732; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_734 = 9'h8b == write_set ? state_vec_139 : _GEN_733; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_735 = 9'h8c == write_set ? state_vec_140 : _GEN_734; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_736 = 9'h8d == write_set ? state_vec_141 : _GEN_735; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_737 = 9'h8e == write_set ? state_vec_142 : _GEN_736; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_738 = 9'h8f == write_set ? state_vec_143 : _GEN_737; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_739 = 9'h90 == write_set ? state_vec_144 : _GEN_738; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_740 = 9'h91 == write_set ? state_vec_145 : _GEN_739; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_741 = 9'h92 == write_set ? state_vec_146 : _GEN_740; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_742 = 9'h93 == write_set ? state_vec_147 : _GEN_741; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_743 = 9'h94 == write_set ? state_vec_148 : _GEN_742; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_744 = 9'h95 == write_set ? state_vec_149 : _GEN_743; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_745 = 9'h96 == write_set ? state_vec_150 : _GEN_744; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_746 = 9'h97 == write_set ? state_vec_151 : _GEN_745; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_747 = 9'h98 == write_set ? state_vec_152 : _GEN_746; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_748 = 9'h99 == write_set ? state_vec_153 : _GEN_747; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_749 = 9'h9a == write_set ? state_vec_154 : _GEN_748; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_750 = 9'h9b == write_set ? state_vec_155 : _GEN_749; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_751 = 9'h9c == write_set ? state_vec_156 : _GEN_750; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_752 = 9'h9d == write_set ? state_vec_157 : _GEN_751; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_753 = 9'h9e == write_set ? state_vec_158 : _GEN_752; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_754 = 9'h9f == write_set ? state_vec_159 : _GEN_753; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_755 = 9'ha0 == write_set ? state_vec_160 : _GEN_754; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_756 = 9'ha1 == write_set ? state_vec_161 : _GEN_755; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_757 = 9'ha2 == write_set ? state_vec_162 : _GEN_756; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_758 = 9'ha3 == write_set ? state_vec_163 : _GEN_757; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_759 = 9'ha4 == write_set ? state_vec_164 : _GEN_758; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_760 = 9'ha5 == write_set ? state_vec_165 : _GEN_759; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_761 = 9'ha6 == write_set ? state_vec_166 : _GEN_760; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_762 = 9'ha7 == write_set ? state_vec_167 : _GEN_761; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_763 = 9'ha8 == write_set ? state_vec_168 : _GEN_762; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_764 = 9'ha9 == write_set ? state_vec_169 : _GEN_763; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_765 = 9'haa == write_set ? state_vec_170 : _GEN_764; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_766 = 9'hab == write_set ? state_vec_171 : _GEN_765; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_767 = 9'hac == write_set ? state_vec_172 : _GEN_766; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_768 = 9'had == write_set ? state_vec_173 : _GEN_767; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_769 = 9'hae == write_set ? state_vec_174 : _GEN_768; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_770 = 9'haf == write_set ? state_vec_175 : _GEN_769; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_771 = 9'hb0 == write_set ? state_vec_176 : _GEN_770; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_772 = 9'hb1 == write_set ? state_vec_177 : _GEN_771; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_773 = 9'hb2 == write_set ? state_vec_178 : _GEN_772; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_774 = 9'hb3 == write_set ? state_vec_179 : _GEN_773; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_775 = 9'hb4 == write_set ? state_vec_180 : _GEN_774; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_776 = 9'hb5 == write_set ? state_vec_181 : _GEN_775; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_777 = 9'hb6 == write_set ? state_vec_182 : _GEN_776; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_778 = 9'hb7 == write_set ? state_vec_183 : _GEN_777; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_779 = 9'hb8 == write_set ? state_vec_184 : _GEN_778; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_780 = 9'hb9 == write_set ? state_vec_185 : _GEN_779; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_781 = 9'hba == write_set ? state_vec_186 : _GEN_780; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_782 = 9'hbb == write_set ? state_vec_187 : _GEN_781; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_783 = 9'hbc == write_set ? state_vec_188 : _GEN_782; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_784 = 9'hbd == write_set ? state_vec_189 : _GEN_783; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_785 = 9'hbe == write_set ? state_vec_190 : _GEN_784; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_786 = 9'hbf == write_set ? state_vec_191 : _GEN_785; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_787 = 9'hc0 == write_set ? state_vec_192 : _GEN_786; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_788 = 9'hc1 == write_set ? state_vec_193 : _GEN_787; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_789 = 9'hc2 == write_set ? state_vec_194 : _GEN_788; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_790 = 9'hc3 == write_set ? state_vec_195 : _GEN_789; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_791 = 9'hc4 == write_set ? state_vec_196 : _GEN_790; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_792 = 9'hc5 == write_set ? state_vec_197 : _GEN_791; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_793 = 9'hc6 == write_set ? state_vec_198 : _GEN_792; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_794 = 9'hc7 == write_set ? state_vec_199 : _GEN_793; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_795 = 9'hc8 == write_set ? state_vec_200 : _GEN_794; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_796 = 9'hc9 == write_set ? state_vec_201 : _GEN_795; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_797 = 9'hca == write_set ? state_vec_202 : _GEN_796; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_798 = 9'hcb == write_set ? state_vec_203 : _GEN_797; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_799 = 9'hcc == write_set ? state_vec_204 : _GEN_798; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_800 = 9'hcd == write_set ? state_vec_205 : _GEN_799; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_801 = 9'hce == write_set ? state_vec_206 : _GEN_800; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_802 = 9'hcf == write_set ? state_vec_207 : _GEN_801; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_803 = 9'hd0 == write_set ? state_vec_208 : _GEN_802; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_804 = 9'hd1 == write_set ? state_vec_209 : _GEN_803; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_805 = 9'hd2 == write_set ? state_vec_210 : _GEN_804; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_806 = 9'hd3 == write_set ? state_vec_211 : _GEN_805; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_807 = 9'hd4 == write_set ? state_vec_212 : _GEN_806; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_808 = 9'hd5 == write_set ? state_vec_213 : _GEN_807; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_809 = 9'hd6 == write_set ? state_vec_214 : _GEN_808; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_810 = 9'hd7 == write_set ? state_vec_215 : _GEN_809; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_811 = 9'hd8 == write_set ? state_vec_216 : _GEN_810; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_812 = 9'hd9 == write_set ? state_vec_217 : _GEN_811; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_813 = 9'hda == write_set ? state_vec_218 : _GEN_812; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_814 = 9'hdb == write_set ? state_vec_219 : _GEN_813; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_815 = 9'hdc == write_set ? state_vec_220 : _GEN_814; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_816 = 9'hdd == write_set ? state_vec_221 : _GEN_815; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_817 = 9'hde == write_set ? state_vec_222 : _GEN_816; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_818 = 9'hdf == write_set ? state_vec_223 : _GEN_817; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_819 = 9'he0 == write_set ? state_vec_224 : _GEN_818; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_820 = 9'he1 == write_set ? state_vec_225 : _GEN_819; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_821 = 9'he2 == write_set ? state_vec_226 : _GEN_820; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_822 = 9'he3 == write_set ? state_vec_227 : _GEN_821; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_823 = 9'he4 == write_set ? state_vec_228 : _GEN_822; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_824 = 9'he5 == write_set ? state_vec_229 : _GEN_823; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_825 = 9'he6 == write_set ? state_vec_230 : _GEN_824; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_826 = 9'he7 == write_set ? state_vec_231 : _GEN_825; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_827 = 9'he8 == write_set ? state_vec_232 : _GEN_826; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_828 = 9'he9 == write_set ? state_vec_233 : _GEN_827; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_829 = 9'hea == write_set ? state_vec_234 : _GEN_828; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_830 = 9'heb == write_set ? state_vec_235 : _GEN_829; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_831 = 9'hec == write_set ? state_vec_236 : _GEN_830; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_832 = 9'hed == write_set ? state_vec_237 : _GEN_831; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_833 = 9'hee == write_set ? state_vec_238 : _GEN_832; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_834 = 9'hef == write_set ? state_vec_239 : _GEN_833; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_835 = 9'hf0 == write_set ? state_vec_240 : _GEN_834; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_836 = 9'hf1 == write_set ? state_vec_241 : _GEN_835; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_837 = 9'hf2 == write_set ? state_vec_242 : _GEN_836; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_838 = 9'hf3 == write_set ? state_vec_243 : _GEN_837; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_839 = 9'hf4 == write_set ? state_vec_244 : _GEN_838; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_840 = 9'hf5 == write_set ? state_vec_245 : _GEN_839; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_841 = 9'hf6 == write_set ? state_vec_246 : _GEN_840; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_842 = 9'hf7 == write_set ? state_vec_247 : _GEN_841; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_843 = 9'hf8 == write_set ? state_vec_248 : _GEN_842; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_844 = 9'hf9 == write_set ? state_vec_249 : _GEN_843; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_845 = 9'hfa == write_set ? state_vec_250 : _GEN_844; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_846 = 9'hfb == write_set ? state_vec_251 : _GEN_845; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_847 = 9'hfc == write_set ? state_vec_252 : _GEN_846; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_848 = 9'hfd == write_set ? state_vec_253 : _GEN_847; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_849 = 9'hfe == write_set ? state_vec_254 : _GEN_848; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_850 = 9'hff == write_set ? state_vec_255 : _GEN_849; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_851 = 9'h100 == write_set ? state_vec_256 : _GEN_850; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_852 = 9'h101 == write_set ? state_vec_257 : _GEN_851; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_853 = 9'h102 == write_set ? state_vec_258 : _GEN_852; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_854 = 9'h103 == write_set ? state_vec_259 : _GEN_853; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_855 = 9'h104 == write_set ? state_vec_260 : _GEN_854; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_856 = 9'h105 == write_set ? state_vec_261 : _GEN_855; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_857 = 9'h106 == write_set ? state_vec_262 : _GEN_856; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_858 = 9'h107 == write_set ? state_vec_263 : _GEN_857; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_859 = 9'h108 == write_set ? state_vec_264 : _GEN_858; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_860 = 9'h109 == write_set ? state_vec_265 : _GEN_859; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_861 = 9'h10a == write_set ? state_vec_266 : _GEN_860; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_862 = 9'h10b == write_set ? state_vec_267 : _GEN_861; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_863 = 9'h10c == write_set ? state_vec_268 : _GEN_862; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_864 = 9'h10d == write_set ? state_vec_269 : _GEN_863; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_865 = 9'h10e == write_set ? state_vec_270 : _GEN_864; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_866 = 9'h10f == write_set ? state_vec_271 : _GEN_865; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_867 = 9'h110 == write_set ? state_vec_272 : _GEN_866; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_868 = 9'h111 == write_set ? state_vec_273 : _GEN_867; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_869 = 9'h112 == write_set ? state_vec_274 : _GEN_868; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_870 = 9'h113 == write_set ? state_vec_275 : _GEN_869; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_871 = 9'h114 == write_set ? state_vec_276 : _GEN_870; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_872 = 9'h115 == write_set ? state_vec_277 : _GEN_871; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_873 = 9'h116 == write_set ? state_vec_278 : _GEN_872; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_874 = 9'h117 == write_set ? state_vec_279 : _GEN_873; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_875 = 9'h118 == write_set ? state_vec_280 : _GEN_874; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_876 = 9'h119 == write_set ? state_vec_281 : _GEN_875; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_877 = 9'h11a == write_set ? state_vec_282 : _GEN_876; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_878 = 9'h11b == write_set ? state_vec_283 : _GEN_877; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_879 = 9'h11c == write_set ? state_vec_284 : _GEN_878; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_880 = 9'h11d == write_set ? state_vec_285 : _GEN_879; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_881 = 9'h11e == write_set ? state_vec_286 : _GEN_880; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_882 = 9'h11f == write_set ? state_vec_287 : _GEN_881; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_883 = 9'h120 == write_set ? state_vec_288 : _GEN_882; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_884 = 9'h121 == write_set ? state_vec_289 : _GEN_883; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_885 = 9'h122 == write_set ? state_vec_290 : _GEN_884; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_886 = 9'h123 == write_set ? state_vec_291 : _GEN_885; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_887 = 9'h124 == write_set ? state_vec_292 : _GEN_886; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_888 = 9'h125 == write_set ? state_vec_293 : _GEN_887; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_889 = 9'h126 == write_set ? state_vec_294 : _GEN_888; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_890 = 9'h127 == write_set ? state_vec_295 : _GEN_889; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_891 = 9'h128 == write_set ? state_vec_296 : _GEN_890; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_892 = 9'h129 == write_set ? state_vec_297 : _GEN_891; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_893 = 9'h12a == write_set ? state_vec_298 : _GEN_892; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_894 = 9'h12b == write_set ? state_vec_299 : _GEN_893; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_895 = 9'h12c == write_set ? state_vec_300 : _GEN_894; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_896 = 9'h12d == write_set ? state_vec_301 : _GEN_895; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_897 = 9'h12e == write_set ? state_vec_302 : _GEN_896; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_898 = 9'h12f == write_set ? state_vec_303 : _GEN_897; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_899 = 9'h130 == write_set ? state_vec_304 : _GEN_898; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_900 = 9'h131 == write_set ? state_vec_305 : _GEN_899; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_901 = 9'h132 == write_set ? state_vec_306 : _GEN_900; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_902 = 9'h133 == write_set ? state_vec_307 : _GEN_901; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_903 = 9'h134 == write_set ? state_vec_308 : _GEN_902; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_904 = 9'h135 == write_set ? state_vec_309 : _GEN_903; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_905 = 9'h136 == write_set ? state_vec_310 : _GEN_904; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_906 = 9'h137 == write_set ? state_vec_311 : _GEN_905; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_907 = 9'h138 == write_set ? state_vec_312 : _GEN_906; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_908 = 9'h139 == write_set ? state_vec_313 : _GEN_907; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_909 = 9'h13a == write_set ? state_vec_314 : _GEN_908; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_910 = 9'h13b == write_set ? state_vec_315 : _GEN_909; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_911 = 9'h13c == write_set ? state_vec_316 : _GEN_910; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_912 = 9'h13d == write_set ? state_vec_317 : _GEN_911; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_913 = 9'h13e == write_set ? state_vec_318 : _GEN_912; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_914 = 9'h13f == write_set ? state_vec_319 : _GEN_913; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_915 = 9'h140 == write_set ? state_vec_320 : _GEN_914; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_916 = 9'h141 == write_set ? state_vec_321 : _GEN_915; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_917 = 9'h142 == write_set ? state_vec_322 : _GEN_916; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_918 = 9'h143 == write_set ? state_vec_323 : _GEN_917; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_919 = 9'h144 == write_set ? state_vec_324 : _GEN_918; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_920 = 9'h145 == write_set ? state_vec_325 : _GEN_919; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_921 = 9'h146 == write_set ? state_vec_326 : _GEN_920; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_922 = 9'h147 == write_set ? state_vec_327 : _GEN_921; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_923 = 9'h148 == write_set ? state_vec_328 : _GEN_922; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_924 = 9'h149 == write_set ? state_vec_329 : _GEN_923; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_925 = 9'h14a == write_set ? state_vec_330 : _GEN_924; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_926 = 9'h14b == write_set ? state_vec_331 : _GEN_925; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_927 = 9'h14c == write_set ? state_vec_332 : _GEN_926; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_928 = 9'h14d == write_set ? state_vec_333 : _GEN_927; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_929 = 9'h14e == write_set ? state_vec_334 : _GEN_928; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_930 = 9'h14f == write_set ? state_vec_335 : _GEN_929; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_931 = 9'h150 == write_set ? state_vec_336 : _GEN_930; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_932 = 9'h151 == write_set ? state_vec_337 : _GEN_931; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_933 = 9'h152 == write_set ? state_vec_338 : _GEN_932; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_934 = 9'h153 == write_set ? state_vec_339 : _GEN_933; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_935 = 9'h154 == write_set ? state_vec_340 : _GEN_934; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_936 = 9'h155 == write_set ? state_vec_341 : _GEN_935; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_937 = 9'h156 == write_set ? state_vec_342 : _GEN_936; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_938 = 9'h157 == write_set ? state_vec_343 : _GEN_937; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_939 = 9'h158 == write_set ? state_vec_344 : _GEN_938; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_940 = 9'h159 == write_set ? state_vec_345 : _GEN_939; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_941 = 9'h15a == write_set ? state_vec_346 : _GEN_940; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_942 = 9'h15b == write_set ? state_vec_347 : _GEN_941; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_943 = 9'h15c == write_set ? state_vec_348 : _GEN_942; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_944 = 9'h15d == write_set ? state_vec_349 : _GEN_943; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_945 = 9'h15e == write_set ? state_vec_350 : _GEN_944; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_946 = 9'h15f == write_set ? state_vec_351 : _GEN_945; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_947 = 9'h160 == write_set ? state_vec_352 : _GEN_946; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_948 = 9'h161 == write_set ? state_vec_353 : _GEN_947; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_949 = 9'h162 == write_set ? state_vec_354 : _GEN_948; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_950 = 9'h163 == write_set ? state_vec_355 : _GEN_949; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_951 = 9'h164 == write_set ? state_vec_356 : _GEN_950; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_952 = 9'h165 == write_set ? state_vec_357 : _GEN_951; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_953 = 9'h166 == write_set ? state_vec_358 : _GEN_952; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_954 = 9'h167 == write_set ? state_vec_359 : _GEN_953; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_955 = 9'h168 == write_set ? state_vec_360 : _GEN_954; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_956 = 9'h169 == write_set ? state_vec_361 : _GEN_955; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_957 = 9'h16a == write_set ? state_vec_362 : _GEN_956; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_958 = 9'h16b == write_set ? state_vec_363 : _GEN_957; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_959 = 9'h16c == write_set ? state_vec_364 : _GEN_958; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_960 = 9'h16d == write_set ? state_vec_365 : _GEN_959; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_961 = 9'h16e == write_set ? state_vec_366 : _GEN_960; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_962 = 9'h16f == write_set ? state_vec_367 : _GEN_961; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_963 = 9'h170 == write_set ? state_vec_368 : _GEN_962; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_964 = 9'h171 == write_set ? state_vec_369 : _GEN_963; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_965 = 9'h172 == write_set ? state_vec_370 : _GEN_964; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_966 = 9'h173 == write_set ? state_vec_371 : _GEN_965; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_967 = 9'h174 == write_set ? state_vec_372 : _GEN_966; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_968 = 9'h175 == write_set ? state_vec_373 : _GEN_967; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_969 = 9'h176 == write_set ? state_vec_374 : _GEN_968; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_970 = 9'h177 == write_set ? state_vec_375 : _GEN_969; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_971 = 9'h178 == write_set ? state_vec_376 : _GEN_970; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_972 = 9'h179 == write_set ? state_vec_377 : _GEN_971; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_973 = 9'h17a == write_set ? state_vec_378 : _GEN_972; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_974 = 9'h17b == write_set ? state_vec_379 : _GEN_973; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_975 = 9'h17c == write_set ? state_vec_380 : _GEN_974; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_976 = 9'h17d == write_set ? state_vec_381 : _GEN_975; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_977 = 9'h17e == write_set ? state_vec_382 : _GEN_976; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_978 = 9'h17f == write_set ? state_vec_383 : _GEN_977; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_979 = 9'h180 == write_set ? state_vec_384 : _GEN_978; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_980 = 9'h181 == write_set ? state_vec_385 : _GEN_979; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_981 = 9'h182 == write_set ? state_vec_386 : _GEN_980; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_982 = 9'h183 == write_set ? state_vec_387 : _GEN_981; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_983 = 9'h184 == write_set ? state_vec_388 : _GEN_982; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_984 = 9'h185 == write_set ? state_vec_389 : _GEN_983; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_985 = 9'h186 == write_set ? state_vec_390 : _GEN_984; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_986 = 9'h187 == write_set ? state_vec_391 : _GEN_985; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_987 = 9'h188 == write_set ? state_vec_392 : _GEN_986; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_988 = 9'h189 == write_set ? state_vec_393 : _GEN_987; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_989 = 9'h18a == write_set ? state_vec_394 : _GEN_988; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_990 = 9'h18b == write_set ? state_vec_395 : _GEN_989; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_991 = 9'h18c == write_set ? state_vec_396 : _GEN_990; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_992 = 9'h18d == write_set ? state_vec_397 : _GEN_991; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_993 = 9'h18e == write_set ? state_vec_398 : _GEN_992; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_994 = 9'h18f == write_set ? state_vec_399 : _GEN_993; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_995 = 9'h190 == write_set ? state_vec_400 : _GEN_994; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_996 = 9'h191 == write_set ? state_vec_401 : _GEN_995; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_997 = 9'h192 == write_set ? state_vec_402 : _GEN_996; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_998 = 9'h193 == write_set ? state_vec_403 : _GEN_997; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_999 = 9'h194 == write_set ? state_vec_404 : _GEN_998; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1000 = 9'h195 == write_set ? state_vec_405 : _GEN_999; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1001 = 9'h196 == write_set ? state_vec_406 : _GEN_1000; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1002 = 9'h197 == write_set ? state_vec_407 : _GEN_1001; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1003 = 9'h198 == write_set ? state_vec_408 : _GEN_1002; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1004 = 9'h199 == write_set ? state_vec_409 : _GEN_1003; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1005 = 9'h19a == write_set ? state_vec_410 : _GEN_1004; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1006 = 9'h19b == write_set ? state_vec_411 : _GEN_1005; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1007 = 9'h19c == write_set ? state_vec_412 : _GEN_1006; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1008 = 9'h19d == write_set ? state_vec_413 : _GEN_1007; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1009 = 9'h19e == write_set ? state_vec_414 : _GEN_1008; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1010 = 9'h19f == write_set ? state_vec_415 : _GEN_1009; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1011 = 9'h1a0 == write_set ? state_vec_416 : _GEN_1010; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1012 = 9'h1a1 == write_set ? state_vec_417 : _GEN_1011; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1013 = 9'h1a2 == write_set ? state_vec_418 : _GEN_1012; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1014 = 9'h1a3 == write_set ? state_vec_419 : _GEN_1013; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1015 = 9'h1a4 == write_set ? state_vec_420 : _GEN_1014; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1016 = 9'h1a5 == write_set ? state_vec_421 : _GEN_1015; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1017 = 9'h1a6 == write_set ? state_vec_422 : _GEN_1016; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1018 = 9'h1a7 == write_set ? state_vec_423 : _GEN_1017; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1019 = 9'h1a8 == write_set ? state_vec_424 : _GEN_1018; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1020 = 9'h1a9 == write_set ? state_vec_425 : _GEN_1019; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1021 = 9'h1aa == write_set ? state_vec_426 : _GEN_1020; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1022 = 9'h1ab == write_set ? state_vec_427 : _GEN_1021; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1023 = 9'h1ac == write_set ? state_vec_428 : _GEN_1022; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1024 = 9'h1ad == write_set ? state_vec_429 : _GEN_1023; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1025 = 9'h1ae == write_set ? state_vec_430 : _GEN_1024; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1026 = 9'h1af == write_set ? state_vec_431 : _GEN_1025; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1027 = 9'h1b0 == write_set ? state_vec_432 : _GEN_1026; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1028 = 9'h1b1 == write_set ? state_vec_433 : _GEN_1027; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1029 = 9'h1b2 == write_set ? state_vec_434 : _GEN_1028; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1030 = 9'h1b3 == write_set ? state_vec_435 : _GEN_1029; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1031 = 9'h1b4 == write_set ? state_vec_436 : _GEN_1030; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1032 = 9'h1b5 == write_set ? state_vec_437 : _GEN_1031; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1033 = 9'h1b6 == write_set ? state_vec_438 : _GEN_1032; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1034 = 9'h1b7 == write_set ? state_vec_439 : _GEN_1033; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1035 = 9'h1b8 == write_set ? state_vec_440 : _GEN_1034; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1036 = 9'h1b9 == write_set ? state_vec_441 : _GEN_1035; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1037 = 9'h1ba == write_set ? state_vec_442 : _GEN_1036; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1038 = 9'h1bb == write_set ? state_vec_443 : _GEN_1037; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1039 = 9'h1bc == write_set ? state_vec_444 : _GEN_1038; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1040 = 9'h1bd == write_set ? state_vec_445 : _GEN_1039; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1041 = 9'h1be == write_set ? state_vec_446 : _GEN_1040; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1042 = 9'h1bf == write_set ? state_vec_447 : _GEN_1041; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1043 = 9'h1c0 == write_set ? state_vec_448 : _GEN_1042; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1044 = 9'h1c1 == write_set ? state_vec_449 : _GEN_1043; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1045 = 9'h1c2 == write_set ? state_vec_450 : _GEN_1044; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1046 = 9'h1c3 == write_set ? state_vec_451 : _GEN_1045; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1047 = 9'h1c4 == write_set ? state_vec_452 : _GEN_1046; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1048 = 9'h1c5 == write_set ? state_vec_453 : _GEN_1047; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1049 = 9'h1c6 == write_set ? state_vec_454 : _GEN_1048; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1050 = 9'h1c7 == write_set ? state_vec_455 : _GEN_1049; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1051 = 9'h1c8 == write_set ? state_vec_456 : _GEN_1050; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1052 = 9'h1c9 == write_set ? state_vec_457 : _GEN_1051; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1053 = 9'h1ca == write_set ? state_vec_458 : _GEN_1052; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1054 = 9'h1cb == write_set ? state_vec_459 : _GEN_1053; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1055 = 9'h1cc == write_set ? state_vec_460 : _GEN_1054; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1056 = 9'h1cd == write_set ? state_vec_461 : _GEN_1055; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1057 = 9'h1ce == write_set ? state_vec_462 : _GEN_1056; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1058 = 9'h1cf == write_set ? state_vec_463 : _GEN_1057; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1059 = 9'h1d0 == write_set ? state_vec_464 : _GEN_1058; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1060 = 9'h1d1 == write_set ? state_vec_465 : _GEN_1059; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1061 = 9'h1d2 == write_set ? state_vec_466 : _GEN_1060; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1062 = 9'h1d3 == write_set ? state_vec_467 : _GEN_1061; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1063 = 9'h1d4 == write_set ? state_vec_468 : _GEN_1062; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1064 = 9'h1d5 == write_set ? state_vec_469 : _GEN_1063; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1065 = 9'h1d6 == write_set ? state_vec_470 : _GEN_1064; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1066 = 9'h1d7 == write_set ? state_vec_471 : _GEN_1065; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1067 = 9'h1d8 == write_set ? state_vec_472 : _GEN_1066; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1068 = 9'h1d9 == write_set ? state_vec_473 : _GEN_1067; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1069 = 9'h1da == write_set ? state_vec_474 : _GEN_1068; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1070 = 9'h1db == write_set ? state_vec_475 : _GEN_1069; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1071 = 9'h1dc == write_set ? state_vec_476 : _GEN_1070; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1072 = 9'h1dd == write_set ? state_vec_477 : _GEN_1071; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1073 = 9'h1de == write_set ? state_vec_478 : _GEN_1072; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1074 = 9'h1df == write_set ? state_vec_479 : _GEN_1073; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1075 = 9'h1e0 == write_set ? state_vec_480 : _GEN_1074; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1076 = 9'h1e1 == write_set ? state_vec_481 : _GEN_1075; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1077 = 9'h1e2 == write_set ? state_vec_482 : _GEN_1076; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1078 = 9'h1e3 == write_set ? state_vec_483 : _GEN_1077; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1079 = 9'h1e4 == write_set ? state_vec_484 : _GEN_1078; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1080 = 9'h1e5 == write_set ? state_vec_485 : _GEN_1079; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1081 = 9'h1e6 == write_set ? state_vec_486 : _GEN_1080; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1082 = 9'h1e7 == write_set ? state_vec_487 : _GEN_1081; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1083 = 9'h1e8 == write_set ? state_vec_488 : _GEN_1082; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1084 = 9'h1e9 == write_set ? state_vec_489 : _GEN_1083; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1085 = 9'h1ea == write_set ? state_vec_490 : _GEN_1084; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1086 = 9'h1eb == write_set ? state_vec_491 : _GEN_1085; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1087 = 9'h1ec == write_set ? state_vec_492 : _GEN_1086; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1088 = 9'h1ed == write_set ? state_vec_493 : _GEN_1087; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1089 = 9'h1ee == write_set ? state_vec_494 : _GEN_1088; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1090 = 9'h1ef == write_set ? state_vec_495 : _GEN_1089; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1091 = 9'h1f0 == write_set ? state_vec_496 : _GEN_1090; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1092 = 9'h1f1 == write_set ? state_vec_497 : _GEN_1091; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1093 = 9'h1f2 == write_set ? state_vec_498 : _GEN_1092; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1094 = 9'h1f3 == write_set ? state_vec_499 : _GEN_1093; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1095 = 9'h1f4 == write_set ? state_vec_500 : _GEN_1094; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1096 = 9'h1f5 == write_set ? state_vec_501 : _GEN_1095; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1097 = 9'h1f6 == write_set ? state_vec_502 : _GEN_1096; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1098 = 9'h1f7 == write_set ? state_vec_503 : _GEN_1097; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1099 = 9'h1f8 == write_set ? state_vec_504 : _GEN_1098; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1100 = 9'h1f9 == write_set ? state_vec_505 : _GEN_1099; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1101 = 9'h1fa == write_set ? state_vec_506 : _GEN_1100; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1102 = 9'h1fb == write_set ? state_vec_507 : _GEN_1101; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1103 = 9'h1fc == write_set ? state_vec_508 : _GEN_1102; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1104 = 9'h1fd == write_set ? state_vec_509 : _GEN_1103; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1105 = 9'h1fe == write_set ? state_vec_510 : _GEN_1104; // @[Replacement.scala 243:{38,38}]
  wire [2:0] _GEN_1106 = 9'h1ff == write_set ? state_vec_511 : _GEN_1105; // @[Replacement.scala 243:{38,38}]
  wire  allocWriteWay_wleft_subtree_older = _GEN_1106[2]; // @[Replacement.scala 243:38]
  wire  allocWriteWay_wleft_subtree_state = _GEN_1106[1]; // @[package.scala 154:13]
  wire  allocWriteWay_wright_subtree_state = _GEN_1106[0]; // @[Replacement.scala 245:38]
  wire  _allocWriteWay_wT_2 = allocWriteWay_wleft_subtree_older ? allocWriteWay_wleft_subtree_state :
    allocWriteWay_wright_subtree_state; // @[Replacement.scala 250:16]
  wire [1:0] _allocWriteWay_wT_3 = {allocWriteWay_wleft_subtree_older,_allocWriteWay_wT_2}; // @[Cat.scala 31:58]
  wire [3:0] _allocWriteWay_wT_4 = ~_allocWriteWay_T; // @[FTB.scala 367:60]
  wire [1:0] _allocWriteWay_wT_9 = _allocWriteWay_wT_4[2] ? 2'h2 : 2'h3; // @[Mux.scala 47:70]
  wire [1:0] _allocWriteWay_wT_10 = _allocWriteWay_wT_4[1] ? 2'h1 : _allocWriteWay_wT_9; // @[Mux.scala 47:70]
  wire [1:0] _allocWriteWay_wT_11 = _allocWriteWay_wT_4[0] ? 2'h0 : _allocWriteWay_wT_10; // @[Mux.scala 47:70]
  wire [1:0] allocWriteWay = allocWriteWay_valid ? _allocWriteWay_wT_3 : _allocWriteWay_wT_11; // @[FTB.scala 367:17]
  wire [1:0] write_way_bits = io_update_write_alloc ? allocWriteWay : io_update_write_way; // @[FTB.scala 401:26]
  wire [1:0] touch_way_0_bits = io_update_write_data_valid ? write_way_bits : hit_way; // @[FTB.scala 359:29]
  wire  set_touch_ways_0_valid = touch_way_0_valid & touch_set_0 == 9'h0; // @[Replacement.scala 315:30]
  wire  state_vec_0_set_left_older = ~touch_way_0_bits[1]; // @[Replacement.scala 196:33]
  wire  state_vec_0_left_subtree_state = state_vec_0[1]; // @[package.scala 154:13]
  wire  state_vec_0_right_subtree_state = state_vec_0[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_0_T_2 = ~touch_way_0_bits[0]; // @[Replacement.scala 218:7]
  wire  _state_vec_0_T_3 = state_vec_0_set_left_older ? state_vec_0_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_0_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_0_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_0_T_8 = {state_vec_0_set_left_older,_state_vec_0_T_3,_state_vec_0_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_1_valid = touch_way_0_valid & touch_set_0 == 9'h1; // @[Replacement.scala 315:30]
  wire  state_vec_1_left_subtree_state = state_vec_1[1]; // @[package.scala 154:13]
  wire  state_vec_1_right_subtree_state = state_vec_1[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_1_T_3 = state_vec_0_set_left_older ? state_vec_1_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_1_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_1_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_1_T_8 = {state_vec_0_set_left_older,_state_vec_1_T_3,_state_vec_1_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_2_valid = touch_way_0_valid & touch_set_0 == 9'h2; // @[Replacement.scala 315:30]
  wire  state_vec_2_left_subtree_state = state_vec_2[1]; // @[package.scala 154:13]
  wire  state_vec_2_right_subtree_state = state_vec_2[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_2_T_3 = state_vec_0_set_left_older ? state_vec_2_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_2_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_2_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_2_T_8 = {state_vec_0_set_left_older,_state_vec_2_T_3,_state_vec_2_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_3_valid = touch_way_0_valid & touch_set_0 == 9'h3; // @[Replacement.scala 315:30]
  wire  state_vec_3_left_subtree_state = state_vec_3[1]; // @[package.scala 154:13]
  wire  state_vec_3_right_subtree_state = state_vec_3[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_3_T_3 = state_vec_0_set_left_older ? state_vec_3_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_3_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_3_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_3_T_8 = {state_vec_0_set_left_older,_state_vec_3_T_3,_state_vec_3_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_4_valid = touch_way_0_valid & touch_set_0 == 9'h4; // @[Replacement.scala 315:30]
  wire  state_vec_4_left_subtree_state = state_vec_4[1]; // @[package.scala 154:13]
  wire  state_vec_4_right_subtree_state = state_vec_4[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_4_T_3 = state_vec_0_set_left_older ? state_vec_4_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_4_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_4_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_4_T_8 = {state_vec_0_set_left_older,_state_vec_4_T_3,_state_vec_4_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_5_valid = touch_way_0_valid & touch_set_0 == 9'h5; // @[Replacement.scala 315:30]
  wire  state_vec_5_left_subtree_state = state_vec_5[1]; // @[package.scala 154:13]
  wire  state_vec_5_right_subtree_state = state_vec_5[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_5_T_3 = state_vec_0_set_left_older ? state_vec_5_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_5_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_5_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_5_T_8 = {state_vec_0_set_left_older,_state_vec_5_T_3,_state_vec_5_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_6_valid = touch_way_0_valid & touch_set_0 == 9'h6; // @[Replacement.scala 315:30]
  wire  state_vec_6_left_subtree_state = state_vec_6[1]; // @[package.scala 154:13]
  wire  state_vec_6_right_subtree_state = state_vec_6[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_6_T_3 = state_vec_0_set_left_older ? state_vec_6_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_6_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_6_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_6_T_8 = {state_vec_0_set_left_older,_state_vec_6_T_3,_state_vec_6_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_7_valid = touch_way_0_valid & touch_set_0 == 9'h7; // @[Replacement.scala 315:30]
  wire  state_vec_7_left_subtree_state = state_vec_7[1]; // @[package.scala 154:13]
  wire  state_vec_7_right_subtree_state = state_vec_7[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_7_T_3 = state_vec_0_set_left_older ? state_vec_7_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_7_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_7_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_7_T_8 = {state_vec_0_set_left_older,_state_vec_7_T_3,_state_vec_7_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_8_valid = touch_way_0_valid & touch_set_0 == 9'h8; // @[Replacement.scala 315:30]
  wire  state_vec_8_left_subtree_state = state_vec_8[1]; // @[package.scala 154:13]
  wire  state_vec_8_right_subtree_state = state_vec_8[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_8_T_3 = state_vec_0_set_left_older ? state_vec_8_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_8_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_8_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_8_T_8 = {state_vec_0_set_left_older,_state_vec_8_T_3,_state_vec_8_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_9_valid = touch_way_0_valid & touch_set_0 == 9'h9; // @[Replacement.scala 315:30]
  wire  state_vec_9_left_subtree_state = state_vec_9[1]; // @[package.scala 154:13]
  wire  state_vec_9_right_subtree_state = state_vec_9[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_9_T_3 = state_vec_0_set_left_older ? state_vec_9_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_9_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_9_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_9_T_8 = {state_vec_0_set_left_older,_state_vec_9_T_3,_state_vec_9_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_10_valid = touch_way_0_valid & touch_set_0 == 9'ha; // @[Replacement.scala 315:30]
  wire  state_vec_10_left_subtree_state = state_vec_10[1]; // @[package.scala 154:13]
  wire  state_vec_10_right_subtree_state = state_vec_10[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_10_T_3 = state_vec_0_set_left_older ? state_vec_10_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_10_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_10_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_10_T_8 = {state_vec_0_set_left_older,_state_vec_10_T_3,_state_vec_10_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_11_valid = touch_way_0_valid & touch_set_0 == 9'hb; // @[Replacement.scala 315:30]
  wire  state_vec_11_left_subtree_state = state_vec_11[1]; // @[package.scala 154:13]
  wire  state_vec_11_right_subtree_state = state_vec_11[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_11_T_3 = state_vec_0_set_left_older ? state_vec_11_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_11_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_11_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_11_T_8 = {state_vec_0_set_left_older,_state_vec_11_T_3,_state_vec_11_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_12_valid = touch_way_0_valid & touch_set_0 == 9'hc; // @[Replacement.scala 315:30]
  wire  state_vec_12_left_subtree_state = state_vec_12[1]; // @[package.scala 154:13]
  wire  state_vec_12_right_subtree_state = state_vec_12[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_12_T_3 = state_vec_0_set_left_older ? state_vec_12_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_12_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_12_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_12_T_8 = {state_vec_0_set_left_older,_state_vec_12_T_3,_state_vec_12_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_13_valid = touch_way_0_valid & touch_set_0 == 9'hd; // @[Replacement.scala 315:30]
  wire  state_vec_13_left_subtree_state = state_vec_13[1]; // @[package.scala 154:13]
  wire  state_vec_13_right_subtree_state = state_vec_13[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_13_T_3 = state_vec_0_set_left_older ? state_vec_13_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_13_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_13_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_13_T_8 = {state_vec_0_set_left_older,_state_vec_13_T_3,_state_vec_13_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_14_valid = touch_way_0_valid & touch_set_0 == 9'he; // @[Replacement.scala 315:30]
  wire  state_vec_14_left_subtree_state = state_vec_14[1]; // @[package.scala 154:13]
  wire  state_vec_14_right_subtree_state = state_vec_14[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_14_T_3 = state_vec_0_set_left_older ? state_vec_14_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_14_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_14_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_14_T_8 = {state_vec_0_set_left_older,_state_vec_14_T_3,_state_vec_14_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_15_valid = touch_way_0_valid & touch_set_0 == 9'hf; // @[Replacement.scala 315:30]
  wire  state_vec_15_left_subtree_state = state_vec_15[1]; // @[package.scala 154:13]
  wire  state_vec_15_right_subtree_state = state_vec_15[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_15_T_3 = state_vec_0_set_left_older ? state_vec_15_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_15_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_15_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_15_T_8 = {state_vec_0_set_left_older,_state_vec_15_T_3,_state_vec_15_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_16_valid = touch_way_0_valid & touch_set_0 == 9'h10; // @[Replacement.scala 315:30]
  wire  state_vec_16_left_subtree_state = state_vec_16[1]; // @[package.scala 154:13]
  wire  state_vec_16_right_subtree_state = state_vec_16[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_16_T_3 = state_vec_0_set_left_older ? state_vec_16_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_16_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_16_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_16_T_8 = {state_vec_0_set_left_older,_state_vec_16_T_3,_state_vec_16_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_17_valid = touch_way_0_valid & touch_set_0 == 9'h11; // @[Replacement.scala 315:30]
  wire  state_vec_17_left_subtree_state = state_vec_17[1]; // @[package.scala 154:13]
  wire  state_vec_17_right_subtree_state = state_vec_17[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_17_T_3 = state_vec_0_set_left_older ? state_vec_17_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_17_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_17_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_17_T_8 = {state_vec_0_set_left_older,_state_vec_17_T_3,_state_vec_17_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_18_valid = touch_way_0_valid & touch_set_0 == 9'h12; // @[Replacement.scala 315:30]
  wire  state_vec_18_left_subtree_state = state_vec_18[1]; // @[package.scala 154:13]
  wire  state_vec_18_right_subtree_state = state_vec_18[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_18_T_3 = state_vec_0_set_left_older ? state_vec_18_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_18_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_18_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_18_T_8 = {state_vec_0_set_left_older,_state_vec_18_T_3,_state_vec_18_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_19_valid = touch_way_0_valid & touch_set_0 == 9'h13; // @[Replacement.scala 315:30]
  wire  state_vec_19_left_subtree_state = state_vec_19[1]; // @[package.scala 154:13]
  wire  state_vec_19_right_subtree_state = state_vec_19[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_19_T_3 = state_vec_0_set_left_older ? state_vec_19_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_19_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_19_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_19_T_8 = {state_vec_0_set_left_older,_state_vec_19_T_3,_state_vec_19_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_20_valid = touch_way_0_valid & touch_set_0 == 9'h14; // @[Replacement.scala 315:30]
  wire  state_vec_20_left_subtree_state = state_vec_20[1]; // @[package.scala 154:13]
  wire  state_vec_20_right_subtree_state = state_vec_20[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_20_T_3 = state_vec_0_set_left_older ? state_vec_20_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_20_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_20_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_20_T_8 = {state_vec_0_set_left_older,_state_vec_20_T_3,_state_vec_20_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_21_valid = touch_way_0_valid & touch_set_0 == 9'h15; // @[Replacement.scala 315:30]
  wire  state_vec_21_left_subtree_state = state_vec_21[1]; // @[package.scala 154:13]
  wire  state_vec_21_right_subtree_state = state_vec_21[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_21_T_3 = state_vec_0_set_left_older ? state_vec_21_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_21_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_21_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_21_T_8 = {state_vec_0_set_left_older,_state_vec_21_T_3,_state_vec_21_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_22_valid = touch_way_0_valid & touch_set_0 == 9'h16; // @[Replacement.scala 315:30]
  wire  state_vec_22_left_subtree_state = state_vec_22[1]; // @[package.scala 154:13]
  wire  state_vec_22_right_subtree_state = state_vec_22[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_22_T_3 = state_vec_0_set_left_older ? state_vec_22_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_22_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_22_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_22_T_8 = {state_vec_0_set_left_older,_state_vec_22_T_3,_state_vec_22_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_23_valid = touch_way_0_valid & touch_set_0 == 9'h17; // @[Replacement.scala 315:30]
  wire  state_vec_23_left_subtree_state = state_vec_23[1]; // @[package.scala 154:13]
  wire  state_vec_23_right_subtree_state = state_vec_23[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_23_T_3 = state_vec_0_set_left_older ? state_vec_23_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_23_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_23_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_23_T_8 = {state_vec_0_set_left_older,_state_vec_23_T_3,_state_vec_23_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_24_valid = touch_way_0_valid & touch_set_0 == 9'h18; // @[Replacement.scala 315:30]
  wire  state_vec_24_left_subtree_state = state_vec_24[1]; // @[package.scala 154:13]
  wire  state_vec_24_right_subtree_state = state_vec_24[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_24_T_3 = state_vec_0_set_left_older ? state_vec_24_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_24_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_24_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_24_T_8 = {state_vec_0_set_left_older,_state_vec_24_T_3,_state_vec_24_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_25_valid = touch_way_0_valid & touch_set_0 == 9'h19; // @[Replacement.scala 315:30]
  wire  state_vec_25_left_subtree_state = state_vec_25[1]; // @[package.scala 154:13]
  wire  state_vec_25_right_subtree_state = state_vec_25[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_25_T_3 = state_vec_0_set_left_older ? state_vec_25_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_25_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_25_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_25_T_8 = {state_vec_0_set_left_older,_state_vec_25_T_3,_state_vec_25_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_26_valid = touch_way_0_valid & touch_set_0 == 9'h1a; // @[Replacement.scala 315:30]
  wire  state_vec_26_left_subtree_state = state_vec_26[1]; // @[package.scala 154:13]
  wire  state_vec_26_right_subtree_state = state_vec_26[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_26_T_3 = state_vec_0_set_left_older ? state_vec_26_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_26_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_26_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_26_T_8 = {state_vec_0_set_left_older,_state_vec_26_T_3,_state_vec_26_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_27_valid = touch_way_0_valid & touch_set_0 == 9'h1b; // @[Replacement.scala 315:30]
  wire  state_vec_27_left_subtree_state = state_vec_27[1]; // @[package.scala 154:13]
  wire  state_vec_27_right_subtree_state = state_vec_27[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_27_T_3 = state_vec_0_set_left_older ? state_vec_27_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_27_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_27_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_27_T_8 = {state_vec_0_set_left_older,_state_vec_27_T_3,_state_vec_27_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_28_valid = touch_way_0_valid & touch_set_0 == 9'h1c; // @[Replacement.scala 315:30]
  wire  state_vec_28_left_subtree_state = state_vec_28[1]; // @[package.scala 154:13]
  wire  state_vec_28_right_subtree_state = state_vec_28[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_28_T_3 = state_vec_0_set_left_older ? state_vec_28_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_28_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_28_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_28_T_8 = {state_vec_0_set_left_older,_state_vec_28_T_3,_state_vec_28_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_29_valid = touch_way_0_valid & touch_set_0 == 9'h1d; // @[Replacement.scala 315:30]
  wire  state_vec_29_left_subtree_state = state_vec_29[1]; // @[package.scala 154:13]
  wire  state_vec_29_right_subtree_state = state_vec_29[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_29_T_3 = state_vec_0_set_left_older ? state_vec_29_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_29_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_29_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_29_T_8 = {state_vec_0_set_left_older,_state_vec_29_T_3,_state_vec_29_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_30_valid = touch_way_0_valid & touch_set_0 == 9'h1e; // @[Replacement.scala 315:30]
  wire  state_vec_30_left_subtree_state = state_vec_30[1]; // @[package.scala 154:13]
  wire  state_vec_30_right_subtree_state = state_vec_30[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_30_T_3 = state_vec_0_set_left_older ? state_vec_30_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_30_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_30_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_30_T_8 = {state_vec_0_set_left_older,_state_vec_30_T_3,_state_vec_30_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_31_valid = touch_way_0_valid & touch_set_0 == 9'h1f; // @[Replacement.scala 315:30]
  wire  state_vec_31_left_subtree_state = state_vec_31[1]; // @[package.scala 154:13]
  wire  state_vec_31_right_subtree_state = state_vec_31[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_31_T_3 = state_vec_0_set_left_older ? state_vec_31_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_31_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_31_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_31_T_8 = {state_vec_0_set_left_older,_state_vec_31_T_3,_state_vec_31_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_32_valid = touch_way_0_valid & touch_set_0 == 9'h20; // @[Replacement.scala 315:30]
  wire  state_vec_32_left_subtree_state = state_vec_32[1]; // @[package.scala 154:13]
  wire  state_vec_32_right_subtree_state = state_vec_32[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_32_T_3 = state_vec_0_set_left_older ? state_vec_32_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_32_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_32_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_32_T_8 = {state_vec_0_set_left_older,_state_vec_32_T_3,_state_vec_32_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_33_valid = touch_way_0_valid & touch_set_0 == 9'h21; // @[Replacement.scala 315:30]
  wire  state_vec_33_left_subtree_state = state_vec_33[1]; // @[package.scala 154:13]
  wire  state_vec_33_right_subtree_state = state_vec_33[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_33_T_3 = state_vec_0_set_left_older ? state_vec_33_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_33_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_33_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_33_T_8 = {state_vec_0_set_left_older,_state_vec_33_T_3,_state_vec_33_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_34_valid = touch_way_0_valid & touch_set_0 == 9'h22; // @[Replacement.scala 315:30]
  wire  state_vec_34_left_subtree_state = state_vec_34[1]; // @[package.scala 154:13]
  wire  state_vec_34_right_subtree_state = state_vec_34[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_34_T_3 = state_vec_0_set_left_older ? state_vec_34_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_34_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_34_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_34_T_8 = {state_vec_0_set_left_older,_state_vec_34_T_3,_state_vec_34_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_35_valid = touch_way_0_valid & touch_set_0 == 9'h23; // @[Replacement.scala 315:30]
  wire  state_vec_35_left_subtree_state = state_vec_35[1]; // @[package.scala 154:13]
  wire  state_vec_35_right_subtree_state = state_vec_35[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_35_T_3 = state_vec_0_set_left_older ? state_vec_35_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_35_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_35_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_35_T_8 = {state_vec_0_set_left_older,_state_vec_35_T_3,_state_vec_35_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_36_valid = touch_way_0_valid & touch_set_0 == 9'h24; // @[Replacement.scala 315:30]
  wire  state_vec_36_left_subtree_state = state_vec_36[1]; // @[package.scala 154:13]
  wire  state_vec_36_right_subtree_state = state_vec_36[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_36_T_3 = state_vec_0_set_left_older ? state_vec_36_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_36_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_36_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_36_T_8 = {state_vec_0_set_left_older,_state_vec_36_T_3,_state_vec_36_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_37_valid = touch_way_0_valid & touch_set_0 == 9'h25; // @[Replacement.scala 315:30]
  wire  state_vec_37_left_subtree_state = state_vec_37[1]; // @[package.scala 154:13]
  wire  state_vec_37_right_subtree_state = state_vec_37[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_37_T_3 = state_vec_0_set_left_older ? state_vec_37_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_37_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_37_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_37_T_8 = {state_vec_0_set_left_older,_state_vec_37_T_3,_state_vec_37_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_38_valid = touch_way_0_valid & touch_set_0 == 9'h26; // @[Replacement.scala 315:30]
  wire  state_vec_38_left_subtree_state = state_vec_38[1]; // @[package.scala 154:13]
  wire  state_vec_38_right_subtree_state = state_vec_38[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_38_T_3 = state_vec_0_set_left_older ? state_vec_38_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_38_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_38_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_38_T_8 = {state_vec_0_set_left_older,_state_vec_38_T_3,_state_vec_38_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_39_valid = touch_way_0_valid & touch_set_0 == 9'h27; // @[Replacement.scala 315:30]
  wire  state_vec_39_left_subtree_state = state_vec_39[1]; // @[package.scala 154:13]
  wire  state_vec_39_right_subtree_state = state_vec_39[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_39_T_3 = state_vec_0_set_left_older ? state_vec_39_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_39_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_39_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_39_T_8 = {state_vec_0_set_left_older,_state_vec_39_T_3,_state_vec_39_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_40_valid = touch_way_0_valid & touch_set_0 == 9'h28; // @[Replacement.scala 315:30]
  wire  state_vec_40_left_subtree_state = state_vec_40[1]; // @[package.scala 154:13]
  wire  state_vec_40_right_subtree_state = state_vec_40[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_40_T_3 = state_vec_0_set_left_older ? state_vec_40_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_40_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_40_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_40_T_8 = {state_vec_0_set_left_older,_state_vec_40_T_3,_state_vec_40_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_41_valid = touch_way_0_valid & touch_set_0 == 9'h29; // @[Replacement.scala 315:30]
  wire  state_vec_41_left_subtree_state = state_vec_41[1]; // @[package.scala 154:13]
  wire  state_vec_41_right_subtree_state = state_vec_41[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_41_T_3 = state_vec_0_set_left_older ? state_vec_41_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_41_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_41_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_41_T_8 = {state_vec_0_set_left_older,_state_vec_41_T_3,_state_vec_41_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_42_valid = touch_way_0_valid & touch_set_0 == 9'h2a; // @[Replacement.scala 315:30]
  wire  state_vec_42_left_subtree_state = state_vec_42[1]; // @[package.scala 154:13]
  wire  state_vec_42_right_subtree_state = state_vec_42[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_42_T_3 = state_vec_0_set_left_older ? state_vec_42_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_42_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_42_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_42_T_8 = {state_vec_0_set_left_older,_state_vec_42_T_3,_state_vec_42_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_43_valid = touch_way_0_valid & touch_set_0 == 9'h2b; // @[Replacement.scala 315:30]
  wire  state_vec_43_left_subtree_state = state_vec_43[1]; // @[package.scala 154:13]
  wire  state_vec_43_right_subtree_state = state_vec_43[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_43_T_3 = state_vec_0_set_left_older ? state_vec_43_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_43_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_43_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_43_T_8 = {state_vec_0_set_left_older,_state_vec_43_T_3,_state_vec_43_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_44_valid = touch_way_0_valid & touch_set_0 == 9'h2c; // @[Replacement.scala 315:30]
  wire  state_vec_44_left_subtree_state = state_vec_44[1]; // @[package.scala 154:13]
  wire  state_vec_44_right_subtree_state = state_vec_44[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_44_T_3 = state_vec_0_set_left_older ? state_vec_44_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_44_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_44_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_44_T_8 = {state_vec_0_set_left_older,_state_vec_44_T_3,_state_vec_44_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_45_valid = touch_way_0_valid & touch_set_0 == 9'h2d; // @[Replacement.scala 315:30]
  wire  state_vec_45_left_subtree_state = state_vec_45[1]; // @[package.scala 154:13]
  wire  state_vec_45_right_subtree_state = state_vec_45[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_45_T_3 = state_vec_0_set_left_older ? state_vec_45_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_45_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_45_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_45_T_8 = {state_vec_0_set_left_older,_state_vec_45_T_3,_state_vec_45_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_46_valid = touch_way_0_valid & touch_set_0 == 9'h2e; // @[Replacement.scala 315:30]
  wire  state_vec_46_left_subtree_state = state_vec_46[1]; // @[package.scala 154:13]
  wire  state_vec_46_right_subtree_state = state_vec_46[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_46_T_3 = state_vec_0_set_left_older ? state_vec_46_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_46_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_46_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_46_T_8 = {state_vec_0_set_left_older,_state_vec_46_T_3,_state_vec_46_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_47_valid = touch_way_0_valid & touch_set_0 == 9'h2f; // @[Replacement.scala 315:30]
  wire  state_vec_47_left_subtree_state = state_vec_47[1]; // @[package.scala 154:13]
  wire  state_vec_47_right_subtree_state = state_vec_47[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_47_T_3 = state_vec_0_set_left_older ? state_vec_47_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_47_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_47_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_47_T_8 = {state_vec_0_set_left_older,_state_vec_47_T_3,_state_vec_47_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_48_valid = touch_way_0_valid & touch_set_0 == 9'h30; // @[Replacement.scala 315:30]
  wire  state_vec_48_left_subtree_state = state_vec_48[1]; // @[package.scala 154:13]
  wire  state_vec_48_right_subtree_state = state_vec_48[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_48_T_3 = state_vec_0_set_left_older ? state_vec_48_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_48_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_48_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_48_T_8 = {state_vec_0_set_left_older,_state_vec_48_T_3,_state_vec_48_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_49_valid = touch_way_0_valid & touch_set_0 == 9'h31; // @[Replacement.scala 315:30]
  wire  state_vec_49_left_subtree_state = state_vec_49[1]; // @[package.scala 154:13]
  wire  state_vec_49_right_subtree_state = state_vec_49[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_49_T_3 = state_vec_0_set_left_older ? state_vec_49_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_49_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_49_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_49_T_8 = {state_vec_0_set_left_older,_state_vec_49_T_3,_state_vec_49_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_50_valid = touch_way_0_valid & touch_set_0 == 9'h32; // @[Replacement.scala 315:30]
  wire  state_vec_50_left_subtree_state = state_vec_50[1]; // @[package.scala 154:13]
  wire  state_vec_50_right_subtree_state = state_vec_50[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_50_T_3 = state_vec_0_set_left_older ? state_vec_50_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_50_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_50_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_50_T_8 = {state_vec_0_set_left_older,_state_vec_50_T_3,_state_vec_50_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_51_valid = touch_way_0_valid & touch_set_0 == 9'h33; // @[Replacement.scala 315:30]
  wire  state_vec_51_left_subtree_state = state_vec_51[1]; // @[package.scala 154:13]
  wire  state_vec_51_right_subtree_state = state_vec_51[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_51_T_3 = state_vec_0_set_left_older ? state_vec_51_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_51_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_51_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_51_T_8 = {state_vec_0_set_left_older,_state_vec_51_T_3,_state_vec_51_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_52_valid = touch_way_0_valid & touch_set_0 == 9'h34; // @[Replacement.scala 315:30]
  wire  state_vec_52_left_subtree_state = state_vec_52[1]; // @[package.scala 154:13]
  wire  state_vec_52_right_subtree_state = state_vec_52[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_52_T_3 = state_vec_0_set_left_older ? state_vec_52_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_52_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_52_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_52_T_8 = {state_vec_0_set_left_older,_state_vec_52_T_3,_state_vec_52_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_53_valid = touch_way_0_valid & touch_set_0 == 9'h35; // @[Replacement.scala 315:30]
  wire  state_vec_53_left_subtree_state = state_vec_53[1]; // @[package.scala 154:13]
  wire  state_vec_53_right_subtree_state = state_vec_53[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_53_T_3 = state_vec_0_set_left_older ? state_vec_53_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_53_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_53_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_53_T_8 = {state_vec_0_set_left_older,_state_vec_53_T_3,_state_vec_53_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_54_valid = touch_way_0_valid & touch_set_0 == 9'h36; // @[Replacement.scala 315:30]
  wire  state_vec_54_left_subtree_state = state_vec_54[1]; // @[package.scala 154:13]
  wire  state_vec_54_right_subtree_state = state_vec_54[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_54_T_3 = state_vec_0_set_left_older ? state_vec_54_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_54_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_54_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_54_T_8 = {state_vec_0_set_left_older,_state_vec_54_T_3,_state_vec_54_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_55_valid = touch_way_0_valid & touch_set_0 == 9'h37; // @[Replacement.scala 315:30]
  wire  state_vec_55_left_subtree_state = state_vec_55[1]; // @[package.scala 154:13]
  wire  state_vec_55_right_subtree_state = state_vec_55[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_55_T_3 = state_vec_0_set_left_older ? state_vec_55_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_55_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_55_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_55_T_8 = {state_vec_0_set_left_older,_state_vec_55_T_3,_state_vec_55_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_56_valid = touch_way_0_valid & touch_set_0 == 9'h38; // @[Replacement.scala 315:30]
  wire  state_vec_56_left_subtree_state = state_vec_56[1]; // @[package.scala 154:13]
  wire  state_vec_56_right_subtree_state = state_vec_56[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_56_T_3 = state_vec_0_set_left_older ? state_vec_56_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_56_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_56_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_56_T_8 = {state_vec_0_set_left_older,_state_vec_56_T_3,_state_vec_56_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_57_valid = touch_way_0_valid & touch_set_0 == 9'h39; // @[Replacement.scala 315:30]
  wire  state_vec_57_left_subtree_state = state_vec_57[1]; // @[package.scala 154:13]
  wire  state_vec_57_right_subtree_state = state_vec_57[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_57_T_3 = state_vec_0_set_left_older ? state_vec_57_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_57_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_57_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_57_T_8 = {state_vec_0_set_left_older,_state_vec_57_T_3,_state_vec_57_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_58_valid = touch_way_0_valid & touch_set_0 == 9'h3a; // @[Replacement.scala 315:30]
  wire  state_vec_58_left_subtree_state = state_vec_58[1]; // @[package.scala 154:13]
  wire  state_vec_58_right_subtree_state = state_vec_58[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_58_T_3 = state_vec_0_set_left_older ? state_vec_58_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_58_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_58_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_58_T_8 = {state_vec_0_set_left_older,_state_vec_58_T_3,_state_vec_58_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_59_valid = touch_way_0_valid & touch_set_0 == 9'h3b; // @[Replacement.scala 315:30]
  wire  state_vec_59_left_subtree_state = state_vec_59[1]; // @[package.scala 154:13]
  wire  state_vec_59_right_subtree_state = state_vec_59[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_59_T_3 = state_vec_0_set_left_older ? state_vec_59_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_59_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_59_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_59_T_8 = {state_vec_0_set_left_older,_state_vec_59_T_3,_state_vec_59_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_60_valid = touch_way_0_valid & touch_set_0 == 9'h3c; // @[Replacement.scala 315:30]
  wire  state_vec_60_left_subtree_state = state_vec_60[1]; // @[package.scala 154:13]
  wire  state_vec_60_right_subtree_state = state_vec_60[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_60_T_3 = state_vec_0_set_left_older ? state_vec_60_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_60_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_60_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_60_T_8 = {state_vec_0_set_left_older,_state_vec_60_T_3,_state_vec_60_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_61_valid = touch_way_0_valid & touch_set_0 == 9'h3d; // @[Replacement.scala 315:30]
  wire  state_vec_61_left_subtree_state = state_vec_61[1]; // @[package.scala 154:13]
  wire  state_vec_61_right_subtree_state = state_vec_61[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_61_T_3 = state_vec_0_set_left_older ? state_vec_61_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_61_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_61_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_61_T_8 = {state_vec_0_set_left_older,_state_vec_61_T_3,_state_vec_61_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_62_valid = touch_way_0_valid & touch_set_0 == 9'h3e; // @[Replacement.scala 315:30]
  wire  state_vec_62_left_subtree_state = state_vec_62[1]; // @[package.scala 154:13]
  wire  state_vec_62_right_subtree_state = state_vec_62[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_62_T_3 = state_vec_0_set_left_older ? state_vec_62_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_62_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_62_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_62_T_8 = {state_vec_0_set_left_older,_state_vec_62_T_3,_state_vec_62_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_63_valid = touch_way_0_valid & touch_set_0 == 9'h3f; // @[Replacement.scala 315:30]
  wire  state_vec_63_left_subtree_state = state_vec_63[1]; // @[package.scala 154:13]
  wire  state_vec_63_right_subtree_state = state_vec_63[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_63_T_3 = state_vec_0_set_left_older ? state_vec_63_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_63_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_63_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_63_T_8 = {state_vec_0_set_left_older,_state_vec_63_T_3,_state_vec_63_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_64_valid = touch_way_0_valid & touch_set_0 == 9'h40; // @[Replacement.scala 315:30]
  wire  state_vec_64_left_subtree_state = state_vec_64[1]; // @[package.scala 154:13]
  wire  state_vec_64_right_subtree_state = state_vec_64[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_64_T_3 = state_vec_0_set_left_older ? state_vec_64_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_64_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_64_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_64_T_8 = {state_vec_0_set_left_older,_state_vec_64_T_3,_state_vec_64_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_65_valid = touch_way_0_valid & touch_set_0 == 9'h41; // @[Replacement.scala 315:30]
  wire  state_vec_65_left_subtree_state = state_vec_65[1]; // @[package.scala 154:13]
  wire  state_vec_65_right_subtree_state = state_vec_65[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_65_T_3 = state_vec_0_set_left_older ? state_vec_65_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_65_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_65_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_65_T_8 = {state_vec_0_set_left_older,_state_vec_65_T_3,_state_vec_65_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_66_valid = touch_way_0_valid & touch_set_0 == 9'h42; // @[Replacement.scala 315:30]
  wire  state_vec_66_left_subtree_state = state_vec_66[1]; // @[package.scala 154:13]
  wire  state_vec_66_right_subtree_state = state_vec_66[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_66_T_3 = state_vec_0_set_left_older ? state_vec_66_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_66_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_66_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_66_T_8 = {state_vec_0_set_left_older,_state_vec_66_T_3,_state_vec_66_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_67_valid = touch_way_0_valid & touch_set_0 == 9'h43; // @[Replacement.scala 315:30]
  wire  state_vec_67_left_subtree_state = state_vec_67[1]; // @[package.scala 154:13]
  wire  state_vec_67_right_subtree_state = state_vec_67[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_67_T_3 = state_vec_0_set_left_older ? state_vec_67_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_67_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_67_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_67_T_8 = {state_vec_0_set_left_older,_state_vec_67_T_3,_state_vec_67_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_68_valid = touch_way_0_valid & touch_set_0 == 9'h44; // @[Replacement.scala 315:30]
  wire  state_vec_68_left_subtree_state = state_vec_68[1]; // @[package.scala 154:13]
  wire  state_vec_68_right_subtree_state = state_vec_68[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_68_T_3 = state_vec_0_set_left_older ? state_vec_68_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_68_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_68_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_68_T_8 = {state_vec_0_set_left_older,_state_vec_68_T_3,_state_vec_68_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_69_valid = touch_way_0_valid & touch_set_0 == 9'h45; // @[Replacement.scala 315:30]
  wire  state_vec_69_left_subtree_state = state_vec_69[1]; // @[package.scala 154:13]
  wire  state_vec_69_right_subtree_state = state_vec_69[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_69_T_3 = state_vec_0_set_left_older ? state_vec_69_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_69_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_69_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_69_T_8 = {state_vec_0_set_left_older,_state_vec_69_T_3,_state_vec_69_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_70_valid = touch_way_0_valid & touch_set_0 == 9'h46; // @[Replacement.scala 315:30]
  wire  state_vec_70_left_subtree_state = state_vec_70[1]; // @[package.scala 154:13]
  wire  state_vec_70_right_subtree_state = state_vec_70[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_70_T_3 = state_vec_0_set_left_older ? state_vec_70_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_70_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_70_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_70_T_8 = {state_vec_0_set_left_older,_state_vec_70_T_3,_state_vec_70_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_71_valid = touch_way_0_valid & touch_set_0 == 9'h47; // @[Replacement.scala 315:30]
  wire  state_vec_71_left_subtree_state = state_vec_71[1]; // @[package.scala 154:13]
  wire  state_vec_71_right_subtree_state = state_vec_71[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_71_T_3 = state_vec_0_set_left_older ? state_vec_71_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_71_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_71_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_71_T_8 = {state_vec_0_set_left_older,_state_vec_71_T_3,_state_vec_71_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_72_valid = touch_way_0_valid & touch_set_0 == 9'h48; // @[Replacement.scala 315:30]
  wire  state_vec_72_left_subtree_state = state_vec_72[1]; // @[package.scala 154:13]
  wire  state_vec_72_right_subtree_state = state_vec_72[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_72_T_3 = state_vec_0_set_left_older ? state_vec_72_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_72_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_72_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_72_T_8 = {state_vec_0_set_left_older,_state_vec_72_T_3,_state_vec_72_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_73_valid = touch_way_0_valid & touch_set_0 == 9'h49; // @[Replacement.scala 315:30]
  wire  state_vec_73_left_subtree_state = state_vec_73[1]; // @[package.scala 154:13]
  wire  state_vec_73_right_subtree_state = state_vec_73[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_73_T_3 = state_vec_0_set_left_older ? state_vec_73_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_73_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_73_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_73_T_8 = {state_vec_0_set_left_older,_state_vec_73_T_3,_state_vec_73_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_74_valid = touch_way_0_valid & touch_set_0 == 9'h4a; // @[Replacement.scala 315:30]
  wire  state_vec_74_left_subtree_state = state_vec_74[1]; // @[package.scala 154:13]
  wire  state_vec_74_right_subtree_state = state_vec_74[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_74_T_3 = state_vec_0_set_left_older ? state_vec_74_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_74_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_74_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_74_T_8 = {state_vec_0_set_left_older,_state_vec_74_T_3,_state_vec_74_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_75_valid = touch_way_0_valid & touch_set_0 == 9'h4b; // @[Replacement.scala 315:30]
  wire  state_vec_75_left_subtree_state = state_vec_75[1]; // @[package.scala 154:13]
  wire  state_vec_75_right_subtree_state = state_vec_75[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_75_T_3 = state_vec_0_set_left_older ? state_vec_75_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_75_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_75_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_75_T_8 = {state_vec_0_set_left_older,_state_vec_75_T_3,_state_vec_75_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_76_valid = touch_way_0_valid & touch_set_0 == 9'h4c; // @[Replacement.scala 315:30]
  wire  state_vec_76_left_subtree_state = state_vec_76[1]; // @[package.scala 154:13]
  wire  state_vec_76_right_subtree_state = state_vec_76[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_76_T_3 = state_vec_0_set_left_older ? state_vec_76_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_76_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_76_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_76_T_8 = {state_vec_0_set_left_older,_state_vec_76_T_3,_state_vec_76_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_77_valid = touch_way_0_valid & touch_set_0 == 9'h4d; // @[Replacement.scala 315:30]
  wire  state_vec_77_left_subtree_state = state_vec_77[1]; // @[package.scala 154:13]
  wire  state_vec_77_right_subtree_state = state_vec_77[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_77_T_3 = state_vec_0_set_left_older ? state_vec_77_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_77_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_77_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_77_T_8 = {state_vec_0_set_left_older,_state_vec_77_T_3,_state_vec_77_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_78_valid = touch_way_0_valid & touch_set_0 == 9'h4e; // @[Replacement.scala 315:30]
  wire  state_vec_78_left_subtree_state = state_vec_78[1]; // @[package.scala 154:13]
  wire  state_vec_78_right_subtree_state = state_vec_78[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_78_T_3 = state_vec_0_set_left_older ? state_vec_78_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_78_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_78_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_78_T_8 = {state_vec_0_set_left_older,_state_vec_78_T_3,_state_vec_78_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_79_valid = touch_way_0_valid & touch_set_0 == 9'h4f; // @[Replacement.scala 315:30]
  wire  state_vec_79_left_subtree_state = state_vec_79[1]; // @[package.scala 154:13]
  wire  state_vec_79_right_subtree_state = state_vec_79[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_79_T_3 = state_vec_0_set_left_older ? state_vec_79_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_79_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_79_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_79_T_8 = {state_vec_0_set_left_older,_state_vec_79_T_3,_state_vec_79_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_80_valid = touch_way_0_valid & touch_set_0 == 9'h50; // @[Replacement.scala 315:30]
  wire  state_vec_80_left_subtree_state = state_vec_80[1]; // @[package.scala 154:13]
  wire  state_vec_80_right_subtree_state = state_vec_80[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_80_T_3 = state_vec_0_set_left_older ? state_vec_80_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_80_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_80_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_80_T_8 = {state_vec_0_set_left_older,_state_vec_80_T_3,_state_vec_80_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_81_valid = touch_way_0_valid & touch_set_0 == 9'h51; // @[Replacement.scala 315:30]
  wire  state_vec_81_left_subtree_state = state_vec_81[1]; // @[package.scala 154:13]
  wire  state_vec_81_right_subtree_state = state_vec_81[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_81_T_3 = state_vec_0_set_left_older ? state_vec_81_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_81_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_81_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_81_T_8 = {state_vec_0_set_left_older,_state_vec_81_T_3,_state_vec_81_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_82_valid = touch_way_0_valid & touch_set_0 == 9'h52; // @[Replacement.scala 315:30]
  wire  state_vec_82_left_subtree_state = state_vec_82[1]; // @[package.scala 154:13]
  wire  state_vec_82_right_subtree_state = state_vec_82[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_82_T_3 = state_vec_0_set_left_older ? state_vec_82_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_82_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_82_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_82_T_8 = {state_vec_0_set_left_older,_state_vec_82_T_3,_state_vec_82_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_83_valid = touch_way_0_valid & touch_set_0 == 9'h53; // @[Replacement.scala 315:30]
  wire  state_vec_83_left_subtree_state = state_vec_83[1]; // @[package.scala 154:13]
  wire  state_vec_83_right_subtree_state = state_vec_83[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_83_T_3 = state_vec_0_set_left_older ? state_vec_83_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_83_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_83_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_83_T_8 = {state_vec_0_set_left_older,_state_vec_83_T_3,_state_vec_83_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_84_valid = touch_way_0_valid & touch_set_0 == 9'h54; // @[Replacement.scala 315:30]
  wire  state_vec_84_left_subtree_state = state_vec_84[1]; // @[package.scala 154:13]
  wire  state_vec_84_right_subtree_state = state_vec_84[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_84_T_3 = state_vec_0_set_left_older ? state_vec_84_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_84_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_84_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_84_T_8 = {state_vec_0_set_left_older,_state_vec_84_T_3,_state_vec_84_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_85_valid = touch_way_0_valid & touch_set_0 == 9'h55; // @[Replacement.scala 315:30]
  wire  state_vec_85_left_subtree_state = state_vec_85[1]; // @[package.scala 154:13]
  wire  state_vec_85_right_subtree_state = state_vec_85[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_85_T_3 = state_vec_0_set_left_older ? state_vec_85_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_85_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_85_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_85_T_8 = {state_vec_0_set_left_older,_state_vec_85_T_3,_state_vec_85_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_86_valid = touch_way_0_valid & touch_set_0 == 9'h56; // @[Replacement.scala 315:30]
  wire  state_vec_86_left_subtree_state = state_vec_86[1]; // @[package.scala 154:13]
  wire  state_vec_86_right_subtree_state = state_vec_86[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_86_T_3 = state_vec_0_set_left_older ? state_vec_86_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_86_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_86_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_86_T_8 = {state_vec_0_set_left_older,_state_vec_86_T_3,_state_vec_86_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_87_valid = touch_way_0_valid & touch_set_0 == 9'h57; // @[Replacement.scala 315:30]
  wire  state_vec_87_left_subtree_state = state_vec_87[1]; // @[package.scala 154:13]
  wire  state_vec_87_right_subtree_state = state_vec_87[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_87_T_3 = state_vec_0_set_left_older ? state_vec_87_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_87_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_87_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_87_T_8 = {state_vec_0_set_left_older,_state_vec_87_T_3,_state_vec_87_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_88_valid = touch_way_0_valid & touch_set_0 == 9'h58; // @[Replacement.scala 315:30]
  wire  state_vec_88_left_subtree_state = state_vec_88[1]; // @[package.scala 154:13]
  wire  state_vec_88_right_subtree_state = state_vec_88[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_88_T_3 = state_vec_0_set_left_older ? state_vec_88_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_88_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_88_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_88_T_8 = {state_vec_0_set_left_older,_state_vec_88_T_3,_state_vec_88_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_89_valid = touch_way_0_valid & touch_set_0 == 9'h59; // @[Replacement.scala 315:30]
  wire  state_vec_89_left_subtree_state = state_vec_89[1]; // @[package.scala 154:13]
  wire  state_vec_89_right_subtree_state = state_vec_89[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_89_T_3 = state_vec_0_set_left_older ? state_vec_89_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_89_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_89_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_89_T_8 = {state_vec_0_set_left_older,_state_vec_89_T_3,_state_vec_89_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_90_valid = touch_way_0_valid & touch_set_0 == 9'h5a; // @[Replacement.scala 315:30]
  wire  state_vec_90_left_subtree_state = state_vec_90[1]; // @[package.scala 154:13]
  wire  state_vec_90_right_subtree_state = state_vec_90[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_90_T_3 = state_vec_0_set_left_older ? state_vec_90_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_90_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_90_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_90_T_8 = {state_vec_0_set_left_older,_state_vec_90_T_3,_state_vec_90_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_91_valid = touch_way_0_valid & touch_set_0 == 9'h5b; // @[Replacement.scala 315:30]
  wire  state_vec_91_left_subtree_state = state_vec_91[1]; // @[package.scala 154:13]
  wire  state_vec_91_right_subtree_state = state_vec_91[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_91_T_3 = state_vec_0_set_left_older ? state_vec_91_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_91_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_91_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_91_T_8 = {state_vec_0_set_left_older,_state_vec_91_T_3,_state_vec_91_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_92_valid = touch_way_0_valid & touch_set_0 == 9'h5c; // @[Replacement.scala 315:30]
  wire  state_vec_92_left_subtree_state = state_vec_92[1]; // @[package.scala 154:13]
  wire  state_vec_92_right_subtree_state = state_vec_92[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_92_T_3 = state_vec_0_set_left_older ? state_vec_92_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_92_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_92_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_92_T_8 = {state_vec_0_set_left_older,_state_vec_92_T_3,_state_vec_92_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_93_valid = touch_way_0_valid & touch_set_0 == 9'h5d; // @[Replacement.scala 315:30]
  wire  state_vec_93_left_subtree_state = state_vec_93[1]; // @[package.scala 154:13]
  wire  state_vec_93_right_subtree_state = state_vec_93[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_93_T_3 = state_vec_0_set_left_older ? state_vec_93_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_93_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_93_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_93_T_8 = {state_vec_0_set_left_older,_state_vec_93_T_3,_state_vec_93_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_94_valid = touch_way_0_valid & touch_set_0 == 9'h5e; // @[Replacement.scala 315:30]
  wire  state_vec_94_left_subtree_state = state_vec_94[1]; // @[package.scala 154:13]
  wire  state_vec_94_right_subtree_state = state_vec_94[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_94_T_3 = state_vec_0_set_left_older ? state_vec_94_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_94_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_94_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_94_T_8 = {state_vec_0_set_left_older,_state_vec_94_T_3,_state_vec_94_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_95_valid = touch_way_0_valid & touch_set_0 == 9'h5f; // @[Replacement.scala 315:30]
  wire  state_vec_95_left_subtree_state = state_vec_95[1]; // @[package.scala 154:13]
  wire  state_vec_95_right_subtree_state = state_vec_95[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_95_T_3 = state_vec_0_set_left_older ? state_vec_95_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_95_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_95_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_95_T_8 = {state_vec_0_set_left_older,_state_vec_95_T_3,_state_vec_95_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_96_valid = touch_way_0_valid & touch_set_0 == 9'h60; // @[Replacement.scala 315:30]
  wire  state_vec_96_left_subtree_state = state_vec_96[1]; // @[package.scala 154:13]
  wire  state_vec_96_right_subtree_state = state_vec_96[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_96_T_3 = state_vec_0_set_left_older ? state_vec_96_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_96_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_96_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_96_T_8 = {state_vec_0_set_left_older,_state_vec_96_T_3,_state_vec_96_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_97_valid = touch_way_0_valid & touch_set_0 == 9'h61; // @[Replacement.scala 315:30]
  wire  state_vec_97_left_subtree_state = state_vec_97[1]; // @[package.scala 154:13]
  wire  state_vec_97_right_subtree_state = state_vec_97[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_97_T_3 = state_vec_0_set_left_older ? state_vec_97_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_97_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_97_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_97_T_8 = {state_vec_0_set_left_older,_state_vec_97_T_3,_state_vec_97_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_98_valid = touch_way_0_valid & touch_set_0 == 9'h62; // @[Replacement.scala 315:30]
  wire  state_vec_98_left_subtree_state = state_vec_98[1]; // @[package.scala 154:13]
  wire  state_vec_98_right_subtree_state = state_vec_98[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_98_T_3 = state_vec_0_set_left_older ? state_vec_98_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_98_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_98_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_98_T_8 = {state_vec_0_set_left_older,_state_vec_98_T_3,_state_vec_98_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_99_valid = touch_way_0_valid & touch_set_0 == 9'h63; // @[Replacement.scala 315:30]
  wire  state_vec_99_left_subtree_state = state_vec_99[1]; // @[package.scala 154:13]
  wire  state_vec_99_right_subtree_state = state_vec_99[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_99_T_3 = state_vec_0_set_left_older ? state_vec_99_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_99_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_99_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_99_T_8 = {state_vec_0_set_left_older,_state_vec_99_T_3,_state_vec_99_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_100_valid = touch_way_0_valid & touch_set_0 == 9'h64; // @[Replacement.scala 315:30]
  wire  state_vec_100_left_subtree_state = state_vec_100[1]; // @[package.scala 154:13]
  wire  state_vec_100_right_subtree_state = state_vec_100[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_100_T_3 = state_vec_0_set_left_older ? state_vec_100_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_100_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_100_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_100_T_8 = {state_vec_0_set_left_older,_state_vec_100_T_3,_state_vec_100_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_101_valid = touch_way_0_valid & touch_set_0 == 9'h65; // @[Replacement.scala 315:30]
  wire  state_vec_101_left_subtree_state = state_vec_101[1]; // @[package.scala 154:13]
  wire  state_vec_101_right_subtree_state = state_vec_101[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_101_T_3 = state_vec_0_set_left_older ? state_vec_101_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_101_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_101_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_101_T_8 = {state_vec_0_set_left_older,_state_vec_101_T_3,_state_vec_101_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_102_valid = touch_way_0_valid & touch_set_0 == 9'h66; // @[Replacement.scala 315:30]
  wire  state_vec_102_left_subtree_state = state_vec_102[1]; // @[package.scala 154:13]
  wire  state_vec_102_right_subtree_state = state_vec_102[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_102_T_3 = state_vec_0_set_left_older ? state_vec_102_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_102_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_102_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_102_T_8 = {state_vec_0_set_left_older,_state_vec_102_T_3,_state_vec_102_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_103_valid = touch_way_0_valid & touch_set_0 == 9'h67; // @[Replacement.scala 315:30]
  wire  state_vec_103_left_subtree_state = state_vec_103[1]; // @[package.scala 154:13]
  wire  state_vec_103_right_subtree_state = state_vec_103[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_103_T_3 = state_vec_0_set_left_older ? state_vec_103_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_103_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_103_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_103_T_8 = {state_vec_0_set_left_older,_state_vec_103_T_3,_state_vec_103_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_104_valid = touch_way_0_valid & touch_set_0 == 9'h68; // @[Replacement.scala 315:30]
  wire  state_vec_104_left_subtree_state = state_vec_104[1]; // @[package.scala 154:13]
  wire  state_vec_104_right_subtree_state = state_vec_104[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_104_T_3 = state_vec_0_set_left_older ? state_vec_104_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_104_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_104_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_104_T_8 = {state_vec_0_set_left_older,_state_vec_104_T_3,_state_vec_104_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_105_valid = touch_way_0_valid & touch_set_0 == 9'h69; // @[Replacement.scala 315:30]
  wire  state_vec_105_left_subtree_state = state_vec_105[1]; // @[package.scala 154:13]
  wire  state_vec_105_right_subtree_state = state_vec_105[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_105_T_3 = state_vec_0_set_left_older ? state_vec_105_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_105_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_105_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_105_T_8 = {state_vec_0_set_left_older,_state_vec_105_T_3,_state_vec_105_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_106_valid = touch_way_0_valid & touch_set_0 == 9'h6a; // @[Replacement.scala 315:30]
  wire  state_vec_106_left_subtree_state = state_vec_106[1]; // @[package.scala 154:13]
  wire  state_vec_106_right_subtree_state = state_vec_106[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_106_T_3 = state_vec_0_set_left_older ? state_vec_106_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_106_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_106_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_106_T_8 = {state_vec_0_set_left_older,_state_vec_106_T_3,_state_vec_106_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_107_valid = touch_way_0_valid & touch_set_0 == 9'h6b; // @[Replacement.scala 315:30]
  wire  state_vec_107_left_subtree_state = state_vec_107[1]; // @[package.scala 154:13]
  wire  state_vec_107_right_subtree_state = state_vec_107[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_107_T_3 = state_vec_0_set_left_older ? state_vec_107_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_107_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_107_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_107_T_8 = {state_vec_0_set_left_older,_state_vec_107_T_3,_state_vec_107_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_108_valid = touch_way_0_valid & touch_set_0 == 9'h6c; // @[Replacement.scala 315:30]
  wire  state_vec_108_left_subtree_state = state_vec_108[1]; // @[package.scala 154:13]
  wire  state_vec_108_right_subtree_state = state_vec_108[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_108_T_3 = state_vec_0_set_left_older ? state_vec_108_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_108_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_108_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_108_T_8 = {state_vec_0_set_left_older,_state_vec_108_T_3,_state_vec_108_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_109_valid = touch_way_0_valid & touch_set_0 == 9'h6d; // @[Replacement.scala 315:30]
  wire  state_vec_109_left_subtree_state = state_vec_109[1]; // @[package.scala 154:13]
  wire  state_vec_109_right_subtree_state = state_vec_109[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_109_T_3 = state_vec_0_set_left_older ? state_vec_109_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_109_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_109_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_109_T_8 = {state_vec_0_set_left_older,_state_vec_109_T_3,_state_vec_109_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_110_valid = touch_way_0_valid & touch_set_0 == 9'h6e; // @[Replacement.scala 315:30]
  wire  state_vec_110_left_subtree_state = state_vec_110[1]; // @[package.scala 154:13]
  wire  state_vec_110_right_subtree_state = state_vec_110[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_110_T_3 = state_vec_0_set_left_older ? state_vec_110_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_110_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_110_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_110_T_8 = {state_vec_0_set_left_older,_state_vec_110_T_3,_state_vec_110_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_111_valid = touch_way_0_valid & touch_set_0 == 9'h6f; // @[Replacement.scala 315:30]
  wire  state_vec_111_left_subtree_state = state_vec_111[1]; // @[package.scala 154:13]
  wire  state_vec_111_right_subtree_state = state_vec_111[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_111_T_3 = state_vec_0_set_left_older ? state_vec_111_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_111_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_111_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_111_T_8 = {state_vec_0_set_left_older,_state_vec_111_T_3,_state_vec_111_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_112_valid = touch_way_0_valid & touch_set_0 == 9'h70; // @[Replacement.scala 315:30]
  wire  state_vec_112_left_subtree_state = state_vec_112[1]; // @[package.scala 154:13]
  wire  state_vec_112_right_subtree_state = state_vec_112[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_112_T_3 = state_vec_0_set_left_older ? state_vec_112_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_112_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_112_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_112_T_8 = {state_vec_0_set_left_older,_state_vec_112_T_3,_state_vec_112_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_113_valid = touch_way_0_valid & touch_set_0 == 9'h71; // @[Replacement.scala 315:30]
  wire  state_vec_113_left_subtree_state = state_vec_113[1]; // @[package.scala 154:13]
  wire  state_vec_113_right_subtree_state = state_vec_113[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_113_T_3 = state_vec_0_set_left_older ? state_vec_113_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_113_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_113_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_113_T_8 = {state_vec_0_set_left_older,_state_vec_113_T_3,_state_vec_113_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_114_valid = touch_way_0_valid & touch_set_0 == 9'h72; // @[Replacement.scala 315:30]
  wire  state_vec_114_left_subtree_state = state_vec_114[1]; // @[package.scala 154:13]
  wire  state_vec_114_right_subtree_state = state_vec_114[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_114_T_3 = state_vec_0_set_left_older ? state_vec_114_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_114_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_114_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_114_T_8 = {state_vec_0_set_left_older,_state_vec_114_T_3,_state_vec_114_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_115_valid = touch_way_0_valid & touch_set_0 == 9'h73; // @[Replacement.scala 315:30]
  wire  state_vec_115_left_subtree_state = state_vec_115[1]; // @[package.scala 154:13]
  wire  state_vec_115_right_subtree_state = state_vec_115[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_115_T_3 = state_vec_0_set_left_older ? state_vec_115_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_115_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_115_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_115_T_8 = {state_vec_0_set_left_older,_state_vec_115_T_3,_state_vec_115_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_116_valid = touch_way_0_valid & touch_set_0 == 9'h74; // @[Replacement.scala 315:30]
  wire  state_vec_116_left_subtree_state = state_vec_116[1]; // @[package.scala 154:13]
  wire  state_vec_116_right_subtree_state = state_vec_116[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_116_T_3 = state_vec_0_set_left_older ? state_vec_116_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_116_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_116_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_116_T_8 = {state_vec_0_set_left_older,_state_vec_116_T_3,_state_vec_116_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_117_valid = touch_way_0_valid & touch_set_0 == 9'h75; // @[Replacement.scala 315:30]
  wire  state_vec_117_left_subtree_state = state_vec_117[1]; // @[package.scala 154:13]
  wire  state_vec_117_right_subtree_state = state_vec_117[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_117_T_3 = state_vec_0_set_left_older ? state_vec_117_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_117_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_117_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_117_T_8 = {state_vec_0_set_left_older,_state_vec_117_T_3,_state_vec_117_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_118_valid = touch_way_0_valid & touch_set_0 == 9'h76; // @[Replacement.scala 315:30]
  wire  state_vec_118_left_subtree_state = state_vec_118[1]; // @[package.scala 154:13]
  wire  state_vec_118_right_subtree_state = state_vec_118[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_118_T_3 = state_vec_0_set_left_older ? state_vec_118_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_118_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_118_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_118_T_8 = {state_vec_0_set_left_older,_state_vec_118_T_3,_state_vec_118_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_119_valid = touch_way_0_valid & touch_set_0 == 9'h77; // @[Replacement.scala 315:30]
  wire  state_vec_119_left_subtree_state = state_vec_119[1]; // @[package.scala 154:13]
  wire  state_vec_119_right_subtree_state = state_vec_119[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_119_T_3 = state_vec_0_set_left_older ? state_vec_119_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_119_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_119_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_119_T_8 = {state_vec_0_set_left_older,_state_vec_119_T_3,_state_vec_119_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_120_valid = touch_way_0_valid & touch_set_0 == 9'h78; // @[Replacement.scala 315:30]
  wire  state_vec_120_left_subtree_state = state_vec_120[1]; // @[package.scala 154:13]
  wire  state_vec_120_right_subtree_state = state_vec_120[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_120_T_3 = state_vec_0_set_left_older ? state_vec_120_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_120_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_120_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_120_T_8 = {state_vec_0_set_left_older,_state_vec_120_T_3,_state_vec_120_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_121_valid = touch_way_0_valid & touch_set_0 == 9'h79; // @[Replacement.scala 315:30]
  wire  state_vec_121_left_subtree_state = state_vec_121[1]; // @[package.scala 154:13]
  wire  state_vec_121_right_subtree_state = state_vec_121[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_121_T_3 = state_vec_0_set_left_older ? state_vec_121_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_121_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_121_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_121_T_8 = {state_vec_0_set_left_older,_state_vec_121_T_3,_state_vec_121_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_122_valid = touch_way_0_valid & touch_set_0 == 9'h7a; // @[Replacement.scala 315:30]
  wire  state_vec_122_left_subtree_state = state_vec_122[1]; // @[package.scala 154:13]
  wire  state_vec_122_right_subtree_state = state_vec_122[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_122_T_3 = state_vec_0_set_left_older ? state_vec_122_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_122_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_122_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_122_T_8 = {state_vec_0_set_left_older,_state_vec_122_T_3,_state_vec_122_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_123_valid = touch_way_0_valid & touch_set_0 == 9'h7b; // @[Replacement.scala 315:30]
  wire  state_vec_123_left_subtree_state = state_vec_123[1]; // @[package.scala 154:13]
  wire  state_vec_123_right_subtree_state = state_vec_123[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_123_T_3 = state_vec_0_set_left_older ? state_vec_123_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_123_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_123_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_123_T_8 = {state_vec_0_set_left_older,_state_vec_123_T_3,_state_vec_123_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_124_valid = touch_way_0_valid & touch_set_0 == 9'h7c; // @[Replacement.scala 315:30]
  wire  state_vec_124_left_subtree_state = state_vec_124[1]; // @[package.scala 154:13]
  wire  state_vec_124_right_subtree_state = state_vec_124[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_124_T_3 = state_vec_0_set_left_older ? state_vec_124_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_124_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_124_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_124_T_8 = {state_vec_0_set_left_older,_state_vec_124_T_3,_state_vec_124_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_125_valid = touch_way_0_valid & touch_set_0 == 9'h7d; // @[Replacement.scala 315:30]
  wire  state_vec_125_left_subtree_state = state_vec_125[1]; // @[package.scala 154:13]
  wire  state_vec_125_right_subtree_state = state_vec_125[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_125_T_3 = state_vec_0_set_left_older ? state_vec_125_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_125_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_125_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_125_T_8 = {state_vec_0_set_left_older,_state_vec_125_T_3,_state_vec_125_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_126_valid = touch_way_0_valid & touch_set_0 == 9'h7e; // @[Replacement.scala 315:30]
  wire  state_vec_126_left_subtree_state = state_vec_126[1]; // @[package.scala 154:13]
  wire  state_vec_126_right_subtree_state = state_vec_126[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_126_T_3 = state_vec_0_set_left_older ? state_vec_126_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_126_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_126_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_126_T_8 = {state_vec_0_set_left_older,_state_vec_126_T_3,_state_vec_126_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_127_valid = touch_way_0_valid & touch_set_0 == 9'h7f; // @[Replacement.scala 315:30]
  wire  state_vec_127_left_subtree_state = state_vec_127[1]; // @[package.scala 154:13]
  wire  state_vec_127_right_subtree_state = state_vec_127[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_127_T_3 = state_vec_0_set_left_older ? state_vec_127_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_127_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_127_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_127_T_8 = {state_vec_0_set_left_older,_state_vec_127_T_3,_state_vec_127_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_128_valid = touch_way_0_valid & touch_set_0 == 9'h80; // @[Replacement.scala 315:30]
  wire  state_vec_128_left_subtree_state = state_vec_128[1]; // @[package.scala 154:13]
  wire  state_vec_128_right_subtree_state = state_vec_128[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_128_T_3 = state_vec_0_set_left_older ? state_vec_128_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_128_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_128_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_128_T_8 = {state_vec_0_set_left_older,_state_vec_128_T_3,_state_vec_128_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_129_valid = touch_way_0_valid & touch_set_0 == 9'h81; // @[Replacement.scala 315:30]
  wire  state_vec_129_left_subtree_state = state_vec_129[1]; // @[package.scala 154:13]
  wire  state_vec_129_right_subtree_state = state_vec_129[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_129_T_3 = state_vec_0_set_left_older ? state_vec_129_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_129_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_129_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_129_T_8 = {state_vec_0_set_left_older,_state_vec_129_T_3,_state_vec_129_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_130_valid = touch_way_0_valid & touch_set_0 == 9'h82; // @[Replacement.scala 315:30]
  wire  state_vec_130_left_subtree_state = state_vec_130[1]; // @[package.scala 154:13]
  wire  state_vec_130_right_subtree_state = state_vec_130[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_130_T_3 = state_vec_0_set_left_older ? state_vec_130_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_130_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_130_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_130_T_8 = {state_vec_0_set_left_older,_state_vec_130_T_3,_state_vec_130_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_131_valid = touch_way_0_valid & touch_set_0 == 9'h83; // @[Replacement.scala 315:30]
  wire  state_vec_131_left_subtree_state = state_vec_131[1]; // @[package.scala 154:13]
  wire  state_vec_131_right_subtree_state = state_vec_131[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_131_T_3 = state_vec_0_set_left_older ? state_vec_131_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_131_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_131_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_131_T_8 = {state_vec_0_set_left_older,_state_vec_131_T_3,_state_vec_131_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_132_valid = touch_way_0_valid & touch_set_0 == 9'h84; // @[Replacement.scala 315:30]
  wire  state_vec_132_left_subtree_state = state_vec_132[1]; // @[package.scala 154:13]
  wire  state_vec_132_right_subtree_state = state_vec_132[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_132_T_3 = state_vec_0_set_left_older ? state_vec_132_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_132_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_132_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_132_T_8 = {state_vec_0_set_left_older,_state_vec_132_T_3,_state_vec_132_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_133_valid = touch_way_0_valid & touch_set_0 == 9'h85; // @[Replacement.scala 315:30]
  wire  state_vec_133_left_subtree_state = state_vec_133[1]; // @[package.scala 154:13]
  wire  state_vec_133_right_subtree_state = state_vec_133[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_133_T_3 = state_vec_0_set_left_older ? state_vec_133_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_133_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_133_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_133_T_8 = {state_vec_0_set_left_older,_state_vec_133_T_3,_state_vec_133_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_134_valid = touch_way_0_valid & touch_set_0 == 9'h86; // @[Replacement.scala 315:30]
  wire  state_vec_134_left_subtree_state = state_vec_134[1]; // @[package.scala 154:13]
  wire  state_vec_134_right_subtree_state = state_vec_134[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_134_T_3 = state_vec_0_set_left_older ? state_vec_134_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_134_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_134_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_134_T_8 = {state_vec_0_set_left_older,_state_vec_134_T_3,_state_vec_134_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_135_valid = touch_way_0_valid & touch_set_0 == 9'h87; // @[Replacement.scala 315:30]
  wire  state_vec_135_left_subtree_state = state_vec_135[1]; // @[package.scala 154:13]
  wire  state_vec_135_right_subtree_state = state_vec_135[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_135_T_3 = state_vec_0_set_left_older ? state_vec_135_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_135_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_135_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_135_T_8 = {state_vec_0_set_left_older,_state_vec_135_T_3,_state_vec_135_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_136_valid = touch_way_0_valid & touch_set_0 == 9'h88; // @[Replacement.scala 315:30]
  wire  state_vec_136_left_subtree_state = state_vec_136[1]; // @[package.scala 154:13]
  wire  state_vec_136_right_subtree_state = state_vec_136[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_136_T_3 = state_vec_0_set_left_older ? state_vec_136_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_136_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_136_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_136_T_8 = {state_vec_0_set_left_older,_state_vec_136_T_3,_state_vec_136_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_137_valid = touch_way_0_valid & touch_set_0 == 9'h89; // @[Replacement.scala 315:30]
  wire  state_vec_137_left_subtree_state = state_vec_137[1]; // @[package.scala 154:13]
  wire  state_vec_137_right_subtree_state = state_vec_137[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_137_T_3 = state_vec_0_set_left_older ? state_vec_137_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_137_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_137_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_137_T_8 = {state_vec_0_set_left_older,_state_vec_137_T_3,_state_vec_137_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_138_valid = touch_way_0_valid & touch_set_0 == 9'h8a; // @[Replacement.scala 315:30]
  wire  state_vec_138_left_subtree_state = state_vec_138[1]; // @[package.scala 154:13]
  wire  state_vec_138_right_subtree_state = state_vec_138[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_138_T_3 = state_vec_0_set_left_older ? state_vec_138_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_138_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_138_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_138_T_8 = {state_vec_0_set_left_older,_state_vec_138_T_3,_state_vec_138_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_139_valid = touch_way_0_valid & touch_set_0 == 9'h8b; // @[Replacement.scala 315:30]
  wire  state_vec_139_left_subtree_state = state_vec_139[1]; // @[package.scala 154:13]
  wire  state_vec_139_right_subtree_state = state_vec_139[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_139_T_3 = state_vec_0_set_left_older ? state_vec_139_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_139_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_139_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_139_T_8 = {state_vec_0_set_left_older,_state_vec_139_T_3,_state_vec_139_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_140_valid = touch_way_0_valid & touch_set_0 == 9'h8c; // @[Replacement.scala 315:30]
  wire  state_vec_140_left_subtree_state = state_vec_140[1]; // @[package.scala 154:13]
  wire  state_vec_140_right_subtree_state = state_vec_140[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_140_T_3 = state_vec_0_set_left_older ? state_vec_140_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_140_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_140_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_140_T_8 = {state_vec_0_set_left_older,_state_vec_140_T_3,_state_vec_140_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_141_valid = touch_way_0_valid & touch_set_0 == 9'h8d; // @[Replacement.scala 315:30]
  wire  state_vec_141_left_subtree_state = state_vec_141[1]; // @[package.scala 154:13]
  wire  state_vec_141_right_subtree_state = state_vec_141[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_141_T_3 = state_vec_0_set_left_older ? state_vec_141_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_141_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_141_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_141_T_8 = {state_vec_0_set_left_older,_state_vec_141_T_3,_state_vec_141_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_142_valid = touch_way_0_valid & touch_set_0 == 9'h8e; // @[Replacement.scala 315:30]
  wire  state_vec_142_left_subtree_state = state_vec_142[1]; // @[package.scala 154:13]
  wire  state_vec_142_right_subtree_state = state_vec_142[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_142_T_3 = state_vec_0_set_left_older ? state_vec_142_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_142_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_142_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_142_T_8 = {state_vec_0_set_left_older,_state_vec_142_T_3,_state_vec_142_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_143_valid = touch_way_0_valid & touch_set_0 == 9'h8f; // @[Replacement.scala 315:30]
  wire  state_vec_143_left_subtree_state = state_vec_143[1]; // @[package.scala 154:13]
  wire  state_vec_143_right_subtree_state = state_vec_143[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_143_T_3 = state_vec_0_set_left_older ? state_vec_143_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_143_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_143_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_143_T_8 = {state_vec_0_set_left_older,_state_vec_143_T_3,_state_vec_143_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_144_valid = touch_way_0_valid & touch_set_0 == 9'h90; // @[Replacement.scala 315:30]
  wire  state_vec_144_left_subtree_state = state_vec_144[1]; // @[package.scala 154:13]
  wire  state_vec_144_right_subtree_state = state_vec_144[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_144_T_3 = state_vec_0_set_left_older ? state_vec_144_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_144_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_144_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_144_T_8 = {state_vec_0_set_left_older,_state_vec_144_T_3,_state_vec_144_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_145_valid = touch_way_0_valid & touch_set_0 == 9'h91; // @[Replacement.scala 315:30]
  wire  state_vec_145_left_subtree_state = state_vec_145[1]; // @[package.scala 154:13]
  wire  state_vec_145_right_subtree_state = state_vec_145[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_145_T_3 = state_vec_0_set_left_older ? state_vec_145_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_145_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_145_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_145_T_8 = {state_vec_0_set_left_older,_state_vec_145_T_3,_state_vec_145_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_146_valid = touch_way_0_valid & touch_set_0 == 9'h92; // @[Replacement.scala 315:30]
  wire  state_vec_146_left_subtree_state = state_vec_146[1]; // @[package.scala 154:13]
  wire  state_vec_146_right_subtree_state = state_vec_146[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_146_T_3 = state_vec_0_set_left_older ? state_vec_146_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_146_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_146_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_146_T_8 = {state_vec_0_set_left_older,_state_vec_146_T_3,_state_vec_146_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_147_valid = touch_way_0_valid & touch_set_0 == 9'h93; // @[Replacement.scala 315:30]
  wire  state_vec_147_left_subtree_state = state_vec_147[1]; // @[package.scala 154:13]
  wire  state_vec_147_right_subtree_state = state_vec_147[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_147_T_3 = state_vec_0_set_left_older ? state_vec_147_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_147_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_147_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_147_T_8 = {state_vec_0_set_left_older,_state_vec_147_T_3,_state_vec_147_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_148_valid = touch_way_0_valid & touch_set_0 == 9'h94; // @[Replacement.scala 315:30]
  wire  state_vec_148_left_subtree_state = state_vec_148[1]; // @[package.scala 154:13]
  wire  state_vec_148_right_subtree_state = state_vec_148[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_148_T_3 = state_vec_0_set_left_older ? state_vec_148_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_148_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_148_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_148_T_8 = {state_vec_0_set_left_older,_state_vec_148_T_3,_state_vec_148_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_149_valid = touch_way_0_valid & touch_set_0 == 9'h95; // @[Replacement.scala 315:30]
  wire  state_vec_149_left_subtree_state = state_vec_149[1]; // @[package.scala 154:13]
  wire  state_vec_149_right_subtree_state = state_vec_149[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_149_T_3 = state_vec_0_set_left_older ? state_vec_149_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_149_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_149_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_149_T_8 = {state_vec_0_set_left_older,_state_vec_149_T_3,_state_vec_149_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_150_valid = touch_way_0_valid & touch_set_0 == 9'h96; // @[Replacement.scala 315:30]
  wire  state_vec_150_left_subtree_state = state_vec_150[1]; // @[package.scala 154:13]
  wire  state_vec_150_right_subtree_state = state_vec_150[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_150_T_3 = state_vec_0_set_left_older ? state_vec_150_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_150_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_150_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_150_T_8 = {state_vec_0_set_left_older,_state_vec_150_T_3,_state_vec_150_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_151_valid = touch_way_0_valid & touch_set_0 == 9'h97; // @[Replacement.scala 315:30]
  wire  state_vec_151_left_subtree_state = state_vec_151[1]; // @[package.scala 154:13]
  wire  state_vec_151_right_subtree_state = state_vec_151[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_151_T_3 = state_vec_0_set_left_older ? state_vec_151_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_151_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_151_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_151_T_8 = {state_vec_0_set_left_older,_state_vec_151_T_3,_state_vec_151_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_152_valid = touch_way_0_valid & touch_set_0 == 9'h98; // @[Replacement.scala 315:30]
  wire  state_vec_152_left_subtree_state = state_vec_152[1]; // @[package.scala 154:13]
  wire  state_vec_152_right_subtree_state = state_vec_152[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_152_T_3 = state_vec_0_set_left_older ? state_vec_152_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_152_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_152_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_152_T_8 = {state_vec_0_set_left_older,_state_vec_152_T_3,_state_vec_152_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_153_valid = touch_way_0_valid & touch_set_0 == 9'h99; // @[Replacement.scala 315:30]
  wire  state_vec_153_left_subtree_state = state_vec_153[1]; // @[package.scala 154:13]
  wire  state_vec_153_right_subtree_state = state_vec_153[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_153_T_3 = state_vec_0_set_left_older ? state_vec_153_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_153_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_153_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_153_T_8 = {state_vec_0_set_left_older,_state_vec_153_T_3,_state_vec_153_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_154_valid = touch_way_0_valid & touch_set_0 == 9'h9a; // @[Replacement.scala 315:30]
  wire  state_vec_154_left_subtree_state = state_vec_154[1]; // @[package.scala 154:13]
  wire  state_vec_154_right_subtree_state = state_vec_154[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_154_T_3 = state_vec_0_set_left_older ? state_vec_154_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_154_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_154_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_154_T_8 = {state_vec_0_set_left_older,_state_vec_154_T_3,_state_vec_154_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_155_valid = touch_way_0_valid & touch_set_0 == 9'h9b; // @[Replacement.scala 315:30]
  wire  state_vec_155_left_subtree_state = state_vec_155[1]; // @[package.scala 154:13]
  wire  state_vec_155_right_subtree_state = state_vec_155[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_155_T_3 = state_vec_0_set_left_older ? state_vec_155_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_155_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_155_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_155_T_8 = {state_vec_0_set_left_older,_state_vec_155_T_3,_state_vec_155_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_156_valid = touch_way_0_valid & touch_set_0 == 9'h9c; // @[Replacement.scala 315:30]
  wire  state_vec_156_left_subtree_state = state_vec_156[1]; // @[package.scala 154:13]
  wire  state_vec_156_right_subtree_state = state_vec_156[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_156_T_3 = state_vec_0_set_left_older ? state_vec_156_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_156_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_156_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_156_T_8 = {state_vec_0_set_left_older,_state_vec_156_T_3,_state_vec_156_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_157_valid = touch_way_0_valid & touch_set_0 == 9'h9d; // @[Replacement.scala 315:30]
  wire  state_vec_157_left_subtree_state = state_vec_157[1]; // @[package.scala 154:13]
  wire  state_vec_157_right_subtree_state = state_vec_157[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_157_T_3 = state_vec_0_set_left_older ? state_vec_157_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_157_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_157_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_157_T_8 = {state_vec_0_set_left_older,_state_vec_157_T_3,_state_vec_157_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_158_valid = touch_way_0_valid & touch_set_0 == 9'h9e; // @[Replacement.scala 315:30]
  wire  state_vec_158_left_subtree_state = state_vec_158[1]; // @[package.scala 154:13]
  wire  state_vec_158_right_subtree_state = state_vec_158[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_158_T_3 = state_vec_0_set_left_older ? state_vec_158_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_158_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_158_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_158_T_8 = {state_vec_0_set_left_older,_state_vec_158_T_3,_state_vec_158_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_159_valid = touch_way_0_valid & touch_set_0 == 9'h9f; // @[Replacement.scala 315:30]
  wire  state_vec_159_left_subtree_state = state_vec_159[1]; // @[package.scala 154:13]
  wire  state_vec_159_right_subtree_state = state_vec_159[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_159_T_3 = state_vec_0_set_left_older ? state_vec_159_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_159_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_159_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_159_T_8 = {state_vec_0_set_left_older,_state_vec_159_T_3,_state_vec_159_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_160_valid = touch_way_0_valid & touch_set_0 == 9'ha0; // @[Replacement.scala 315:30]
  wire  state_vec_160_left_subtree_state = state_vec_160[1]; // @[package.scala 154:13]
  wire  state_vec_160_right_subtree_state = state_vec_160[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_160_T_3 = state_vec_0_set_left_older ? state_vec_160_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_160_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_160_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_160_T_8 = {state_vec_0_set_left_older,_state_vec_160_T_3,_state_vec_160_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_161_valid = touch_way_0_valid & touch_set_0 == 9'ha1; // @[Replacement.scala 315:30]
  wire  state_vec_161_left_subtree_state = state_vec_161[1]; // @[package.scala 154:13]
  wire  state_vec_161_right_subtree_state = state_vec_161[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_161_T_3 = state_vec_0_set_left_older ? state_vec_161_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_161_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_161_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_161_T_8 = {state_vec_0_set_left_older,_state_vec_161_T_3,_state_vec_161_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_162_valid = touch_way_0_valid & touch_set_0 == 9'ha2; // @[Replacement.scala 315:30]
  wire  state_vec_162_left_subtree_state = state_vec_162[1]; // @[package.scala 154:13]
  wire  state_vec_162_right_subtree_state = state_vec_162[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_162_T_3 = state_vec_0_set_left_older ? state_vec_162_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_162_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_162_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_162_T_8 = {state_vec_0_set_left_older,_state_vec_162_T_3,_state_vec_162_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_163_valid = touch_way_0_valid & touch_set_0 == 9'ha3; // @[Replacement.scala 315:30]
  wire  state_vec_163_left_subtree_state = state_vec_163[1]; // @[package.scala 154:13]
  wire  state_vec_163_right_subtree_state = state_vec_163[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_163_T_3 = state_vec_0_set_left_older ? state_vec_163_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_163_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_163_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_163_T_8 = {state_vec_0_set_left_older,_state_vec_163_T_3,_state_vec_163_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_164_valid = touch_way_0_valid & touch_set_0 == 9'ha4; // @[Replacement.scala 315:30]
  wire  state_vec_164_left_subtree_state = state_vec_164[1]; // @[package.scala 154:13]
  wire  state_vec_164_right_subtree_state = state_vec_164[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_164_T_3 = state_vec_0_set_left_older ? state_vec_164_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_164_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_164_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_164_T_8 = {state_vec_0_set_left_older,_state_vec_164_T_3,_state_vec_164_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_165_valid = touch_way_0_valid & touch_set_0 == 9'ha5; // @[Replacement.scala 315:30]
  wire  state_vec_165_left_subtree_state = state_vec_165[1]; // @[package.scala 154:13]
  wire  state_vec_165_right_subtree_state = state_vec_165[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_165_T_3 = state_vec_0_set_left_older ? state_vec_165_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_165_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_165_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_165_T_8 = {state_vec_0_set_left_older,_state_vec_165_T_3,_state_vec_165_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_166_valid = touch_way_0_valid & touch_set_0 == 9'ha6; // @[Replacement.scala 315:30]
  wire  state_vec_166_left_subtree_state = state_vec_166[1]; // @[package.scala 154:13]
  wire  state_vec_166_right_subtree_state = state_vec_166[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_166_T_3 = state_vec_0_set_left_older ? state_vec_166_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_166_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_166_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_166_T_8 = {state_vec_0_set_left_older,_state_vec_166_T_3,_state_vec_166_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_167_valid = touch_way_0_valid & touch_set_0 == 9'ha7; // @[Replacement.scala 315:30]
  wire  state_vec_167_left_subtree_state = state_vec_167[1]; // @[package.scala 154:13]
  wire  state_vec_167_right_subtree_state = state_vec_167[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_167_T_3 = state_vec_0_set_left_older ? state_vec_167_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_167_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_167_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_167_T_8 = {state_vec_0_set_left_older,_state_vec_167_T_3,_state_vec_167_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_168_valid = touch_way_0_valid & touch_set_0 == 9'ha8; // @[Replacement.scala 315:30]
  wire  state_vec_168_left_subtree_state = state_vec_168[1]; // @[package.scala 154:13]
  wire  state_vec_168_right_subtree_state = state_vec_168[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_168_T_3 = state_vec_0_set_left_older ? state_vec_168_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_168_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_168_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_168_T_8 = {state_vec_0_set_left_older,_state_vec_168_T_3,_state_vec_168_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_169_valid = touch_way_0_valid & touch_set_0 == 9'ha9; // @[Replacement.scala 315:30]
  wire  state_vec_169_left_subtree_state = state_vec_169[1]; // @[package.scala 154:13]
  wire  state_vec_169_right_subtree_state = state_vec_169[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_169_T_3 = state_vec_0_set_left_older ? state_vec_169_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_169_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_169_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_169_T_8 = {state_vec_0_set_left_older,_state_vec_169_T_3,_state_vec_169_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_170_valid = touch_way_0_valid & touch_set_0 == 9'haa; // @[Replacement.scala 315:30]
  wire  state_vec_170_left_subtree_state = state_vec_170[1]; // @[package.scala 154:13]
  wire  state_vec_170_right_subtree_state = state_vec_170[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_170_T_3 = state_vec_0_set_left_older ? state_vec_170_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_170_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_170_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_170_T_8 = {state_vec_0_set_left_older,_state_vec_170_T_3,_state_vec_170_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_171_valid = touch_way_0_valid & touch_set_0 == 9'hab; // @[Replacement.scala 315:30]
  wire  state_vec_171_left_subtree_state = state_vec_171[1]; // @[package.scala 154:13]
  wire  state_vec_171_right_subtree_state = state_vec_171[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_171_T_3 = state_vec_0_set_left_older ? state_vec_171_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_171_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_171_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_171_T_8 = {state_vec_0_set_left_older,_state_vec_171_T_3,_state_vec_171_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_172_valid = touch_way_0_valid & touch_set_0 == 9'hac; // @[Replacement.scala 315:30]
  wire  state_vec_172_left_subtree_state = state_vec_172[1]; // @[package.scala 154:13]
  wire  state_vec_172_right_subtree_state = state_vec_172[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_172_T_3 = state_vec_0_set_left_older ? state_vec_172_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_172_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_172_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_172_T_8 = {state_vec_0_set_left_older,_state_vec_172_T_3,_state_vec_172_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_173_valid = touch_way_0_valid & touch_set_0 == 9'had; // @[Replacement.scala 315:30]
  wire  state_vec_173_left_subtree_state = state_vec_173[1]; // @[package.scala 154:13]
  wire  state_vec_173_right_subtree_state = state_vec_173[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_173_T_3 = state_vec_0_set_left_older ? state_vec_173_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_173_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_173_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_173_T_8 = {state_vec_0_set_left_older,_state_vec_173_T_3,_state_vec_173_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_174_valid = touch_way_0_valid & touch_set_0 == 9'hae; // @[Replacement.scala 315:30]
  wire  state_vec_174_left_subtree_state = state_vec_174[1]; // @[package.scala 154:13]
  wire  state_vec_174_right_subtree_state = state_vec_174[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_174_T_3 = state_vec_0_set_left_older ? state_vec_174_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_174_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_174_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_174_T_8 = {state_vec_0_set_left_older,_state_vec_174_T_3,_state_vec_174_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_175_valid = touch_way_0_valid & touch_set_0 == 9'haf; // @[Replacement.scala 315:30]
  wire  state_vec_175_left_subtree_state = state_vec_175[1]; // @[package.scala 154:13]
  wire  state_vec_175_right_subtree_state = state_vec_175[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_175_T_3 = state_vec_0_set_left_older ? state_vec_175_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_175_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_175_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_175_T_8 = {state_vec_0_set_left_older,_state_vec_175_T_3,_state_vec_175_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_176_valid = touch_way_0_valid & touch_set_0 == 9'hb0; // @[Replacement.scala 315:30]
  wire  state_vec_176_left_subtree_state = state_vec_176[1]; // @[package.scala 154:13]
  wire  state_vec_176_right_subtree_state = state_vec_176[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_176_T_3 = state_vec_0_set_left_older ? state_vec_176_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_176_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_176_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_176_T_8 = {state_vec_0_set_left_older,_state_vec_176_T_3,_state_vec_176_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_177_valid = touch_way_0_valid & touch_set_0 == 9'hb1; // @[Replacement.scala 315:30]
  wire  state_vec_177_left_subtree_state = state_vec_177[1]; // @[package.scala 154:13]
  wire  state_vec_177_right_subtree_state = state_vec_177[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_177_T_3 = state_vec_0_set_left_older ? state_vec_177_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_177_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_177_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_177_T_8 = {state_vec_0_set_left_older,_state_vec_177_T_3,_state_vec_177_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_178_valid = touch_way_0_valid & touch_set_0 == 9'hb2; // @[Replacement.scala 315:30]
  wire  state_vec_178_left_subtree_state = state_vec_178[1]; // @[package.scala 154:13]
  wire  state_vec_178_right_subtree_state = state_vec_178[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_178_T_3 = state_vec_0_set_left_older ? state_vec_178_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_178_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_178_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_178_T_8 = {state_vec_0_set_left_older,_state_vec_178_T_3,_state_vec_178_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_179_valid = touch_way_0_valid & touch_set_0 == 9'hb3; // @[Replacement.scala 315:30]
  wire  state_vec_179_left_subtree_state = state_vec_179[1]; // @[package.scala 154:13]
  wire  state_vec_179_right_subtree_state = state_vec_179[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_179_T_3 = state_vec_0_set_left_older ? state_vec_179_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_179_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_179_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_179_T_8 = {state_vec_0_set_left_older,_state_vec_179_T_3,_state_vec_179_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_180_valid = touch_way_0_valid & touch_set_0 == 9'hb4; // @[Replacement.scala 315:30]
  wire  state_vec_180_left_subtree_state = state_vec_180[1]; // @[package.scala 154:13]
  wire  state_vec_180_right_subtree_state = state_vec_180[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_180_T_3 = state_vec_0_set_left_older ? state_vec_180_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_180_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_180_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_180_T_8 = {state_vec_0_set_left_older,_state_vec_180_T_3,_state_vec_180_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_181_valid = touch_way_0_valid & touch_set_0 == 9'hb5; // @[Replacement.scala 315:30]
  wire  state_vec_181_left_subtree_state = state_vec_181[1]; // @[package.scala 154:13]
  wire  state_vec_181_right_subtree_state = state_vec_181[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_181_T_3 = state_vec_0_set_left_older ? state_vec_181_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_181_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_181_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_181_T_8 = {state_vec_0_set_left_older,_state_vec_181_T_3,_state_vec_181_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_182_valid = touch_way_0_valid & touch_set_0 == 9'hb6; // @[Replacement.scala 315:30]
  wire  state_vec_182_left_subtree_state = state_vec_182[1]; // @[package.scala 154:13]
  wire  state_vec_182_right_subtree_state = state_vec_182[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_182_T_3 = state_vec_0_set_left_older ? state_vec_182_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_182_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_182_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_182_T_8 = {state_vec_0_set_left_older,_state_vec_182_T_3,_state_vec_182_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_183_valid = touch_way_0_valid & touch_set_0 == 9'hb7; // @[Replacement.scala 315:30]
  wire  state_vec_183_left_subtree_state = state_vec_183[1]; // @[package.scala 154:13]
  wire  state_vec_183_right_subtree_state = state_vec_183[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_183_T_3 = state_vec_0_set_left_older ? state_vec_183_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_183_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_183_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_183_T_8 = {state_vec_0_set_left_older,_state_vec_183_T_3,_state_vec_183_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_184_valid = touch_way_0_valid & touch_set_0 == 9'hb8; // @[Replacement.scala 315:30]
  wire  state_vec_184_left_subtree_state = state_vec_184[1]; // @[package.scala 154:13]
  wire  state_vec_184_right_subtree_state = state_vec_184[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_184_T_3 = state_vec_0_set_left_older ? state_vec_184_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_184_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_184_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_184_T_8 = {state_vec_0_set_left_older,_state_vec_184_T_3,_state_vec_184_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_185_valid = touch_way_0_valid & touch_set_0 == 9'hb9; // @[Replacement.scala 315:30]
  wire  state_vec_185_left_subtree_state = state_vec_185[1]; // @[package.scala 154:13]
  wire  state_vec_185_right_subtree_state = state_vec_185[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_185_T_3 = state_vec_0_set_left_older ? state_vec_185_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_185_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_185_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_185_T_8 = {state_vec_0_set_left_older,_state_vec_185_T_3,_state_vec_185_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_186_valid = touch_way_0_valid & touch_set_0 == 9'hba; // @[Replacement.scala 315:30]
  wire  state_vec_186_left_subtree_state = state_vec_186[1]; // @[package.scala 154:13]
  wire  state_vec_186_right_subtree_state = state_vec_186[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_186_T_3 = state_vec_0_set_left_older ? state_vec_186_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_186_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_186_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_186_T_8 = {state_vec_0_set_left_older,_state_vec_186_T_3,_state_vec_186_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_187_valid = touch_way_0_valid & touch_set_0 == 9'hbb; // @[Replacement.scala 315:30]
  wire  state_vec_187_left_subtree_state = state_vec_187[1]; // @[package.scala 154:13]
  wire  state_vec_187_right_subtree_state = state_vec_187[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_187_T_3 = state_vec_0_set_left_older ? state_vec_187_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_187_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_187_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_187_T_8 = {state_vec_0_set_left_older,_state_vec_187_T_3,_state_vec_187_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_188_valid = touch_way_0_valid & touch_set_0 == 9'hbc; // @[Replacement.scala 315:30]
  wire  state_vec_188_left_subtree_state = state_vec_188[1]; // @[package.scala 154:13]
  wire  state_vec_188_right_subtree_state = state_vec_188[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_188_T_3 = state_vec_0_set_left_older ? state_vec_188_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_188_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_188_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_188_T_8 = {state_vec_0_set_left_older,_state_vec_188_T_3,_state_vec_188_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_189_valid = touch_way_0_valid & touch_set_0 == 9'hbd; // @[Replacement.scala 315:30]
  wire  state_vec_189_left_subtree_state = state_vec_189[1]; // @[package.scala 154:13]
  wire  state_vec_189_right_subtree_state = state_vec_189[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_189_T_3 = state_vec_0_set_left_older ? state_vec_189_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_189_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_189_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_189_T_8 = {state_vec_0_set_left_older,_state_vec_189_T_3,_state_vec_189_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_190_valid = touch_way_0_valid & touch_set_0 == 9'hbe; // @[Replacement.scala 315:30]
  wire  state_vec_190_left_subtree_state = state_vec_190[1]; // @[package.scala 154:13]
  wire  state_vec_190_right_subtree_state = state_vec_190[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_190_T_3 = state_vec_0_set_left_older ? state_vec_190_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_190_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_190_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_190_T_8 = {state_vec_0_set_left_older,_state_vec_190_T_3,_state_vec_190_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_191_valid = touch_way_0_valid & touch_set_0 == 9'hbf; // @[Replacement.scala 315:30]
  wire  state_vec_191_left_subtree_state = state_vec_191[1]; // @[package.scala 154:13]
  wire  state_vec_191_right_subtree_state = state_vec_191[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_191_T_3 = state_vec_0_set_left_older ? state_vec_191_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_191_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_191_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_191_T_8 = {state_vec_0_set_left_older,_state_vec_191_T_3,_state_vec_191_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_192_valid = touch_way_0_valid & touch_set_0 == 9'hc0; // @[Replacement.scala 315:30]
  wire  state_vec_192_left_subtree_state = state_vec_192[1]; // @[package.scala 154:13]
  wire  state_vec_192_right_subtree_state = state_vec_192[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_192_T_3 = state_vec_0_set_left_older ? state_vec_192_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_192_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_192_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_192_T_8 = {state_vec_0_set_left_older,_state_vec_192_T_3,_state_vec_192_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_193_valid = touch_way_0_valid & touch_set_0 == 9'hc1; // @[Replacement.scala 315:30]
  wire  state_vec_193_left_subtree_state = state_vec_193[1]; // @[package.scala 154:13]
  wire  state_vec_193_right_subtree_state = state_vec_193[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_193_T_3 = state_vec_0_set_left_older ? state_vec_193_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_193_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_193_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_193_T_8 = {state_vec_0_set_left_older,_state_vec_193_T_3,_state_vec_193_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_194_valid = touch_way_0_valid & touch_set_0 == 9'hc2; // @[Replacement.scala 315:30]
  wire  state_vec_194_left_subtree_state = state_vec_194[1]; // @[package.scala 154:13]
  wire  state_vec_194_right_subtree_state = state_vec_194[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_194_T_3 = state_vec_0_set_left_older ? state_vec_194_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_194_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_194_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_194_T_8 = {state_vec_0_set_left_older,_state_vec_194_T_3,_state_vec_194_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_195_valid = touch_way_0_valid & touch_set_0 == 9'hc3; // @[Replacement.scala 315:30]
  wire  state_vec_195_left_subtree_state = state_vec_195[1]; // @[package.scala 154:13]
  wire  state_vec_195_right_subtree_state = state_vec_195[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_195_T_3 = state_vec_0_set_left_older ? state_vec_195_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_195_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_195_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_195_T_8 = {state_vec_0_set_left_older,_state_vec_195_T_3,_state_vec_195_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_196_valid = touch_way_0_valid & touch_set_0 == 9'hc4; // @[Replacement.scala 315:30]
  wire  state_vec_196_left_subtree_state = state_vec_196[1]; // @[package.scala 154:13]
  wire  state_vec_196_right_subtree_state = state_vec_196[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_196_T_3 = state_vec_0_set_left_older ? state_vec_196_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_196_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_196_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_196_T_8 = {state_vec_0_set_left_older,_state_vec_196_T_3,_state_vec_196_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_197_valid = touch_way_0_valid & touch_set_0 == 9'hc5; // @[Replacement.scala 315:30]
  wire  state_vec_197_left_subtree_state = state_vec_197[1]; // @[package.scala 154:13]
  wire  state_vec_197_right_subtree_state = state_vec_197[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_197_T_3 = state_vec_0_set_left_older ? state_vec_197_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_197_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_197_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_197_T_8 = {state_vec_0_set_left_older,_state_vec_197_T_3,_state_vec_197_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_198_valid = touch_way_0_valid & touch_set_0 == 9'hc6; // @[Replacement.scala 315:30]
  wire  state_vec_198_left_subtree_state = state_vec_198[1]; // @[package.scala 154:13]
  wire  state_vec_198_right_subtree_state = state_vec_198[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_198_T_3 = state_vec_0_set_left_older ? state_vec_198_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_198_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_198_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_198_T_8 = {state_vec_0_set_left_older,_state_vec_198_T_3,_state_vec_198_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_199_valid = touch_way_0_valid & touch_set_0 == 9'hc7; // @[Replacement.scala 315:30]
  wire  state_vec_199_left_subtree_state = state_vec_199[1]; // @[package.scala 154:13]
  wire  state_vec_199_right_subtree_state = state_vec_199[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_199_T_3 = state_vec_0_set_left_older ? state_vec_199_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_199_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_199_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_199_T_8 = {state_vec_0_set_left_older,_state_vec_199_T_3,_state_vec_199_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_200_valid = touch_way_0_valid & touch_set_0 == 9'hc8; // @[Replacement.scala 315:30]
  wire  state_vec_200_left_subtree_state = state_vec_200[1]; // @[package.scala 154:13]
  wire  state_vec_200_right_subtree_state = state_vec_200[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_200_T_3 = state_vec_0_set_left_older ? state_vec_200_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_200_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_200_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_200_T_8 = {state_vec_0_set_left_older,_state_vec_200_T_3,_state_vec_200_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_201_valid = touch_way_0_valid & touch_set_0 == 9'hc9; // @[Replacement.scala 315:30]
  wire  state_vec_201_left_subtree_state = state_vec_201[1]; // @[package.scala 154:13]
  wire  state_vec_201_right_subtree_state = state_vec_201[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_201_T_3 = state_vec_0_set_left_older ? state_vec_201_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_201_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_201_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_201_T_8 = {state_vec_0_set_left_older,_state_vec_201_T_3,_state_vec_201_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_202_valid = touch_way_0_valid & touch_set_0 == 9'hca; // @[Replacement.scala 315:30]
  wire  state_vec_202_left_subtree_state = state_vec_202[1]; // @[package.scala 154:13]
  wire  state_vec_202_right_subtree_state = state_vec_202[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_202_T_3 = state_vec_0_set_left_older ? state_vec_202_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_202_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_202_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_202_T_8 = {state_vec_0_set_left_older,_state_vec_202_T_3,_state_vec_202_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_203_valid = touch_way_0_valid & touch_set_0 == 9'hcb; // @[Replacement.scala 315:30]
  wire  state_vec_203_left_subtree_state = state_vec_203[1]; // @[package.scala 154:13]
  wire  state_vec_203_right_subtree_state = state_vec_203[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_203_T_3 = state_vec_0_set_left_older ? state_vec_203_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_203_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_203_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_203_T_8 = {state_vec_0_set_left_older,_state_vec_203_T_3,_state_vec_203_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_204_valid = touch_way_0_valid & touch_set_0 == 9'hcc; // @[Replacement.scala 315:30]
  wire  state_vec_204_left_subtree_state = state_vec_204[1]; // @[package.scala 154:13]
  wire  state_vec_204_right_subtree_state = state_vec_204[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_204_T_3 = state_vec_0_set_left_older ? state_vec_204_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_204_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_204_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_204_T_8 = {state_vec_0_set_left_older,_state_vec_204_T_3,_state_vec_204_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_205_valid = touch_way_0_valid & touch_set_0 == 9'hcd; // @[Replacement.scala 315:30]
  wire  state_vec_205_left_subtree_state = state_vec_205[1]; // @[package.scala 154:13]
  wire  state_vec_205_right_subtree_state = state_vec_205[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_205_T_3 = state_vec_0_set_left_older ? state_vec_205_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_205_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_205_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_205_T_8 = {state_vec_0_set_left_older,_state_vec_205_T_3,_state_vec_205_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_206_valid = touch_way_0_valid & touch_set_0 == 9'hce; // @[Replacement.scala 315:30]
  wire  state_vec_206_left_subtree_state = state_vec_206[1]; // @[package.scala 154:13]
  wire  state_vec_206_right_subtree_state = state_vec_206[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_206_T_3 = state_vec_0_set_left_older ? state_vec_206_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_206_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_206_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_206_T_8 = {state_vec_0_set_left_older,_state_vec_206_T_3,_state_vec_206_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_207_valid = touch_way_0_valid & touch_set_0 == 9'hcf; // @[Replacement.scala 315:30]
  wire  state_vec_207_left_subtree_state = state_vec_207[1]; // @[package.scala 154:13]
  wire  state_vec_207_right_subtree_state = state_vec_207[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_207_T_3 = state_vec_0_set_left_older ? state_vec_207_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_207_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_207_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_207_T_8 = {state_vec_0_set_left_older,_state_vec_207_T_3,_state_vec_207_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_208_valid = touch_way_0_valid & touch_set_0 == 9'hd0; // @[Replacement.scala 315:30]
  wire  state_vec_208_left_subtree_state = state_vec_208[1]; // @[package.scala 154:13]
  wire  state_vec_208_right_subtree_state = state_vec_208[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_208_T_3 = state_vec_0_set_left_older ? state_vec_208_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_208_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_208_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_208_T_8 = {state_vec_0_set_left_older,_state_vec_208_T_3,_state_vec_208_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_209_valid = touch_way_0_valid & touch_set_0 == 9'hd1; // @[Replacement.scala 315:30]
  wire  state_vec_209_left_subtree_state = state_vec_209[1]; // @[package.scala 154:13]
  wire  state_vec_209_right_subtree_state = state_vec_209[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_209_T_3 = state_vec_0_set_left_older ? state_vec_209_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_209_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_209_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_209_T_8 = {state_vec_0_set_left_older,_state_vec_209_T_3,_state_vec_209_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_210_valid = touch_way_0_valid & touch_set_0 == 9'hd2; // @[Replacement.scala 315:30]
  wire  state_vec_210_left_subtree_state = state_vec_210[1]; // @[package.scala 154:13]
  wire  state_vec_210_right_subtree_state = state_vec_210[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_210_T_3 = state_vec_0_set_left_older ? state_vec_210_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_210_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_210_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_210_T_8 = {state_vec_0_set_left_older,_state_vec_210_T_3,_state_vec_210_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_211_valid = touch_way_0_valid & touch_set_0 == 9'hd3; // @[Replacement.scala 315:30]
  wire  state_vec_211_left_subtree_state = state_vec_211[1]; // @[package.scala 154:13]
  wire  state_vec_211_right_subtree_state = state_vec_211[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_211_T_3 = state_vec_0_set_left_older ? state_vec_211_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_211_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_211_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_211_T_8 = {state_vec_0_set_left_older,_state_vec_211_T_3,_state_vec_211_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_212_valid = touch_way_0_valid & touch_set_0 == 9'hd4; // @[Replacement.scala 315:30]
  wire  state_vec_212_left_subtree_state = state_vec_212[1]; // @[package.scala 154:13]
  wire  state_vec_212_right_subtree_state = state_vec_212[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_212_T_3 = state_vec_0_set_left_older ? state_vec_212_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_212_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_212_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_212_T_8 = {state_vec_0_set_left_older,_state_vec_212_T_3,_state_vec_212_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_213_valid = touch_way_0_valid & touch_set_0 == 9'hd5; // @[Replacement.scala 315:30]
  wire  state_vec_213_left_subtree_state = state_vec_213[1]; // @[package.scala 154:13]
  wire  state_vec_213_right_subtree_state = state_vec_213[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_213_T_3 = state_vec_0_set_left_older ? state_vec_213_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_213_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_213_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_213_T_8 = {state_vec_0_set_left_older,_state_vec_213_T_3,_state_vec_213_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_214_valid = touch_way_0_valid & touch_set_0 == 9'hd6; // @[Replacement.scala 315:30]
  wire  state_vec_214_left_subtree_state = state_vec_214[1]; // @[package.scala 154:13]
  wire  state_vec_214_right_subtree_state = state_vec_214[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_214_T_3 = state_vec_0_set_left_older ? state_vec_214_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_214_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_214_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_214_T_8 = {state_vec_0_set_left_older,_state_vec_214_T_3,_state_vec_214_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_215_valid = touch_way_0_valid & touch_set_0 == 9'hd7; // @[Replacement.scala 315:30]
  wire  state_vec_215_left_subtree_state = state_vec_215[1]; // @[package.scala 154:13]
  wire  state_vec_215_right_subtree_state = state_vec_215[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_215_T_3 = state_vec_0_set_left_older ? state_vec_215_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_215_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_215_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_215_T_8 = {state_vec_0_set_left_older,_state_vec_215_T_3,_state_vec_215_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_216_valid = touch_way_0_valid & touch_set_0 == 9'hd8; // @[Replacement.scala 315:30]
  wire  state_vec_216_left_subtree_state = state_vec_216[1]; // @[package.scala 154:13]
  wire  state_vec_216_right_subtree_state = state_vec_216[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_216_T_3 = state_vec_0_set_left_older ? state_vec_216_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_216_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_216_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_216_T_8 = {state_vec_0_set_left_older,_state_vec_216_T_3,_state_vec_216_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_217_valid = touch_way_0_valid & touch_set_0 == 9'hd9; // @[Replacement.scala 315:30]
  wire  state_vec_217_left_subtree_state = state_vec_217[1]; // @[package.scala 154:13]
  wire  state_vec_217_right_subtree_state = state_vec_217[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_217_T_3 = state_vec_0_set_left_older ? state_vec_217_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_217_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_217_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_217_T_8 = {state_vec_0_set_left_older,_state_vec_217_T_3,_state_vec_217_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_218_valid = touch_way_0_valid & touch_set_0 == 9'hda; // @[Replacement.scala 315:30]
  wire  state_vec_218_left_subtree_state = state_vec_218[1]; // @[package.scala 154:13]
  wire  state_vec_218_right_subtree_state = state_vec_218[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_218_T_3 = state_vec_0_set_left_older ? state_vec_218_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_218_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_218_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_218_T_8 = {state_vec_0_set_left_older,_state_vec_218_T_3,_state_vec_218_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_219_valid = touch_way_0_valid & touch_set_0 == 9'hdb; // @[Replacement.scala 315:30]
  wire  state_vec_219_left_subtree_state = state_vec_219[1]; // @[package.scala 154:13]
  wire  state_vec_219_right_subtree_state = state_vec_219[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_219_T_3 = state_vec_0_set_left_older ? state_vec_219_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_219_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_219_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_219_T_8 = {state_vec_0_set_left_older,_state_vec_219_T_3,_state_vec_219_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_220_valid = touch_way_0_valid & touch_set_0 == 9'hdc; // @[Replacement.scala 315:30]
  wire  state_vec_220_left_subtree_state = state_vec_220[1]; // @[package.scala 154:13]
  wire  state_vec_220_right_subtree_state = state_vec_220[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_220_T_3 = state_vec_0_set_left_older ? state_vec_220_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_220_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_220_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_220_T_8 = {state_vec_0_set_left_older,_state_vec_220_T_3,_state_vec_220_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_221_valid = touch_way_0_valid & touch_set_0 == 9'hdd; // @[Replacement.scala 315:30]
  wire  state_vec_221_left_subtree_state = state_vec_221[1]; // @[package.scala 154:13]
  wire  state_vec_221_right_subtree_state = state_vec_221[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_221_T_3 = state_vec_0_set_left_older ? state_vec_221_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_221_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_221_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_221_T_8 = {state_vec_0_set_left_older,_state_vec_221_T_3,_state_vec_221_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_222_valid = touch_way_0_valid & touch_set_0 == 9'hde; // @[Replacement.scala 315:30]
  wire  state_vec_222_left_subtree_state = state_vec_222[1]; // @[package.scala 154:13]
  wire  state_vec_222_right_subtree_state = state_vec_222[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_222_T_3 = state_vec_0_set_left_older ? state_vec_222_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_222_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_222_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_222_T_8 = {state_vec_0_set_left_older,_state_vec_222_T_3,_state_vec_222_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_223_valid = touch_way_0_valid & touch_set_0 == 9'hdf; // @[Replacement.scala 315:30]
  wire  state_vec_223_left_subtree_state = state_vec_223[1]; // @[package.scala 154:13]
  wire  state_vec_223_right_subtree_state = state_vec_223[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_223_T_3 = state_vec_0_set_left_older ? state_vec_223_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_223_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_223_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_223_T_8 = {state_vec_0_set_left_older,_state_vec_223_T_3,_state_vec_223_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_224_valid = touch_way_0_valid & touch_set_0 == 9'he0; // @[Replacement.scala 315:30]
  wire  state_vec_224_left_subtree_state = state_vec_224[1]; // @[package.scala 154:13]
  wire  state_vec_224_right_subtree_state = state_vec_224[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_224_T_3 = state_vec_0_set_left_older ? state_vec_224_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_224_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_224_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_224_T_8 = {state_vec_0_set_left_older,_state_vec_224_T_3,_state_vec_224_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_225_valid = touch_way_0_valid & touch_set_0 == 9'he1; // @[Replacement.scala 315:30]
  wire  state_vec_225_left_subtree_state = state_vec_225[1]; // @[package.scala 154:13]
  wire  state_vec_225_right_subtree_state = state_vec_225[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_225_T_3 = state_vec_0_set_left_older ? state_vec_225_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_225_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_225_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_225_T_8 = {state_vec_0_set_left_older,_state_vec_225_T_3,_state_vec_225_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_226_valid = touch_way_0_valid & touch_set_0 == 9'he2; // @[Replacement.scala 315:30]
  wire  state_vec_226_left_subtree_state = state_vec_226[1]; // @[package.scala 154:13]
  wire  state_vec_226_right_subtree_state = state_vec_226[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_226_T_3 = state_vec_0_set_left_older ? state_vec_226_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_226_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_226_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_226_T_8 = {state_vec_0_set_left_older,_state_vec_226_T_3,_state_vec_226_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_227_valid = touch_way_0_valid & touch_set_0 == 9'he3; // @[Replacement.scala 315:30]
  wire  state_vec_227_left_subtree_state = state_vec_227[1]; // @[package.scala 154:13]
  wire  state_vec_227_right_subtree_state = state_vec_227[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_227_T_3 = state_vec_0_set_left_older ? state_vec_227_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_227_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_227_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_227_T_8 = {state_vec_0_set_left_older,_state_vec_227_T_3,_state_vec_227_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_228_valid = touch_way_0_valid & touch_set_0 == 9'he4; // @[Replacement.scala 315:30]
  wire  state_vec_228_left_subtree_state = state_vec_228[1]; // @[package.scala 154:13]
  wire  state_vec_228_right_subtree_state = state_vec_228[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_228_T_3 = state_vec_0_set_left_older ? state_vec_228_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_228_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_228_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_228_T_8 = {state_vec_0_set_left_older,_state_vec_228_T_3,_state_vec_228_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_229_valid = touch_way_0_valid & touch_set_0 == 9'he5; // @[Replacement.scala 315:30]
  wire  state_vec_229_left_subtree_state = state_vec_229[1]; // @[package.scala 154:13]
  wire  state_vec_229_right_subtree_state = state_vec_229[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_229_T_3 = state_vec_0_set_left_older ? state_vec_229_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_229_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_229_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_229_T_8 = {state_vec_0_set_left_older,_state_vec_229_T_3,_state_vec_229_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_230_valid = touch_way_0_valid & touch_set_0 == 9'he6; // @[Replacement.scala 315:30]
  wire  state_vec_230_left_subtree_state = state_vec_230[1]; // @[package.scala 154:13]
  wire  state_vec_230_right_subtree_state = state_vec_230[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_230_T_3 = state_vec_0_set_left_older ? state_vec_230_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_230_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_230_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_230_T_8 = {state_vec_0_set_left_older,_state_vec_230_T_3,_state_vec_230_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_231_valid = touch_way_0_valid & touch_set_0 == 9'he7; // @[Replacement.scala 315:30]
  wire  state_vec_231_left_subtree_state = state_vec_231[1]; // @[package.scala 154:13]
  wire  state_vec_231_right_subtree_state = state_vec_231[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_231_T_3 = state_vec_0_set_left_older ? state_vec_231_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_231_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_231_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_231_T_8 = {state_vec_0_set_left_older,_state_vec_231_T_3,_state_vec_231_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_232_valid = touch_way_0_valid & touch_set_0 == 9'he8; // @[Replacement.scala 315:30]
  wire  state_vec_232_left_subtree_state = state_vec_232[1]; // @[package.scala 154:13]
  wire  state_vec_232_right_subtree_state = state_vec_232[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_232_T_3 = state_vec_0_set_left_older ? state_vec_232_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_232_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_232_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_232_T_8 = {state_vec_0_set_left_older,_state_vec_232_T_3,_state_vec_232_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_233_valid = touch_way_0_valid & touch_set_0 == 9'he9; // @[Replacement.scala 315:30]
  wire  state_vec_233_left_subtree_state = state_vec_233[1]; // @[package.scala 154:13]
  wire  state_vec_233_right_subtree_state = state_vec_233[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_233_T_3 = state_vec_0_set_left_older ? state_vec_233_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_233_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_233_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_233_T_8 = {state_vec_0_set_left_older,_state_vec_233_T_3,_state_vec_233_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_234_valid = touch_way_0_valid & touch_set_0 == 9'hea; // @[Replacement.scala 315:30]
  wire  state_vec_234_left_subtree_state = state_vec_234[1]; // @[package.scala 154:13]
  wire  state_vec_234_right_subtree_state = state_vec_234[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_234_T_3 = state_vec_0_set_left_older ? state_vec_234_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_234_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_234_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_234_T_8 = {state_vec_0_set_left_older,_state_vec_234_T_3,_state_vec_234_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_235_valid = touch_way_0_valid & touch_set_0 == 9'heb; // @[Replacement.scala 315:30]
  wire  state_vec_235_left_subtree_state = state_vec_235[1]; // @[package.scala 154:13]
  wire  state_vec_235_right_subtree_state = state_vec_235[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_235_T_3 = state_vec_0_set_left_older ? state_vec_235_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_235_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_235_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_235_T_8 = {state_vec_0_set_left_older,_state_vec_235_T_3,_state_vec_235_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_236_valid = touch_way_0_valid & touch_set_0 == 9'hec; // @[Replacement.scala 315:30]
  wire  state_vec_236_left_subtree_state = state_vec_236[1]; // @[package.scala 154:13]
  wire  state_vec_236_right_subtree_state = state_vec_236[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_236_T_3 = state_vec_0_set_left_older ? state_vec_236_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_236_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_236_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_236_T_8 = {state_vec_0_set_left_older,_state_vec_236_T_3,_state_vec_236_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_237_valid = touch_way_0_valid & touch_set_0 == 9'hed; // @[Replacement.scala 315:30]
  wire  state_vec_237_left_subtree_state = state_vec_237[1]; // @[package.scala 154:13]
  wire  state_vec_237_right_subtree_state = state_vec_237[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_237_T_3 = state_vec_0_set_left_older ? state_vec_237_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_237_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_237_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_237_T_8 = {state_vec_0_set_left_older,_state_vec_237_T_3,_state_vec_237_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_238_valid = touch_way_0_valid & touch_set_0 == 9'hee; // @[Replacement.scala 315:30]
  wire  state_vec_238_left_subtree_state = state_vec_238[1]; // @[package.scala 154:13]
  wire  state_vec_238_right_subtree_state = state_vec_238[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_238_T_3 = state_vec_0_set_left_older ? state_vec_238_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_238_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_238_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_238_T_8 = {state_vec_0_set_left_older,_state_vec_238_T_3,_state_vec_238_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_239_valid = touch_way_0_valid & touch_set_0 == 9'hef; // @[Replacement.scala 315:30]
  wire  state_vec_239_left_subtree_state = state_vec_239[1]; // @[package.scala 154:13]
  wire  state_vec_239_right_subtree_state = state_vec_239[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_239_T_3 = state_vec_0_set_left_older ? state_vec_239_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_239_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_239_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_239_T_8 = {state_vec_0_set_left_older,_state_vec_239_T_3,_state_vec_239_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_240_valid = touch_way_0_valid & touch_set_0 == 9'hf0; // @[Replacement.scala 315:30]
  wire  state_vec_240_left_subtree_state = state_vec_240[1]; // @[package.scala 154:13]
  wire  state_vec_240_right_subtree_state = state_vec_240[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_240_T_3 = state_vec_0_set_left_older ? state_vec_240_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_240_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_240_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_240_T_8 = {state_vec_0_set_left_older,_state_vec_240_T_3,_state_vec_240_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_241_valid = touch_way_0_valid & touch_set_0 == 9'hf1; // @[Replacement.scala 315:30]
  wire  state_vec_241_left_subtree_state = state_vec_241[1]; // @[package.scala 154:13]
  wire  state_vec_241_right_subtree_state = state_vec_241[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_241_T_3 = state_vec_0_set_left_older ? state_vec_241_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_241_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_241_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_241_T_8 = {state_vec_0_set_left_older,_state_vec_241_T_3,_state_vec_241_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_242_valid = touch_way_0_valid & touch_set_0 == 9'hf2; // @[Replacement.scala 315:30]
  wire  state_vec_242_left_subtree_state = state_vec_242[1]; // @[package.scala 154:13]
  wire  state_vec_242_right_subtree_state = state_vec_242[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_242_T_3 = state_vec_0_set_left_older ? state_vec_242_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_242_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_242_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_242_T_8 = {state_vec_0_set_left_older,_state_vec_242_T_3,_state_vec_242_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_243_valid = touch_way_0_valid & touch_set_0 == 9'hf3; // @[Replacement.scala 315:30]
  wire  state_vec_243_left_subtree_state = state_vec_243[1]; // @[package.scala 154:13]
  wire  state_vec_243_right_subtree_state = state_vec_243[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_243_T_3 = state_vec_0_set_left_older ? state_vec_243_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_243_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_243_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_243_T_8 = {state_vec_0_set_left_older,_state_vec_243_T_3,_state_vec_243_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_244_valid = touch_way_0_valid & touch_set_0 == 9'hf4; // @[Replacement.scala 315:30]
  wire  state_vec_244_left_subtree_state = state_vec_244[1]; // @[package.scala 154:13]
  wire  state_vec_244_right_subtree_state = state_vec_244[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_244_T_3 = state_vec_0_set_left_older ? state_vec_244_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_244_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_244_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_244_T_8 = {state_vec_0_set_left_older,_state_vec_244_T_3,_state_vec_244_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_245_valid = touch_way_0_valid & touch_set_0 == 9'hf5; // @[Replacement.scala 315:30]
  wire  state_vec_245_left_subtree_state = state_vec_245[1]; // @[package.scala 154:13]
  wire  state_vec_245_right_subtree_state = state_vec_245[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_245_T_3 = state_vec_0_set_left_older ? state_vec_245_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_245_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_245_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_245_T_8 = {state_vec_0_set_left_older,_state_vec_245_T_3,_state_vec_245_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_246_valid = touch_way_0_valid & touch_set_0 == 9'hf6; // @[Replacement.scala 315:30]
  wire  state_vec_246_left_subtree_state = state_vec_246[1]; // @[package.scala 154:13]
  wire  state_vec_246_right_subtree_state = state_vec_246[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_246_T_3 = state_vec_0_set_left_older ? state_vec_246_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_246_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_246_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_246_T_8 = {state_vec_0_set_left_older,_state_vec_246_T_3,_state_vec_246_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_247_valid = touch_way_0_valid & touch_set_0 == 9'hf7; // @[Replacement.scala 315:30]
  wire  state_vec_247_left_subtree_state = state_vec_247[1]; // @[package.scala 154:13]
  wire  state_vec_247_right_subtree_state = state_vec_247[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_247_T_3 = state_vec_0_set_left_older ? state_vec_247_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_247_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_247_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_247_T_8 = {state_vec_0_set_left_older,_state_vec_247_T_3,_state_vec_247_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_248_valid = touch_way_0_valid & touch_set_0 == 9'hf8; // @[Replacement.scala 315:30]
  wire  state_vec_248_left_subtree_state = state_vec_248[1]; // @[package.scala 154:13]
  wire  state_vec_248_right_subtree_state = state_vec_248[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_248_T_3 = state_vec_0_set_left_older ? state_vec_248_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_248_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_248_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_248_T_8 = {state_vec_0_set_left_older,_state_vec_248_T_3,_state_vec_248_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_249_valid = touch_way_0_valid & touch_set_0 == 9'hf9; // @[Replacement.scala 315:30]
  wire  state_vec_249_left_subtree_state = state_vec_249[1]; // @[package.scala 154:13]
  wire  state_vec_249_right_subtree_state = state_vec_249[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_249_T_3 = state_vec_0_set_left_older ? state_vec_249_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_249_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_249_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_249_T_8 = {state_vec_0_set_left_older,_state_vec_249_T_3,_state_vec_249_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_250_valid = touch_way_0_valid & touch_set_0 == 9'hfa; // @[Replacement.scala 315:30]
  wire  state_vec_250_left_subtree_state = state_vec_250[1]; // @[package.scala 154:13]
  wire  state_vec_250_right_subtree_state = state_vec_250[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_250_T_3 = state_vec_0_set_left_older ? state_vec_250_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_250_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_250_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_250_T_8 = {state_vec_0_set_left_older,_state_vec_250_T_3,_state_vec_250_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_251_valid = touch_way_0_valid & touch_set_0 == 9'hfb; // @[Replacement.scala 315:30]
  wire  state_vec_251_left_subtree_state = state_vec_251[1]; // @[package.scala 154:13]
  wire  state_vec_251_right_subtree_state = state_vec_251[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_251_T_3 = state_vec_0_set_left_older ? state_vec_251_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_251_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_251_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_251_T_8 = {state_vec_0_set_left_older,_state_vec_251_T_3,_state_vec_251_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_252_valid = touch_way_0_valid & touch_set_0 == 9'hfc; // @[Replacement.scala 315:30]
  wire  state_vec_252_left_subtree_state = state_vec_252[1]; // @[package.scala 154:13]
  wire  state_vec_252_right_subtree_state = state_vec_252[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_252_T_3 = state_vec_0_set_left_older ? state_vec_252_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_252_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_252_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_252_T_8 = {state_vec_0_set_left_older,_state_vec_252_T_3,_state_vec_252_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_253_valid = touch_way_0_valid & touch_set_0 == 9'hfd; // @[Replacement.scala 315:30]
  wire  state_vec_253_left_subtree_state = state_vec_253[1]; // @[package.scala 154:13]
  wire  state_vec_253_right_subtree_state = state_vec_253[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_253_T_3 = state_vec_0_set_left_older ? state_vec_253_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_253_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_253_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_253_T_8 = {state_vec_0_set_left_older,_state_vec_253_T_3,_state_vec_253_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_254_valid = touch_way_0_valid & touch_set_0 == 9'hfe; // @[Replacement.scala 315:30]
  wire  state_vec_254_left_subtree_state = state_vec_254[1]; // @[package.scala 154:13]
  wire  state_vec_254_right_subtree_state = state_vec_254[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_254_T_3 = state_vec_0_set_left_older ? state_vec_254_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_254_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_254_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_254_T_8 = {state_vec_0_set_left_older,_state_vec_254_T_3,_state_vec_254_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_255_valid = touch_way_0_valid & touch_set_0 == 9'hff; // @[Replacement.scala 315:30]
  wire  state_vec_255_left_subtree_state = state_vec_255[1]; // @[package.scala 154:13]
  wire  state_vec_255_right_subtree_state = state_vec_255[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_255_T_3 = state_vec_0_set_left_older ? state_vec_255_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_255_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_255_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_255_T_8 = {state_vec_0_set_left_older,_state_vec_255_T_3,_state_vec_255_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_256_valid = touch_way_0_valid & touch_set_0 == 9'h100; // @[Replacement.scala 315:30]
  wire  state_vec_256_left_subtree_state = state_vec_256[1]; // @[package.scala 154:13]
  wire  state_vec_256_right_subtree_state = state_vec_256[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_256_T_3 = state_vec_0_set_left_older ? state_vec_256_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_256_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_256_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_256_T_8 = {state_vec_0_set_left_older,_state_vec_256_T_3,_state_vec_256_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_257_valid = touch_way_0_valid & touch_set_0 == 9'h101; // @[Replacement.scala 315:30]
  wire  state_vec_257_left_subtree_state = state_vec_257[1]; // @[package.scala 154:13]
  wire  state_vec_257_right_subtree_state = state_vec_257[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_257_T_3 = state_vec_0_set_left_older ? state_vec_257_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_257_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_257_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_257_T_8 = {state_vec_0_set_left_older,_state_vec_257_T_3,_state_vec_257_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_258_valid = touch_way_0_valid & touch_set_0 == 9'h102; // @[Replacement.scala 315:30]
  wire  state_vec_258_left_subtree_state = state_vec_258[1]; // @[package.scala 154:13]
  wire  state_vec_258_right_subtree_state = state_vec_258[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_258_T_3 = state_vec_0_set_left_older ? state_vec_258_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_258_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_258_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_258_T_8 = {state_vec_0_set_left_older,_state_vec_258_T_3,_state_vec_258_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_259_valid = touch_way_0_valid & touch_set_0 == 9'h103; // @[Replacement.scala 315:30]
  wire  state_vec_259_left_subtree_state = state_vec_259[1]; // @[package.scala 154:13]
  wire  state_vec_259_right_subtree_state = state_vec_259[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_259_T_3 = state_vec_0_set_left_older ? state_vec_259_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_259_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_259_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_259_T_8 = {state_vec_0_set_left_older,_state_vec_259_T_3,_state_vec_259_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_260_valid = touch_way_0_valid & touch_set_0 == 9'h104; // @[Replacement.scala 315:30]
  wire  state_vec_260_left_subtree_state = state_vec_260[1]; // @[package.scala 154:13]
  wire  state_vec_260_right_subtree_state = state_vec_260[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_260_T_3 = state_vec_0_set_left_older ? state_vec_260_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_260_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_260_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_260_T_8 = {state_vec_0_set_left_older,_state_vec_260_T_3,_state_vec_260_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_261_valid = touch_way_0_valid & touch_set_0 == 9'h105; // @[Replacement.scala 315:30]
  wire  state_vec_261_left_subtree_state = state_vec_261[1]; // @[package.scala 154:13]
  wire  state_vec_261_right_subtree_state = state_vec_261[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_261_T_3 = state_vec_0_set_left_older ? state_vec_261_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_261_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_261_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_261_T_8 = {state_vec_0_set_left_older,_state_vec_261_T_3,_state_vec_261_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_262_valid = touch_way_0_valid & touch_set_0 == 9'h106; // @[Replacement.scala 315:30]
  wire  state_vec_262_left_subtree_state = state_vec_262[1]; // @[package.scala 154:13]
  wire  state_vec_262_right_subtree_state = state_vec_262[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_262_T_3 = state_vec_0_set_left_older ? state_vec_262_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_262_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_262_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_262_T_8 = {state_vec_0_set_left_older,_state_vec_262_T_3,_state_vec_262_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_263_valid = touch_way_0_valid & touch_set_0 == 9'h107; // @[Replacement.scala 315:30]
  wire  state_vec_263_left_subtree_state = state_vec_263[1]; // @[package.scala 154:13]
  wire  state_vec_263_right_subtree_state = state_vec_263[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_263_T_3 = state_vec_0_set_left_older ? state_vec_263_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_263_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_263_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_263_T_8 = {state_vec_0_set_left_older,_state_vec_263_T_3,_state_vec_263_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_264_valid = touch_way_0_valid & touch_set_0 == 9'h108; // @[Replacement.scala 315:30]
  wire  state_vec_264_left_subtree_state = state_vec_264[1]; // @[package.scala 154:13]
  wire  state_vec_264_right_subtree_state = state_vec_264[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_264_T_3 = state_vec_0_set_left_older ? state_vec_264_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_264_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_264_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_264_T_8 = {state_vec_0_set_left_older,_state_vec_264_T_3,_state_vec_264_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_265_valid = touch_way_0_valid & touch_set_0 == 9'h109; // @[Replacement.scala 315:30]
  wire  state_vec_265_left_subtree_state = state_vec_265[1]; // @[package.scala 154:13]
  wire  state_vec_265_right_subtree_state = state_vec_265[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_265_T_3 = state_vec_0_set_left_older ? state_vec_265_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_265_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_265_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_265_T_8 = {state_vec_0_set_left_older,_state_vec_265_T_3,_state_vec_265_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_266_valid = touch_way_0_valid & touch_set_0 == 9'h10a; // @[Replacement.scala 315:30]
  wire  state_vec_266_left_subtree_state = state_vec_266[1]; // @[package.scala 154:13]
  wire  state_vec_266_right_subtree_state = state_vec_266[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_266_T_3 = state_vec_0_set_left_older ? state_vec_266_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_266_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_266_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_266_T_8 = {state_vec_0_set_left_older,_state_vec_266_T_3,_state_vec_266_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_267_valid = touch_way_0_valid & touch_set_0 == 9'h10b; // @[Replacement.scala 315:30]
  wire  state_vec_267_left_subtree_state = state_vec_267[1]; // @[package.scala 154:13]
  wire  state_vec_267_right_subtree_state = state_vec_267[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_267_T_3 = state_vec_0_set_left_older ? state_vec_267_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_267_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_267_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_267_T_8 = {state_vec_0_set_left_older,_state_vec_267_T_3,_state_vec_267_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_268_valid = touch_way_0_valid & touch_set_0 == 9'h10c; // @[Replacement.scala 315:30]
  wire  state_vec_268_left_subtree_state = state_vec_268[1]; // @[package.scala 154:13]
  wire  state_vec_268_right_subtree_state = state_vec_268[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_268_T_3 = state_vec_0_set_left_older ? state_vec_268_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_268_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_268_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_268_T_8 = {state_vec_0_set_left_older,_state_vec_268_T_3,_state_vec_268_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_269_valid = touch_way_0_valid & touch_set_0 == 9'h10d; // @[Replacement.scala 315:30]
  wire  state_vec_269_left_subtree_state = state_vec_269[1]; // @[package.scala 154:13]
  wire  state_vec_269_right_subtree_state = state_vec_269[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_269_T_3 = state_vec_0_set_left_older ? state_vec_269_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_269_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_269_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_269_T_8 = {state_vec_0_set_left_older,_state_vec_269_T_3,_state_vec_269_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_270_valid = touch_way_0_valid & touch_set_0 == 9'h10e; // @[Replacement.scala 315:30]
  wire  state_vec_270_left_subtree_state = state_vec_270[1]; // @[package.scala 154:13]
  wire  state_vec_270_right_subtree_state = state_vec_270[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_270_T_3 = state_vec_0_set_left_older ? state_vec_270_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_270_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_270_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_270_T_8 = {state_vec_0_set_left_older,_state_vec_270_T_3,_state_vec_270_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_271_valid = touch_way_0_valid & touch_set_0 == 9'h10f; // @[Replacement.scala 315:30]
  wire  state_vec_271_left_subtree_state = state_vec_271[1]; // @[package.scala 154:13]
  wire  state_vec_271_right_subtree_state = state_vec_271[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_271_T_3 = state_vec_0_set_left_older ? state_vec_271_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_271_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_271_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_271_T_8 = {state_vec_0_set_left_older,_state_vec_271_T_3,_state_vec_271_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_272_valid = touch_way_0_valid & touch_set_0 == 9'h110; // @[Replacement.scala 315:30]
  wire  state_vec_272_left_subtree_state = state_vec_272[1]; // @[package.scala 154:13]
  wire  state_vec_272_right_subtree_state = state_vec_272[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_272_T_3 = state_vec_0_set_left_older ? state_vec_272_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_272_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_272_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_272_T_8 = {state_vec_0_set_left_older,_state_vec_272_T_3,_state_vec_272_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_273_valid = touch_way_0_valid & touch_set_0 == 9'h111; // @[Replacement.scala 315:30]
  wire  state_vec_273_left_subtree_state = state_vec_273[1]; // @[package.scala 154:13]
  wire  state_vec_273_right_subtree_state = state_vec_273[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_273_T_3 = state_vec_0_set_left_older ? state_vec_273_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_273_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_273_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_273_T_8 = {state_vec_0_set_left_older,_state_vec_273_T_3,_state_vec_273_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_274_valid = touch_way_0_valid & touch_set_0 == 9'h112; // @[Replacement.scala 315:30]
  wire  state_vec_274_left_subtree_state = state_vec_274[1]; // @[package.scala 154:13]
  wire  state_vec_274_right_subtree_state = state_vec_274[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_274_T_3 = state_vec_0_set_left_older ? state_vec_274_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_274_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_274_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_274_T_8 = {state_vec_0_set_left_older,_state_vec_274_T_3,_state_vec_274_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_275_valid = touch_way_0_valid & touch_set_0 == 9'h113; // @[Replacement.scala 315:30]
  wire  state_vec_275_left_subtree_state = state_vec_275[1]; // @[package.scala 154:13]
  wire  state_vec_275_right_subtree_state = state_vec_275[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_275_T_3 = state_vec_0_set_left_older ? state_vec_275_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_275_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_275_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_275_T_8 = {state_vec_0_set_left_older,_state_vec_275_T_3,_state_vec_275_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_276_valid = touch_way_0_valid & touch_set_0 == 9'h114; // @[Replacement.scala 315:30]
  wire  state_vec_276_left_subtree_state = state_vec_276[1]; // @[package.scala 154:13]
  wire  state_vec_276_right_subtree_state = state_vec_276[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_276_T_3 = state_vec_0_set_left_older ? state_vec_276_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_276_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_276_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_276_T_8 = {state_vec_0_set_left_older,_state_vec_276_T_3,_state_vec_276_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_277_valid = touch_way_0_valid & touch_set_0 == 9'h115; // @[Replacement.scala 315:30]
  wire  state_vec_277_left_subtree_state = state_vec_277[1]; // @[package.scala 154:13]
  wire  state_vec_277_right_subtree_state = state_vec_277[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_277_T_3 = state_vec_0_set_left_older ? state_vec_277_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_277_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_277_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_277_T_8 = {state_vec_0_set_left_older,_state_vec_277_T_3,_state_vec_277_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_278_valid = touch_way_0_valid & touch_set_0 == 9'h116; // @[Replacement.scala 315:30]
  wire  state_vec_278_left_subtree_state = state_vec_278[1]; // @[package.scala 154:13]
  wire  state_vec_278_right_subtree_state = state_vec_278[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_278_T_3 = state_vec_0_set_left_older ? state_vec_278_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_278_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_278_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_278_T_8 = {state_vec_0_set_left_older,_state_vec_278_T_3,_state_vec_278_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_279_valid = touch_way_0_valid & touch_set_0 == 9'h117; // @[Replacement.scala 315:30]
  wire  state_vec_279_left_subtree_state = state_vec_279[1]; // @[package.scala 154:13]
  wire  state_vec_279_right_subtree_state = state_vec_279[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_279_T_3 = state_vec_0_set_left_older ? state_vec_279_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_279_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_279_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_279_T_8 = {state_vec_0_set_left_older,_state_vec_279_T_3,_state_vec_279_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_280_valid = touch_way_0_valid & touch_set_0 == 9'h118; // @[Replacement.scala 315:30]
  wire  state_vec_280_left_subtree_state = state_vec_280[1]; // @[package.scala 154:13]
  wire  state_vec_280_right_subtree_state = state_vec_280[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_280_T_3 = state_vec_0_set_left_older ? state_vec_280_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_280_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_280_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_280_T_8 = {state_vec_0_set_left_older,_state_vec_280_T_3,_state_vec_280_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_281_valid = touch_way_0_valid & touch_set_0 == 9'h119; // @[Replacement.scala 315:30]
  wire  state_vec_281_left_subtree_state = state_vec_281[1]; // @[package.scala 154:13]
  wire  state_vec_281_right_subtree_state = state_vec_281[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_281_T_3 = state_vec_0_set_left_older ? state_vec_281_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_281_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_281_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_281_T_8 = {state_vec_0_set_left_older,_state_vec_281_T_3,_state_vec_281_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_282_valid = touch_way_0_valid & touch_set_0 == 9'h11a; // @[Replacement.scala 315:30]
  wire  state_vec_282_left_subtree_state = state_vec_282[1]; // @[package.scala 154:13]
  wire  state_vec_282_right_subtree_state = state_vec_282[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_282_T_3 = state_vec_0_set_left_older ? state_vec_282_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_282_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_282_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_282_T_8 = {state_vec_0_set_left_older,_state_vec_282_T_3,_state_vec_282_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_283_valid = touch_way_0_valid & touch_set_0 == 9'h11b; // @[Replacement.scala 315:30]
  wire  state_vec_283_left_subtree_state = state_vec_283[1]; // @[package.scala 154:13]
  wire  state_vec_283_right_subtree_state = state_vec_283[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_283_T_3 = state_vec_0_set_left_older ? state_vec_283_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_283_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_283_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_283_T_8 = {state_vec_0_set_left_older,_state_vec_283_T_3,_state_vec_283_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_284_valid = touch_way_0_valid & touch_set_0 == 9'h11c; // @[Replacement.scala 315:30]
  wire  state_vec_284_left_subtree_state = state_vec_284[1]; // @[package.scala 154:13]
  wire  state_vec_284_right_subtree_state = state_vec_284[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_284_T_3 = state_vec_0_set_left_older ? state_vec_284_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_284_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_284_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_284_T_8 = {state_vec_0_set_left_older,_state_vec_284_T_3,_state_vec_284_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_285_valid = touch_way_0_valid & touch_set_0 == 9'h11d; // @[Replacement.scala 315:30]
  wire  state_vec_285_left_subtree_state = state_vec_285[1]; // @[package.scala 154:13]
  wire  state_vec_285_right_subtree_state = state_vec_285[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_285_T_3 = state_vec_0_set_left_older ? state_vec_285_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_285_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_285_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_285_T_8 = {state_vec_0_set_left_older,_state_vec_285_T_3,_state_vec_285_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_286_valid = touch_way_0_valid & touch_set_0 == 9'h11e; // @[Replacement.scala 315:30]
  wire  state_vec_286_left_subtree_state = state_vec_286[1]; // @[package.scala 154:13]
  wire  state_vec_286_right_subtree_state = state_vec_286[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_286_T_3 = state_vec_0_set_left_older ? state_vec_286_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_286_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_286_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_286_T_8 = {state_vec_0_set_left_older,_state_vec_286_T_3,_state_vec_286_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_287_valid = touch_way_0_valid & touch_set_0 == 9'h11f; // @[Replacement.scala 315:30]
  wire  state_vec_287_left_subtree_state = state_vec_287[1]; // @[package.scala 154:13]
  wire  state_vec_287_right_subtree_state = state_vec_287[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_287_T_3 = state_vec_0_set_left_older ? state_vec_287_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_287_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_287_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_287_T_8 = {state_vec_0_set_left_older,_state_vec_287_T_3,_state_vec_287_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_288_valid = touch_way_0_valid & touch_set_0 == 9'h120; // @[Replacement.scala 315:30]
  wire  state_vec_288_left_subtree_state = state_vec_288[1]; // @[package.scala 154:13]
  wire  state_vec_288_right_subtree_state = state_vec_288[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_288_T_3 = state_vec_0_set_left_older ? state_vec_288_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_288_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_288_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_288_T_8 = {state_vec_0_set_left_older,_state_vec_288_T_3,_state_vec_288_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_289_valid = touch_way_0_valid & touch_set_0 == 9'h121; // @[Replacement.scala 315:30]
  wire  state_vec_289_left_subtree_state = state_vec_289[1]; // @[package.scala 154:13]
  wire  state_vec_289_right_subtree_state = state_vec_289[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_289_T_3 = state_vec_0_set_left_older ? state_vec_289_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_289_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_289_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_289_T_8 = {state_vec_0_set_left_older,_state_vec_289_T_3,_state_vec_289_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_290_valid = touch_way_0_valid & touch_set_0 == 9'h122; // @[Replacement.scala 315:30]
  wire  state_vec_290_left_subtree_state = state_vec_290[1]; // @[package.scala 154:13]
  wire  state_vec_290_right_subtree_state = state_vec_290[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_290_T_3 = state_vec_0_set_left_older ? state_vec_290_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_290_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_290_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_290_T_8 = {state_vec_0_set_left_older,_state_vec_290_T_3,_state_vec_290_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_291_valid = touch_way_0_valid & touch_set_0 == 9'h123; // @[Replacement.scala 315:30]
  wire  state_vec_291_left_subtree_state = state_vec_291[1]; // @[package.scala 154:13]
  wire  state_vec_291_right_subtree_state = state_vec_291[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_291_T_3 = state_vec_0_set_left_older ? state_vec_291_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_291_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_291_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_291_T_8 = {state_vec_0_set_left_older,_state_vec_291_T_3,_state_vec_291_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_292_valid = touch_way_0_valid & touch_set_0 == 9'h124; // @[Replacement.scala 315:30]
  wire  state_vec_292_left_subtree_state = state_vec_292[1]; // @[package.scala 154:13]
  wire  state_vec_292_right_subtree_state = state_vec_292[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_292_T_3 = state_vec_0_set_left_older ? state_vec_292_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_292_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_292_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_292_T_8 = {state_vec_0_set_left_older,_state_vec_292_T_3,_state_vec_292_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_293_valid = touch_way_0_valid & touch_set_0 == 9'h125; // @[Replacement.scala 315:30]
  wire  state_vec_293_left_subtree_state = state_vec_293[1]; // @[package.scala 154:13]
  wire  state_vec_293_right_subtree_state = state_vec_293[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_293_T_3 = state_vec_0_set_left_older ? state_vec_293_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_293_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_293_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_293_T_8 = {state_vec_0_set_left_older,_state_vec_293_T_3,_state_vec_293_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_294_valid = touch_way_0_valid & touch_set_0 == 9'h126; // @[Replacement.scala 315:30]
  wire  state_vec_294_left_subtree_state = state_vec_294[1]; // @[package.scala 154:13]
  wire  state_vec_294_right_subtree_state = state_vec_294[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_294_T_3 = state_vec_0_set_left_older ? state_vec_294_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_294_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_294_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_294_T_8 = {state_vec_0_set_left_older,_state_vec_294_T_3,_state_vec_294_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_295_valid = touch_way_0_valid & touch_set_0 == 9'h127; // @[Replacement.scala 315:30]
  wire  state_vec_295_left_subtree_state = state_vec_295[1]; // @[package.scala 154:13]
  wire  state_vec_295_right_subtree_state = state_vec_295[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_295_T_3 = state_vec_0_set_left_older ? state_vec_295_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_295_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_295_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_295_T_8 = {state_vec_0_set_left_older,_state_vec_295_T_3,_state_vec_295_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_296_valid = touch_way_0_valid & touch_set_0 == 9'h128; // @[Replacement.scala 315:30]
  wire  state_vec_296_left_subtree_state = state_vec_296[1]; // @[package.scala 154:13]
  wire  state_vec_296_right_subtree_state = state_vec_296[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_296_T_3 = state_vec_0_set_left_older ? state_vec_296_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_296_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_296_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_296_T_8 = {state_vec_0_set_left_older,_state_vec_296_T_3,_state_vec_296_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_297_valid = touch_way_0_valid & touch_set_0 == 9'h129; // @[Replacement.scala 315:30]
  wire  state_vec_297_left_subtree_state = state_vec_297[1]; // @[package.scala 154:13]
  wire  state_vec_297_right_subtree_state = state_vec_297[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_297_T_3 = state_vec_0_set_left_older ? state_vec_297_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_297_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_297_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_297_T_8 = {state_vec_0_set_left_older,_state_vec_297_T_3,_state_vec_297_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_298_valid = touch_way_0_valid & touch_set_0 == 9'h12a; // @[Replacement.scala 315:30]
  wire  state_vec_298_left_subtree_state = state_vec_298[1]; // @[package.scala 154:13]
  wire  state_vec_298_right_subtree_state = state_vec_298[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_298_T_3 = state_vec_0_set_left_older ? state_vec_298_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_298_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_298_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_298_T_8 = {state_vec_0_set_left_older,_state_vec_298_T_3,_state_vec_298_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_299_valid = touch_way_0_valid & touch_set_0 == 9'h12b; // @[Replacement.scala 315:30]
  wire  state_vec_299_left_subtree_state = state_vec_299[1]; // @[package.scala 154:13]
  wire  state_vec_299_right_subtree_state = state_vec_299[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_299_T_3 = state_vec_0_set_left_older ? state_vec_299_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_299_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_299_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_299_T_8 = {state_vec_0_set_left_older,_state_vec_299_T_3,_state_vec_299_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_300_valid = touch_way_0_valid & touch_set_0 == 9'h12c; // @[Replacement.scala 315:30]
  wire  state_vec_300_left_subtree_state = state_vec_300[1]; // @[package.scala 154:13]
  wire  state_vec_300_right_subtree_state = state_vec_300[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_300_T_3 = state_vec_0_set_left_older ? state_vec_300_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_300_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_300_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_300_T_8 = {state_vec_0_set_left_older,_state_vec_300_T_3,_state_vec_300_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_301_valid = touch_way_0_valid & touch_set_0 == 9'h12d; // @[Replacement.scala 315:30]
  wire  state_vec_301_left_subtree_state = state_vec_301[1]; // @[package.scala 154:13]
  wire  state_vec_301_right_subtree_state = state_vec_301[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_301_T_3 = state_vec_0_set_left_older ? state_vec_301_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_301_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_301_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_301_T_8 = {state_vec_0_set_left_older,_state_vec_301_T_3,_state_vec_301_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_302_valid = touch_way_0_valid & touch_set_0 == 9'h12e; // @[Replacement.scala 315:30]
  wire  state_vec_302_left_subtree_state = state_vec_302[1]; // @[package.scala 154:13]
  wire  state_vec_302_right_subtree_state = state_vec_302[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_302_T_3 = state_vec_0_set_left_older ? state_vec_302_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_302_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_302_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_302_T_8 = {state_vec_0_set_left_older,_state_vec_302_T_3,_state_vec_302_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_303_valid = touch_way_0_valid & touch_set_0 == 9'h12f; // @[Replacement.scala 315:30]
  wire  state_vec_303_left_subtree_state = state_vec_303[1]; // @[package.scala 154:13]
  wire  state_vec_303_right_subtree_state = state_vec_303[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_303_T_3 = state_vec_0_set_left_older ? state_vec_303_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_303_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_303_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_303_T_8 = {state_vec_0_set_left_older,_state_vec_303_T_3,_state_vec_303_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_304_valid = touch_way_0_valid & touch_set_0 == 9'h130; // @[Replacement.scala 315:30]
  wire  state_vec_304_left_subtree_state = state_vec_304[1]; // @[package.scala 154:13]
  wire  state_vec_304_right_subtree_state = state_vec_304[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_304_T_3 = state_vec_0_set_left_older ? state_vec_304_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_304_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_304_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_304_T_8 = {state_vec_0_set_left_older,_state_vec_304_T_3,_state_vec_304_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_305_valid = touch_way_0_valid & touch_set_0 == 9'h131; // @[Replacement.scala 315:30]
  wire  state_vec_305_left_subtree_state = state_vec_305[1]; // @[package.scala 154:13]
  wire  state_vec_305_right_subtree_state = state_vec_305[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_305_T_3 = state_vec_0_set_left_older ? state_vec_305_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_305_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_305_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_305_T_8 = {state_vec_0_set_left_older,_state_vec_305_T_3,_state_vec_305_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_306_valid = touch_way_0_valid & touch_set_0 == 9'h132; // @[Replacement.scala 315:30]
  wire  state_vec_306_left_subtree_state = state_vec_306[1]; // @[package.scala 154:13]
  wire  state_vec_306_right_subtree_state = state_vec_306[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_306_T_3 = state_vec_0_set_left_older ? state_vec_306_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_306_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_306_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_306_T_8 = {state_vec_0_set_left_older,_state_vec_306_T_3,_state_vec_306_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_307_valid = touch_way_0_valid & touch_set_0 == 9'h133; // @[Replacement.scala 315:30]
  wire  state_vec_307_left_subtree_state = state_vec_307[1]; // @[package.scala 154:13]
  wire  state_vec_307_right_subtree_state = state_vec_307[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_307_T_3 = state_vec_0_set_left_older ? state_vec_307_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_307_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_307_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_307_T_8 = {state_vec_0_set_left_older,_state_vec_307_T_3,_state_vec_307_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_308_valid = touch_way_0_valid & touch_set_0 == 9'h134; // @[Replacement.scala 315:30]
  wire  state_vec_308_left_subtree_state = state_vec_308[1]; // @[package.scala 154:13]
  wire  state_vec_308_right_subtree_state = state_vec_308[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_308_T_3 = state_vec_0_set_left_older ? state_vec_308_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_308_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_308_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_308_T_8 = {state_vec_0_set_left_older,_state_vec_308_T_3,_state_vec_308_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_309_valid = touch_way_0_valid & touch_set_0 == 9'h135; // @[Replacement.scala 315:30]
  wire  state_vec_309_left_subtree_state = state_vec_309[1]; // @[package.scala 154:13]
  wire  state_vec_309_right_subtree_state = state_vec_309[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_309_T_3 = state_vec_0_set_left_older ? state_vec_309_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_309_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_309_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_309_T_8 = {state_vec_0_set_left_older,_state_vec_309_T_3,_state_vec_309_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_310_valid = touch_way_0_valid & touch_set_0 == 9'h136; // @[Replacement.scala 315:30]
  wire  state_vec_310_left_subtree_state = state_vec_310[1]; // @[package.scala 154:13]
  wire  state_vec_310_right_subtree_state = state_vec_310[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_310_T_3 = state_vec_0_set_left_older ? state_vec_310_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_310_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_310_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_310_T_8 = {state_vec_0_set_left_older,_state_vec_310_T_3,_state_vec_310_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_311_valid = touch_way_0_valid & touch_set_0 == 9'h137; // @[Replacement.scala 315:30]
  wire  state_vec_311_left_subtree_state = state_vec_311[1]; // @[package.scala 154:13]
  wire  state_vec_311_right_subtree_state = state_vec_311[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_311_T_3 = state_vec_0_set_left_older ? state_vec_311_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_311_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_311_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_311_T_8 = {state_vec_0_set_left_older,_state_vec_311_T_3,_state_vec_311_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_312_valid = touch_way_0_valid & touch_set_0 == 9'h138; // @[Replacement.scala 315:30]
  wire  state_vec_312_left_subtree_state = state_vec_312[1]; // @[package.scala 154:13]
  wire  state_vec_312_right_subtree_state = state_vec_312[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_312_T_3 = state_vec_0_set_left_older ? state_vec_312_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_312_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_312_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_312_T_8 = {state_vec_0_set_left_older,_state_vec_312_T_3,_state_vec_312_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_313_valid = touch_way_0_valid & touch_set_0 == 9'h139; // @[Replacement.scala 315:30]
  wire  state_vec_313_left_subtree_state = state_vec_313[1]; // @[package.scala 154:13]
  wire  state_vec_313_right_subtree_state = state_vec_313[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_313_T_3 = state_vec_0_set_left_older ? state_vec_313_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_313_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_313_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_313_T_8 = {state_vec_0_set_left_older,_state_vec_313_T_3,_state_vec_313_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_314_valid = touch_way_0_valid & touch_set_0 == 9'h13a; // @[Replacement.scala 315:30]
  wire  state_vec_314_left_subtree_state = state_vec_314[1]; // @[package.scala 154:13]
  wire  state_vec_314_right_subtree_state = state_vec_314[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_314_T_3 = state_vec_0_set_left_older ? state_vec_314_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_314_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_314_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_314_T_8 = {state_vec_0_set_left_older,_state_vec_314_T_3,_state_vec_314_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_315_valid = touch_way_0_valid & touch_set_0 == 9'h13b; // @[Replacement.scala 315:30]
  wire  state_vec_315_left_subtree_state = state_vec_315[1]; // @[package.scala 154:13]
  wire  state_vec_315_right_subtree_state = state_vec_315[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_315_T_3 = state_vec_0_set_left_older ? state_vec_315_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_315_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_315_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_315_T_8 = {state_vec_0_set_left_older,_state_vec_315_T_3,_state_vec_315_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_316_valid = touch_way_0_valid & touch_set_0 == 9'h13c; // @[Replacement.scala 315:30]
  wire  state_vec_316_left_subtree_state = state_vec_316[1]; // @[package.scala 154:13]
  wire  state_vec_316_right_subtree_state = state_vec_316[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_316_T_3 = state_vec_0_set_left_older ? state_vec_316_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_316_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_316_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_316_T_8 = {state_vec_0_set_left_older,_state_vec_316_T_3,_state_vec_316_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_317_valid = touch_way_0_valid & touch_set_0 == 9'h13d; // @[Replacement.scala 315:30]
  wire  state_vec_317_left_subtree_state = state_vec_317[1]; // @[package.scala 154:13]
  wire  state_vec_317_right_subtree_state = state_vec_317[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_317_T_3 = state_vec_0_set_left_older ? state_vec_317_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_317_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_317_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_317_T_8 = {state_vec_0_set_left_older,_state_vec_317_T_3,_state_vec_317_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_318_valid = touch_way_0_valid & touch_set_0 == 9'h13e; // @[Replacement.scala 315:30]
  wire  state_vec_318_left_subtree_state = state_vec_318[1]; // @[package.scala 154:13]
  wire  state_vec_318_right_subtree_state = state_vec_318[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_318_T_3 = state_vec_0_set_left_older ? state_vec_318_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_318_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_318_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_318_T_8 = {state_vec_0_set_left_older,_state_vec_318_T_3,_state_vec_318_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_319_valid = touch_way_0_valid & touch_set_0 == 9'h13f; // @[Replacement.scala 315:30]
  wire  state_vec_319_left_subtree_state = state_vec_319[1]; // @[package.scala 154:13]
  wire  state_vec_319_right_subtree_state = state_vec_319[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_319_T_3 = state_vec_0_set_left_older ? state_vec_319_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_319_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_319_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_319_T_8 = {state_vec_0_set_left_older,_state_vec_319_T_3,_state_vec_319_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_320_valid = touch_way_0_valid & touch_set_0 == 9'h140; // @[Replacement.scala 315:30]
  wire  state_vec_320_left_subtree_state = state_vec_320[1]; // @[package.scala 154:13]
  wire  state_vec_320_right_subtree_state = state_vec_320[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_320_T_3 = state_vec_0_set_left_older ? state_vec_320_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_320_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_320_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_320_T_8 = {state_vec_0_set_left_older,_state_vec_320_T_3,_state_vec_320_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_321_valid = touch_way_0_valid & touch_set_0 == 9'h141; // @[Replacement.scala 315:30]
  wire  state_vec_321_left_subtree_state = state_vec_321[1]; // @[package.scala 154:13]
  wire  state_vec_321_right_subtree_state = state_vec_321[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_321_T_3 = state_vec_0_set_left_older ? state_vec_321_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_321_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_321_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_321_T_8 = {state_vec_0_set_left_older,_state_vec_321_T_3,_state_vec_321_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_322_valid = touch_way_0_valid & touch_set_0 == 9'h142; // @[Replacement.scala 315:30]
  wire  state_vec_322_left_subtree_state = state_vec_322[1]; // @[package.scala 154:13]
  wire  state_vec_322_right_subtree_state = state_vec_322[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_322_T_3 = state_vec_0_set_left_older ? state_vec_322_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_322_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_322_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_322_T_8 = {state_vec_0_set_left_older,_state_vec_322_T_3,_state_vec_322_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_323_valid = touch_way_0_valid & touch_set_0 == 9'h143; // @[Replacement.scala 315:30]
  wire  state_vec_323_left_subtree_state = state_vec_323[1]; // @[package.scala 154:13]
  wire  state_vec_323_right_subtree_state = state_vec_323[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_323_T_3 = state_vec_0_set_left_older ? state_vec_323_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_323_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_323_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_323_T_8 = {state_vec_0_set_left_older,_state_vec_323_T_3,_state_vec_323_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_324_valid = touch_way_0_valid & touch_set_0 == 9'h144; // @[Replacement.scala 315:30]
  wire  state_vec_324_left_subtree_state = state_vec_324[1]; // @[package.scala 154:13]
  wire  state_vec_324_right_subtree_state = state_vec_324[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_324_T_3 = state_vec_0_set_left_older ? state_vec_324_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_324_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_324_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_324_T_8 = {state_vec_0_set_left_older,_state_vec_324_T_3,_state_vec_324_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_325_valid = touch_way_0_valid & touch_set_0 == 9'h145; // @[Replacement.scala 315:30]
  wire  state_vec_325_left_subtree_state = state_vec_325[1]; // @[package.scala 154:13]
  wire  state_vec_325_right_subtree_state = state_vec_325[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_325_T_3 = state_vec_0_set_left_older ? state_vec_325_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_325_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_325_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_325_T_8 = {state_vec_0_set_left_older,_state_vec_325_T_3,_state_vec_325_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_326_valid = touch_way_0_valid & touch_set_0 == 9'h146; // @[Replacement.scala 315:30]
  wire  state_vec_326_left_subtree_state = state_vec_326[1]; // @[package.scala 154:13]
  wire  state_vec_326_right_subtree_state = state_vec_326[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_326_T_3 = state_vec_0_set_left_older ? state_vec_326_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_326_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_326_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_326_T_8 = {state_vec_0_set_left_older,_state_vec_326_T_3,_state_vec_326_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_327_valid = touch_way_0_valid & touch_set_0 == 9'h147; // @[Replacement.scala 315:30]
  wire  state_vec_327_left_subtree_state = state_vec_327[1]; // @[package.scala 154:13]
  wire  state_vec_327_right_subtree_state = state_vec_327[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_327_T_3 = state_vec_0_set_left_older ? state_vec_327_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_327_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_327_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_327_T_8 = {state_vec_0_set_left_older,_state_vec_327_T_3,_state_vec_327_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_328_valid = touch_way_0_valid & touch_set_0 == 9'h148; // @[Replacement.scala 315:30]
  wire  state_vec_328_left_subtree_state = state_vec_328[1]; // @[package.scala 154:13]
  wire  state_vec_328_right_subtree_state = state_vec_328[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_328_T_3 = state_vec_0_set_left_older ? state_vec_328_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_328_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_328_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_328_T_8 = {state_vec_0_set_left_older,_state_vec_328_T_3,_state_vec_328_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_329_valid = touch_way_0_valid & touch_set_0 == 9'h149; // @[Replacement.scala 315:30]
  wire  state_vec_329_left_subtree_state = state_vec_329[1]; // @[package.scala 154:13]
  wire  state_vec_329_right_subtree_state = state_vec_329[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_329_T_3 = state_vec_0_set_left_older ? state_vec_329_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_329_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_329_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_329_T_8 = {state_vec_0_set_left_older,_state_vec_329_T_3,_state_vec_329_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_330_valid = touch_way_0_valid & touch_set_0 == 9'h14a; // @[Replacement.scala 315:30]
  wire  state_vec_330_left_subtree_state = state_vec_330[1]; // @[package.scala 154:13]
  wire  state_vec_330_right_subtree_state = state_vec_330[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_330_T_3 = state_vec_0_set_left_older ? state_vec_330_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_330_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_330_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_330_T_8 = {state_vec_0_set_left_older,_state_vec_330_T_3,_state_vec_330_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_331_valid = touch_way_0_valid & touch_set_0 == 9'h14b; // @[Replacement.scala 315:30]
  wire  state_vec_331_left_subtree_state = state_vec_331[1]; // @[package.scala 154:13]
  wire  state_vec_331_right_subtree_state = state_vec_331[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_331_T_3 = state_vec_0_set_left_older ? state_vec_331_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_331_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_331_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_331_T_8 = {state_vec_0_set_left_older,_state_vec_331_T_3,_state_vec_331_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_332_valid = touch_way_0_valid & touch_set_0 == 9'h14c; // @[Replacement.scala 315:30]
  wire  state_vec_332_left_subtree_state = state_vec_332[1]; // @[package.scala 154:13]
  wire  state_vec_332_right_subtree_state = state_vec_332[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_332_T_3 = state_vec_0_set_left_older ? state_vec_332_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_332_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_332_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_332_T_8 = {state_vec_0_set_left_older,_state_vec_332_T_3,_state_vec_332_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_333_valid = touch_way_0_valid & touch_set_0 == 9'h14d; // @[Replacement.scala 315:30]
  wire  state_vec_333_left_subtree_state = state_vec_333[1]; // @[package.scala 154:13]
  wire  state_vec_333_right_subtree_state = state_vec_333[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_333_T_3 = state_vec_0_set_left_older ? state_vec_333_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_333_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_333_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_333_T_8 = {state_vec_0_set_left_older,_state_vec_333_T_3,_state_vec_333_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_334_valid = touch_way_0_valid & touch_set_0 == 9'h14e; // @[Replacement.scala 315:30]
  wire  state_vec_334_left_subtree_state = state_vec_334[1]; // @[package.scala 154:13]
  wire  state_vec_334_right_subtree_state = state_vec_334[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_334_T_3 = state_vec_0_set_left_older ? state_vec_334_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_334_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_334_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_334_T_8 = {state_vec_0_set_left_older,_state_vec_334_T_3,_state_vec_334_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_335_valid = touch_way_0_valid & touch_set_0 == 9'h14f; // @[Replacement.scala 315:30]
  wire  state_vec_335_left_subtree_state = state_vec_335[1]; // @[package.scala 154:13]
  wire  state_vec_335_right_subtree_state = state_vec_335[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_335_T_3 = state_vec_0_set_left_older ? state_vec_335_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_335_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_335_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_335_T_8 = {state_vec_0_set_left_older,_state_vec_335_T_3,_state_vec_335_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_336_valid = touch_way_0_valid & touch_set_0 == 9'h150; // @[Replacement.scala 315:30]
  wire  state_vec_336_left_subtree_state = state_vec_336[1]; // @[package.scala 154:13]
  wire  state_vec_336_right_subtree_state = state_vec_336[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_336_T_3 = state_vec_0_set_left_older ? state_vec_336_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_336_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_336_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_336_T_8 = {state_vec_0_set_left_older,_state_vec_336_T_3,_state_vec_336_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_337_valid = touch_way_0_valid & touch_set_0 == 9'h151; // @[Replacement.scala 315:30]
  wire  state_vec_337_left_subtree_state = state_vec_337[1]; // @[package.scala 154:13]
  wire  state_vec_337_right_subtree_state = state_vec_337[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_337_T_3 = state_vec_0_set_left_older ? state_vec_337_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_337_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_337_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_337_T_8 = {state_vec_0_set_left_older,_state_vec_337_T_3,_state_vec_337_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_338_valid = touch_way_0_valid & touch_set_0 == 9'h152; // @[Replacement.scala 315:30]
  wire  state_vec_338_left_subtree_state = state_vec_338[1]; // @[package.scala 154:13]
  wire  state_vec_338_right_subtree_state = state_vec_338[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_338_T_3 = state_vec_0_set_left_older ? state_vec_338_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_338_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_338_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_338_T_8 = {state_vec_0_set_left_older,_state_vec_338_T_3,_state_vec_338_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_339_valid = touch_way_0_valid & touch_set_0 == 9'h153; // @[Replacement.scala 315:30]
  wire  state_vec_339_left_subtree_state = state_vec_339[1]; // @[package.scala 154:13]
  wire  state_vec_339_right_subtree_state = state_vec_339[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_339_T_3 = state_vec_0_set_left_older ? state_vec_339_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_339_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_339_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_339_T_8 = {state_vec_0_set_left_older,_state_vec_339_T_3,_state_vec_339_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_340_valid = touch_way_0_valid & touch_set_0 == 9'h154; // @[Replacement.scala 315:30]
  wire  state_vec_340_left_subtree_state = state_vec_340[1]; // @[package.scala 154:13]
  wire  state_vec_340_right_subtree_state = state_vec_340[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_340_T_3 = state_vec_0_set_left_older ? state_vec_340_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_340_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_340_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_340_T_8 = {state_vec_0_set_left_older,_state_vec_340_T_3,_state_vec_340_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_341_valid = touch_way_0_valid & touch_set_0 == 9'h155; // @[Replacement.scala 315:30]
  wire  state_vec_341_left_subtree_state = state_vec_341[1]; // @[package.scala 154:13]
  wire  state_vec_341_right_subtree_state = state_vec_341[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_341_T_3 = state_vec_0_set_left_older ? state_vec_341_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_341_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_341_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_341_T_8 = {state_vec_0_set_left_older,_state_vec_341_T_3,_state_vec_341_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_342_valid = touch_way_0_valid & touch_set_0 == 9'h156; // @[Replacement.scala 315:30]
  wire  state_vec_342_left_subtree_state = state_vec_342[1]; // @[package.scala 154:13]
  wire  state_vec_342_right_subtree_state = state_vec_342[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_342_T_3 = state_vec_0_set_left_older ? state_vec_342_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_342_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_342_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_342_T_8 = {state_vec_0_set_left_older,_state_vec_342_T_3,_state_vec_342_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_343_valid = touch_way_0_valid & touch_set_0 == 9'h157; // @[Replacement.scala 315:30]
  wire  state_vec_343_left_subtree_state = state_vec_343[1]; // @[package.scala 154:13]
  wire  state_vec_343_right_subtree_state = state_vec_343[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_343_T_3 = state_vec_0_set_left_older ? state_vec_343_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_343_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_343_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_343_T_8 = {state_vec_0_set_left_older,_state_vec_343_T_3,_state_vec_343_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_344_valid = touch_way_0_valid & touch_set_0 == 9'h158; // @[Replacement.scala 315:30]
  wire  state_vec_344_left_subtree_state = state_vec_344[1]; // @[package.scala 154:13]
  wire  state_vec_344_right_subtree_state = state_vec_344[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_344_T_3 = state_vec_0_set_left_older ? state_vec_344_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_344_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_344_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_344_T_8 = {state_vec_0_set_left_older,_state_vec_344_T_3,_state_vec_344_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_345_valid = touch_way_0_valid & touch_set_0 == 9'h159; // @[Replacement.scala 315:30]
  wire  state_vec_345_left_subtree_state = state_vec_345[1]; // @[package.scala 154:13]
  wire  state_vec_345_right_subtree_state = state_vec_345[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_345_T_3 = state_vec_0_set_left_older ? state_vec_345_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_345_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_345_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_345_T_8 = {state_vec_0_set_left_older,_state_vec_345_T_3,_state_vec_345_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_346_valid = touch_way_0_valid & touch_set_0 == 9'h15a; // @[Replacement.scala 315:30]
  wire  state_vec_346_left_subtree_state = state_vec_346[1]; // @[package.scala 154:13]
  wire  state_vec_346_right_subtree_state = state_vec_346[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_346_T_3 = state_vec_0_set_left_older ? state_vec_346_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_346_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_346_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_346_T_8 = {state_vec_0_set_left_older,_state_vec_346_T_3,_state_vec_346_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_347_valid = touch_way_0_valid & touch_set_0 == 9'h15b; // @[Replacement.scala 315:30]
  wire  state_vec_347_left_subtree_state = state_vec_347[1]; // @[package.scala 154:13]
  wire  state_vec_347_right_subtree_state = state_vec_347[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_347_T_3 = state_vec_0_set_left_older ? state_vec_347_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_347_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_347_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_347_T_8 = {state_vec_0_set_left_older,_state_vec_347_T_3,_state_vec_347_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_348_valid = touch_way_0_valid & touch_set_0 == 9'h15c; // @[Replacement.scala 315:30]
  wire  state_vec_348_left_subtree_state = state_vec_348[1]; // @[package.scala 154:13]
  wire  state_vec_348_right_subtree_state = state_vec_348[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_348_T_3 = state_vec_0_set_left_older ? state_vec_348_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_348_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_348_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_348_T_8 = {state_vec_0_set_left_older,_state_vec_348_T_3,_state_vec_348_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_349_valid = touch_way_0_valid & touch_set_0 == 9'h15d; // @[Replacement.scala 315:30]
  wire  state_vec_349_left_subtree_state = state_vec_349[1]; // @[package.scala 154:13]
  wire  state_vec_349_right_subtree_state = state_vec_349[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_349_T_3 = state_vec_0_set_left_older ? state_vec_349_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_349_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_349_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_349_T_8 = {state_vec_0_set_left_older,_state_vec_349_T_3,_state_vec_349_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_350_valid = touch_way_0_valid & touch_set_0 == 9'h15e; // @[Replacement.scala 315:30]
  wire  state_vec_350_left_subtree_state = state_vec_350[1]; // @[package.scala 154:13]
  wire  state_vec_350_right_subtree_state = state_vec_350[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_350_T_3 = state_vec_0_set_left_older ? state_vec_350_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_350_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_350_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_350_T_8 = {state_vec_0_set_left_older,_state_vec_350_T_3,_state_vec_350_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_351_valid = touch_way_0_valid & touch_set_0 == 9'h15f; // @[Replacement.scala 315:30]
  wire  state_vec_351_left_subtree_state = state_vec_351[1]; // @[package.scala 154:13]
  wire  state_vec_351_right_subtree_state = state_vec_351[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_351_T_3 = state_vec_0_set_left_older ? state_vec_351_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_351_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_351_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_351_T_8 = {state_vec_0_set_left_older,_state_vec_351_T_3,_state_vec_351_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_352_valid = touch_way_0_valid & touch_set_0 == 9'h160; // @[Replacement.scala 315:30]
  wire  state_vec_352_left_subtree_state = state_vec_352[1]; // @[package.scala 154:13]
  wire  state_vec_352_right_subtree_state = state_vec_352[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_352_T_3 = state_vec_0_set_left_older ? state_vec_352_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_352_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_352_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_352_T_8 = {state_vec_0_set_left_older,_state_vec_352_T_3,_state_vec_352_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_353_valid = touch_way_0_valid & touch_set_0 == 9'h161; // @[Replacement.scala 315:30]
  wire  state_vec_353_left_subtree_state = state_vec_353[1]; // @[package.scala 154:13]
  wire  state_vec_353_right_subtree_state = state_vec_353[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_353_T_3 = state_vec_0_set_left_older ? state_vec_353_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_353_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_353_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_353_T_8 = {state_vec_0_set_left_older,_state_vec_353_T_3,_state_vec_353_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_354_valid = touch_way_0_valid & touch_set_0 == 9'h162; // @[Replacement.scala 315:30]
  wire  state_vec_354_left_subtree_state = state_vec_354[1]; // @[package.scala 154:13]
  wire  state_vec_354_right_subtree_state = state_vec_354[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_354_T_3 = state_vec_0_set_left_older ? state_vec_354_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_354_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_354_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_354_T_8 = {state_vec_0_set_left_older,_state_vec_354_T_3,_state_vec_354_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_355_valid = touch_way_0_valid & touch_set_0 == 9'h163; // @[Replacement.scala 315:30]
  wire  state_vec_355_left_subtree_state = state_vec_355[1]; // @[package.scala 154:13]
  wire  state_vec_355_right_subtree_state = state_vec_355[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_355_T_3 = state_vec_0_set_left_older ? state_vec_355_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_355_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_355_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_355_T_8 = {state_vec_0_set_left_older,_state_vec_355_T_3,_state_vec_355_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_356_valid = touch_way_0_valid & touch_set_0 == 9'h164; // @[Replacement.scala 315:30]
  wire  state_vec_356_left_subtree_state = state_vec_356[1]; // @[package.scala 154:13]
  wire  state_vec_356_right_subtree_state = state_vec_356[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_356_T_3 = state_vec_0_set_left_older ? state_vec_356_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_356_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_356_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_356_T_8 = {state_vec_0_set_left_older,_state_vec_356_T_3,_state_vec_356_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_357_valid = touch_way_0_valid & touch_set_0 == 9'h165; // @[Replacement.scala 315:30]
  wire  state_vec_357_left_subtree_state = state_vec_357[1]; // @[package.scala 154:13]
  wire  state_vec_357_right_subtree_state = state_vec_357[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_357_T_3 = state_vec_0_set_left_older ? state_vec_357_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_357_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_357_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_357_T_8 = {state_vec_0_set_left_older,_state_vec_357_T_3,_state_vec_357_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_358_valid = touch_way_0_valid & touch_set_0 == 9'h166; // @[Replacement.scala 315:30]
  wire  state_vec_358_left_subtree_state = state_vec_358[1]; // @[package.scala 154:13]
  wire  state_vec_358_right_subtree_state = state_vec_358[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_358_T_3 = state_vec_0_set_left_older ? state_vec_358_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_358_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_358_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_358_T_8 = {state_vec_0_set_left_older,_state_vec_358_T_3,_state_vec_358_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_359_valid = touch_way_0_valid & touch_set_0 == 9'h167; // @[Replacement.scala 315:30]
  wire  state_vec_359_left_subtree_state = state_vec_359[1]; // @[package.scala 154:13]
  wire  state_vec_359_right_subtree_state = state_vec_359[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_359_T_3 = state_vec_0_set_left_older ? state_vec_359_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_359_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_359_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_359_T_8 = {state_vec_0_set_left_older,_state_vec_359_T_3,_state_vec_359_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_360_valid = touch_way_0_valid & touch_set_0 == 9'h168; // @[Replacement.scala 315:30]
  wire  state_vec_360_left_subtree_state = state_vec_360[1]; // @[package.scala 154:13]
  wire  state_vec_360_right_subtree_state = state_vec_360[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_360_T_3 = state_vec_0_set_left_older ? state_vec_360_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_360_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_360_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_360_T_8 = {state_vec_0_set_left_older,_state_vec_360_T_3,_state_vec_360_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_361_valid = touch_way_0_valid & touch_set_0 == 9'h169; // @[Replacement.scala 315:30]
  wire  state_vec_361_left_subtree_state = state_vec_361[1]; // @[package.scala 154:13]
  wire  state_vec_361_right_subtree_state = state_vec_361[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_361_T_3 = state_vec_0_set_left_older ? state_vec_361_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_361_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_361_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_361_T_8 = {state_vec_0_set_left_older,_state_vec_361_T_3,_state_vec_361_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_362_valid = touch_way_0_valid & touch_set_0 == 9'h16a; // @[Replacement.scala 315:30]
  wire  state_vec_362_left_subtree_state = state_vec_362[1]; // @[package.scala 154:13]
  wire  state_vec_362_right_subtree_state = state_vec_362[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_362_T_3 = state_vec_0_set_left_older ? state_vec_362_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_362_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_362_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_362_T_8 = {state_vec_0_set_left_older,_state_vec_362_T_3,_state_vec_362_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_363_valid = touch_way_0_valid & touch_set_0 == 9'h16b; // @[Replacement.scala 315:30]
  wire  state_vec_363_left_subtree_state = state_vec_363[1]; // @[package.scala 154:13]
  wire  state_vec_363_right_subtree_state = state_vec_363[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_363_T_3 = state_vec_0_set_left_older ? state_vec_363_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_363_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_363_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_363_T_8 = {state_vec_0_set_left_older,_state_vec_363_T_3,_state_vec_363_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_364_valid = touch_way_0_valid & touch_set_0 == 9'h16c; // @[Replacement.scala 315:30]
  wire  state_vec_364_left_subtree_state = state_vec_364[1]; // @[package.scala 154:13]
  wire  state_vec_364_right_subtree_state = state_vec_364[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_364_T_3 = state_vec_0_set_left_older ? state_vec_364_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_364_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_364_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_364_T_8 = {state_vec_0_set_left_older,_state_vec_364_T_3,_state_vec_364_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_365_valid = touch_way_0_valid & touch_set_0 == 9'h16d; // @[Replacement.scala 315:30]
  wire  state_vec_365_left_subtree_state = state_vec_365[1]; // @[package.scala 154:13]
  wire  state_vec_365_right_subtree_state = state_vec_365[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_365_T_3 = state_vec_0_set_left_older ? state_vec_365_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_365_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_365_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_365_T_8 = {state_vec_0_set_left_older,_state_vec_365_T_3,_state_vec_365_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_366_valid = touch_way_0_valid & touch_set_0 == 9'h16e; // @[Replacement.scala 315:30]
  wire  state_vec_366_left_subtree_state = state_vec_366[1]; // @[package.scala 154:13]
  wire  state_vec_366_right_subtree_state = state_vec_366[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_366_T_3 = state_vec_0_set_left_older ? state_vec_366_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_366_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_366_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_366_T_8 = {state_vec_0_set_left_older,_state_vec_366_T_3,_state_vec_366_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_367_valid = touch_way_0_valid & touch_set_0 == 9'h16f; // @[Replacement.scala 315:30]
  wire  state_vec_367_left_subtree_state = state_vec_367[1]; // @[package.scala 154:13]
  wire  state_vec_367_right_subtree_state = state_vec_367[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_367_T_3 = state_vec_0_set_left_older ? state_vec_367_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_367_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_367_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_367_T_8 = {state_vec_0_set_left_older,_state_vec_367_T_3,_state_vec_367_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_368_valid = touch_way_0_valid & touch_set_0 == 9'h170; // @[Replacement.scala 315:30]
  wire  state_vec_368_left_subtree_state = state_vec_368[1]; // @[package.scala 154:13]
  wire  state_vec_368_right_subtree_state = state_vec_368[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_368_T_3 = state_vec_0_set_left_older ? state_vec_368_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_368_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_368_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_368_T_8 = {state_vec_0_set_left_older,_state_vec_368_T_3,_state_vec_368_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_369_valid = touch_way_0_valid & touch_set_0 == 9'h171; // @[Replacement.scala 315:30]
  wire  state_vec_369_left_subtree_state = state_vec_369[1]; // @[package.scala 154:13]
  wire  state_vec_369_right_subtree_state = state_vec_369[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_369_T_3 = state_vec_0_set_left_older ? state_vec_369_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_369_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_369_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_369_T_8 = {state_vec_0_set_left_older,_state_vec_369_T_3,_state_vec_369_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_370_valid = touch_way_0_valid & touch_set_0 == 9'h172; // @[Replacement.scala 315:30]
  wire  state_vec_370_left_subtree_state = state_vec_370[1]; // @[package.scala 154:13]
  wire  state_vec_370_right_subtree_state = state_vec_370[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_370_T_3 = state_vec_0_set_left_older ? state_vec_370_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_370_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_370_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_370_T_8 = {state_vec_0_set_left_older,_state_vec_370_T_3,_state_vec_370_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_371_valid = touch_way_0_valid & touch_set_0 == 9'h173; // @[Replacement.scala 315:30]
  wire  state_vec_371_left_subtree_state = state_vec_371[1]; // @[package.scala 154:13]
  wire  state_vec_371_right_subtree_state = state_vec_371[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_371_T_3 = state_vec_0_set_left_older ? state_vec_371_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_371_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_371_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_371_T_8 = {state_vec_0_set_left_older,_state_vec_371_T_3,_state_vec_371_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_372_valid = touch_way_0_valid & touch_set_0 == 9'h174; // @[Replacement.scala 315:30]
  wire  state_vec_372_left_subtree_state = state_vec_372[1]; // @[package.scala 154:13]
  wire  state_vec_372_right_subtree_state = state_vec_372[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_372_T_3 = state_vec_0_set_left_older ? state_vec_372_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_372_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_372_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_372_T_8 = {state_vec_0_set_left_older,_state_vec_372_T_3,_state_vec_372_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_373_valid = touch_way_0_valid & touch_set_0 == 9'h175; // @[Replacement.scala 315:30]
  wire  state_vec_373_left_subtree_state = state_vec_373[1]; // @[package.scala 154:13]
  wire  state_vec_373_right_subtree_state = state_vec_373[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_373_T_3 = state_vec_0_set_left_older ? state_vec_373_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_373_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_373_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_373_T_8 = {state_vec_0_set_left_older,_state_vec_373_T_3,_state_vec_373_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_374_valid = touch_way_0_valid & touch_set_0 == 9'h176; // @[Replacement.scala 315:30]
  wire  state_vec_374_left_subtree_state = state_vec_374[1]; // @[package.scala 154:13]
  wire  state_vec_374_right_subtree_state = state_vec_374[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_374_T_3 = state_vec_0_set_left_older ? state_vec_374_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_374_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_374_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_374_T_8 = {state_vec_0_set_left_older,_state_vec_374_T_3,_state_vec_374_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_375_valid = touch_way_0_valid & touch_set_0 == 9'h177; // @[Replacement.scala 315:30]
  wire  state_vec_375_left_subtree_state = state_vec_375[1]; // @[package.scala 154:13]
  wire  state_vec_375_right_subtree_state = state_vec_375[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_375_T_3 = state_vec_0_set_left_older ? state_vec_375_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_375_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_375_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_375_T_8 = {state_vec_0_set_left_older,_state_vec_375_T_3,_state_vec_375_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_376_valid = touch_way_0_valid & touch_set_0 == 9'h178; // @[Replacement.scala 315:30]
  wire  state_vec_376_left_subtree_state = state_vec_376[1]; // @[package.scala 154:13]
  wire  state_vec_376_right_subtree_state = state_vec_376[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_376_T_3 = state_vec_0_set_left_older ? state_vec_376_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_376_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_376_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_376_T_8 = {state_vec_0_set_left_older,_state_vec_376_T_3,_state_vec_376_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_377_valid = touch_way_0_valid & touch_set_0 == 9'h179; // @[Replacement.scala 315:30]
  wire  state_vec_377_left_subtree_state = state_vec_377[1]; // @[package.scala 154:13]
  wire  state_vec_377_right_subtree_state = state_vec_377[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_377_T_3 = state_vec_0_set_left_older ? state_vec_377_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_377_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_377_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_377_T_8 = {state_vec_0_set_left_older,_state_vec_377_T_3,_state_vec_377_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_378_valid = touch_way_0_valid & touch_set_0 == 9'h17a; // @[Replacement.scala 315:30]
  wire  state_vec_378_left_subtree_state = state_vec_378[1]; // @[package.scala 154:13]
  wire  state_vec_378_right_subtree_state = state_vec_378[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_378_T_3 = state_vec_0_set_left_older ? state_vec_378_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_378_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_378_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_378_T_8 = {state_vec_0_set_left_older,_state_vec_378_T_3,_state_vec_378_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_379_valid = touch_way_0_valid & touch_set_0 == 9'h17b; // @[Replacement.scala 315:30]
  wire  state_vec_379_left_subtree_state = state_vec_379[1]; // @[package.scala 154:13]
  wire  state_vec_379_right_subtree_state = state_vec_379[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_379_T_3 = state_vec_0_set_left_older ? state_vec_379_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_379_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_379_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_379_T_8 = {state_vec_0_set_left_older,_state_vec_379_T_3,_state_vec_379_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_380_valid = touch_way_0_valid & touch_set_0 == 9'h17c; // @[Replacement.scala 315:30]
  wire  state_vec_380_left_subtree_state = state_vec_380[1]; // @[package.scala 154:13]
  wire  state_vec_380_right_subtree_state = state_vec_380[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_380_T_3 = state_vec_0_set_left_older ? state_vec_380_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_380_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_380_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_380_T_8 = {state_vec_0_set_left_older,_state_vec_380_T_3,_state_vec_380_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_381_valid = touch_way_0_valid & touch_set_0 == 9'h17d; // @[Replacement.scala 315:30]
  wire  state_vec_381_left_subtree_state = state_vec_381[1]; // @[package.scala 154:13]
  wire  state_vec_381_right_subtree_state = state_vec_381[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_381_T_3 = state_vec_0_set_left_older ? state_vec_381_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_381_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_381_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_381_T_8 = {state_vec_0_set_left_older,_state_vec_381_T_3,_state_vec_381_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_382_valid = touch_way_0_valid & touch_set_0 == 9'h17e; // @[Replacement.scala 315:30]
  wire  state_vec_382_left_subtree_state = state_vec_382[1]; // @[package.scala 154:13]
  wire  state_vec_382_right_subtree_state = state_vec_382[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_382_T_3 = state_vec_0_set_left_older ? state_vec_382_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_382_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_382_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_382_T_8 = {state_vec_0_set_left_older,_state_vec_382_T_3,_state_vec_382_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_383_valid = touch_way_0_valid & touch_set_0 == 9'h17f; // @[Replacement.scala 315:30]
  wire  state_vec_383_left_subtree_state = state_vec_383[1]; // @[package.scala 154:13]
  wire  state_vec_383_right_subtree_state = state_vec_383[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_383_T_3 = state_vec_0_set_left_older ? state_vec_383_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_383_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_383_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_383_T_8 = {state_vec_0_set_left_older,_state_vec_383_T_3,_state_vec_383_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_384_valid = touch_way_0_valid & touch_set_0 == 9'h180; // @[Replacement.scala 315:30]
  wire  state_vec_384_left_subtree_state = state_vec_384[1]; // @[package.scala 154:13]
  wire  state_vec_384_right_subtree_state = state_vec_384[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_384_T_3 = state_vec_0_set_left_older ? state_vec_384_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_384_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_384_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_384_T_8 = {state_vec_0_set_left_older,_state_vec_384_T_3,_state_vec_384_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_385_valid = touch_way_0_valid & touch_set_0 == 9'h181; // @[Replacement.scala 315:30]
  wire  state_vec_385_left_subtree_state = state_vec_385[1]; // @[package.scala 154:13]
  wire  state_vec_385_right_subtree_state = state_vec_385[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_385_T_3 = state_vec_0_set_left_older ? state_vec_385_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_385_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_385_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_385_T_8 = {state_vec_0_set_left_older,_state_vec_385_T_3,_state_vec_385_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_386_valid = touch_way_0_valid & touch_set_0 == 9'h182; // @[Replacement.scala 315:30]
  wire  state_vec_386_left_subtree_state = state_vec_386[1]; // @[package.scala 154:13]
  wire  state_vec_386_right_subtree_state = state_vec_386[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_386_T_3 = state_vec_0_set_left_older ? state_vec_386_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_386_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_386_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_386_T_8 = {state_vec_0_set_left_older,_state_vec_386_T_3,_state_vec_386_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_387_valid = touch_way_0_valid & touch_set_0 == 9'h183; // @[Replacement.scala 315:30]
  wire  state_vec_387_left_subtree_state = state_vec_387[1]; // @[package.scala 154:13]
  wire  state_vec_387_right_subtree_state = state_vec_387[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_387_T_3 = state_vec_0_set_left_older ? state_vec_387_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_387_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_387_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_387_T_8 = {state_vec_0_set_left_older,_state_vec_387_T_3,_state_vec_387_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_388_valid = touch_way_0_valid & touch_set_0 == 9'h184; // @[Replacement.scala 315:30]
  wire  state_vec_388_left_subtree_state = state_vec_388[1]; // @[package.scala 154:13]
  wire  state_vec_388_right_subtree_state = state_vec_388[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_388_T_3 = state_vec_0_set_left_older ? state_vec_388_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_388_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_388_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_388_T_8 = {state_vec_0_set_left_older,_state_vec_388_T_3,_state_vec_388_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_389_valid = touch_way_0_valid & touch_set_0 == 9'h185; // @[Replacement.scala 315:30]
  wire  state_vec_389_left_subtree_state = state_vec_389[1]; // @[package.scala 154:13]
  wire  state_vec_389_right_subtree_state = state_vec_389[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_389_T_3 = state_vec_0_set_left_older ? state_vec_389_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_389_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_389_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_389_T_8 = {state_vec_0_set_left_older,_state_vec_389_T_3,_state_vec_389_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_390_valid = touch_way_0_valid & touch_set_0 == 9'h186; // @[Replacement.scala 315:30]
  wire  state_vec_390_left_subtree_state = state_vec_390[1]; // @[package.scala 154:13]
  wire  state_vec_390_right_subtree_state = state_vec_390[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_390_T_3 = state_vec_0_set_left_older ? state_vec_390_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_390_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_390_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_390_T_8 = {state_vec_0_set_left_older,_state_vec_390_T_3,_state_vec_390_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_391_valid = touch_way_0_valid & touch_set_0 == 9'h187; // @[Replacement.scala 315:30]
  wire  state_vec_391_left_subtree_state = state_vec_391[1]; // @[package.scala 154:13]
  wire  state_vec_391_right_subtree_state = state_vec_391[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_391_T_3 = state_vec_0_set_left_older ? state_vec_391_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_391_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_391_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_391_T_8 = {state_vec_0_set_left_older,_state_vec_391_T_3,_state_vec_391_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_392_valid = touch_way_0_valid & touch_set_0 == 9'h188; // @[Replacement.scala 315:30]
  wire  state_vec_392_left_subtree_state = state_vec_392[1]; // @[package.scala 154:13]
  wire  state_vec_392_right_subtree_state = state_vec_392[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_392_T_3 = state_vec_0_set_left_older ? state_vec_392_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_392_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_392_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_392_T_8 = {state_vec_0_set_left_older,_state_vec_392_T_3,_state_vec_392_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_393_valid = touch_way_0_valid & touch_set_0 == 9'h189; // @[Replacement.scala 315:30]
  wire  state_vec_393_left_subtree_state = state_vec_393[1]; // @[package.scala 154:13]
  wire  state_vec_393_right_subtree_state = state_vec_393[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_393_T_3 = state_vec_0_set_left_older ? state_vec_393_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_393_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_393_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_393_T_8 = {state_vec_0_set_left_older,_state_vec_393_T_3,_state_vec_393_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_394_valid = touch_way_0_valid & touch_set_0 == 9'h18a; // @[Replacement.scala 315:30]
  wire  state_vec_394_left_subtree_state = state_vec_394[1]; // @[package.scala 154:13]
  wire  state_vec_394_right_subtree_state = state_vec_394[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_394_T_3 = state_vec_0_set_left_older ? state_vec_394_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_394_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_394_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_394_T_8 = {state_vec_0_set_left_older,_state_vec_394_T_3,_state_vec_394_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_395_valid = touch_way_0_valid & touch_set_0 == 9'h18b; // @[Replacement.scala 315:30]
  wire  state_vec_395_left_subtree_state = state_vec_395[1]; // @[package.scala 154:13]
  wire  state_vec_395_right_subtree_state = state_vec_395[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_395_T_3 = state_vec_0_set_left_older ? state_vec_395_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_395_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_395_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_395_T_8 = {state_vec_0_set_left_older,_state_vec_395_T_3,_state_vec_395_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_396_valid = touch_way_0_valid & touch_set_0 == 9'h18c; // @[Replacement.scala 315:30]
  wire  state_vec_396_left_subtree_state = state_vec_396[1]; // @[package.scala 154:13]
  wire  state_vec_396_right_subtree_state = state_vec_396[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_396_T_3 = state_vec_0_set_left_older ? state_vec_396_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_396_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_396_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_396_T_8 = {state_vec_0_set_left_older,_state_vec_396_T_3,_state_vec_396_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_397_valid = touch_way_0_valid & touch_set_0 == 9'h18d; // @[Replacement.scala 315:30]
  wire  state_vec_397_left_subtree_state = state_vec_397[1]; // @[package.scala 154:13]
  wire  state_vec_397_right_subtree_state = state_vec_397[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_397_T_3 = state_vec_0_set_left_older ? state_vec_397_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_397_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_397_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_397_T_8 = {state_vec_0_set_left_older,_state_vec_397_T_3,_state_vec_397_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_398_valid = touch_way_0_valid & touch_set_0 == 9'h18e; // @[Replacement.scala 315:30]
  wire  state_vec_398_left_subtree_state = state_vec_398[1]; // @[package.scala 154:13]
  wire  state_vec_398_right_subtree_state = state_vec_398[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_398_T_3 = state_vec_0_set_left_older ? state_vec_398_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_398_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_398_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_398_T_8 = {state_vec_0_set_left_older,_state_vec_398_T_3,_state_vec_398_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_399_valid = touch_way_0_valid & touch_set_0 == 9'h18f; // @[Replacement.scala 315:30]
  wire  state_vec_399_left_subtree_state = state_vec_399[1]; // @[package.scala 154:13]
  wire  state_vec_399_right_subtree_state = state_vec_399[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_399_T_3 = state_vec_0_set_left_older ? state_vec_399_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_399_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_399_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_399_T_8 = {state_vec_0_set_left_older,_state_vec_399_T_3,_state_vec_399_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_400_valid = touch_way_0_valid & touch_set_0 == 9'h190; // @[Replacement.scala 315:30]
  wire  state_vec_400_left_subtree_state = state_vec_400[1]; // @[package.scala 154:13]
  wire  state_vec_400_right_subtree_state = state_vec_400[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_400_T_3 = state_vec_0_set_left_older ? state_vec_400_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_400_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_400_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_400_T_8 = {state_vec_0_set_left_older,_state_vec_400_T_3,_state_vec_400_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_401_valid = touch_way_0_valid & touch_set_0 == 9'h191; // @[Replacement.scala 315:30]
  wire  state_vec_401_left_subtree_state = state_vec_401[1]; // @[package.scala 154:13]
  wire  state_vec_401_right_subtree_state = state_vec_401[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_401_T_3 = state_vec_0_set_left_older ? state_vec_401_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_401_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_401_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_401_T_8 = {state_vec_0_set_left_older,_state_vec_401_T_3,_state_vec_401_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_402_valid = touch_way_0_valid & touch_set_0 == 9'h192; // @[Replacement.scala 315:30]
  wire  state_vec_402_left_subtree_state = state_vec_402[1]; // @[package.scala 154:13]
  wire  state_vec_402_right_subtree_state = state_vec_402[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_402_T_3 = state_vec_0_set_left_older ? state_vec_402_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_402_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_402_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_402_T_8 = {state_vec_0_set_left_older,_state_vec_402_T_3,_state_vec_402_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_403_valid = touch_way_0_valid & touch_set_0 == 9'h193; // @[Replacement.scala 315:30]
  wire  state_vec_403_left_subtree_state = state_vec_403[1]; // @[package.scala 154:13]
  wire  state_vec_403_right_subtree_state = state_vec_403[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_403_T_3 = state_vec_0_set_left_older ? state_vec_403_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_403_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_403_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_403_T_8 = {state_vec_0_set_left_older,_state_vec_403_T_3,_state_vec_403_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_404_valid = touch_way_0_valid & touch_set_0 == 9'h194; // @[Replacement.scala 315:30]
  wire  state_vec_404_left_subtree_state = state_vec_404[1]; // @[package.scala 154:13]
  wire  state_vec_404_right_subtree_state = state_vec_404[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_404_T_3 = state_vec_0_set_left_older ? state_vec_404_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_404_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_404_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_404_T_8 = {state_vec_0_set_left_older,_state_vec_404_T_3,_state_vec_404_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_405_valid = touch_way_0_valid & touch_set_0 == 9'h195; // @[Replacement.scala 315:30]
  wire  state_vec_405_left_subtree_state = state_vec_405[1]; // @[package.scala 154:13]
  wire  state_vec_405_right_subtree_state = state_vec_405[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_405_T_3 = state_vec_0_set_left_older ? state_vec_405_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_405_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_405_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_405_T_8 = {state_vec_0_set_left_older,_state_vec_405_T_3,_state_vec_405_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_406_valid = touch_way_0_valid & touch_set_0 == 9'h196; // @[Replacement.scala 315:30]
  wire  state_vec_406_left_subtree_state = state_vec_406[1]; // @[package.scala 154:13]
  wire  state_vec_406_right_subtree_state = state_vec_406[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_406_T_3 = state_vec_0_set_left_older ? state_vec_406_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_406_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_406_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_406_T_8 = {state_vec_0_set_left_older,_state_vec_406_T_3,_state_vec_406_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_407_valid = touch_way_0_valid & touch_set_0 == 9'h197; // @[Replacement.scala 315:30]
  wire  state_vec_407_left_subtree_state = state_vec_407[1]; // @[package.scala 154:13]
  wire  state_vec_407_right_subtree_state = state_vec_407[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_407_T_3 = state_vec_0_set_left_older ? state_vec_407_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_407_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_407_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_407_T_8 = {state_vec_0_set_left_older,_state_vec_407_T_3,_state_vec_407_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_408_valid = touch_way_0_valid & touch_set_0 == 9'h198; // @[Replacement.scala 315:30]
  wire  state_vec_408_left_subtree_state = state_vec_408[1]; // @[package.scala 154:13]
  wire  state_vec_408_right_subtree_state = state_vec_408[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_408_T_3 = state_vec_0_set_left_older ? state_vec_408_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_408_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_408_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_408_T_8 = {state_vec_0_set_left_older,_state_vec_408_T_3,_state_vec_408_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_409_valid = touch_way_0_valid & touch_set_0 == 9'h199; // @[Replacement.scala 315:30]
  wire  state_vec_409_left_subtree_state = state_vec_409[1]; // @[package.scala 154:13]
  wire  state_vec_409_right_subtree_state = state_vec_409[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_409_T_3 = state_vec_0_set_left_older ? state_vec_409_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_409_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_409_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_409_T_8 = {state_vec_0_set_left_older,_state_vec_409_T_3,_state_vec_409_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_410_valid = touch_way_0_valid & touch_set_0 == 9'h19a; // @[Replacement.scala 315:30]
  wire  state_vec_410_left_subtree_state = state_vec_410[1]; // @[package.scala 154:13]
  wire  state_vec_410_right_subtree_state = state_vec_410[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_410_T_3 = state_vec_0_set_left_older ? state_vec_410_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_410_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_410_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_410_T_8 = {state_vec_0_set_left_older,_state_vec_410_T_3,_state_vec_410_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_411_valid = touch_way_0_valid & touch_set_0 == 9'h19b; // @[Replacement.scala 315:30]
  wire  state_vec_411_left_subtree_state = state_vec_411[1]; // @[package.scala 154:13]
  wire  state_vec_411_right_subtree_state = state_vec_411[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_411_T_3 = state_vec_0_set_left_older ? state_vec_411_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_411_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_411_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_411_T_8 = {state_vec_0_set_left_older,_state_vec_411_T_3,_state_vec_411_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_412_valid = touch_way_0_valid & touch_set_0 == 9'h19c; // @[Replacement.scala 315:30]
  wire  state_vec_412_left_subtree_state = state_vec_412[1]; // @[package.scala 154:13]
  wire  state_vec_412_right_subtree_state = state_vec_412[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_412_T_3 = state_vec_0_set_left_older ? state_vec_412_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_412_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_412_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_412_T_8 = {state_vec_0_set_left_older,_state_vec_412_T_3,_state_vec_412_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_413_valid = touch_way_0_valid & touch_set_0 == 9'h19d; // @[Replacement.scala 315:30]
  wire  state_vec_413_left_subtree_state = state_vec_413[1]; // @[package.scala 154:13]
  wire  state_vec_413_right_subtree_state = state_vec_413[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_413_T_3 = state_vec_0_set_left_older ? state_vec_413_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_413_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_413_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_413_T_8 = {state_vec_0_set_left_older,_state_vec_413_T_3,_state_vec_413_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_414_valid = touch_way_0_valid & touch_set_0 == 9'h19e; // @[Replacement.scala 315:30]
  wire  state_vec_414_left_subtree_state = state_vec_414[1]; // @[package.scala 154:13]
  wire  state_vec_414_right_subtree_state = state_vec_414[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_414_T_3 = state_vec_0_set_left_older ? state_vec_414_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_414_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_414_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_414_T_8 = {state_vec_0_set_left_older,_state_vec_414_T_3,_state_vec_414_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_415_valid = touch_way_0_valid & touch_set_0 == 9'h19f; // @[Replacement.scala 315:30]
  wire  state_vec_415_left_subtree_state = state_vec_415[1]; // @[package.scala 154:13]
  wire  state_vec_415_right_subtree_state = state_vec_415[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_415_T_3 = state_vec_0_set_left_older ? state_vec_415_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_415_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_415_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_415_T_8 = {state_vec_0_set_left_older,_state_vec_415_T_3,_state_vec_415_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_416_valid = touch_way_0_valid & touch_set_0 == 9'h1a0; // @[Replacement.scala 315:30]
  wire  state_vec_416_left_subtree_state = state_vec_416[1]; // @[package.scala 154:13]
  wire  state_vec_416_right_subtree_state = state_vec_416[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_416_T_3 = state_vec_0_set_left_older ? state_vec_416_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_416_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_416_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_416_T_8 = {state_vec_0_set_left_older,_state_vec_416_T_3,_state_vec_416_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_417_valid = touch_way_0_valid & touch_set_0 == 9'h1a1; // @[Replacement.scala 315:30]
  wire  state_vec_417_left_subtree_state = state_vec_417[1]; // @[package.scala 154:13]
  wire  state_vec_417_right_subtree_state = state_vec_417[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_417_T_3 = state_vec_0_set_left_older ? state_vec_417_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_417_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_417_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_417_T_8 = {state_vec_0_set_left_older,_state_vec_417_T_3,_state_vec_417_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_418_valid = touch_way_0_valid & touch_set_0 == 9'h1a2; // @[Replacement.scala 315:30]
  wire  state_vec_418_left_subtree_state = state_vec_418[1]; // @[package.scala 154:13]
  wire  state_vec_418_right_subtree_state = state_vec_418[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_418_T_3 = state_vec_0_set_left_older ? state_vec_418_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_418_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_418_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_418_T_8 = {state_vec_0_set_left_older,_state_vec_418_T_3,_state_vec_418_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_419_valid = touch_way_0_valid & touch_set_0 == 9'h1a3; // @[Replacement.scala 315:30]
  wire  state_vec_419_left_subtree_state = state_vec_419[1]; // @[package.scala 154:13]
  wire  state_vec_419_right_subtree_state = state_vec_419[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_419_T_3 = state_vec_0_set_left_older ? state_vec_419_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_419_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_419_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_419_T_8 = {state_vec_0_set_left_older,_state_vec_419_T_3,_state_vec_419_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_420_valid = touch_way_0_valid & touch_set_0 == 9'h1a4; // @[Replacement.scala 315:30]
  wire  state_vec_420_left_subtree_state = state_vec_420[1]; // @[package.scala 154:13]
  wire  state_vec_420_right_subtree_state = state_vec_420[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_420_T_3 = state_vec_0_set_left_older ? state_vec_420_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_420_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_420_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_420_T_8 = {state_vec_0_set_left_older,_state_vec_420_T_3,_state_vec_420_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_421_valid = touch_way_0_valid & touch_set_0 == 9'h1a5; // @[Replacement.scala 315:30]
  wire  state_vec_421_left_subtree_state = state_vec_421[1]; // @[package.scala 154:13]
  wire  state_vec_421_right_subtree_state = state_vec_421[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_421_T_3 = state_vec_0_set_left_older ? state_vec_421_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_421_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_421_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_421_T_8 = {state_vec_0_set_left_older,_state_vec_421_T_3,_state_vec_421_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_422_valid = touch_way_0_valid & touch_set_0 == 9'h1a6; // @[Replacement.scala 315:30]
  wire  state_vec_422_left_subtree_state = state_vec_422[1]; // @[package.scala 154:13]
  wire  state_vec_422_right_subtree_state = state_vec_422[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_422_T_3 = state_vec_0_set_left_older ? state_vec_422_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_422_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_422_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_422_T_8 = {state_vec_0_set_left_older,_state_vec_422_T_3,_state_vec_422_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_423_valid = touch_way_0_valid & touch_set_0 == 9'h1a7; // @[Replacement.scala 315:30]
  wire  state_vec_423_left_subtree_state = state_vec_423[1]; // @[package.scala 154:13]
  wire  state_vec_423_right_subtree_state = state_vec_423[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_423_T_3 = state_vec_0_set_left_older ? state_vec_423_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_423_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_423_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_423_T_8 = {state_vec_0_set_left_older,_state_vec_423_T_3,_state_vec_423_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_424_valid = touch_way_0_valid & touch_set_0 == 9'h1a8; // @[Replacement.scala 315:30]
  wire  state_vec_424_left_subtree_state = state_vec_424[1]; // @[package.scala 154:13]
  wire  state_vec_424_right_subtree_state = state_vec_424[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_424_T_3 = state_vec_0_set_left_older ? state_vec_424_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_424_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_424_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_424_T_8 = {state_vec_0_set_left_older,_state_vec_424_T_3,_state_vec_424_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_425_valid = touch_way_0_valid & touch_set_0 == 9'h1a9; // @[Replacement.scala 315:30]
  wire  state_vec_425_left_subtree_state = state_vec_425[1]; // @[package.scala 154:13]
  wire  state_vec_425_right_subtree_state = state_vec_425[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_425_T_3 = state_vec_0_set_left_older ? state_vec_425_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_425_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_425_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_425_T_8 = {state_vec_0_set_left_older,_state_vec_425_T_3,_state_vec_425_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_426_valid = touch_way_0_valid & touch_set_0 == 9'h1aa; // @[Replacement.scala 315:30]
  wire  state_vec_426_left_subtree_state = state_vec_426[1]; // @[package.scala 154:13]
  wire  state_vec_426_right_subtree_state = state_vec_426[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_426_T_3 = state_vec_0_set_left_older ? state_vec_426_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_426_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_426_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_426_T_8 = {state_vec_0_set_left_older,_state_vec_426_T_3,_state_vec_426_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_427_valid = touch_way_0_valid & touch_set_0 == 9'h1ab; // @[Replacement.scala 315:30]
  wire  state_vec_427_left_subtree_state = state_vec_427[1]; // @[package.scala 154:13]
  wire  state_vec_427_right_subtree_state = state_vec_427[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_427_T_3 = state_vec_0_set_left_older ? state_vec_427_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_427_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_427_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_427_T_8 = {state_vec_0_set_left_older,_state_vec_427_T_3,_state_vec_427_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_428_valid = touch_way_0_valid & touch_set_0 == 9'h1ac; // @[Replacement.scala 315:30]
  wire  state_vec_428_left_subtree_state = state_vec_428[1]; // @[package.scala 154:13]
  wire  state_vec_428_right_subtree_state = state_vec_428[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_428_T_3 = state_vec_0_set_left_older ? state_vec_428_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_428_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_428_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_428_T_8 = {state_vec_0_set_left_older,_state_vec_428_T_3,_state_vec_428_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_429_valid = touch_way_0_valid & touch_set_0 == 9'h1ad; // @[Replacement.scala 315:30]
  wire  state_vec_429_left_subtree_state = state_vec_429[1]; // @[package.scala 154:13]
  wire  state_vec_429_right_subtree_state = state_vec_429[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_429_T_3 = state_vec_0_set_left_older ? state_vec_429_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_429_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_429_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_429_T_8 = {state_vec_0_set_left_older,_state_vec_429_T_3,_state_vec_429_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_430_valid = touch_way_0_valid & touch_set_0 == 9'h1ae; // @[Replacement.scala 315:30]
  wire  state_vec_430_left_subtree_state = state_vec_430[1]; // @[package.scala 154:13]
  wire  state_vec_430_right_subtree_state = state_vec_430[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_430_T_3 = state_vec_0_set_left_older ? state_vec_430_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_430_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_430_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_430_T_8 = {state_vec_0_set_left_older,_state_vec_430_T_3,_state_vec_430_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_431_valid = touch_way_0_valid & touch_set_0 == 9'h1af; // @[Replacement.scala 315:30]
  wire  state_vec_431_left_subtree_state = state_vec_431[1]; // @[package.scala 154:13]
  wire  state_vec_431_right_subtree_state = state_vec_431[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_431_T_3 = state_vec_0_set_left_older ? state_vec_431_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_431_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_431_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_431_T_8 = {state_vec_0_set_left_older,_state_vec_431_T_3,_state_vec_431_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_432_valid = touch_way_0_valid & touch_set_0 == 9'h1b0; // @[Replacement.scala 315:30]
  wire  state_vec_432_left_subtree_state = state_vec_432[1]; // @[package.scala 154:13]
  wire  state_vec_432_right_subtree_state = state_vec_432[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_432_T_3 = state_vec_0_set_left_older ? state_vec_432_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_432_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_432_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_432_T_8 = {state_vec_0_set_left_older,_state_vec_432_T_3,_state_vec_432_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_433_valid = touch_way_0_valid & touch_set_0 == 9'h1b1; // @[Replacement.scala 315:30]
  wire  state_vec_433_left_subtree_state = state_vec_433[1]; // @[package.scala 154:13]
  wire  state_vec_433_right_subtree_state = state_vec_433[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_433_T_3 = state_vec_0_set_left_older ? state_vec_433_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_433_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_433_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_433_T_8 = {state_vec_0_set_left_older,_state_vec_433_T_3,_state_vec_433_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_434_valid = touch_way_0_valid & touch_set_0 == 9'h1b2; // @[Replacement.scala 315:30]
  wire  state_vec_434_left_subtree_state = state_vec_434[1]; // @[package.scala 154:13]
  wire  state_vec_434_right_subtree_state = state_vec_434[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_434_T_3 = state_vec_0_set_left_older ? state_vec_434_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_434_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_434_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_434_T_8 = {state_vec_0_set_left_older,_state_vec_434_T_3,_state_vec_434_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_435_valid = touch_way_0_valid & touch_set_0 == 9'h1b3; // @[Replacement.scala 315:30]
  wire  state_vec_435_left_subtree_state = state_vec_435[1]; // @[package.scala 154:13]
  wire  state_vec_435_right_subtree_state = state_vec_435[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_435_T_3 = state_vec_0_set_left_older ? state_vec_435_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_435_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_435_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_435_T_8 = {state_vec_0_set_left_older,_state_vec_435_T_3,_state_vec_435_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_436_valid = touch_way_0_valid & touch_set_0 == 9'h1b4; // @[Replacement.scala 315:30]
  wire  state_vec_436_left_subtree_state = state_vec_436[1]; // @[package.scala 154:13]
  wire  state_vec_436_right_subtree_state = state_vec_436[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_436_T_3 = state_vec_0_set_left_older ? state_vec_436_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_436_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_436_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_436_T_8 = {state_vec_0_set_left_older,_state_vec_436_T_3,_state_vec_436_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_437_valid = touch_way_0_valid & touch_set_0 == 9'h1b5; // @[Replacement.scala 315:30]
  wire  state_vec_437_left_subtree_state = state_vec_437[1]; // @[package.scala 154:13]
  wire  state_vec_437_right_subtree_state = state_vec_437[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_437_T_3 = state_vec_0_set_left_older ? state_vec_437_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_437_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_437_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_437_T_8 = {state_vec_0_set_left_older,_state_vec_437_T_3,_state_vec_437_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_438_valid = touch_way_0_valid & touch_set_0 == 9'h1b6; // @[Replacement.scala 315:30]
  wire  state_vec_438_left_subtree_state = state_vec_438[1]; // @[package.scala 154:13]
  wire  state_vec_438_right_subtree_state = state_vec_438[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_438_T_3 = state_vec_0_set_left_older ? state_vec_438_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_438_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_438_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_438_T_8 = {state_vec_0_set_left_older,_state_vec_438_T_3,_state_vec_438_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_439_valid = touch_way_0_valid & touch_set_0 == 9'h1b7; // @[Replacement.scala 315:30]
  wire  state_vec_439_left_subtree_state = state_vec_439[1]; // @[package.scala 154:13]
  wire  state_vec_439_right_subtree_state = state_vec_439[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_439_T_3 = state_vec_0_set_left_older ? state_vec_439_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_439_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_439_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_439_T_8 = {state_vec_0_set_left_older,_state_vec_439_T_3,_state_vec_439_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_440_valid = touch_way_0_valid & touch_set_0 == 9'h1b8; // @[Replacement.scala 315:30]
  wire  state_vec_440_left_subtree_state = state_vec_440[1]; // @[package.scala 154:13]
  wire  state_vec_440_right_subtree_state = state_vec_440[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_440_T_3 = state_vec_0_set_left_older ? state_vec_440_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_440_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_440_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_440_T_8 = {state_vec_0_set_left_older,_state_vec_440_T_3,_state_vec_440_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_441_valid = touch_way_0_valid & touch_set_0 == 9'h1b9; // @[Replacement.scala 315:30]
  wire  state_vec_441_left_subtree_state = state_vec_441[1]; // @[package.scala 154:13]
  wire  state_vec_441_right_subtree_state = state_vec_441[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_441_T_3 = state_vec_0_set_left_older ? state_vec_441_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_441_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_441_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_441_T_8 = {state_vec_0_set_left_older,_state_vec_441_T_3,_state_vec_441_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_442_valid = touch_way_0_valid & touch_set_0 == 9'h1ba; // @[Replacement.scala 315:30]
  wire  state_vec_442_left_subtree_state = state_vec_442[1]; // @[package.scala 154:13]
  wire  state_vec_442_right_subtree_state = state_vec_442[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_442_T_3 = state_vec_0_set_left_older ? state_vec_442_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_442_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_442_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_442_T_8 = {state_vec_0_set_left_older,_state_vec_442_T_3,_state_vec_442_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_443_valid = touch_way_0_valid & touch_set_0 == 9'h1bb; // @[Replacement.scala 315:30]
  wire  state_vec_443_left_subtree_state = state_vec_443[1]; // @[package.scala 154:13]
  wire  state_vec_443_right_subtree_state = state_vec_443[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_443_T_3 = state_vec_0_set_left_older ? state_vec_443_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_443_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_443_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_443_T_8 = {state_vec_0_set_left_older,_state_vec_443_T_3,_state_vec_443_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_444_valid = touch_way_0_valid & touch_set_0 == 9'h1bc; // @[Replacement.scala 315:30]
  wire  state_vec_444_left_subtree_state = state_vec_444[1]; // @[package.scala 154:13]
  wire  state_vec_444_right_subtree_state = state_vec_444[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_444_T_3 = state_vec_0_set_left_older ? state_vec_444_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_444_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_444_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_444_T_8 = {state_vec_0_set_left_older,_state_vec_444_T_3,_state_vec_444_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_445_valid = touch_way_0_valid & touch_set_0 == 9'h1bd; // @[Replacement.scala 315:30]
  wire  state_vec_445_left_subtree_state = state_vec_445[1]; // @[package.scala 154:13]
  wire  state_vec_445_right_subtree_state = state_vec_445[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_445_T_3 = state_vec_0_set_left_older ? state_vec_445_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_445_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_445_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_445_T_8 = {state_vec_0_set_left_older,_state_vec_445_T_3,_state_vec_445_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_446_valid = touch_way_0_valid & touch_set_0 == 9'h1be; // @[Replacement.scala 315:30]
  wire  state_vec_446_left_subtree_state = state_vec_446[1]; // @[package.scala 154:13]
  wire  state_vec_446_right_subtree_state = state_vec_446[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_446_T_3 = state_vec_0_set_left_older ? state_vec_446_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_446_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_446_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_446_T_8 = {state_vec_0_set_left_older,_state_vec_446_T_3,_state_vec_446_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_447_valid = touch_way_0_valid & touch_set_0 == 9'h1bf; // @[Replacement.scala 315:30]
  wire  state_vec_447_left_subtree_state = state_vec_447[1]; // @[package.scala 154:13]
  wire  state_vec_447_right_subtree_state = state_vec_447[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_447_T_3 = state_vec_0_set_left_older ? state_vec_447_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_447_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_447_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_447_T_8 = {state_vec_0_set_left_older,_state_vec_447_T_3,_state_vec_447_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_448_valid = touch_way_0_valid & touch_set_0 == 9'h1c0; // @[Replacement.scala 315:30]
  wire  state_vec_448_left_subtree_state = state_vec_448[1]; // @[package.scala 154:13]
  wire  state_vec_448_right_subtree_state = state_vec_448[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_448_T_3 = state_vec_0_set_left_older ? state_vec_448_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_448_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_448_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_448_T_8 = {state_vec_0_set_left_older,_state_vec_448_T_3,_state_vec_448_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_449_valid = touch_way_0_valid & touch_set_0 == 9'h1c1; // @[Replacement.scala 315:30]
  wire  state_vec_449_left_subtree_state = state_vec_449[1]; // @[package.scala 154:13]
  wire  state_vec_449_right_subtree_state = state_vec_449[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_449_T_3 = state_vec_0_set_left_older ? state_vec_449_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_449_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_449_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_449_T_8 = {state_vec_0_set_left_older,_state_vec_449_T_3,_state_vec_449_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_450_valid = touch_way_0_valid & touch_set_0 == 9'h1c2; // @[Replacement.scala 315:30]
  wire  state_vec_450_left_subtree_state = state_vec_450[1]; // @[package.scala 154:13]
  wire  state_vec_450_right_subtree_state = state_vec_450[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_450_T_3 = state_vec_0_set_left_older ? state_vec_450_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_450_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_450_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_450_T_8 = {state_vec_0_set_left_older,_state_vec_450_T_3,_state_vec_450_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_451_valid = touch_way_0_valid & touch_set_0 == 9'h1c3; // @[Replacement.scala 315:30]
  wire  state_vec_451_left_subtree_state = state_vec_451[1]; // @[package.scala 154:13]
  wire  state_vec_451_right_subtree_state = state_vec_451[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_451_T_3 = state_vec_0_set_left_older ? state_vec_451_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_451_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_451_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_451_T_8 = {state_vec_0_set_left_older,_state_vec_451_T_3,_state_vec_451_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_452_valid = touch_way_0_valid & touch_set_0 == 9'h1c4; // @[Replacement.scala 315:30]
  wire  state_vec_452_left_subtree_state = state_vec_452[1]; // @[package.scala 154:13]
  wire  state_vec_452_right_subtree_state = state_vec_452[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_452_T_3 = state_vec_0_set_left_older ? state_vec_452_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_452_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_452_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_452_T_8 = {state_vec_0_set_left_older,_state_vec_452_T_3,_state_vec_452_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_453_valid = touch_way_0_valid & touch_set_0 == 9'h1c5; // @[Replacement.scala 315:30]
  wire  state_vec_453_left_subtree_state = state_vec_453[1]; // @[package.scala 154:13]
  wire  state_vec_453_right_subtree_state = state_vec_453[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_453_T_3 = state_vec_0_set_left_older ? state_vec_453_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_453_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_453_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_453_T_8 = {state_vec_0_set_left_older,_state_vec_453_T_3,_state_vec_453_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_454_valid = touch_way_0_valid & touch_set_0 == 9'h1c6; // @[Replacement.scala 315:30]
  wire  state_vec_454_left_subtree_state = state_vec_454[1]; // @[package.scala 154:13]
  wire  state_vec_454_right_subtree_state = state_vec_454[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_454_T_3 = state_vec_0_set_left_older ? state_vec_454_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_454_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_454_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_454_T_8 = {state_vec_0_set_left_older,_state_vec_454_T_3,_state_vec_454_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_455_valid = touch_way_0_valid & touch_set_0 == 9'h1c7; // @[Replacement.scala 315:30]
  wire  state_vec_455_left_subtree_state = state_vec_455[1]; // @[package.scala 154:13]
  wire  state_vec_455_right_subtree_state = state_vec_455[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_455_T_3 = state_vec_0_set_left_older ? state_vec_455_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_455_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_455_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_455_T_8 = {state_vec_0_set_left_older,_state_vec_455_T_3,_state_vec_455_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_456_valid = touch_way_0_valid & touch_set_0 == 9'h1c8; // @[Replacement.scala 315:30]
  wire  state_vec_456_left_subtree_state = state_vec_456[1]; // @[package.scala 154:13]
  wire  state_vec_456_right_subtree_state = state_vec_456[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_456_T_3 = state_vec_0_set_left_older ? state_vec_456_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_456_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_456_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_456_T_8 = {state_vec_0_set_left_older,_state_vec_456_T_3,_state_vec_456_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_457_valid = touch_way_0_valid & touch_set_0 == 9'h1c9; // @[Replacement.scala 315:30]
  wire  state_vec_457_left_subtree_state = state_vec_457[1]; // @[package.scala 154:13]
  wire  state_vec_457_right_subtree_state = state_vec_457[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_457_T_3 = state_vec_0_set_left_older ? state_vec_457_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_457_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_457_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_457_T_8 = {state_vec_0_set_left_older,_state_vec_457_T_3,_state_vec_457_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_458_valid = touch_way_0_valid & touch_set_0 == 9'h1ca; // @[Replacement.scala 315:30]
  wire  state_vec_458_left_subtree_state = state_vec_458[1]; // @[package.scala 154:13]
  wire  state_vec_458_right_subtree_state = state_vec_458[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_458_T_3 = state_vec_0_set_left_older ? state_vec_458_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_458_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_458_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_458_T_8 = {state_vec_0_set_left_older,_state_vec_458_T_3,_state_vec_458_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_459_valid = touch_way_0_valid & touch_set_0 == 9'h1cb; // @[Replacement.scala 315:30]
  wire  state_vec_459_left_subtree_state = state_vec_459[1]; // @[package.scala 154:13]
  wire  state_vec_459_right_subtree_state = state_vec_459[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_459_T_3 = state_vec_0_set_left_older ? state_vec_459_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_459_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_459_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_459_T_8 = {state_vec_0_set_left_older,_state_vec_459_T_3,_state_vec_459_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_460_valid = touch_way_0_valid & touch_set_0 == 9'h1cc; // @[Replacement.scala 315:30]
  wire  state_vec_460_left_subtree_state = state_vec_460[1]; // @[package.scala 154:13]
  wire  state_vec_460_right_subtree_state = state_vec_460[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_460_T_3 = state_vec_0_set_left_older ? state_vec_460_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_460_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_460_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_460_T_8 = {state_vec_0_set_left_older,_state_vec_460_T_3,_state_vec_460_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_461_valid = touch_way_0_valid & touch_set_0 == 9'h1cd; // @[Replacement.scala 315:30]
  wire  state_vec_461_left_subtree_state = state_vec_461[1]; // @[package.scala 154:13]
  wire  state_vec_461_right_subtree_state = state_vec_461[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_461_T_3 = state_vec_0_set_left_older ? state_vec_461_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_461_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_461_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_461_T_8 = {state_vec_0_set_left_older,_state_vec_461_T_3,_state_vec_461_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_462_valid = touch_way_0_valid & touch_set_0 == 9'h1ce; // @[Replacement.scala 315:30]
  wire  state_vec_462_left_subtree_state = state_vec_462[1]; // @[package.scala 154:13]
  wire  state_vec_462_right_subtree_state = state_vec_462[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_462_T_3 = state_vec_0_set_left_older ? state_vec_462_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_462_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_462_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_462_T_8 = {state_vec_0_set_left_older,_state_vec_462_T_3,_state_vec_462_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_463_valid = touch_way_0_valid & touch_set_0 == 9'h1cf; // @[Replacement.scala 315:30]
  wire  state_vec_463_left_subtree_state = state_vec_463[1]; // @[package.scala 154:13]
  wire  state_vec_463_right_subtree_state = state_vec_463[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_463_T_3 = state_vec_0_set_left_older ? state_vec_463_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_463_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_463_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_463_T_8 = {state_vec_0_set_left_older,_state_vec_463_T_3,_state_vec_463_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_464_valid = touch_way_0_valid & touch_set_0 == 9'h1d0; // @[Replacement.scala 315:30]
  wire  state_vec_464_left_subtree_state = state_vec_464[1]; // @[package.scala 154:13]
  wire  state_vec_464_right_subtree_state = state_vec_464[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_464_T_3 = state_vec_0_set_left_older ? state_vec_464_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_464_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_464_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_464_T_8 = {state_vec_0_set_left_older,_state_vec_464_T_3,_state_vec_464_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_465_valid = touch_way_0_valid & touch_set_0 == 9'h1d1; // @[Replacement.scala 315:30]
  wire  state_vec_465_left_subtree_state = state_vec_465[1]; // @[package.scala 154:13]
  wire  state_vec_465_right_subtree_state = state_vec_465[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_465_T_3 = state_vec_0_set_left_older ? state_vec_465_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_465_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_465_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_465_T_8 = {state_vec_0_set_left_older,_state_vec_465_T_3,_state_vec_465_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_466_valid = touch_way_0_valid & touch_set_0 == 9'h1d2; // @[Replacement.scala 315:30]
  wire  state_vec_466_left_subtree_state = state_vec_466[1]; // @[package.scala 154:13]
  wire  state_vec_466_right_subtree_state = state_vec_466[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_466_T_3 = state_vec_0_set_left_older ? state_vec_466_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_466_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_466_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_466_T_8 = {state_vec_0_set_left_older,_state_vec_466_T_3,_state_vec_466_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_467_valid = touch_way_0_valid & touch_set_0 == 9'h1d3; // @[Replacement.scala 315:30]
  wire  state_vec_467_left_subtree_state = state_vec_467[1]; // @[package.scala 154:13]
  wire  state_vec_467_right_subtree_state = state_vec_467[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_467_T_3 = state_vec_0_set_left_older ? state_vec_467_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_467_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_467_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_467_T_8 = {state_vec_0_set_left_older,_state_vec_467_T_3,_state_vec_467_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_468_valid = touch_way_0_valid & touch_set_0 == 9'h1d4; // @[Replacement.scala 315:30]
  wire  state_vec_468_left_subtree_state = state_vec_468[1]; // @[package.scala 154:13]
  wire  state_vec_468_right_subtree_state = state_vec_468[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_468_T_3 = state_vec_0_set_left_older ? state_vec_468_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_468_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_468_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_468_T_8 = {state_vec_0_set_left_older,_state_vec_468_T_3,_state_vec_468_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_469_valid = touch_way_0_valid & touch_set_0 == 9'h1d5; // @[Replacement.scala 315:30]
  wire  state_vec_469_left_subtree_state = state_vec_469[1]; // @[package.scala 154:13]
  wire  state_vec_469_right_subtree_state = state_vec_469[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_469_T_3 = state_vec_0_set_left_older ? state_vec_469_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_469_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_469_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_469_T_8 = {state_vec_0_set_left_older,_state_vec_469_T_3,_state_vec_469_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_470_valid = touch_way_0_valid & touch_set_0 == 9'h1d6; // @[Replacement.scala 315:30]
  wire  state_vec_470_left_subtree_state = state_vec_470[1]; // @[package.scala 154:13]
  wire  state_vec_470_right_subtree_state = state_vec_470[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_470_T_3 = state_vec_0_set_left_older ? state_vec_470_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_470_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_470_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_470_T_8 = {state_vec_0_set_left_older,_state_vec_470_T_3,_state_vec_470_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_471_valid = touch_way_0_valid & touch_set_0 == 9'h1d7; // @[Replacement.scala 315:30]
  wire  state_vec_471_left_subtree_state = state_vec_471[1]; // @[package.scala 154:13]
  wire  state_vec_471_right_subtree_state = state_vec_471[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_471_T_3 = state_vec_0_set_left_older ? state_vec_471_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_471_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_471_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_471_T_8 = {state_vec_0_set_left_older,_state_vec_471_T_3,_state_vec_471_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_472_valid = touch_way_0_valid & touch_set_0 == 9'h1d8; // @[Replacement.scala 315:30]
  wire  state_vec_472_left_subtree_state = state_vec_472[1]; // @[package.scala 154:13]
  wire  state_vec_472_right_subtree_state = state_vec_472[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_472_T_3 = state_vec_0_set_left_older ? state_vec_472_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_472_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_472_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_472_T_8 = {state_vec_0_set_left_older,_state_vec_472_T_3,_state_vec_472_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_473_valid = touch_way_0_valid & touch_set_0 == 9'h1d9; // @[Replacement.scala 315:30]
  wire  state_vec_473_left_subtree_state = state_vec_473[1]; // @[package.scala 154:13]
  wire  state_vec_473_right_subtree_state = state_vec_473[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_473_T_3 = state_vec_0_set_left_older ? state_vec_473_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_473_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_473_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_473_T_8 = {state_vec_0_set_left_older,_state_vec_473_T_3,_state_vec_473_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_474_valid = touch_way_0_valid & touch_set_0 == 9'h1da; // @[Replacement.scala 315:30]
  wire  state_vec_474_left_subtree_state = state_vec_474[1]; // @[package.scala 154:13]
  wire  state_vec_474_right_subtree_state = state_vec_474[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_474_T_3 = state_vec_0_set_left_older ? state_vec_474_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_474_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_474_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_474_T_8 = {state_vec_0_set_left_older,_state_vec_474_T_3,_state_vec_474_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_475_valid = touch_way_0_valid & touch_set_0 == 9'h1db; // @[Replacement.scala 315:30]
  wire  state_vec_475_left_subtree_state = state_vec_475[1]; // @[package.scala 154:13]
  wire  state_vec_475_right_subtree_state = state_vec_475[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_475_T_3 = state_vec_0_set_left_older ? state_vec_475_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_475_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_475_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_475_T_8 = {state_vec_0_set_left_older,_state_vec_475_T_3,_state_vec_475_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_476_valid = touch_way_0_valid & touch_set_0 == 9'h1dc; // @[Replacement.scala 315:30]
  wire  state_vec_476_left_subtree_state = state_vec_476[1]; // @[package.scala 154:13]
  wire  state_vec_476_right_subtree_state = state_vec_476[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_476_T_3 = state_vec_0_set_left_older ? state_vec_476_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_476_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_476_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_476_T_8 = {state_vec_0_set_left_older,_state_vec_476_T_3,_state_vec_476_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_477_valid = touch_way_0_valid & touch_set_0 == 9'h1dd; // @[Replacement.scala 315:30]
  wire  state_vec_477_left_subtree_state = state_vec_477[1]; // @[package.scala 154:13]
  wire  state_vec_477_right_subtree_state = state_vec_477[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_477_T_3 = state_vec_0_set_left_older ? state_vec_477_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_477_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_477_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_477_T_8 = {state_vec_0_set_left_older,_state_vec_477_T_3,_state_vec_477_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_478_valid = touch_way_0_valid & touch_set_0 == 9'h1de; // @[Replacement.scala 315:30]
  wire  state_vec_478_left_subtree_state = state_vec_478[1]; // @[package.scala 154:13]
  wire  state_vec_478_right_subtree_state = state_vec_478[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_478_T_3 = state_vec_0_set_left_older ? state_vec_478_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_478_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_478_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_478_T_8 = {state_vec_0_set_left_older,_state_vec_478_T_3,_state_vec_478_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_479_valid = touch_way_0_valid & touch_set_0 == 9'h1df; // @[Replacement.scala 315:30]
  wire  state_vec_479_left_subtree_state = state_vec_479[1]; // @[package.scala 154:13]
  wire  state_vec_479_right_subtree_state = state_vec_479[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_479_T_3 = state_vec_0_set_left_older ? state_vec_479_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_479_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_479_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_479_T_8 = {state_vec_0_set_left_older,_state_vec_479_T_3,_state_vec_479_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_480_valid = touch_way_0_valid & touch_set_0 == 9'h1e0; // @[Replacement.scala 315:30]
  wire  state_vec_480_left_subtree_state = state_vec_480[1]; // @[package.scala 154:13]
  wire  state_vec_480_right_subtree_state = state_vec_480[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_480_T_3 = state_vec_0_set_left_older ? state_vec_480_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_480_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_480_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_480_T_8 = {state_vec_0_set_left_older,_state_vec_480_T_3,_state_vec_480_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_481_valid = touch_way_0_valid & touch_set_0 == 9'h1e1; // @[Replacement.scala 315:30]
  wire  state_vec_481_left_subtree_state = state_vec_481[1]; // @[package.scala 154:13]
  wire  state_vec_481_right_subtree_state = state_vec_481[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_481_T_3 = state_vec_0_set_left_older ? state_vec_481_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_481_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_481_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_481_T_8 = {state_vec_0_set_left_older,_state_vec_481_T_3,_state_vec_481_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_482_valid = touch_way_0_valid & touch_set_0 == 9'h1e2; // @[Replacement.scala 315:30]
  wire  state_vec_482_left_subtree_state = state_vec_482[1]; // @[package.scala 154:13]
  wire  state_vec_482_right_subtree_state = state_vec_482[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_482_T_3 = state_vec_0_set_left_older ? state_vec_482_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_482_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_482_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_482_T_8 = {state_vec_0_set_left_older,_state_vec_482_T_3,_state_vec_482_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_483_valid = touch_way_0_valid & touch_set_0 == 9'h1e3; // @[Replacement.scala 315:30]
  wire  state_vec_483_left_subtree_state = state_vec_483[1]; // @[package.scala 154:13]
  wire  state_vec_483_right_subtree_state = state_vec_483[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_483_T_3 = state_vec_0_set_left_older ? state_vec_483_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_483_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_483_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_483_T_8 = {state_vec_0_set_left_older,_state_vec_483_T_3,_state_vec_483_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_484_valid = touch_way_0_valid & touch_set_0 == 9'h1e4; // @[Replacement.scala 315:30]
  wire  state_vec_484_left_subtree_state = state_vec_484[1]; // @[package.scala 154:13]
  wire  state_vec_484_right_subtree_state = state_vec_484[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_484_T_3 = state_vec_0_set_left_older ? state_vec_484_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_484_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_484_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_484_T_8 = {state_vec_0_set_left_older,_state_vec_484_T_3,_state_vec_484_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_485_valid = touch_way_0_valid & touch_set_0 == 9'h1e5; // @[Replacement.scala 315:30]
  wire  state_vec_485_left_subtree_state = state_vec_485[1]; // @[package.scala 154:13]
  wire  state_vec_485_right_subtree_state = state_vec_485[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_485_T_3 = state_vec_0_set_left_older ? state_vec_485_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_485_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_485_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_485_T_8 = {state_vec_0_set_left_older,_state_vec_485_T_3,_state_vec_485_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_486_valid = touch_way_0_valid & touch_set_0 == 9'h1e6; // @[Replacement.scala 315:30]
  wire  state_vec_486_left_subtree_state = state_vec_486[1]; // @[package.scala 154:13]
  wire  state_vec_486_right_subtree_state = state_vec_486[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_486_T_3 = state_vec_0_set_left_older ? state_vec_486_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_486_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_486_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_486_T_8 = {state_vec_0_set_left_older,_state_vec_486_T_3,_state_vec_486_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_487_valid = touch_way_0_valid & touch_set_0 == 9'h1e7; // @[Replacement.scala 315:30]
  wire  state_vec_487_left_subtree_state = state_vec_487[1]; // @[package.scala 154:13]
  wire  state_vec_487_right_subtree_state = state_vec_487[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_487_T_3 = state_vec_0_set_left_older ? state_vec_487_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_487_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_487_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_487_T_8 = {state_vec_0_set_left_older,_state_vec_487_T_3,_state_vec_487_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_488_valid = touch_way_0_valid & touch_set_0 == 9'h1e8; // @[Replacement.scala 315:30]
  wire  state_vec_488_left_subtree_state = state_vec_488[1]; // @[package.scala 154:13]
  wire  state_vec_488_right_subtree_state = state_vec_488[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_488_T_3 = state_vec_0_set_left_older ? state_vec_488_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_488_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_488_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_488_T_8 = {state_vec_0_set_left_older,_state_vec_488_T_3,_state_vec_488_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_489_valid = touch_way_0_valid & touch_set_0 == 9'h1e9; // @[Replacement.scala 315:30]
  wire  state_vec_489_left_subtree_state = state_vec_489[1]; // @[package.scala 154:13]
  wire  state_vec_489_right_subtree_state = state_vec_489[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_489_T_3 = state_vec_0_set_left_older ? state_vec_489_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_489_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_489_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_489_T_8 = {state_vec_0_set_left_older,_state_vec_489_T_3,_state_vec_489_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_490_valid = touch_way_0_valid & touch_set_0 == 9'h1ea; // @[Replacement.scala 315:30]
  wire  state_vec_490_left_subtree_state = state_vec_490[1]; // @[package.scala 154:13]
  wire  state_vec_490_right_subtree_state = state_vec_490[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_490_T_3 = state_vec_0_set_left_older ? state_vec_490_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_490_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_490_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_490_T_8 = {state_vec_0_set_left_older,_state_vec_490_T_3,_state_vec_490_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_491_valid = touch_way_0_valid & touch_set_0 == 9'h1eb; // @[Replacement.scala 315:30]
  wire  state_vec_491_left_subtree_state = state_vec_491[1]; // @[package.scala 154:13]
  wire  state_vec_491_right_subtree_state = state_vec_491[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_491_T_3 = state_vec_0_set_left_older ? state_vec_491_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_491_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_491_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_491_T_8 = {state_vec_0_set_left_older,_state_vec_491_T_3,_state_vec_491_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_492_valid = touch_way_0_valid & touch_set_0 == 9'h1ec; // @[Replacement.scala 315:30]
  wire  state_vec_492_left_subtree_state = state_vec_492[1]; // @[package.scala 154:13]
  wire  state_vec_492_right_subtree_state = state_vec_492[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_492_T_3 = state_vec_0_set_left_older ? state_vec_492_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_492_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_492_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_492_T_8 = {state_vec_0_set_left_older,_state_vec_492_T_3,_state_vec_492_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_493_valid = touch_way_0_valid & touch_set_0 == 9'h1ed; // @[Replacement.scala 315:30]
  wire  state_vec_493_left_subtree_state = state_vec_493[1]; // @[package.scala 154:13]
  wire  state_vec_493_right_subtree_state = state_vec_493[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_493_T_3 = state_vec_0_set_left_older ? state_vec_493_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_493_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_493_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_493_T_8 = {state_vec_0_set_left_older,_state_vec_493_T_3,_state_vec_493_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_494_valid = touch_way_0_valid & touch_set_0 == 9'h1ee; // @[Replacement.scala 315:30]
  wire  state_vec_494_left_subtree_state = state_vec_494[1]; // @[package.scala 154:13]
  wire  state_vec_494_right_subtree_state = state_vec_494[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_494_T_3 = state_vec_0_set_left_older ? state_vec_494_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_494_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_494_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_494_T_8 = {state_vec_0_set_left_older,_state_vec_494_T_3,_state_vec_494_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_495_valid = touch_way_0_valid & touch_set_0 == 9'h1ef; // @[Replacement.scala 315:30]
  wire  state_vec_495_left_subtree_state = state_vec_495[1]; // @[package.scala 154:13]
  wire  state_vec_495_right_subtree_state = state_vec_495[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_495_T_3 = state_vec_0_set_left_older ? state_vec_495_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_495_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_495_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_495_T_8 = {state_vec_0_set_left_older,_state_vec_495_T_3,_state_vec_495_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_496_valid = touch_way_0_valid & touch_set_0 == 9'h1f0; // @[Replacement.scala 315:30]
  wire  state_vec_496_left_subtree_state = state_vec_496[1]; // @[package.scala 154:13]
  wire  state_vec_496_right_subtree_state = state_vec_496[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_496_T_3 = state_vec_0_set_left_older ? state_vec_496_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_496_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_496_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_496_T_8 = {state_vec_0_set_left_older,_state_vec_496_T_3,_state_vec_496_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_497_valid = touch_way_0_valid & touch_set_0 == 9'h1f1; // @[Replacement.scala 315:30]
  wire  state_vec_497_left_subtree_state = state_vec_497[1]; // @[package.scala 154:13]
  wire  state_vec_497_right_subtree_state = state_vec_497[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_497_T_3 = state_vec_0_set_left_older ? state_vec_497_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_497_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_497_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_497_T_8 = {state_vec_0_set_left_older,_state_vec_497_T_3,_state_vec_497_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_498_valid = touch_way_0_valid & touch_set_0 == 9'h1f2; // @[Replacement.scala 315:30]
  wire  state_vec_498_left_subtree_state = state_vec_498[1]; // @[package.scala 154:13]
  wire  state_vec_498_right_subtree_state = state_vec_498[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_498_T_3 = state_vec_0_set_left_older ? state_vec_498_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_498_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_498_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_498_T_8 = {state_vec_0_set_left_older,_state_vec_498_T_3,_state_vec_498_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_499_valid = touch_way_0_valid & touch_set_0 == 9'h1f3; // @[Replacement.scala 315:30]
  wire  state_vec_499_left_subtree_state = state_vec_499[1]; // @[package.scala 154:13]
  wire  state_vec_499_right_subtree_state = state_vec_499[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_499_T_3 = state_vec_0_set_left_older ? state_vec_499_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_499_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_499_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_499_T_8 = {state_vec_0_set_left_older,_state_vec_499_T_3,_state_vec_499_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_500_valid = touch_way_0_valid & touch_set_0 == 9'h1f4; // @[Replacement.scala 315:30]
  wire  state_vec_500_left_subtree_state = state_vec_500[1]; // @[package.scala 154:13]
  wire  state_vec_500_right_subtree_state = state_vec_500[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_500_T_3 = state_vec_0_set_left_older ? state_vec_500_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_500_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_500_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_500_T_8 = {state_vec_0_set_left_older,_state_vec_500_T_3,_state_vec_500_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_501_valid = touch_way_0_valid & touch_set_0 == 9'h1f5; // @[Replacement.scala 315:30]
  wire  state_vec_501_left_subtree_state = state_vec_501[1]; // @[package.scala 154:13]
  wire  state_vec_501_right_subtree_state = state_vec_501[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_501_T_3 = state_vec_0_set_left_older ? state_vec_501_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_501_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_501_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_501_T_8 = {state_vec_0_set_left_older,_state_vec_501_T_3,_state_vec_501_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_502_valid = touch_way_0_valid & touch_set_0 == 9'h1f6; // @[Replacement.scala 315:30]
  wire  state_vec_502_left_subtree_state = state_vec_502[1]; // @[package.scala 154:13]
  wire  state_vec_502_right_subtree_state = state_vec_502[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_502_T_3 = state_vec_0_set_left_older ? state_vec_502_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_502_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_502_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_502_T_8 = {state_vec_0_set_left_older,_state_vec_502_T_3,_state_vec_502_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_503_valid = touch_way_0_valid & touch_set_0 == 9'h1f7; // @[Replacement.scala 315:30]
  wire  state_vec_503_left_subtree_state = state_vec_503[1]; // @[package.scala 154:13]
  wire  state_vec_503_right_subtree_state = state_vec_503[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_503_T_3 = state_vec_0_set_left_older ? state_vec_503_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_503_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_503_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_503_T_8 = {state_vec_0_set_left_older,_state_vec_503_T_3,_state_vec_503_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_504_valid = touch_way_0_valid & touch_set_0 == 9'h1f8; // @[Replacement.scala 315:30]
  wire  state_vec_504_left_subtree_state = state_vec_504[1]; // @[package.scala 154:13]
  wire  state_vec_504_right_subtree_state = state_vec_504[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_504_T_3 = state_vec_0_set_left_older ? state_vec_504_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_504_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_504_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_504_T_8 = {state_vec_0_set_left_older,_state_vec_504_T_3,_state_vec_504_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_505_valid = touch_way_0_valid & touch_set_0 == 9'h1f9; // @[Replacement.scala 315:30]
  wire  state_vec_505_left_subtree_state = state_vec_505[1]; // @[package.scala 154:13]
  wire  state_vec_505_right_subtree_state = state_vec_505[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_505_T_3 = state_vec_0_set_left_older ? state_vec_505_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_505_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_505_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_505_T_8 = {state_vec_0_set_left_older,_state_vec_505_T_3,_state_vec_505_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_506_valid = touch_way_0_valid & touch_set_0 == 9'h1fa; // @[Replacement.scala 315:30]
  wire  state_vec_506_left_subtree_state = state_vec_506[1]; // @[package.scala 154:13]
  wire  state_vec_506_right_subtree_state = state_vec_506[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_506_T_3 = state_vec_0_set_left_older ? state_vec_506_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_506_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_506_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_506_T_8 = {state_vec_0_set_left_older,_state_vec_506_T_3,_state_vec_506_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_507_valid = touch_way_0_valid & touch_set_0 == 9'h1fb; // @[Replacement.scala 315:30]
  wire  state_vec_507_left_subtree_state = state_vec_507[1]; // @[package.scala 154:13]
  wire  state_vec_507_right_subtree_state = state_vec_507[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_507_T_3 = state_vec_0_set_left_older ? state_vec_507_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_507_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_507_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_507_T_8 = {state_vec_0_set_left_older,_state_vec_507_T_3,_state_vec_507_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_508_valid = touch_way_0_valid & touch_set_0 == 9'h1fc; // @[Replacement.scala 315:30]
  wire  state_vec_508_left_subtree_state = state_vec_508[1]; // @[package.scala 154:13]
  wire  state_vec_508_right_subtree_state = state_vec_508[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_508_T_3 = state_vec_0_set_left_older ? state_vec_508_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_508_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_508_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_508_T_8 = {state_vec_0_set_left_older,_state_vec_508_T_3,_state_vec_508_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_509_valid = touch_way_0_valid & touch_set_0 == 9'h1fd; // @[Replacement.scala 315:30]
  wire  state_vec_509_left_subtree_state = state_vec_509[1]; // @[package.scala 154:13]
  wire  state_vec_509_right_subtree_state = state_vec_509[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_509_T_3 = state_vec_0_set_left_older ? state_vec_509_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_509_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_509_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_509_T_8 = {state_vec_0_set_left_older,_state_vec_509_T_3,_state_vec_509_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_510_valid = touch_way_0_valid & touch_set_0 == 9'h1fe; // @[Replacement.scala 315:30]
  wire  state_vec_510_left_subtree_state = state_vec_510[1]; // @[package.scala 154:13]
  wire  state_vec_510_right_subtree_state = state_vec_510[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_510_T_3 = state_vec_0_set_left_older ? state_vec_510_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_510_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_510_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_510_T_8 = {state_vec_0_set_left_older,_state_vec_510_T_3,_state_vec_510_T_7}; // @[Cat.scala 31:58]
  wire  set_touch_ways_0_511_valid = touch_way_0_valid & touch_set_0 == 9'h1ff; // @[Replacement.scala 315:30]
  wire  state_vec_511_left_subtree_state = state_vec_511[1]; // @[package.scala 154:13]
  wire  state_vec_511_right_subtree_state = state_vec_511[0]; // @[Replacement.scala 198:38]
  wire  _state_vec_511_T_3 = state_vec_0_set_left_older ? state_vec_511_left_subtree_state : _state_vec_0_T_2; // @[Replacement.scala 203:16]
  wire  _state_vec_511_T_7 = state_vec_0_set_left_older ? _state_vec_0_T_2 : state_vec_511_right_subtree_state; // @[Replacement.scala 206:16]
  wire [2:0] _state_vec_511_T_8 = {state_vec_0_set_left_older,_state_vec_511_T_3,_state_vec_511_T_7}; // @[Cat.scala 31:58]
  wire [2:0] _io_read_resp_T_49 = total_hits_0 ? _GEN_11 : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_resp_T_50 = total_hits_1 ? _GEN_31 : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_resp_T_51 = total_hits_2 ? _GEN_51 : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_resp_T_52 = total_hits_3 ? _GEN_71 : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_resp_T_53 = _io_read_resp_T_49 | _io_read_resp_T_50; // @[Mux.scala 27:73]
  wire [2:0] _io_read_resp_T_54 = _io_read_resp_T_53 | _io_read_resp_T_51; // @[Mux.scala 27:73]
  wire [1:0] _io_read_resp_T_70 = total_hits_0 ? _GEN_8 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_resp_T_71 = total_hits_1 ? _GEN_28 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_resp_T_72 = total_hits_2 ? _GEN_48 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_resp_T_73 = total_hits_3 ? _GEN_68 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_resp_T_74 = _io_read_resp_T_70 | _io_read_resp_T_71; // @[Mux.scala 27:73]
  wire [1:0] _io_read_resp_T_75 = _io_read_resp_T_74 | _io_read_resp_T_72; // @[Mux.scala 27:73]
  wire [19:0] _io_read_resp_T_77 = total_hits_0 ? _GEN_7 : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _io_read_resp_T_78 = total_hits_1 ? _GEN_27 : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _io_read_resp_T_79 = total_hits_2 ? _GEN_47 : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _io_read_resp_T_80 = total_hits_3 ? _GEN_67 : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _io_read_resp_T_81 = _io_read_resp_T_77 | _io_read_resp_T_78; // @[Mux.scala 27:73]
  wire [19:0] _io_read_resp_T_82 = _io_read_resp_T_81 | _io_read_resp_T_79; // @[Mux.scala 27:73]
  wire [2:0] _io_read_resp_T_84 = total_hits_0 ? _GEN_6 : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_resp_T_85 = total_hits_1 ? _GEN_26 : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_resp_T_86 = total_hits_2 ? _GEN_46 : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_resp_T_87 = total_hits_3 ? _GEN_66 : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_resp_T_88 = _io_read_resp_T_84 | _io_read_resp_T_85; // @[Mux.scala 27:73]
  wire [2:0] _io_read_resp_T_89 = _io_read_resp_T_88 | _io_read_resp_T_86; // @[Mux.scala 27:73]
  wire [1:0] _io_read_resp_T_105 = total_hits_0 ? _GEN_3 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_resp_T_106 = total_hits_1 ? _GEN_23 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_resp_T_107 = total_hits_2 ? _GEN_43 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_resp_T_108 = total_hits_3 ? _GEN_63 : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_resp_T_109 = _io_read_resp_T_105 | _io_read_resp_T_106; // @[Mux.scala 27:73]
  wire [1:0] _io_read_resp_T_110 = _io_read_resp_T_109 | _io_read_resp_T_107; // @[Mux.scala 27:73]
  wire [11:0] _io_read_resp_T_112 = total_hits_0 ? _GEN_2 : 12'h0; // @[Mux.scala 27:73]
  wire [11:0] _io_read_resp_T_113 = total_hits_1 ? _GEN_22 : 12'h0; // @[Mux.scala 27:73]
  wire [11:0] _io_read_resp_T_114 = total_hits_2 ? _GEN_42 : 12'h0; // @[Mux.scala 27:73]
  wire [11:0] _io_read_resp_T_115 = total_hits_3 ? _GEN_62 : 12'h0; // @[Mux.scala 27:73]
  wire [11:0] _io_read_resp_T_116 = _io_read_resp_T_112 | _io_read_resp_T_113; // @[Mux.scala 27:73]
  wire [11:0] _io_read_resp_T_117 = _io_read_resp_T_116 | _io_read_resp_T_114; // @[Mux.scala 27:73]
  wire [2:0] _io_read_resp_T_119 = total_hits_0 ? _GEN_1 : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_resp_T_120 = total_hits_1 ? _GEN_21 : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_resp_T_121 = total_hits_2 ? _GEN_41 : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_resp_T_122 = total_hits_3 ? _GEN_61 : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_resp_T_123 = _io_read_resp_T_119 | _io_read_resp_T_120; // @[Mux.scala 27:73]
  wire [2:0] _io_read_resp_T_124 = _io_read_resp_T_123 | _io_read_resp_T_121; // @[Mux.scala 27:73]
  SRAMTemplate_12 ftb ( // @[FTB.scala 302:21]
    .clock(ftb_clock),
    .reset(ftb_reset),
    .io_rreq_ready(ftb_io_rreq_ready),
    .io_rreq_valid(ftb_io_rreq_valid),
    .io_rreq_bits_setIdx(ftb_io_rreq_bits_setIdx),
    .io_rresp_data_0_entry_valid(ftb_io_rresp_data_0_entry_valid),
    .io_rresp_data_0_entry_brSlots_0_offset(ftb_io_rresp_data_0_entry_brSlots_0_offset),
    .io_rresp_data_0_entry_brSlots_0_lower(ftb_io_rresp_data_0_entry_brSlots_0_lower),
    .io_rresp_data_0_entry_brSlots_0_tarStat(ftb_io_rresp_data_0_entry_brSlots_0_tarStat),
    .io_rresp_data_0_entry_brSlots_0_sharing(ftb_io_rresp_data_0_entry_brSlots_0_sharing),
    .io_rresp_data_0_entry_brSlots_0_valid(ftb_io_rresp_data_0_entry_brSlots_0_valid),
    .io_rresp_data_0_entry_tailSlot_offset(ftb_io_rresp_data_0_entry_tailSlot_offset),
    .io_rresp_data_0_entry_tailSlot_lower(ftb_io_rresp_data_0_entry_tailSlot_lower),
    .io_rresp_data_0_entry_tailSlot_tarStat(ftb_io_rresp_data_0_entry_tailSlot_tarStat),
    .io_rresp_data_0_entry_tailSlot_sharing(ftb_io_rresp_data_0_entry_tailSlot_sharing),
    .io_rresp_data_0_entry_tailSlot_valid(ftb_io_rresp_data_0_entry_tailSlot_valid),
    .io_rresp_data_0_entry_pftAddr(ftb_io_rresp_data_0_entry_pftAddr),
    .io_rresp_data_0_entry_carry(ftb_io_rresp_data_0_entry_carry),
    .io_rresp_data_0_entry_isCall(ftb_io_rresp_data_0_entry_isCall),
    .io_rresp_data_0_entry_isRet(ftb_io_rresp_data_0_entry_isRet),
    .io_rresp_data_0_entry_isJalr(ftb_io_rresp_data_0_entry_isJalr),
    .io_rresp_data_0_entry_last_may_be_rvi_call(ftb_io_rresp_data_0_entry_last_may_be_rvi_call),
    .io_rresp_data_0_entry_always_taken_0(ftb_io_rresp_data_0_entry_always_taken_0),
    .io_rresp_data_0_entry_always_taken_1(ftb_io_rresp_data_0_entry_always_taken_1),
    .io_rresp_data_0_tag(ftb_io_rresp_data_0_tag),
    .io_rresp_data_1_entry_valid(ftb_io_rresp_data_1_entry_valid),
    .io_rresp_data_1_entry_brSlots_0_offset(ftb_io_rresp_data_1_entry_brSlots_0_offset),
    .io_rresp_data_1_entry_brSlots_0_lower(ftb_io_rresp_data_1_entry_brSlots_0_lower),
    .io_rresp_data_1_entry_brSlots_0_tarStat(ftb_io_rresp_data_1_entry_brSlots_0_tarStat),
    .io_rresp_data_1_entry_brSlots_0_sharing(ftb_io_rresp_data_1_entry_brSlots_0_sharing),
    .io_rresp_data_1_entry_brSlots_0_valid(ftb_io_rresp_data_1_entry_brSlots_0_valid),
    .io_rresp_data_1_entry_tailSlot_offset(ftb_io_rresp_data_1_entry_tailSlot_offset),
    .io_rresp_data_1_entry_tailSlot_lower(ftb_io_rresp_data_1_entry_tailSlot_lower),
    .io_rresp_data_1_entry_tailSlot_tarStat(ftb_io_rresp_data_1_entry_tailSlot_tarStat),
    .io_rresp_data_1_entry_tailSlot_sharing(ftb_io_rresp_data_1_entry_tailSlot_sharing),
    .io_rresp_data_1_entry_tailSlot_valid(ftb_io_rresp_data_1_entry_tailSlot_valid),
    .io_rresp_data_1_entry_pftAddr(ftb_io_rresp_data_1_entry_pftAddr),
    .io_rresp_data_1_entry_carry(ftb_io_rresp_data_1_entry_carry),
    .io_rresp_data_1_entry_isCall(ftb_io_rresp_data_1_entry_isCall),
    .io_rresp_data_1_entry_isRet(ftb_io_rresp_data_1_entry_isRet),
    .io_rresp_data_1_entry_isJalr(ftb_io_rresp_data_1_entry_isJalr),
    .io_rresp_data_1_entry_last_may_be_rvi_call(ftb_io_rresp_data_1_entry_last_may_be_rvi_call),
    .io_rresp_data_1_entry_always_taken_0(ftb_io_rresp_data_1_entry_always_taken_0),
    .io_rresp_data_1_entry_always_taken_1(ftb_io_rresp_data_1_entry_always_taken_1),
    .io_rresp_data_1_tag(ftb_io_rresp_data_1_tag),
    .io_rresp_data_2_entry_valid(ftb_io_rresp_data_2_entry_valid),
    .io_rresp_data_2_entry_brSlots_0_offset(ftb_io_rresp_data_2_entry_brSlots_0_offset),
    .io_rresp_data_2_entry_brSlots_0_lower(ftb_io_rresp_data_2_entry_brSlots_0_lower),
    .io_rresp_data_2_entry_brSlots_0_tarStat(ftb_io_rresp_data_2_entry_brSlots_0_tarStat),
    .io_rresp_data_2_entry_brSlots_0_sharing(ftb_io_rresp_data_2_entry_brSlots_0_sharing),
    .io_rresp_data_2_entry_brSlots_0_valid(ftb_io_rresp_data_2_entry_brSlots_0_valid),
    .io_rresp_data_2_entry_tailSlot_offset(ftb_io_rresp_data_2_entry_tailSlot_offset),
    .io_rresp_data_2_entry_tailSlot_lower(ftb_io_rresp_data_2_entry_tailSlot_lower),
    .io_rresp_data_2_entry_tailSlot_tarStat(ftb_io_rresp_data_2_entry_tailSlot_tarStat),
    .io_rresp_data_2_entry_tailSlot_sharing(ftb_io_rresp_data_2_entry_tailSlot_sharing),
    .io_rresp_data_2_entry_tailSlot_valid(ftb_io_rresp_data_2_entry_tailSlot_valid),
    .io_rresp_data_2_entry_pftAddr(ftb_io_rresp_data_2_entry_pftAddr),
    .io_rresp_data_2_entry_carry(ftb_io_rresp_data_2_entry_carry),
    .io_rresp_data_2_entry_isCall(ftb_io_rresp_data_2_entry_isCall),
    .io_rresp_data_2_entry_isRet(ftb_io_rresp_data_2_entry_isRet),
    .io_rresp_data_2_entry_isJalr(ftb_io_rresp_data_2_entry_isJalr),
    .io_rresp_data_2_entry_last_may_be_rvi_call(ftb_io_rresp_data_2_entry_last_may_be_rvi_call),
    .io_rresp_data_2_entry_always_taken_0(ftb_io_rresp_data_2_entry_always_taken_0),
    .io_rresp_data_2_entry_always_taken_1(ftb_io_rresp_data_2_entry_always_taken_1),
    .io_rresp_data_2_tag(ftb_io_rresp_data_2_tag),
    .io_rresp_data_3_entry_valid(ftb_io_rresp_data_3_entry_valid),
    .io_rresp_data_3_entry_brSlots_0_offset(ftb_io_rresp_data_3_entry_brSlots_0_offset),
    .io_rresp_data_3_entry_brSlots_0_lower(ftb_io_rresp_data_3_entry_brSlots_0_lower),
    .io_rresp_data_3_entry_brSlots_0_tarStat(ftb_io_rresp_data_3_entry_brSlots_0_tarStat),
    .io_rresp_data_3_entry_brSlots_0_sharing(ftb_io_rresp_data_3_entry_brSlots_0_sharing),
    .io_rresp_data_3_entry_brSlots_0_valid(ftb_io_rresp_data_3_entry_brSlots_0_valid),
    .io_rresp_data_3_entry_tailSlot_offset(ftb_io_rresp_data_3_entry_tailSlot_offset),
    .io_rresp_data_3_entry_tailSlot_lower(ftb_io_rresp_data_3_entry_tailSlot_lower),
    .io_rresp_data_3_entry_tailSlot_tarStat(ftb_io_rresp_data_3_entry_tailSlot_tarStat),
    .io_rresp_data_3_entry_tailSlot_sharing(ftb_io_rresp_data_3_entry_tailSlot_sharing),
    .io_rresp_data_3_entry_tailSlot_valid(ftb_io_rresp_data_3_entry_tailSlot_valid),
    .io_rresp_data_3_entry_pftAddr(ftb_io_rresp_data_3_entry_pftAddr),
    .io_rresp_data_3_entry_carry(ftb_io_rresp_data_3_entry_carry),
    .io_rresp_data_3_entry_isCall(ftb_io_rresp_data_3_entry_isCall),
    .io_rresp_data_3_entry_isRet(ftb_io_rresp_data_3_entry_isRet),
    .io_rresp_data_3_entry_isJalr(ftb_io_rresp_data_3_entry_isJalr),
    .io_rresp_data_3_entry_last_may_be_rvi_call(ftb_io_rresp_data_3_entry_last_may_be_rvi_call),
    .io_rresp_data_3_entry_always_taken_0(ftb_io_rresp_data_3_entry_always_taken_0),
    .io_rresp_data_3_entry_always_taken_1(ftb_io_rresp_data_3_entry_always_taken_1),
    .io_rresp_data_3_tag(ftb_io_rresp_data_3_tag),
    .io_wreq_valid(ftb_io_wreq_valid),
    .io_wreq_bits_setIdx(ftb_io_wreq_bits_setIdx),
    .io_wreq_bits_data_0_entry_valid(ftb_io_wreq_bits_data_0_entry_valid),
    .io_wreq_bits_data_0_entry_brSlots_0_offset(ftb_io_wreq_bits_data_0_entry_brSlots_0_offset),
    .io_wreq_bits_data_0_entry_brSlots_0_lower(ftb_io_wreq_bits_data_0_entry_brSlots_0_lower),
    .io_wreq_bits_data_0_entry_brSlots_0_tarStat(ftb_io_wreq_bits_data_0_entry_brSlots_0_tarStat),
    .io_wreq_bits_data_0_entry_brSlots_0_sharing(ftb_io_wreq_bits_data_0_entry_brSlots_0_sharing),
    .io_wreq_bits_data_0_entry_brSlots_0_valid(ftb_io_wreq_bits_data_0_entry_brSlots_0_valid),
    .io_wreq_bits_data_0_entry_tailSlot_offset(ftb_io_wreq_bits_data_0_entry_tailSlot_offset),
    .io_wreq_bits_data_0_entry_tailSlot_lower(ftb_io_wreq_bits_data_0_entry_tailSlot_lower),
    .io_wreq_bits_data_0_entry_tailSlot_tarStat(ftb_io_wreq_bits_data_0_entry_tailSlot_tarStat),
    .io_wreq_bits_data_0_entry_tailSlot_sharing(ftb_io_wreq_bits_data_0_entry_tailSlot_sharing),
    .io_wreq_bits_data_0_entry_tailSlot_valid(ftb_io_wreq_bits_data_0_entry_tailSlot_valid),
    .io_wreq_bits_data_0_entry_pftAddr(ftb_io_wreq_bits_data_0_entry_pftAddr),
    .io_wreq_bits_data_0_entry_carry(ftb_io_wreq_bits_data_0_entry_carry),
    .io_wreq_bits_data_0_entry_isCall(ftb_io_wreq_bits_data_0_entry_isCall),
    .io_wreq_bits_data_0_entry_isRet(ftb_io_wreq_bits_data_0_entry_isRet),
    .io_wreq_bits_data_0_entry_isJalr(ftb_io_wreq_bits_data_0_entry_isJalr),
    .io_wreq_bits_data_0_entry_last_may_be_rvi_call(ftb_io_wreq_bits_data_0_entry_last_may_be_rvi_call),
    .io_wreq_bits_data_0_entry_always_taken_0(ftb_io_wreq_bits_data_0_entry_always_taken_0),
    .io_wreq_bits_data_0_entry_always_taken_1(ftb_io_wreq_bits_data_0_entry_always_taken_1),
    .io_wreq_bits_data_0_tag(ftb_io_wreq_bits_data_0_tag),
    .io_wreq_bits_data_1_entry_valid(ftb_io_wreq_bits_data_1_entry_valid),
    .io_wreq_bits_data_1_entry_brSlots_0_offset(ftb_io_wreq_bits_data_1_entry_brSlots_0_offset),
    .io_wreq_bits_data_1_entry_brSlots_0_lower(ftb_io_wreq_bits_data_1_entry_brSlots_0_lower),
    .io_wreq_bits_data_1_entry_brSlots_0_tarStat(ftb_io_wreq_bits_data_1_entry_brSlots_0_tarStat),
    .io_wreq_bits_data_1_entry_brSlots_0_sharing(ftb_io_wreq_bits_data_1_entry_brSlots_0_sharing),
    .io_wreq_bits_data_1_entry_brSlots_0_valid(ftb_io_wreq_bits_data_1_entry_brSlots_0_valid),
    .io_wreq_bits_data_1_entry_tailSlot_offset(ftb_io_wreq_bits_data_1_entry_tailSlot_offset),
    .io_wreq_bits_data_1_entry_tailSlot_lower(ftb_io_wreq_bits_data_1_entry_tailSlot_lower),
    .io_wreq_bits_data_1_entry_tailSlot_tarStat(ftb_io_wreq_bits_data_1_entry_tailSlot_tarStat),
    .io_wreq_bits_data_1_entry_tailSlot_sharing(ftb_io_wreq_bits_data_1_entry_tailSlot_sharing),
    .io_wreq_bits_data_1_entry_tailSlot_valid(ftb_io_wreq_bits_data_1_entry_tailSlot_valid),
    .io_wreq_bits_data_1_entry_pftAddr(ftb_io_wreq_bits_data_1_entry_pftAddr),
    .io_wreq_bits_data_1_entry_carry(ftb_io_wreq_bits_data_1_entry_carry),
    .io_wreq_bits_data_1_entry_isCall(ftb_io_wreq_bits_data_1_entry_isCall),
    .io_wreq_bits_data_1_entry_isRet(ftb_io_wreq_bits_data_1_entry_isRet),
    .io_wreq_bits_data_1_entry_isJalr(ftb_io_wreq_bits_data_1_entry_isJalr),
    .io_wreq_bits_data_1_entry_last_may_be_rvi_call(ftb_io_wreq_bits_data_1_entry_last_may_be_rvi_call),
    .io_wreq_bits_data_1_entry_always_taken_0(ftb_io_wreq_bits_data_1_entry_always_taken_0),
    .io_wreq_bits_data_1_entry_always_taken_1(ftb_io_wreq_bits_data_1_entry_always_taken_1),
    .io_wreq_bits_data_1_tag(ftb_io_wreq_bits_data_1_tag),
    .io_wreq_bits_data_2_entry_valid(ftb_io_wreq_bits_data_2_entry_valid),
    .io_wreq_bits_data_2_entry_brSlots_0_offset(ftb_io_wreq_bits_data_2_entry_brSlots_0_offset),
    .io_wreq_bits_data_2_entry_brSlots_0_lower(ftb_io_wreq_bits_data_2_entry_brSlots_0_lower),
    .io_wreq_bits_data_2_entry_brSlots_0_tarStat(ftb_io_wreq_bits_data_2_entry_brSlots_0_tarStat),
    .io_wreq_bits_data_2_entry_brSlots_0_sharing(ftb_io_wreq_bits_data_2_entry_brSlots_0_sharing),
    .io_wreq_bits_data_2_entry_brSlots_0_valid(ftb_io_wreq_bits_data_2_entry_brSlots_0_valid),
    .io_wreq_bits_data_2_entry_tailSlot_offset(ftb_io_wreq_bits_data_2_entry_tailSlot_offset),
    .io_wreq_bits_data_2_entry_tailSlot_lower(ftb_io_wreq_bits_data_2_entry_tailSlot_lower),
    .io_wreq_bits_data_2_entry_tailSlot_tarStat(ftb_io_wreq_bits_data_2_entry_tailSlot_tarStat),
    .io_wreq_bits_data_2_entry_tailSlot_sharing(ftb_io_wreq_bits_data_2_entry_tailSlot_sharing),
    .io_wreq_bits_data_2_entry_tailSlot_valid(ftb_io_wreq_bits_data_2_entry_tailSlot_valid),
    .io_wreq_bits_data_2_entry_pftAddr(ftb_io_wreq_bits_data_2_entry_pftAddr),
    .io_wreq_bits_data_2_entry_carry(ftb_io_wreq_bits_data_2_entry_carry),
    .io_wreq_bits_data_2_entry_isCall(ftb_io_wreq_bits_data_2_entry_isCall),
    .io_wreq_bits_data_2_entry_isRet(ftb_io_wreq_bits_data_2_entry_isRet),
    .io_wreq_bits_data_2_entry_isJalr(ftb_io_wreq_bits_data_2_entry_isJalr),
    .io_wreq_bits_data_2_entry_last_may_be_rvi_call(ftb_io_wreq_bits_data_2_entry_last_may_be_rvi_call),
    .io_wreq_bits_data_2_entry_always_taken_0(ftb_io_wreq_bits_data_2_entry_always_taken_0),
    .io_wreq_bits_data_2_entry_always_taken_1(ftb_io_wreq_bits_data_2_entry_always_taken_1),
    .io_wreq_bits_data_2_tag(ftb_io_wreq_bits_data_2_tag),
    .io_wreq_bits_data_3_entry_valid(ftb_io_wreq_bits_data_3_entry_valid),
    .io_wreq_bits_data_3_entry_brSlots_0_offset(ftb_io_wreq_bits_data_3_entry_brSlots_0_offset),
    .io_wreq_bits_data_3_entry_brSlots_0_lower(ftb_io_wreq_bits_data_3_entry_brSlots_0_lower),
    .io_wreq_bits_data_3_entry_brSlots_0_tarStat(ftb_io_wreq_bits_data_3_entry_brSlots_0_tarStat),
    .io_wreq_bits_data_3_entry_brSlots_0_sharing(ftb_io_wreq_bits_data_3_entry_brSlots_0_sharing),
    .io_wreq_bits_data_3_entry_brSlots_0_valid(ftb_io_wreq_bits_data_3_entry_brSlots_0_valid),
    .io_wreq_bits_data_3_entry_tailSlot_offset(ftb_io_wreq_bits_data_3_entry_tailSlot_offset),
    .io_wreq_bits_data_3_entry_tailSlot_lower(ftb_io_wreq_bits_data_3_entry_tailSlot_lower),
    .io_wreq_bits_data_3_entry_tailSlot_tarStat(ftb_io_wreq_bits_data_3_entry_tailSlot_tarStat),
    .io_wreq_bits_data_3_entry_tailSlot_sharing(ftb_io_wreq_bits_data_3_entry_tailSlot_sharing),
    .io_wreq_bits_data_3_entry_tailSlot_valid(ftb_io_wreq_bits_data_3_entry_tailSlot_valid),
    .io_wreq_bits_data_3_entry_pftAddr(ftb_io_wreq_bits_data_3_entry_pftAddr),
    .io_wreq_bits_data_3_entry_carry(ftb_io_wreq_bits_data_3_entry_carry),
    .io_wreq_bits_data_3_entry_isCall(ftb_io_wreq_bits_data_3_entry_isCall),
    .io_wreq_bits_data_3_entry_isRet(ftb_io_wreq_bits_data_3_entry_isRet),
    .io_wreq_bits_data_3_entry_isJalr(ftb_io_wreq_bits_data_3_entry_isJalr),
    .io_wreq_bits_data_3_entry_last_may_be_rvi_call(ftb_io_wreq_bits_data_3_entry_last_may_be_rvi_call),
    .io_wreq_bits_data_3_entry_always_taken_0(ftb_io_wreq_bits_data_3_entry_always_taken_0),
    .io_wreq_bits_data_3_entry_always_taken_1(ftb_io_wreq_bits_data_3_entry_always_taken_1),
    .io_wreq_bits_data_3_tag(ftb_io_wreq_bits_data_3_tag),
    .io_wreq_bits_waymask(ftb_io_wreq_bits_waymask)
  );
  assign io_req_pc_ready = ftb_io_rreq_ready; // @[FTB.scala 311:21]
  assign io_read_resp_valid = total_hits_0 & _GEN_0 | total_hits_1 & _GEN_20 | total_hits_2 & _GEN_40 | total_hits_3 &
    _GEN_60; // @[Mux.scala 27:73]
  assign io_read_resp_brSlots_0_offset = _io_read_resp_T_124 | _io_read_resp_T_122; // @[Mux.scala 27:73]
  assign io_read_resp_brSlots_0_lower = _io_read_resp_T_117 | _io_read_resp_T_115; // @[Mux.scala 27:73]
  assign io_read_resp_brSlots_0_tarStat = _io_read_resp_T_110 | _io_read_resp_T_108; // @[Mux.scala 27:73]
  assign io_read_resp_brSlots_0_sharing = total_hits_0 & _GEN_4 | total_hits_1 & _GEN_24 | total_hits_2 & _GEN_44 |
    total_hits_3 & _GEN_64; // @[Mux.scala 27:73]
  assign io_read_resp_brSlots_0_valid = total_hits_0 & _GEN_5 | total_hits_1 & _GEN_25 | total_hits_2 & _GEN_45 |
    total_hits_3 & _GEN_65; // @[Mux.scala 27:73]
  assign io_read_resp_tailSlot_offset = _io_read_resp_T_89 | _io_read_resp_T_87; // @[Mux.scala 27:73]
  assign io_read_resp_tailSlot_lower = _io_read_resp_T_82 | _io_read_resp_T_80; // @[Mux.scala 27:73]
  assign io_read_resp_tailSlot_tarStat = _io_read_resp_T_75 | _io_read_resp_T_73; // @[Mux.scala 27:73]
  assign io_read_resp_tailSlot_sharing = total_hits_0 & _GEN_9 | total_hits_1 & _GEN_29 | total_hits_2 & _GEN_49 |
    total_hits_3 & _GEN_69; // @[Mux.scala 27:73]
  assign io_read_resp_tailSlot_valid = total_hits_0 & _GEN_10 | total_hits_1 & _GEN_30 | total_hits_2 & _GEN_50 |
    total_hits_3 & _GEN_70; // @[Mux.scala 27:73]
  assign io_read_resp_pftAddr = _io_read_resp_T_54 | _io_read_resp_T_52; // @[Mux.scala 27:73]
  assign io_read_resp_carry = total_hits_0 & _GEN_12 | total_hits_1 & _GEN_32 | total_hits_2 & _GEN_52 | total_hits_3 &
    _GEN_72; // @[Mux.scala 27:73]
  assign io_read_resp_isCall = total_hits_0 & _GEN_13 | total_hits_1 & _GEN_33 | total_hits_2 & _GEN_53 | total_hits_3
     & _GEN_73; // @[Mux.scala 27:73]
  assign io_read_resp_isRet = total_hits_0 & _GEN_14 | total_hits_1 & _GEN_34 | total_hits_2 & _GEN_54 | total_hits_3 &
    _GEN_74; // @[Mux.scala 27:73]
  assign io_read_resp_isJalr = total_hits_0 & _GEN_15 | total_hits_1 & _GEN_35 | total_hits_2 & _GEN_55 | total_hits_3
     & _GEN_75; // @[Mux.scala 27:73]
  assign io_read_resp_last_may_be_rvi_call = total_hits_0 & _GEN_16 | total_hits_1 & _GEN_36 | total_hits_2 & _GEN_56 |
    total_hits_3 & _GEN_76; // @[Mux.scala 27:73]
  assign io_read_resp_always_taken_0 = total_hits_0 & _GEN_17 | total_hits_1 & _GEN_37 | total_hits_2 & _GEN_57 |
    total_hits_3 & _GEN_77; // @[Mux.scala 27:73]
  assign io_read_resp_always_taken_1 = total_hits_0 & _GEN_18 | total_hits_1 & _GEN_38 | total_hits_2 & _GEN_58 |
    total_hits_3 & _GEN_78; // @[Mux.scala 27:73]
  assign io_read_hits_valid = total_hits_0 | total_hits_1 | total_hits_2 | total_hits_3; // @[FTB.scala 323:34]
  assign io_read_hits_bits = {_hit_way_T_1,_hit_way_T_2[1]}; // @[Cat.scala 31:58]
  assign io_update_hits_valid = u_total_hits_0 | u_total_hits_1 | u_total_hits_2 | u_total_hits_3; // @[FTB.scala 329:38]
  assign io_update_hits_bits = {_u_hit_way_T_1,_u_hit_way_T_2[1]}; // @[Cat.scala 31:58]
  assign ftb_clock = clock;
  assign ftb_reset = reset;
  assign ftb_io_rreq_valid = io_req_pc_valid | io_u_req_pc_valid; // @[FTB.scala 306:43]
  assign ftb_io_rreq_bits_setIdx = io_u_req_pc_valid ? io_u_req_pc_bits[9:1] : io_req_pc_bits[9:1]; // @[FTB.scala 307:36]
  assign ftb_io_wreq_valid = io_update_write_data_valid; // @[SRAMTemplate.scala 84:20]
  assign ftb_io_wreq_bits_setIdx = io_update_pc[9:1]; // @[FrontendBundle.scala 389:65]
  assign ftb_io_wreq_bits_data_0_entry_valid = io_update_write_data_bits_entry_valid; // @[SRAMTemplate.scala 88:{25,25}]
  assign ftb_io_wreq_bits_data_0_entry_brSlots_0_offset = io_update_write_data_bits_entry_brSlots_0_offset; // @[SRAMTemplate.scala 88:{25,25}]
  assign ftb_io_wreq_bits_data_0_entry_brSlots_0_lower = io_update_write_data_bits_entry_brSlots_0_lower; // @[SRAMTemplate.scala 88:{25,25}]
  assign ftb_io_wreq_bits_data_0_entry_brSlots_0_tarStat = io_update_write_data_bits_entry_brSlots_0_tarStat; // @[SRAMTemplate.scala 88:{25,25}]
  assign ftb_io_wreq_bits_data_0_entry_brSlots_0_sharing = io_update_write_data_bits_entry_brSlots_0_sharing; // @[SRAMTemplate.scala 88:{25,25}]
  assign ftb_io_wreq_bits_data_0_entry_brSlots_0_valid = io_update_write_data_bits_entry_brSlots_0_valid; // @[SRAMTemplate.scala 88:{25,25}]
  assign ftb_io_wreq_bits_data_0_entry_tailSlot_offset = io_update_write_data_bits_entry_tailSlot_offset; // @[SRAMTemplate.scala 88:{25,25}]
  assign ftb_io_wreq_bits_data_0_entry_tailSlot_lower = io_update_write_data_bits_entry_tailSlot_lower; // @[SRAMTemplate.scala 88:{25,25}]
  assign ftb_io_wreq_bits_data_0_entry_tailSlot_tarStat = io_update_write_data_bits_entry_tailSlot_tarStat; // @[SRAMTemplate.scala 88:{25,25}]
  assign ftb_io_wreq_bits_data_0_entry_tailSlot_sharing = io_update_write_data_bits_entry_tailSlot_sharing; // @[SRAMTemplate.scala 88:{25,25}]
  assign ftb_io_wreq_bits_data_0_entry_tailSlot_valid = io_update_write_data_bits_entry_tailSlot_valid; // @[SRAMTemplate.scala 88:{25,25}]
  assign ftb_io_wreq_bits_data_0_entry_pftAddr = io_update_write_data_bits_entry_pftAddr; // @[SRAMTemplate.scala 88:{25,25}]
  assign ftb_io_wreq_bits_data_0_entry_carry = io_update_write_data_bits_entry_carry; // @[SRAMTemplate.scala 88:{25,25}]
  assign ftb_io_wreq_bits_data_0_entry_isCall = io_update_write_data_bits_entry_isCall; // @[SRAMTemplate.scala 88:{25,25}]
  assign ftb_io_wreq_bits_data_0_entry_isRet = io_update_write_data_bits_entry_isRet; // @[SRAMTemplate.scala 88:{25,25}]
  assign ftb_io_wreq_bits_data_0_entry_isJalr = io_update_write_data_bits_entry_isJalr; // @[SRAMTemplate.scala 88:{25,25}]
  assign ftb_io_wreq_bits_data_0_entry_last_may_be_rvi_call = io_update_write_data_bits_entry_last_may_be_rvi_call; // @[SRAMTemplate.scala 88:{25,25}]
  assign ftb_io_wreq_bits_data_0_entry_always_taken_0 = io_update_write_data_bits_entry_always_taken_0; // @[SRAMTemplate.scala 88:{25,25}]
  assign ftb_io_wreq_bits_data_0_entry_always_taken_1 = io_update_write_data_bits_entry_always_taken_1; // @[SRAMTemplate.scala 88:{25,25}]
  assign ftb_io_wreq_bits_data_0_tag = io_update_write_data_bits_tag; // @[SRAMTemplate.scala 88:{25,25}]
  assign ftb_io_wreq_bits_data_1_entry_valid = io_update_write_data_bits_entry_valid; // @[SRAMTemplate.scala 88:{25,25}]
  assign ftb_io_wreq_bits_data_1_entry_brSlots_0_offset = io_update_write_data_bits_entry_brSlots_0_offset; // @[SRAMTemplate.scala 88:{25,25}]
  assign ftb_io_wreq_bits_data_1_entry_brSlots_0_lower = io_update_write_data_bits_entry_brSlots_0_lower; // @[SRAMTemplate.scala 88:{25,25}]
  assign ftb_io_wreq_bits_data_1_entry_brSlots_0_tarStat = io_update_write_data_bits_entry_brSlots_0_tarStat; // @[SRAMTemplate.scala 88:{25,25}]
  assign ftb_io_wreq_bits_data_1_entry_brSlots_0_sharing = io_update_write_data_bits_entry_brSlots_0_sharing; // @[SRAMTemplate.scala 88:{25,25}]
  assign ftb_io_wreq_bits_data_1_entry_brSlots_0_valid = io_update_write_data_bits_entry_brSlots_0_valid; // @[SRAMTemplate.scala 88:{25,25}]
  assign ftb_io_wreq_bits_data_1_entry_tailSlot_offset = io_update_write_data_bits_entry_tailSlot_offset; // @[SRAMTemplate.scala 88:{25,25}]
  assign ftb_io_wreq_bits_data_1_entry_tailSlot_lower = io_update_write_data_bits_entry_tailSlot_lower; // @[SRAMTemplate.scala 88:{25,25}]
  assign ftb_io_wreq_bits_data_1_entry_tailSlot_tarStat = io_update_write_data_bits_entry_tailSlot_tarStat; // @[SRAMTemplate.scala 88:{25,25}]
  assign ftb_io_wreq_bits_data_1_entry_tailSlot_sharing = io_update_write_data_bits_entry_tailSlot_sharing; // @[SRAMTemplate.scala 88:{25,25}]
  assign ftb_io_wreq_bits_data_1_entry_tailSlot_valid = io_update_write_data_bits_entry_tailSlot_valid; // @[SRAMTemplate.scala 88:{25,25}]
  assign ftb_io_wreq_bits_data_1_entry_pftAddr = io_update_write_data_bits_entry_pftAddr; // @[SRAMTemplate.scala 88:{25,25}]
  assign ftb_io_wreq_bits_data_1_entry_carry = io_update_write_data_bits_entry_carry; // @[SRAMTemplate.scala 88:{25,25}]
  assign ftb_io_wreq_bits_data_1_entry_isCall = io_update_write_data_bits_entry_isCall; // @[SRAMTemplate.scala 88:{25,25}]
  assign ftb_io_wreq_bits_data_1_entry_isRet = io_update_write_data_bits_entry_isRet; // @[SRAMTemplate.scala 88:{25,25}]
  assign ftb_io_wreq_bits_data_1_entry_isJalr = io_update_write_data_bits_entry_isJalr; // @[SRAMTemplate.scala 88:{25,25}]
  assign ftb_io_wreq_bits_data_1_entry_last_may_be_rvi_call = io_update_write_data_bits_entry_last_may_be_rvi_call; // @[SRAMTemplate.scala 88:{25,25}]
  assign ftb_io_wreq_bits_data_1_entry_always_taken_0 = io_update_write_data_bits_entry_always_taken_0; // @[SRAMTemplate.scala 88:{25,25}]
  assign ftb_io_wreq_bits_data_1_entry_always_taken_1 = io_update_write_data_bits_entry_always_taken_1; // @[SRAMTemplate.scala 88:{25,25}]
  assign ftb_io_wreq_bits_data_1_tag = io_update_write_data_bits_tag; // @[SRAMTemplate.scala 88:{25,25}]
  assign ftb_io_wreq_bits_data_2_entry_valid = io_update_write_data_bits_entry_valid; // @[SRAMTemplate.scala 88:{25,25}]
  assign ftb_io_wreq_bits_data_2_entry_brSlots_0_offset = io_update_write_data_bits_entry_brSlots_0_offset; // @[SRAMTemplate.scala 88:{25,25}]
  assign ftb_io_wreq_bits_data_2_entry_brSlots_0_lower = io_update_write_data_bits_entry_brSlots_0_lower; // @[SRAMTemplate.scala 88:{25,25}]
  assign ftb_io_wreq_bits_data_2_entry_brSlots_0_tarStat = io_update_write_data_bits_entry_brSlots_0_tarStat; // @[SRAMTemplate.scala 88:{25,25}]
  assign ftb_io_wreq_bits_data_2_entry_brSlots_0_sharing = io_update_write_data_bits_entry_brSlots_0_sharing; // @[SRAMTemplate.scala 88:{25,25}]
  assign ftb_io_wreq_bits_data_2_entry_brSlots_0_valid = io_update_write_data_bits_entry_brSlots_0_valid; // @[SRAMTemplate.scala 88:{25,25}]
  assign ftb_io_wreq_bits_data_2_entry_tailSlot_offset = io_update_write_data_bits_entry_tailSlot_offset; // @[SRAMTemplate.scala 88:{25,25}]
  assign ftb_io_wreq_bits_data_2_entry_tailSlot_lower = io_update_write_data_bits_entry_tailSlot_lower; // @[SRAMTemplate.scala 88:{25,25}]
  assign ftb_io_wreq_bits_data_2_entry_tailSlot_tarStat = io_update_write_data_bits_entry_tailSlot_tarStat; // @[SRAMTemplate.scala 88:{25,25}]
  assign ftb_io_wreq_bits_data_2_entry_tailSlot_sharing = io_update_write_data_bits_entry_tailSlot_sharing; // @[SRAMTemplate.scala 88:{25,25}]
  assign ftb_io_wreq_bits_data_2_entry_tailSlot_valid = io_update_write_data_bits_entry_tailSlot_valid; // @[SRAMTemplate.scala 88:{25,25}]
  assign ftb_io_wreq_bits_data_2_entry_pftAddr = io_update_write_data_bits_entry_pftAddr; // @[SRAMTemplate.scala 88:{25,25}]
  assign ftb_io_wreq_bits_data_2_entry_carry = io_update_write_data_bits_entry_carry; // @[SRAMTemplate.scala 88:{25,25}]
  assign ftb_io_wreq_bits_data_2_entry_isCall = io_update_write_data_bits_entry_isCall; // @[SRAMTemplate.scala 88:{25,25}]
  assign ftb_io_wreq_bits_data_2_entry_isRet = io_update_write_data_bits_entry_isRet; // @[SRAMTemplate.scala 88:{25,25}]
  assign ftb_io_wreq_bits_data_2_entry_isJalr = io_update_write_data_bits_entry_isJalr; // @[SRAMTemplate.scala 88:{25,25}]
  assign ftb_io_wreq_bits_data_2_entry_last_may_be_rvi_call = io_update_write_data_bits_entry_last_may_be_rvi_call; // @[SRAMTemplate.scala 88:{25,25}]
  assign ftb_io_wreq_bits_data_2_entry_always_taken_0 = io_update_write_data_bits_entry_always_taken_0; // @[SRAMTemplate.scala 88:{25,25}]
  assign ftb_io_wreq_bits_data_2_entry_always_taken_1 = io_update_write_data_bits_entry_always_taken_1; // @[SRAMTemplate.scala 88:{25,25}]
  assign ftb_io_wreq_bits_data_2_tag = io_update_write_data_bits_tag; // @[SRAMTemplate.scala 88:{25,25}]
  assign ftb_io_wreq_bits_data_3_entry_valid = io_update_write_data_bits_entry_valid; // @[SRAMTemplate.scala 88:{25,25}]
  assign ftb_io_wreq_bits_data_3_entry_brSlots_0_offset = io_update_write_data_bits_entry_brSlots_0_offset; // @[SRAMTemplate.scala 88:{25,25}]
  assign ftb_io_wreq_bits_data_3_entry_brSlots_0_lower = io_update_write_data_bits_entry_brSlots_0_lower; // @[SRAMTemplate.scala 88:{25,25}]
  assign ftb_io_wreq_bits_data_3_entry_brSlots_0_tarStat = io_update_write_data_bits_entry_brSlots_0_tarStat; // @[SRAMTemplate.scala 88:{25,25}]
  assign ftb_io_wreq_bits_data_3_entry_brSlots_0_sharing = io_update_write_data_bits_entry_brSlots_0_sharing; // @[SRAMTemplate.scala 88:{25,25}]
  assign ftb_io_wreq_bits_data_3_entry_brSlots_0_valid = io_update_write_data_bits_entry_brSlots_0_valid; // @[SRAMTemplate.scala 88:{25,25}]
  assign ftb_io_wreq_bits_data_3_entry_tailSlot_offset = io_update_write_data_bits_entry_tailSlot_offset; // @[SRAMTemplate.scala 88:{25,25}]
  assign ftb_io_wreq_bits_data_3_entry_tailSlot_lower = io_update_write_data_bits_entry_tailSlot_lower; // @[SRAMTemplate.scala 88:{25,25}]
  assign ftb_io_wreq_bits_data_3_entry_tailSlot_tarStat = io_update_write_data_bits_entry_tailSlot_tarStat; // @[SRAMTemplate.scala 88:{25,25}]
  assign ftb_io_wreq_bits_data_3_entry_tailSlot_sharing = io_update_write_data_bits_entry_tailSlot_sharing; // @[SRAMTemplate.scala 88:{25,25}]
  assign ftb_io_wreq_bits_data_3_entry_tailSlot_valid = io_update_write_data_bits_entry_tailSlot_valid; // @[SRAMTemplate.scala 88:{25,25}]
  assign ftb_io_wreq_bits_data_3_entry_pftAddr = io_update_write_data_bits_entry_pftAddr; // @[SRAMTemplate.scala 88:{25,25}]
  assign ftb_io_wreq_bits_data_3_entry_carry = io_update_write_data_bits_entry_carry; // @[SRAMTemplate.scala 88:{25,25}]
  assign ftb_io_wreq_bits_data_3_entry_isCall = io_update_write_data_bits_entry_isCall; // @[SRAMTemplate.scala 88:{25,25}]
  assign ftb_io_wreq_bits_data_3_entry_isRet = io_update_write_data_bits_entry_isRet; // @[SRAMTemplate.scala 88:{25,25}]
  assign ftb_io_wreq_bits_data_3_entry_isJalr = io_update_write_data_bits_entry_isJalr; // @[SRAMTemplate.scala 88:{25,25}]
  assign ftb_io_wreq_bits_data_3_entry_last_may_be_rvi_call = io_update_write_data_bits_entry_last_may_be_rvi_call; // @[SRAMTemplate.scala 88:{25,25}]
  assign ftb_io_wreq_bits_data_3_entry_always_taken_0 = io_update_write_data_bits_entry_always_taken_0; // @[SRAMTemplate.scala 88:{25,25}]
  assign ftb_io_wreq_bits_data_3_entry_always_taken_1 = io_update_write_data_bits_entry_always_taken_1; // @[SRAMTemplate.scala 88:{25,25}]
  assign ftb_io_wreq_bits_data_3_tag = io_update_write_data_bits_tag; // @[SRAMTemplate.scala 88:{25,25}]
  assign ftb_io_wreq_bits_waymask = 4'h1 << write_way_bits; // @[OneHot.scala 57:35]
  always @(posedge clock) begin
    pred_rdata_REG <= io_req_pc_valid & ~io_update_access; // @[FTB.scala 305:79]
    if (pred_rdata_REG) begin // @[Reg.scala 17:18]
      pred_rdata_hold_data_0_entry_valid <= ftb_io_rresp_data_0_entry_valid; // @[Reg.scala 17:22]
    end
    if (pred_rdata_REG) begin // @[Reg.scala 17:18]
      pred_rdata_hold_data_0_entry_brSlots_0_offset <= ftb_io_rresp_data_0_entry_brSlots_0_offset; // @[Reg.scala 17:22]
    end
    if (pred_rdata_REG) begin // @[Reg.scala 17:18]
      pred_rdata_hold_data_0_entry_brSlots_0_lower <= ftb_io_rresp_data_0_entry_brSlots_0_lower; // @[Reg.scala 17:22]
    end
    if (pred_rdata_REG) begin // @[Reg.scala 17:18]
      pred_rdata_hold_data_0_entry_brSlots_0_tarStat <= ftb_io_rresp_data_0_entry_brSlots_0_tarStat; // @[Reg.scala 17:22]
    end
    if (pred_rdata_REG) begin // @[Reg.scala 17:18]
      pred_rdata_hold_data_0_entry_brSlots_0_sharing <= ftb_io_rresp_data_0_entry_brSlots_0_sharing; // @[Reg.scala 17:22]
    end
    if (pred_rdata_REG) begin // @[Reg.scala 17:18]
      pred_rdata_hold_data_0_entry_brSlots_0_valid <= ftb_io_rresp_data_0_entry_brSlots_0_valid; // @[Reg.scala 17:22]
    end
    if (pred_rdata_REG) begin // @[Reg.scala 17:18]
      pred_rdata_hold_data_0_entry_tailSlot_offset <= ftb_io_rresp_data_0_entry_tailSlot_offset; // @[Reg.scala 17:22]
    end
    if (pred_rdata_REG) begin // @[Reg.scala 17:18]
      pred_rdata_hold_data_0_entry_tailSlot_lower <= ftb_io_rresp_data_0_entry_tailSlot_lower; // @[Reg.scala 17:22]
    end
    if (pred_rdata_REG) begin // @[Reg.scala 17:18]
      pred_rdata_hold_data_0_entry_tailSlot_tarStat <= ftb_io_rresp_data_0_entry_tailSlot_tarStat; // @[Reg.scala 17:22]
    end
    if (pred_rdata_REG) begin // @[Reg.scala 17:18]
      pred_rdata_hold_data_0_entry_tailSlot_sharing <= ftb_io_rresp_data_0_entry_tailSlot_sharing; // @[Reg.scala 17:22]
    end
    if (pred_rdata_REG) begin // @[Reg.scala 17:18]
      pred_rdata_hold_data_0_entry_tailSlot_valid <= ftb_io_rresp_data_0_entry_tailSlot_valid; // @[Reg.scala 17:22]
    end
    if (pred_rdata_REG) begin // @[Reg.scala 17:18]
      pred_rdata_hold_data_0_entry_pftAddr <= ftb_io_rresp_data_0_entry_pftAddr; // @[Reg.scala 17:22]
    end
    if (pred_rdata_REG) begin // @[Reg.scala 17:18]
      pred_rdata_hold_data_0_entry_carry <= ftb_io_rresp_data_0_entry_carry; // @[Reg.scala 17:22]
    end
    if (pred_rdata_REG) begin // @[Reg.scala 17:18]
      pred_rdata_hold_data_0_entry_isCall <= ftb_io_rresp_data_0_entry_isCall; // @[Reg.scala 17:22]
    end
    if (pred_rdata_REG) begin // @[Reg.scala 17:18]
      pred_rdata_hold_data_0_entry_isRet <= ftb_io_rresp_data_0_entry_isRet; // @[Reg.scala 17:22]
    end
    if (pred_rdata_REG) begin // @[Reg.scala 17:18]
      pred_rdata_hold_data_0_entry_isJalr <= ftb_io_rresp_data_0_entry_isJalr; // @[Reg.scala 17:22]
    end
    if (pred_rdata_REG) begin // @[Reg.scala 17:18]
      pred_rdata_hold_data_0_entry_last_may_be_rvi_call <= ftb_io_rresp_data_0_entry_last_may_be_rvi_call; // @[Reg.scala 17:22]
    end
    if (pred_rdata_REG) begin // @[Reg.scala 17:18]
      pred_rdata_hold_data_0_entry_always_taken_0 <= ftb_io_rresp_data_0_entry_always_taken_0; // @[Reg.scala 17:22]
    end
    if (pred_rdata_REG) begin // @[Reg.scala 17:18]
      pred_rdata_hold_data_0_entry_always_taken_1 <= ftb_io_rresp_data_0_entry_always_taken_1; // @[Reg.scala 17:22]
    end
    if (pred_rdata_REG) begin // @[Reg.scala 17:18]
      pred_rdata_hold_data_0_tag <= ftb_io_rresp_data_0_tag; // @[Reg.scala 17:22]
    end
    if (pred_rdata_REG) begin // @[Reg.scala 17:18]
      pred_rdata_hold_data_1_entry_valid <= ftb_io_rresp_data_1_entry_valid; // @[Reg.scala 17:22]
    end
    if (pred_rdata_REG) begin // @[Reg.scala 17:18]
      pred_rdata_hold_data_1_entry_brSlots_0_offset <= ftb_io_rresp_data_1_entry_brSlots_0_offset; // @[Reg.scala 17:22]
    end
    if (pred_rdata_REG) begin // @[Reg.scala 17:18]
      pred_rdata_hold_data_1_entry_brSlots_0_lower <= ftb_io_rresp_data_1_entry_brSlots_0_lower; // @[Reg.scala 17:22]
    end
    if (pred_rdata_REG) begin // @[Reg.scala 17:18]
      pred_rdata_hold_data_1_entry_brSlots_0_tarStat <= ftb_io_rresp_data_1_entry_brSlots_0_tarStat; // @[Reg.scala 17:22]
    end
    if (pred_rdata_REG) begin // @[Reg.scala 17:18]
      pred_rdata_hold_data_1_entry_brSlots_0_sharing <= ftb_io_rresp_data_1_entry_brSlots_0_sharing; // @[Reg.scala 17:22]
    end
    if (pred_rdata_REG) begin // @[Reg.scala 17:18]
      pred_rdata_hold_data_1_entry_brSlots_0_valid <= ftb_io_rresp_data_1_entry_brSlots_0_valid; // @[Reg.scala 17:22]
    end
    if (pred_rdata_REG) begin // @[Reg.scala 17:18]
      pred_rdata_hold_data_1_entry_tailSlot_offset <= ftb_io_rresp_data_1_entry_tailSlot_offset; // @[Reg.scala 17:22]
    end
    if (pred_rdata_REG) begin // @[Reg.scala 17:18]
      pred_rdata_hold_data_1_entry_tailSlot_lower <= ftb_io_rresp_data_1_entry_tailSlot_lower; // @[Reg.scala 17:22]
    end
    if (pred_rdata_REG) begin // @[Reg.scala 17:18]
      pred_rdata_hold_data_1_entry_tailSlot_tarStat <= ftb_io_rresp_data_1_entry_tailSlot_tarStat; // @[Reg.scala 17:22]
    end
    if (pred_rdata_REG) begin // @[Reg.scala 17:18]
      pred_rdata_hold_data_1_entry_tailSlot_sharing <= ftb_io_rresp_data_1_entry_tailSlot_sharing; // @[Reg.scala 17:22]
    end
    if (pred_rdata_REG) begin // @[Reg.scala 17:18]
      pred_rdata_hold_data_1_entry_tailSlot_valid <= ftb_io_rresp_data_1_entry_tailSlot_valid; // @[Reg.scala 17:22]
    end
    if (pred_rdata_REG) begin // @[Reg.scala 17:18]
      pred_rdata_hold_data_1_entry_pftAddr <= ftb_io_rresp_data_1_entry_pftAddr; // @[Reg.scala 17:22]
    end
    if (pred_rdata_REG) begin // @[Reg.scala 17:18]
      pred_rdata_hold_data_1_entry_carry <= ftb_io_rresp_data_1_entry_carry; // @[Reg.scala 17:22]
    end
    if (pred_rdata_REG) begin // @[Reg.scala 17:18]
      pred_rdata_hold_data_1_entry_isCall <= ftb_io_rresp_data_1_entry_isCall; // @[Reg.scala 17:22]
    end
    if (pred_rdata_REG) begin // @[Reg.scala 17:18]
      pred_rdata_hold_data_1_entry_isRet <= ftb_io_rresp_data_1_entry_isRet; // @[Reg.scala 17:22]
    end
    if (pred_rdata_REG) begin // @[Reg.scala 17:18]
      pred_rdata_hold_data_1_entry_isJalr <= ftb_io_rresp_data_1_entry_isJalr; // @[Reg.scala 17:22]
    end
    if (pred_rdata_REG) begin // @[Reg.scala 17:18]
      pred_rdata_hold_data_1_entry_last_may_be_rvi_call <= ftb_io_rresp_data_1_entry_last_may_be_rvi_call; // @[Reg.scala 17:22]
    end
    if (pred_rdata_REG) begin // @[Reg.scala 17:18]
      pred_rdata_hold_data_1_entry_always_taken_0 <= ftb_io_rresp_data_1_entry_always_taken_0; // @[Reg.scala 17:22]
    end
    if (pred_rdata_REG) begin // @[Reg.scala 17:18]
      pred_rdata_hold_data_1_entry_always_taken_1 <= ftb_io_rresp_data_1_entry_always_taken_1; // @[Reg.scala 17:22]
    end
    if (pred_rdata_REG) begin // @[Reg.scala 17:18]
      pred_rdata_hold_data_1_tag <= ftb_io_rresp_data_1_tag; // @[Reg.scala 17:22]
    end
    if (pred_rdata_REG) begin // @[Reg.scala 17:18]
      pred_rdata_hold_data_2_entry_valid <= ftb_io_rresp_data_2_entry_valid; // @[Reg.scala 17:22]
    end
    if (pred_rdata_REG) begin // @[Reg.scala 17:18]
      pred_rdata_hold_data_2_entry_brSlots_0_offset <= ftb_io_rresp_data_2_entry_brSlots_0_offset; // @[Reg.scala 17:22]
    end
    if (pred_rdata_REG) begin // @[Reg.scala 17:18]
      pred_rdata_hold_data_2_entry_brSlots_0_lower <= ftb_io_rresp_data_2_entry_brSlots_0_lower; // @[Reg.scala 17:22]
    end
    if (pred_rdata_REG) begin // @[Reg.scala 17:18]
      pred_rdata_hold_data_2_entry_brSlots_0_tarStat <= ftb_io_rresp_data_2_entry_brSlots_0_tarStat; // @[Reg.scala 17:22]
    end
    if (pred_rdata_REG) begin // @[Reg.scala 17:18]
      pred_rdata_hold_data_2_entry_brSlots_0_sharing <= ftb_io_rresp_data_2_entry_brSlots_0_sharing; // @[Reg.scala 17:22]
    end
    if (pred_rdata_REG) begin // @[Reg.scala 17:18]
      pred_rdata_hold_data_2_entry_brSlots_0_valid <= ftb_io_rresp_data_2_entry_brSlots_0_valid; // @[Reg.scala 17:22]
    end
    if (pred_rdata_REG) begin // @[Reg.scala 17:18]
      pred_rdata_hold_data_2_entry_tailSlot_offset <= ftb_io_rresp_data_2_entry_tailSlot_offset; // @[Reg.scala 17:22]
    end
    if (pred_rdata_REG) begin // @[Reg.scala 17:18]
      pred_rdata_hold_data_2_entry_tailSlot_lower <= ftb_io_rresp_data_2_entry_tailSlot_lower; // @[Reg.scala 17:22]
    end
    if (pred_rdata_REG) begin // @[Reg.scala 17:18]
      pred_rdata_hold_data_2_entry_tailSlot_tarStat <= ftb_io_rresp_data_2_entry_tailSlot_tarStat; // @[Reg.scala 17:22]
    end
    if (pred_rdata_REG) begin // @[Reg.scala 17:18]
      pred_rdata_hold_data_2_entry_tailSlot_sharing <= ftb_io_rresp_data_2_entry_tailSlot_sharing; // @[Reg.scala 17:22]
    end
    if (pred_rdata_REG) begin // @[Reg.scala 17:18]
      pred_rdata_hold_data_2_entry_tailSlot_valid <= ftb_io_rresp_data_2_entry_tailSlot_valid; // @[Reg.scala 17:22]
    end
    if (pred_rdata_REG) begin // @[Reg.scala 17:18]
      pred_rdata_hold_data_2_entry_pftAddr <= ftb_io_rresp_data_2_entry_pftAddr; // @[Reg.scala 17:22]
    end
    if (pred_rdata_REG) begin // @[Reg.scala 17:18]
      pred_rdata_hold_data_2_entry_carry <= ftb_io_rresp_data_2_entry_carry; // @[Reg.scala 17:22]
    end
    if (pred_rdata_REG) begin // @[Reg.scala 17:18]
      pred_rdata_hold_data_2_entry_isCall <= ftb_io_rresp_data_2_entry_isCall; // @[Reg.scala 17:22]
    end
    if (pred_rdata_REG) begin // @[Reg.scala 17:18]
      pred_rdata_hold_data_2_entry_isRet <= ftb_io_rresp_data_2_entry_isRet; // @[Reg.scala 17:22]
    end
    if (pred_rdata_REG) begin // @[Reg.scala 17:18]
      pred_rdata_hold_data_2_entry_isJalr <= ftb_io_rresp_data_2_entry_isJalr; // @[Reg.scala 17:22]
    end
    if (pred_rdata_REG) begin // @[Reg.scala 17:18]
      pred_rdata_hold_data_2_entry_last_may_be_rvi_call <= ftb_io_rresp_data_2_entry_last_may_be_rvi_call; // @[Reg.scala 17:22]
    end
    if (pred_rdata_REG) begin // @[Reg.scala 17:18]
      pred_rdata_hold_data_2_entry_always_taken_0 <= ftb_io_rresp_data_2_entry_always_taken_0; // @[Reg.scala 17:22]
    end
    if (pred_rdata_REG) begin // @[Reg.scala 17:18]
      pred_rdata_hold_data_2_entry_always_taken_1 <= ftb_io_rresp_data_2_entry_always_taken_1; // @[Reg.scala 17:22]
    end
    if (pred_rdata_REG) begin // @[Reg.scala 17:18]
      pred_rdata_hold_data_2_tag <= ftb_io_rresp_data_2_tag; // @[Reg.scala 17:22]
    end
    if (pred_rdata_REG) begin // @[Reg.scala 17:18]
      pred_rdata_hold_data_3_entry_valid <= ftb_io_rresp_data_3_entry_valid; // @[Reg.scala 17:22]
    end
    if (pred_rdata_REG) begin // @[Reg.scala 17:18]
      pred_rdata_hold_data_3_entry_brSlots_0_offset <= ftb_io_rresp_data_3_entry_brSlots_0_offset; // @[Reg.scala 17:22]
    end
    if (pred_rdata_REG) begin // @[Reg.scala 17:18]
      pred_rdata_hold_data_3_entry_brSlots_0_lower <= ftb_io_rresp_data_3_entry_brSlots_0_lower; // @[Reg.scala 17:22]
    end
    if (pred_rdata_REG) begin // @[Reg.scala 17:18]
      pred_rdata_hold_data_3_entry_brSlots_0_tarStat <= ftb_io_rresp_data_3_entry_brSlots_0_tarStat; // @[Reg.scala 17:22]
    end
    if (pred_rdata_REG) begin // @[Reg.scala 17:18]
      pred_rdata_hold_data_3_entry_brSlots_0_sharing <= ftb_io_rresp_data_3_entry_brSlots_0_sharing; // @[Reg.scala 17:22]
    end
    if (pred_rdata_REG) begin // @[Reg.scala 17:18]
      pred_rdata_hold_data_3_entry_brSlots_0_valid <= ftb_io_rresp_data_3_entry_brSlots_0_valid; // @[Reg.scala 17:22]
    end
    if (pred_rdata_REG) begin // @[Reg.scala 17:18]
      pred_rdata_hold_data_3_entry_tailSlot_offset <= ftb_io_rresp_data_3_entry_tailSlot_offset; // @[Reg.scala 17:22]
    end
    if (pred_rdata_REG) begin // @[Reg.scala 17:18]
      pred_rdata_hold_data_3_entry_tailSlot_lower <= ftb_io_rresp_data_3_entry_tailSlot_lower; // @[Reg.scala 17:22]
    end
    if (pred_rdata_REG) begin // @[Reg.scala 17:18]
      pred_rdata_hold_data_3_entry_tailSlot_tarStat <= ftb_io_rresp_data_3_entry_tailSlot_tarStat; // @[Reg.scala 17:22]
    end
    if (pred_rdata_REG) begin // @[Reg.scala 17:18]
      pred_rdata_hold_data_3_entry_tailSlot_sharing <= ftb_io_rresp_data_3_entry_tailSlot_sharing; // @[Reg.scala 17:22]
    end
    if (pred_rdata_REG) begin // @[Reg.scala 17:18]
      pred_rdata_hold_data_3_entry_tailSlot_valid <= ftb_io_rresp_data_3_entry_tailSlot_valid; // @[Reg.scala 17:22]
    end
    if (pred_rdata_REG) begin // @[Reg.scala 17:18]
      pred_rdata_hold_data_3_entry_pftAddr <= ftb_io_rresp_data_3_entry_pftAddr; // @[Reg.scala 17:22]
    end
    if (pred_rdata_REG) begin // @[Reg.scala 17:18]
      pred_rdata_hold_data_3_entry_carry <= ftb_io_rresp_data_3_entry_carry; // @[Reg.scala 17:22]
    end
    if (pred_rdata_REG) begin // @[Reg.scala 17:18]
      pred_rdata_hold_data_3_entry_isCall <= ftb_io_rresp_data_3_entry_isCall; // @[Reg.scala 17:22]
    end
    if (pred_rdata_REG) begin // @[Reg.scala 17:18]
      pred_rdata_hold_data_3_entry_isRet <= ftb_io_rresp_data_3_entry_isRet; // @[Reg.scala 17:22]
    end
    if (pred_rdata_REG) begin // @[Reg.scala 17:18]
      pred_rdata_hold_data_3_entry_isJalr <= ftb_io_rresp_data_3_entry_isJalr; // @[Reg.scala 17:22]
    end
    if (pred_rdata_REG) begin // @[Reg.scala 17:18]
      pred_rdata_hold_data_3_entry_last_may_be_rvi_call <= ftb_io_rresp_data_3_entry_last_may_be_rvi_call; // @[Reg.scala 17:22]
    end
    if (pred_rdata_REG) begin // @[Reg.scala 17:18]
      pred_rdata_hold_data_3_entry_always_taken_0 <= ftb_io_rresp_data_3_entry_always_taken_0; // @[Reg.scala 17:22]
    end
    if (pred_rdata_REG) begin // @[Reg.scala 17:18]
      pred_rdata_hold_data_3_entry_always_taken_1 <= ftb_io_rresp_data_3_entry_always_taken_1; // @[Reg.scala 17:22]
    end
    if (pred_rdata_REG) begin // @[Reg.scala 17:18]
      pred_rdata_hold_data_3_tag <= ftb_io_rresp_data_3_tag; // @[Reg.scala 17:22]
    end
    if (io_req_pc_valid) begin // @[Reg.scala 17:18]
      req_tag <= io_req_pc_bits[29:10]; // @[Reg.scala 17:22]
    end
    if (io_req_pc_valid) begin // @[Reg.scala 17:18]
      req_idx <= io_req_pc_bits[9:1]; // @[Reg.scala 17:22]
    end
    if (io_u_req_pc_valid) begin // @[Reg.scala 17:18]
      u_req_tag <= io_u_req_pc_bits[29:10]; // @[Reg.scala 17:22]
    end
    u_total_hits_REG <= io_update_access; // @[FTB.scala 328:96]
    u_total_hits_REG_1 <= io_update_access; // @[FTB.scala 328:96]
    u_total_hits_REG_2 <= io_update_access; // @[FTB.scala 328:96]
    u_total_hits_REG_3 <= io_update_access; // @[FTB.scala 328:96]
    allocWriteWay_REG_3 <= ftb_io_rresp_data_3_entry_valid; // @[FTB.scala 386:{49,49}]
    allocWriteWay_REG_2 <= ftb_io_rresp_data_2_entry_valid; // @[FTB.scala 386:{49,49}]
    allocWriteWay_REG_1 <= ftb_io_rresp_data_1_entry_valid; // @[FTB.scala 386:{49,49}]
    allocWriteWay_REG_0 <= ftb_io_rresp_data_0_entry_valid; // @[FTB.scala 386:{49,49}]
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_0 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_valid) begin
        state_vec_0 <= _state_vec_0_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_1 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_1_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_1_valid) begin
        state_vec_1 <= _state_vec_1_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_2 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_2_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_2_valid) begin
        state_vec_2 <= _state_vec_2_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_3 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_3_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_3_valid) begin
        state_vec_3 <= _state_vec_3_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_4 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_4_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_4_valid) begin
        state_vec_4 <= _state_vec_4_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_5 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_5_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_5_valid) begin
        state_vec_5 <= _state_vec_5_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_6 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_6_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_6_valid) begin
        state_vec_6 <= _state_vec_6_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_7 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_7_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_7_valid) begin
        state_vec_7 <= _state_vec_7_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_8 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_8_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_8_valid) begin
        state_vec_8 <= _state_vec_8_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_9 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_9_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_9_valid) begin
        state_vec_9 <= _state_vec_9_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_10 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_10_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_10_valid) begin
        state_vec_10 <= _state_vec_10_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_11 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_11_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_11_valid) begin
        state_vec_11 <= _state_vec_11_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_12 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_12_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_12_valid) begin
        state_vec_12 <= _state_vec_12_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_13 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_13_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_13_valid) begin
        state_vec_13 <= _state_vec_13_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_14 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_14_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_14_valid) begin
        state_vec_14 <= _state_vec_14_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_15 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_15_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_15_valid) begin
        state_vec_15 <= _state_vec_15_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_16 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_16_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_16_valid) begin
        state_vec_16 <= _state_vec_16_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_17 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_17_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_17_valid) begin
        state_vec_17 <= _state_vec_17_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_18 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_18_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_18_valid) begin
        state_vec_18 <= _state_vec_18_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_19 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_19_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_19_valid) begin
        state_vec_19 <= _state_vec_19_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_20 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_20_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_20_valid) begin
        state_vec_20 <= _state_vec_20_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_21 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_21_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_21_valid) begin
        state_vec_21 <= _state_vec_21_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_22 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_22_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_22_valid) begin
        state_vec_22 <= _state_vec_22_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_23 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_23_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_23_valid) begin
        state_vec_23 <= _state_vec_23_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_24 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_24_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_24_valid) begin
        state_vec_24 <= _state_vec_24_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_25 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_25_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_25_valid) begin
        state_vec_25 <= _state_vec_25_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_26 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_26_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_26_valid) begin
        state_vec_26 <= _state_vec_26_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_27 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_27_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_27_valid) begin
        state_vec_27 <= _state_vec_27_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_28 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_28_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_28_valid) begin
        state_vec_28 <= _state_vec_28_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_29 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_29_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_29_valid) begin
        state_vec_29 <= _state_vec_29_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_30 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_30_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_30_valid) begin
        state_vec_30 <= _state_vec_30_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_31 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_31_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_31_valid) begin
        state_vec_31 <= _state_vec_31_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_32 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_32_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_32_valid) begin
        state_vec_32 <= _state_vec_32_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_33 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_33_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_33_valid) begin
        state_vec_33 <= _state_vec_33_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_34 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_34_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_34_valid) begin
        state_vec_34 <= _state_vec_34_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_35 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_35_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_35_valid) begin
        state_vec_35 <= _state_vec_35_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_36 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_36_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_36_valid) begin
        state_vec_36 <= _state_vec_36_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_37 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_37_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_37_valid) begin
        state_vec_37 <= _state_vec_37_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_38 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_38_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_38_valid) begin
        state_vec_38 <= _state_vec_38_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_39 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_39_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_39_valid) begin
        state_vec_39 <= _state_vec_39_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_40 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_40_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_40_valid) begin
        state_vec_40 <= _state_vec_40_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_41 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_41_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_41_valid) begin
        state_vec_41 <= _state_vec_41_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_42 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_42_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_42_valid) begin
        state_vec_42 <= _state_vec_42_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_43 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_43_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_43_valid) begin
        state_vec_43 <= _state_vec_43_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_44 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_44_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_44_valid) begin
        state_vec_44 <= _state_vec_44_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_45 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_45_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_45_valid) begin
        state_vec_45 <= _state_vec_45_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_46 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_46_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_46_valid) begin
        state_vec_46 <= _state_vec_46_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_47 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_47_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_47_valid) begin
        state_vec_47 <= _state_vec_47_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_48 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_48_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_48_valid) begin
        state_vec_48 <= _state_vec_48_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_49 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_49_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_49_valid) begin
        state_vec_49 <= _state_vec_49_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_50 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_50_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_50_valid) begin
        state_vec_50 <= _state_vec_50_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_51 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_51_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_51_valid) begin
        state_vec_51 <= _state_vec_51_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_52 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_52_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_52_valid) begin
        state_vec_52 <= _state_vec_52_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_53 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_53_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_53_valid) begin
        state_vec_53 <= _state_vec_53_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_54 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_54_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_54_valid) begin
        state_vec_54 <= _state_vec_54_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_55 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_55_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_55_valid) begin
        state_vec_55 <= _state_vec_55_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_56 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_56_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_56_valid) begin
        state_vec_56 <= _state_vec_56_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_57 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_57_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_57_valid) begin
        state_vec_57 <= _state_vec_57_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_58 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_58_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_58_valid) begin
        state_vec_58 <= _state_vec_58_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_59 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_59_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_59_valid) begin
        state_vec_59 <= _state_vec_59_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_60 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_60_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_60_valid) begin
        state_vec_60 <= _state_vec_60_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_61 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_61_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_61_valid) begin
        state_vec_61 <= _state_vec_61_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_62 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_62_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_62_valid) begin
        state_vec_62 <= _state_vec_62_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_63 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_63_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_63_valid) begin
        state_vec_63 <= _state_vec_63_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_64 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_64_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_64_valid) begin
        state_vec_64 <= _state_vec_64_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_65 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_65_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_65_valid) begin
        state_vec_65 <= _state_vec_65_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_66 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_66_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_66_valid) begin
        state_vec_66 <= _state_vec_66_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_67 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_67_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_67_valid) begin
        state_vec_67 <= _state_vec_67_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_68 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_68_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_68_valid) begin
        state_vec_68 <= _state_vec_68_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_69 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_69_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_69_valid) begin
        state_vec_69 <= _state_vec_69_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_70 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_70_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_70_valid) begin
        state_vec_70 <= _state_vec_70_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_71 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_71_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_71_valid) begin
        state_vec_71 <= _state_vec_71_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_72 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_72_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_72_valid) begin
        state_vec_72 <= _state_vec_72_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_73 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_73_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_73_valid) begin
        state_vec_73 <= _state_vec_73_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_74 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_74_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_74_valid) begin
        state_vec_74 <= _state_vec_74_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_75 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_75_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_75_valid) begin
        state_vec_75 <= _state_vec_75_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_76 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_76_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_76_valid) begin
        state_vec_76 <= _state_vec_76_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_77 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_77_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_77_valid) begin
        state_vec_77 <= _state_vec_77_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_78 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_78_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_78_valid) begin
        state_vec_78 <= _state_vec_78_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_79 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_79_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_79_valid) begin
        state_vec_79 <= _state_vec_79_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_80 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_80_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_80_valid) begin
        state_vec_80 <= _state_vec_80_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_81 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_81_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_81_valid) begin
        state_vec_81 <= _state_vec_81_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_82 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_82_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_82_valid) begin
        state_vec_82 <= _state_vec_82_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_83 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_83_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_83_valid) begin
        state_vec_83 <= _state_vec_83_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_84 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_84_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_84_valid) begin
        state_vec_84 <= _state_vec_84_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_85 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_85_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_85_valid) begin
        state_vec_85 <= _state_vec_85_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_86 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_86_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_86_valid) begin
        state_vec_86 <= _state_vec_86_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_87 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_87_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_87_valid) begin
        state_vec_87 <= _state_vec_87_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_88 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_88_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_88_valid) begin
        state_vec_88 <= _state_vec_88_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_89 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_89_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_89_valid) begin
        state_vec_89 <= _state_vec_89_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_90 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_90_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_90_valid) begin
        state_vec_90 <= _state_vec_90_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_91 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_91_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_91_valid) begin
        state_vec_91 <= _state_vec_91_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_92 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_92_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_92_valid) begin
        state_vec_92 <= _state_vec_92_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_93 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_93_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_93_valid) begin
        state_vec_93 <= _state_vec_93_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_94 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_94_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_94_valid) begin
        state_vec_94 <= _state_vec_94_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_95 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_95_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_95_valid) begin
        state_vec_95 <= _state_vec_95_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_96 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_96_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_96_valid) begin
        state_vec_96 <= _state_vec_96_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_97 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_97_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_97_valid) begin
        state_vec_97 <= _state_vec_97_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_98 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_98_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_98_valid) begin
        state_vec_98 <= _state_vec_98_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_99 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_99_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_99_valid) begin
        state_vec_99 <= _state_vec_99_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_100 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_100_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_100_valid) begin
        state_vec_100 <= _state_vec_100_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_101 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_101_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_101_valid) begin
        state_vec_101 <= _state_vec_101_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_102 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_102_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_102_valid) begin
        state_vec_102 <= _state_vec_102_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_103 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_103_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_103_valid) begin
        state_vec_103 <= _state_vec_103_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_104 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_104_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_104_valid) begin
        state_vec_104 <= _state_vec_104_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_105 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_105_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_105_valid) begin
        state_vec_105 <= _state_vec_105_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_106 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_106_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_106_valid) begin
        state_vec_106 <= _state_vec_106_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_107 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_107_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_107_valid) begin
        state_vec_107 <= _state_vec_107_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_108 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_108_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_108_valid) begin
        state_vec_108 <= _state_vec_108_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_109 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_109_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_109_valid) begin
        state_vec_109 <= _state_vec_109_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_110 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_110_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_110_valid) begin
        state_vec_110 <= _state_vec_110_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_111 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_111_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_111_valid) begin
        state_vec_111 <= _state_vec_111_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_112 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_112_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_112_valid) begin
        state_vec_112 <= _state_vec_112_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_113 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_113_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_113_valid) begin
        state_vec_113 <= _state_vec_113_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_114 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_114_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_114_valid) begin
        state_vec_114 <= _state_vec_114_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_115 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_115_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_115_valid) begin
        state_vec_115 <= _state_vec_115_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_116 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_116_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_116_valid) begin
        state_vec_116 <= _state_vec_116_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_117 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_117_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_117_valid) begin
        state_vec_117 <= _state_vec_117_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_118 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_118_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_118_valid) begin
        state_vec_118 <= _state_vec_118_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_119 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_119_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_119_valid) begin
        state_vec_119 <= _state_vec_119_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_120 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_120_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_120_valid) begin
        state_vec_120 <= _state_vec_120_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_121 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_121_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_121_valid) begin
        state_vec_121 <= _state_vec_121_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_122 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_122_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_122_valid) begin
        state_vec_122 <= _state_vec_122_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_123 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_123_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_123_valid) begin
        state_vec_123 <= _state_vec_123_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_124 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_124_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_124_valid) begin
        state_vec_124 <= _state_vec_124_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_125 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_125_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_125_valid) begin
        state_vec_125 <= _state_vec_125_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_126 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_126_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_126_valid) begin
        state_vec_126 <= _state_vec_126_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_127 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_127_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_127_valid) begin
        state_vec_127 <= _state_vec_127_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_128 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_128_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_128_valid) begin
        state_vec_128 <= _state_vec_128_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_129 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_129_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_129_valid) begin
        state_vec_129 <= _state_vec_129_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_130 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_130_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_130_valid) begin
        state_vec_130 <= _state_vec_130_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_131 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_131_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_131_valid) begin
        state_vec_131 <= _state_vec_131_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_132 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_132_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_132_valid) begin
        state_vec_132 <= _state_vec_132_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_133 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_133_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_133_valid) begin
        state_vec_133 <= _state_vec_133_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_134 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_134_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_134_valid) begin
        state_vec_134 <= _state_vec_134_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_135 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_135_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_135_valid) begin
        state_vec_135 <= _state_vec_135_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_136 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_136_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_136_valid) begin
        state_vec_136 <= _state_vec_136_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_137 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_137_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_137_valid) begin
        state_vec_137 <= _state_vec_137_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_138 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_138_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_138_valid) begin
        state_vec_138 <= _state_vec_138_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_139 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_139_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_139_valid) begin
        state_vec_139 <= _state_vec_139_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_140 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_140_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_140_valid) begin
        state_vec_140 <= _state_vec_140_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_141 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_141_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_141_valid) begin
        state_vec_141 <= _state_vec_141_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_142 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_142_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_142_valid) begin
        state_vec_142 <= _state_vec_142_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_143 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_143_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_143_valid) begin
        state_vec_143 <= _state_vec_143_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_144 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_144_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_144_valid) begin
        state_vec_144 <= _state_vec_144_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_145 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_145_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_145_valid) begin
        state_vec_145 <= _state_vec_145_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_146 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_146_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_146_valid) begin
        state_vec_146 <= _state_vec_146_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_147 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_147_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_147_valid) begin
        state_vec_147 <= _state_vec_147_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_148 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_148_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_148_valid) begin
        state_vec_148 <= _state_vec_148_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_149 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_149_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_149_valid) begin
        state_vec_149 <= _state_vec_149_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_150 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_150_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_150_valid) begin
        state_vec_150 <= _state_vec_150_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_151 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_151_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_151_valid) begin
        state_vec_151 <= _state_vec_151_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_152 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_152_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_152_valid) begin
        state_vec_152 <= _state_vec_152_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_153 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_153_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_153_valid) begin
        state_vec_153 <= _state_vec_153_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_154 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_154_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_154_valid) begin
        state_vec_154 <= _state_vec_154_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_155 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_155_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_155_valid) begin
        state_vec_155 <= _state_vec_155_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_156 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_156_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_156_valid) begin
        state_vec_156 <= _state_vec_156_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_157 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_157_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_157_valid) begin
        state_vec_157 <= _state_vec_157_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_158 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_158_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_158_valid) begin
        state_vec_158 <= _state_vec_158_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_159 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_159_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_159_valid) begin
        state_vec_159 <= _state_vec_159_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_160 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_160_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_160_valid) begin
        state_vec_160 <= _state_vec_160_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_161 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_161_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_161_valid) begin
        state_vec_161 <= _state_vec_161_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_162 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_162_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_162_valid) begin
        state_vec_162 <= _state_vec_162_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_163 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_163_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_163_valid) begin
        state_vec_163 <= _state_vec_163_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_164 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_164_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_164_valid) begin
        state_vec_164 <= _state_vec_164_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_165 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_165_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_165_valid) begin
        state_vec_165 <= _state_vec_165_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_166 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_166_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_166_valid) begin
        state_vec_166 <= _state_vec_166_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_167 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_167_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_167_valid) begin
        state_vec_167 <= _state_vec_167_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_168 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_168_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_168_valid) begin
        state_vec_168 <= _state_vec_168_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_169 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_169_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_169_valid) begin
        state_vec_169 <= _state_vec_169_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_170 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_170_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_170_valid) begin
        state_vec_170 <= _state_vec_170_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_171 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_171_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_171_valid) begin
        state_vec_171 <= _state_vec_171_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_172 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_172_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_172_valid) begin
        state_vec_172 <= _state_vec_172_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_173 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_173_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_173_valid) begin
        state_vec_173 <= _state_vec_173_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_174 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_174_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_174_valid) begin
        state_vec_174 <= _state_vec_174_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_175 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_175_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_175_valid) begin
        state_vec_175 <= _state_vec_175_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_176 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_176_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_176_valid) begin
        state_vec_176 <= _state_vec_176_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_177 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_177_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_177_valid) begin
        state_vec_177 <= _state_vec_177_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_178 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_178_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_178_valid) begin
        state_vec_178 <= _state_vec_178_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_179 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_179_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_179_valid) begin
        state_vec_179 <= _state_vec_179_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_180 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_180_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_180_valid) begin
        state_vec_180 <= _state_vec_180_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_181 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_181_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_181_valid) begin
        state_vec_181 <= _state_vec_181_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_182 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_182_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_182_valid) begin
        state_vec_182 <= _state_vec_182_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_183 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_183_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_183_valid) begin
        state_vec_183 <= _state_vec_183_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_184 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_184_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_184_valid) begin
        state_vec_184 <= _state_vec_184_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_185 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_185_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_185_valid) begin
        state_vec_185 <= _state_vec_185_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_186 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_186_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_186_valid) begin
        state_vec_186 <= _state_vec_186_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_187 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_187_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_187_valid) begin
        state_vec_187 <= _state_vec_187_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_188 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_188_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_188_valid) begin
        state_vec_188 <= _state_vec_188_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_189 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_189_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_189_valid) begin
        state_vec_189 <= _state_vec_189_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_190 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_190_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_190_valid) begin
        state_vec_190 <= _state_vec_190_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_191 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_191_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_191_valid) begin
        state_vec_191 <= _state_vec_191_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_192 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_192_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_192_valid) begin
        state_vec_192 <= _state_vec_192_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_193 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_193_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_193_valid) begin
        state_vec_193 <= _state_vec_193_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_194 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_194_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_194_valid) begin
        state_vec_194 <= _state_vec_194_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_195 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_195_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_195_valid) begin
        state_vec_195 <= _state_vec_195_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_196 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_196_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_196_valid) begin
        state_vec_196 <= _state_vec_196_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_197 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_197_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_197_valid) begin
        state_vec_197 <= _state_vec_197_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_198 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_198_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_198_valid) begin
        state_vec_198 <= _state_vec_198_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_199 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_199_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_199_valid) begin
        state_vec_199 <= _state_vec_199_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_200 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_200_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_200_valid) begin
        state_vec_200 <= _state_vec_200_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_201 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_201_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_201_valid) begin
        state_vec_201 <= _state_vec_201_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_202 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_202_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_202_valid) begin
        state_vec_202 <= _state_vec_202_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_203 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_203_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_203_valid) begin
        state_vec_203 <= _state_vec_203_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_204 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_204_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_204_valid) begin
        state_vec_204 <= _state_vec_204_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_205 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_205_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_205_valid) begin
        state_vec_205 <= _state_vec_205_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_206 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_206_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_206_valid) begin
        state_vec_206 <= _state_vec_206_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_207 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_207_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_207_valid) begin
        state_vec_207 <= _state_vec_207_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_208 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_208_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_208_valid) begin
        state_vec_208 <= _state_vec_208_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_209 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_209_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_209_valid) begin
        state_vec_209 <= _state_vec_209_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_210 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_210_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_210_valid) begin
        state_vec_210 <= _state_vec_210_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_211 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_211_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_211_valid) begin
        state_vec_211 <= _state_vec_211_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_212 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_212_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_212_valid) begin
        state_vec_212 <= _state_vec_212_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_213 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_213_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_213_valid) begin
        state_vec_213 <= _state_vec_213_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_214 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_214_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_214_valid) begin
        state_vec_214 <= _state_vec_214_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_215 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_215_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_215_valid) begin
        state_vec_215 <= _state_vec_215_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_216 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_216_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_216_valid) begin
        state_vec_216 <= _state_vec_216_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_217 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_217_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_217_valid) begin
        state_vec_217 <= _state_vec_217_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_218 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_218_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_218_valid) begin
        state_vec_218 <= _state_vec_218_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_219 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_219_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_219_valid) begin
        state_vec_219 <= _state_vec_219_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_220 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_220_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_220_valid) begin
        state_vec_220 <= _state_vec_220_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_221 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_221_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_221_valid) begin
        state_vec_221 <= _state_vec_221_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_222 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_222_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_222_valid) begin
        state_vec_222 <= _state_vec_222_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_223 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_223_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_223_valid) begin
        state_vec_223 <= _state_vec_223_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_224 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_224_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_224_valid) begin
        state_vec_224 <= _state_vec_224_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_225 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_225_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_225_valid) begin
        state_vec_225 <= _state_vec_225_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_226 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_226_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_226_valid) begin
        state_vec_226 <= _state_vec_226_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_227 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_227_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_227_valid) begin
        state_vec_227 <= _state_vec_227_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_228 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_228_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_228_valid) begin
        state_vec_228 <= _state_vec_228_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_229 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_229_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_229_valid) begin
        state_vec_229 <= _state_vec_229_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_230 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_230_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_230_valid) begin
        state_vec_230 <= _state_vec_230_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_231 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_231_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_231_valid) begin
        state_vec_231 <= _state_vec_231_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_232 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_232_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_232_valid) begin
        state_vec_232 <= _state_vec_232_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_233 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_233_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_233_valid) begin
        state_vec_233 <= _state_vec_233_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_234 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_234_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_234_valid) begin
        state_vec_234 <= _state_vec_234_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_235 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_235_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_235_valid) begin
        state_vec_235 <= _state_vec_235_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_236 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_236_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_236_valid) begin
        state_vec_236 <= _state_vec_236_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_237 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_237_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_237_valid) begin
        state_vec_237 <= _state_vec_237_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_238 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_238_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_238_valid) begin
        state_vec_238 <= _state_vec_238_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_239 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_239_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_239_valid) begin
        state_vec_239 <= _state_vec_239_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_240 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_240_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_240_valid) begin
        state_vec_240 <= _state_vec_240_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_241 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_241_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_241_valid) begin
        state_vec_241 <= _state_vec_241_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_242 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_242_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_242_valid) begin
        state_vec_242 <= _state_vec_242_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_243 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_243_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_243_valid) begin
        state_vec_243 <= _state_vec_243_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_244 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_244_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_244_valid) begin
        state_vec_244 <= _state_vec_244_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_245 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_245_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_245_valid) begin
        state_vec_245 <= _state_vec_245_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_246 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_246_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_246_valid) begin
        state_vec_246 <= _state_vec_246_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_247 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_247_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_247_valid) begin
        state_vec_247 <= _state_vec_247_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_248 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_248_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_248_valid) begin
        state_vec_248 <= _state_vec_248_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_249 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_249_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_249_valid) begin
        state_vec_249 <= _state_vec_249_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_250 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_250_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_250_valid) begin
        state_vec_250 <= _state_vec_250_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_251 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_251_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_251_valid) begin
        state_vec_251 <= _state_vec_251_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_252 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_252_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_252_valid) begin
        state_vec_252 <= _state_vec_252_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_253 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_253_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_253_valid) begin
        state_vec_253 <= _state_vec_253_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_254 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_254_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_254_valid) begin
        state_vec_254 <= _state_vec_254_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_255 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_255_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_255_valid) begin
        state_vec_255 <= _state_vec_255_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_256 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_256_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_256_valid) begin
        state_vec_256 <= _state_vec_256_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_257 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_257_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_257_valid) begin
        state_vec_257 <= _state_vec_257_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_258 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_258_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_258_valid) begin
        state_vec_258 <= _state_vec_258_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_259 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_259_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_259_valid) begin
        state_vec_259 <= _state_vec_259_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_260 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_260_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_260_valid) begin
        state_vec_260 <= _state_vec_260_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_261 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_261_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_261_valid) begin
        state_vec_261 <= _state_vec_261_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_262 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_262_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_262_valid) begin
        state_vec_262 <= _state_vec_262_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_263 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_263_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_263_valid) begin
        state_vec_263 <= _state_vec_263_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_264 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_264_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_264_valid) begin
        state_vec_264 <= _state_vec_264_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_265 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_265_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_265_valid) begin
        state_vec_265 <= _state_vec_265_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_266 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_266_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_266_valid) begin
        state_vec_266 <= _state_vec_266_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_267 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_267_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_267_valid) begin
        state_vec_267 <= _state_vec_267_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_268 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_268_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_268_valid) begin
        state_vec_268 <= _state_vec_268_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_269 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_269_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_269_valid) begin
        state_vec_269 <= _state_vec_269_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_270 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_270_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_270_valid) begin
        state_vec_270 <= _state_vec_270_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_271 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_271_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_271_valid) begin
        state_vec_271 <= _state_vec_271_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_272 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_272_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_272_valid) begin
        state_vec_272 <= _state_vec_272_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_273 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_273_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_273_valid) begin
        state_vec_273 <= _state_vec_273_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_274 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_274_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_274_valid) begin
        state_vec_274 <= _state_vec_274_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_275 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_275_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_275_valid) begin
        state_vec_275 <= _state_vec_275_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_276 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_276_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_276_valid) begin
        state_vec_276 <= _state_vec_276_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_277 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_277_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_277_valid) begin
        state_vec_277 <= _state_vec_277_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_278 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_278_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_278_valid) begin
        state_vec_278 <= _state_vec_278_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_279 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_279_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_279_valid) begin
        state_vec_279 <= _state_vec_279_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_280 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_280_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_280_valid) begin
        state_vec_280 <= _state_vec_280_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_281 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_281_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_281_valid) begin
        state_vec_281 <= _state_vec_281_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_282 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_282_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_282_valid) begin
        state_vec_282 <= _state_vec_282_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_283 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_283_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_283_valid) begin
        state_vec_283 <= _state_vec_283_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_284 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_284_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_284_valid) begin
        state_vec_284 <= _state_vec_284_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_285 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_285_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_285_valid) begin
        state_vec_285 <= _state_vec_285_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_286 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_286_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_286_valid) begin
        state_vec_286 <= _state_vec_286_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_287 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_287_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_287_valid) begin
        state_vec_287 <= _state_vec_287_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_288 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_288_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_288_valid) begin
        state_vec_288 <= _state_vec_288_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_289 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_289_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_289_valid) begin
        state_vec_289 <= _state_vec_289_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_290 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_290_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_290_valid) begin
        state_vec_290 <= _state_vec_290_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_291 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_291_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_291_valid) begin
        state_vec_291 <= _state_vec_291_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_292 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_292_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_292_valid) begin
        state_vec_292 <= _state_vec_292_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_293 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_293_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_293_valid) begin
        state_vec_293 <= _state_vec_293_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_294 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_294_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_294_valid) begin
        state_vec_294 <= _state_vec_294_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_295 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_295_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_295_valid) begin
        state_vec_295 <= _state_vec_295_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_296 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_296_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_296_valid) begin
        state_vec_296 <= _state_vec_296_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_297 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_297_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_297_valid) begin
        state_vec_297 <= _state_vec_297_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_298 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_298_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_298_valid) begin
        state_vec_298 <= _state_vec_298_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_299 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_299_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_299_valid) begin
        state_vec_299 <= _state_vec_299_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_300 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_300_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_300_valid) begin
        state_vec_300 <= _state_vec_300_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_301 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_301_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_301_valid) begin
        state_vec_301 <= _state_vec_301_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_302 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_302_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_302_valid) begin
        state_vec_302 <= _state_vec_302_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_303 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_303_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_303_valid) begin
        state_vec_303 <= _state_vec_303_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_304 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_304_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_304_valid) begin
        state_vec_304 <= _state_vec_304_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_305 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_305_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_305_valid) begin
        state_vec_305 <= _state_vec_305_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_306 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_306_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_306_valid) begin
        state_vec_306 <= _state_vec_306_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_307 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_307_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_307_valid) begin
        state_vec_307 <= _state_vec_307_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_308 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_308_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_308_valid) begin
        state_vec_308 <= _state_vec_308_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_309 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_309_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_309_valid) begin
        state_vec_309 <= _state_vec_309_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_310 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_310_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_310_valid) begin
        state_vec_310 <= _state_vec_310_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_311 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_311_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_311_valid) begin
        state_vec_311 <= _state_vec_311_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_312 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_312_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_312_valid) begin
        state_vec_312 <= _state_vec_312_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_313 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_313_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_313_valid) begin
        state_vec_313 <= _state_vec_313_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_314 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_314_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_314_valid) begin
        state_vec_314 <= _state_vec_314_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_315 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_315_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_315_valid) begin
        state_vec_315 <= _state_vec_315_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_316 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_316_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_316_valid) begin
        state_vec_316 <= _state_vec_316_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_317 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_317_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_317_valid) begin
        state_vec_317 <= _state_vec_317_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_318 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_318_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_318_valid) begin
        state_vec_318 <= _state_vec_318_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_319 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_319_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_319_valid) begin
        state_vec_319 <= _state_vec_319_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_320 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_320_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_320_valid) begin
        state_vec_320 <= _state_vec_320_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_321 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_321_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_321_valid) begin
        state_vec_321 <= _state_vec_321_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_322 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_322_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_322_valid) begin
        state_vec_322 <= _state_vec_322_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_323 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_323_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_323_valid) begin
        state_vec_323 <= _state_vec_323_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_324 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_324_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_324_valid) begin
        state_vec_324 <= _state_vec_324_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_325 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_325_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_325_valid) begin
        state_vec_325 <= _state_vec_325_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_326 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_326_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_326_valid) begin
        state_vec_326 <= _state_vec_326_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_327 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_327_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_327_valid) begin
        state_vec_327 <= _state_vec_327_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_328 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_328_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_328_valid) begin
        state_vec_328 <= _state_vec_328_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_329 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_329_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_329_valid) begin
        state_vec_329 <= _state_vec_329_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_330 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_330_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_330_valid) begin
        state_vec_330 <= _state_vec_330_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_331 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_331_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_331_valid) begin
        state_vec_331 <= _state_vec_331_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_332 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_332_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_332_valid) begin
        state_vec_332 <= _state_vec_332_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_333 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_333_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_333_valid) begin
        state_vec_333 <= _state_vec_333_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_334 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_334_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_334_valid) begin
        state_vec_334 <= _state_vec_334_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_335 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_335_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_335_valid) begin
        state_vec_335 <= _state_vec_335_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_336 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_336_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_336_valid) begin
        state_vec_336 <= _state_vec_336_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_337 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_337_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_337_valid) begin
        state_vec_337 <= _state_vec_337_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_338 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_338_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_338_valid) begin
        state_vec_338 <= _state_vec_338_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_339 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_339_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_339_valid) begin
        state_vec_339 <= _state_vec_339_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_340 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_340_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_340_valid) begin
        state_vec_340 <= _state_vec_340_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_341 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_341_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_341_valid) begin
        state_vec_341 <= _state_vec_341_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_342 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_342_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_342_valid) begin
        state_vec_342 <= _state_vec_342_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_343 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_343_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_343_valid) begin
        state_vec_343 <= _state_vec_343_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_344 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_344_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_344_valid) begin
        state_vec_344 <= _state_vec_344_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_345 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_345_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_345_valid) begin
        state_vec_345 <= _state_vec_345_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_346 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_346_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_346_valid) begin
        state_vec_346 <= _state_vec_346_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_347 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_347_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_347_valid) begin
        state_vec_347 <= _state_vec_347_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_348 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_348_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_348_valid) begin
        state_vec_348 <= _state_vec_348_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_349 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_349_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_349_valid) begin
        state_vec_349 <= _state_vec_349_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_350 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_350_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_350_valid) begin
        state_vec_350 <= _state_vec_350_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_351 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_351_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_351_valid) begin
        state_vec_351 <= _state_vec_351_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_352 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_352_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_352_valid) begin
        state_vec_352 <= _state_vec_352_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_353 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_353_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_353_valid) begin
        state_vec_353 <= _state_vec_353_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_354 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_354_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_354_valid) begin
        state_vec_354 <= _state_vec_354_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_355 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_355_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_355_valid) begin
        state_vec_355 <= _state_vec_355_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_356 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_356_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_356_valid) begin
        state_vec_356 <= _state_vec_356_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_357 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_357_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_357_valid) begin
        state_vec_357 <= _state_vec_357_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_358 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_358_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_358_valid) begin
        state_vec_358 <= _state_vec_358_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_359 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_359_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_359_valid) begin
        state_vec_359 <= _state_vec_359_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_360 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_360_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_360_valid) begin
        state_vec_360 <= _state_vec_360_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_361 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_361_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_361_valid) begin
        state_vec_361 <= _state_vec_361_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_362 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_362_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_362_valid) begin
        state_vec_362 <= _state_vec_362_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_363 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_363_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_363_valid) begin
        state_vec_363 <= _state_vec_363_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_364 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_364_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_364_valid) begin
        state_vec_364 <= _state_vec_364_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_365 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_365_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_365_valid) begin
        state_vec_365 <= _state_vec_365_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_366 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_366_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_366_valid) begin
        state_vec_366 <= _state_vec_366_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_367 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_367_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_367_valid) begin
        state_vec_367 <= _state_vec_367_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_368 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_368_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_368_valid) begin
        state_vec_368 <= _state_vec_368_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_369 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_369_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_369_valid) begin
        state_vec_369 <= _state_vec_369_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_370 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_370_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_370_valid) begin
        state_vec_370 <= _state_vec_370_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_371 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_371_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_371_valid) begin
        state_vec_371 <= _state_vec_371_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_372 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_372_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_372_valid) begin
        state_vec_372 <= _state_vec_372_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_373 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_373_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_373_valid) begin
        state_vec_373 <= _state_vec_373_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_374 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_374_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_374_valid) begin
        state_vec_374 <= _state_vec_374_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_375 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_375_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_375_valid) begin
        state_vec_375 <= _state_vec_375_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_376 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_376_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_376_valid) begin
        state_vec_376 <= _state_vec_376_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_377 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_377_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_377_valid) begin
        state_vec_377 <= _state_vec_377_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_378 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_378_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_378_valid) begin
        state_vec_378 <= _state_vec_378_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_379 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_379_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_379_valid) begin
        state_vec_379 <= _state_vec_379_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_380 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_380_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_380_valid) begin
        state_vec_380 <= _state_vec_380_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_381 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_381_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_381_valid) begin
        state_vec_381 <= _state_vec_381_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_382 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_382_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_382_valid) begin
        state_vec_382 <= _state_vec_382_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_383 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_383_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_383_valid) begin
        state_vec_383 <= _state_vec_383_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_384 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_384_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_384_valid) begin
        state_vec_384 <= _state_vec_384_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_385 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_385_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_385_valid) begin
        state_vec_385 <= _state_vec_385_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_386 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_386_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_386_valid) begin
        state_vec_386 <= _state_vec_386_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_387 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_387_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_387_valid) begin
        state_vec_387 <= _state_vec_387_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_388 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_388_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_388_valid) begin
        state_vec_388 <= _state_vec_388_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_389 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_389_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_389_valid) begin
        state_vec_389 <= _state_vec_389_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_390 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_390_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_390_valid) begin
        state_vec_390 <= _state_vec_390_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_391 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_391_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_391_valid) begin
        state_vec_391 <= _state_vec_391_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_392 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_392_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_392_valid) begin
        state_vec_392 <= _state_vec_392_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_393 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_393_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_393_valid) begin
        state_vec_393 <= _state_vec_393_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_394 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_394_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_394_valid) begin
        state_vec_394 <= _state_vec_394_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_395 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_395_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_395_valid) begin
        state_vec_395 <= _state_vec_395_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_396 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_396_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_396_valid) begin
        state_vec_396 <= _state_vec_396_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_397 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_397_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_397_valid) begin
        state_vec_397 <= _state_vec_397_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_398 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_398_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_398_valid) begin
        state_vec_398 <= _state_vec_398_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_399 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_399_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_399_valid) begin
        state_vec_399 <= _state_vec_399_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_400 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_400_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_400_valid) begin
        state_vec_400 <= _state_vec_400_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_401 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_401_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_401_valid) begin
        state_vec_401 <= _state_vec_401_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_402 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_402_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_402_valid) begin
        state_vec_402 <= _state_vec_402_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_403 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_403_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_403_valid) begin
        state_vec_403 <= _state_vec_403_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_404 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_404_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_404_valid) begin
        state_vec_404 <= _state_vec_404_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_405 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_405_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_405_valid) begin
        state_vec_405 <= _state_vec_405_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_406 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_406_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_406_valid) begin
        state_vec_406 <= _state_vec_406_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_407 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_407_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_407_valid) begin
        state_vec_407 <= _state_vec_407_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_408 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_408_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_408_valid) begin
        state_vec_408 <= _state_vec_408_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_409 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_409_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_409_valid) begin
        state_vec_409 <= _state_vec_409_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_410 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_410_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_410_valid) begin
        state_vec_410 <= _state_vec_410_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_411 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_411_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_411_valid) begin
        state_vec_411 <= _state_vec_411_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_412 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_412_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_412_valid) begin
        state_vec_412 <= _state_vec_412_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_413 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_413_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_413_valid) begin
        state_vec_413 <= _state_vec_413_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_414 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_414_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_414_valid) begin
        state_vec_414 <= _state_vec_414_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_415 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_415_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_415_valid) begin
        state_vec_415 <= _state_vec_415_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_416 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_416_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_416_valid) begin
        state_vec_416 <= _state_vec_416_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_417 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_417_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_417_valid) begin
        state_vec_417 <= _state_vec_417_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_418 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_418_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_418_valid) begin
        state_vec_418 <= _state_vec_418_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_419 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_419_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_419_valid) begin
        state_vec_419 <= _state_vec_419_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_420 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_420_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_420_valid) begin
        state_vec_420 <= _state_vec_420_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_421 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_421_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_421_valid) begin
        state_vec_421 <= _state_vec_421_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_422 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_422_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_422_valid) begin
        state_vec_422 <= _state_vec_422_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_423 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_423_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_423_valid) begin
        state_vec_423 <= _state_vec_423_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_424 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_424_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_424_valid) begin
        state_vec_424 <= _state_vec_424_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_425 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_425_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_425_valid) begin
        state_vec_425 <= _state_vec_425_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_426 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_426_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_426_valid) begin
        state_vec_426 <= _state_vec_426_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_427 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_427_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_427_valid) begin
        state_vec_427 <= _state_vec_427_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_428 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_428_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_428_valid) begin
        state_vec_428 <= _state_vec_428_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_429 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_429_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_429_valid) begin
        state_vec_429 <= _state_vec_429_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_430 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_430_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_430_valid) begin
        state_vec_430 <= _state_vec_430_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_431 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_431_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_431_valid) begin
        state_vec_431 <= _state_vec_431_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_432 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_432_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_432_valid) begin
        state_vec_432 <= _state_vec_432_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_433 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_433_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_433_valid) begin
        state_vec_433 <= _state_vec_433_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_434 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_434_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_434_valid) begin
        state_vec_434 <= _state_vec_434_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_435 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_435_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_435_valid) begin
        state_vec_435 <= _state_vec_435_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_436 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_436_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_436_valid) begin
        state_vec_436 <= _state_vec_436_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_437 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_437_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_437_valid) begin
        state_vec_437 <= _state_vec_437_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_438 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_438_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_438_valid) begin
        state_vec_438 <= _state_vec_438_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_439 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_439_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_439_valid) begin
        state_vec_439 <= _state_vec_439_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_440 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_440_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_440_valid) begin
        state_vec_440 <= _state_vec_440_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_441 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_441_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_441_valid) begin
        state_vec_441 <= _state_vec_441_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_442 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_442_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_442_valid) begin
        state_vec_442 <= _state_vec_442_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_443 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_443_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_443_valid) begin
        state_vec_443 <= _state_vec_443_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_444 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_444_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_444_valid) begin
        state_vec_444 <= _state_vec_444_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_445 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_445_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_445_valid) begin
        state_vec_445 <= _state_vec_445_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_446 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_446_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_446_valid) begin
        state_vec_446 <= _state_vec_446_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_447 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_447_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_447_valid) begin
        state_vec_447 <= _state_vec_447_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_448 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_448_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_448_valid) begin
        state_vec_448 <= _state_vec_448_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_449 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_449_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_449_valid) begin
        state_vec_449 <= _state_vec_449_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_450 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_450_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_450_valid) begin
        state_vec_450 <= _state_vec_450_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_451 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_451_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_451_valid) begin
        state_vec_451 <= _state_vec_451_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_452 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_452_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_452_valid) begin
        state_vec_452 <= _state_vec_452_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_453 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_453_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_453_valid) begin
        state_vec_453 <= _state_vec_453_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_454 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_454_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_454_valid) begin
        state_vec_454 <= _state_vec_454_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_455 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_455_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_455_valid) begin
        state_vec_455 <= _state_vec_455_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_456 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_456_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_456_valid) begin
        state_vec_456 <= _state_vec_456_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_457 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_457_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_457_valid) begin
        state_vec_457 <= _state_vec_457_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_458 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_458_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_458_valid) begin
        state_vec_458 <= _state_vec_458_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_459 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_459_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_459_valid) begin
        state_vec_459 <= _state_vec_459_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_460 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_460_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_460_valid) begin
        state_vec_460 <= _state_vec_460_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_461 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_461_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_461_valid) begin
        state_vec_461 <= _state_vec_461_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_462 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_462_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_462_valid) begin
        state_vec_462 <= _state_vec_462_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_463 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_463_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_463_valid) begin
        state_vec_463 <= _state_vec_463_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_464 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_464_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_464_valid) begin
        state_vec_464 <= _state_vec_464_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_465 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_465_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_465_valid) begin
        state_vec_465 <= _state_vec_465_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_466 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_466_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_466_valid) begin
        state_vec_466 <= _state_vec_466_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_467 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_467_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_467_valid) begin
        state_vec_467 <= _state_vec_467_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_468 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_468_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_468_valid) begin
        state_vec_468 <= _state_vec_468_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_469 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_469_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_469_valid) begin
        state_vec_469 <= _state_vec_469_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_470 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_470_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_470_valid) begin
        state_vec_470 <= _state_vec_470_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_471 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_471_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_471_valid) begin
        state_vec_471 <= _state_vec_471_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_472 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_472_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_472_valid) begin
        state_vec_472 <= _state_vec_472_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_473 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_473_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_473_valid) begin
        state_vec_473 <= _state_vec_473_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_474 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_474_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_474_valid) begin
        state_vec_474 <= _state_vec_474_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_475 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_475_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_475_valid) begin
        state_vec_475 <= _state_vec_475_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_476 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_476_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_476_valid) begin
        state_vec_476 <= _state_vec_476_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_477 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_477_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_477_valid) begin
        state_vec_477 <= _state_vec_477_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_478 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_478_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_478_valid) begin
        state_vec_478 <= _state_vec_478_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_479 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_479_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_479_valid) begin
        state_vec_479 <= _state_vec_479_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_480 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_480_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_480_valid) begin
        state_vec_480 <= _state_vec_480_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_481 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_481_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_481_valid) begin
        state_vec_481 <= _state_vec_481_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_482 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_482_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_482_valid) begin
        state_vec_482 <= _state_vec_482_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_483 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_483_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_483_valid) begin
        state_vec_483 <= _state_vec_483_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_484 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_484_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_484_valid) begin
        state_vec_484 <= _state_vec_484_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_485 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_485_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_485_valid) begin
        state_vec_485 <= _state_vec_485_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_486 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_486_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_486_valid) begin
        state_vec_486 <= _state_vec_486_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_487 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_487_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_487_valid) begin
        state_vec_487 <= _state_vec_487_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_488 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_488_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_488_valid) begin
        state_vec_488 <= _state_vec_488_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_489 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_489_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_489_valid) begin
        state_vec_489 <= _state_vec_489_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_490 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_490_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_490_valid) begin
        state_vec_490 <= _state_vec_490_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_491 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_491_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_491_valid) begin
        state_vec_491 <= _state_vec_491_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_492 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_492_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_492_valid) begin
        state_vec_492 <= _state_vec_492_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_493 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_493_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_493_valid) begin
        state_vec_493 <= _state_vec_493_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_494 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_494_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_494_valid) begin
        state_vec_494 <= _state_vec_494_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_495 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_495_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_495_valid) begin
        state_vec_495 <= _state_vec_495_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_496 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_496_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_496_valid) begin
        state_vec_496 <= _state_vec_496_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_497 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_497_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_497_valid) begin
        state_vec_497 <= _state_vec_497_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_498 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_498_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_498_valid) begin
        state_vec_498 <= _state_vec_498_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_499 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_499_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_499_valid) begin
        state_vec_499 <= _state_vec_499_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_500 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_500_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_500_valid) begin
        state_vec_500 <= _state_vec_500_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_501 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_501_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_501_valid) begin
        state_vec_501 <= _state_vec_501_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_502 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_502_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_502_valid) begin
        state_vec_502 <= _state_vec_502_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_503 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_503_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_503_valid) begin
        state_vec_503 <= _state_vec_503_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_504 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_504_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_504_valid) begin
        state_vec_504 <= _state_vec_504_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_505 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_505_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_505_valid) begin
        state_vec_505 <= _state_vec_505_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_506 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_506_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_506_valid) begin
        state_vec_506 <= _state_vec_506_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_507 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_507_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_507_valid) begin
        state_vec_507 <= _state_vec_507_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_508 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_508_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_508_valid) begin
        state_vec_508 <= _state_vec_508_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_509 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_509_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_509_valid) begin
        state_vec_509 <= _state_vec_509_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_510 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_510_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_510_valid) begin
        state_vec_510 <= _state_vec_510_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Replacement.scala 316:46]
      state_vec_511 <= 3'h0; // @[Replacement.scala 22:56]
    end else if (set_touch_ways_0_511_valid) begin // @[Replacement.scala 305:17]
      if (set_touch_ways_0_511_valid) begin
        state_vec_511 <= _state_vec_511_T_8;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  pred_rdata_REG = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  pred_rdata_hold_data_0_entry_valid = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  pred_rdata_hold_data_0_entry_brSlots_0_offset = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  pred_rdata_hold_data_0_entry_brSlots_0_lower = _RAND_3[11:0];
  _RAND_4 = {1{`RANDOM}};
  pred_rdata_hold_data_0_entry_brSlots_0_tarStat = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  pred_rdata_hold_data_0_entry_brSlots_0_sharing = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  pred_rdata_hold_data_0_entry_brSlots_0_valid = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  pred_rdata_hold_data_0_entry_tailSlot_offset = _RAND_7[2:0];
  _RAND_8 = {1{`RANDOM}};
  pred_rdata_hold_data_0_entry_tailSlot_lower = _RAND_8[19:0];
  _RAND_9 = {1{`RANDOM}};
  pred_rdata_hold_data_0_entry_tailSlot_tarStat = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  pred_rdata_hold_data_0_entry_tailSlot_sharing = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  pred_rdata_hold_data_0_entry_tailSlot_valid = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  pred_rdata_hold_data_0_entry_pftAddr = _RAND_12[2:0];
  _RAND_13 = {1{`RANDOM}};
  pred_rdata_hold_data_0_entry_carry = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  pred_rdata_hold_data_0_entry_isCall = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  pred_rdata_hold_data_0_entry_isRet = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  pred_rdata_hold_data_0_entry_isJalr = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  pred_rdata_hold_data_0_entry_last_may_be_rvi_call = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  pred_rdata_hold_data_0_entry_always_taken_0 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  pred_rdata_hold_data_0_entry_always_taken_1 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  pred_rdata_hold_data_0_tag = _RAND_20[19:0];
  _RAND_21 = {1{`RANDOM}};
  pred_rdata_hold_data_1_entry_valid = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  pred_rdata_hold_data_1_entry_brSlots_0_offset = _RAND_22[2:0];
  _RAND_23 = {1{`RANDOM}};
  pred_rdata_hold_data_1_entry_brSlots_0_lower = _RAND_23[11:0];
  _RAND_24 = {1{`RANDOM}};
  pred_rdata_hold_data_1_entry_brSlots_0_tarStat = _RAND_24[1:0];
  _RAND_25 = {1{`RANDOM}};
  pred_rdata_hold_data_1_entry_brSlots_0_sharing = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  pred_rdata_hold_data_1_entry_brSlots_0_valid = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  pred_rdata_hold_data_1_entry_tailSlot_offset = _RAND_27[2:0];
  _RAND_28 = {1{`RANDOM}};
  pred_rdata_hold_data_1_entry_tailSlot_lower = _RAND_28[19:0];
  _RAND_29 = {1{`RANDOM}};
  pred_rdata_hold_data_1_entry_tailSlot_tarStat = _RAND_29[1:0];
  _RAND_30 = {1{`RANDOM}};
  pred_rdata_hold_data_1_entry_tailSlot_sharing = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  pred_rdata_hold_data_1_entry_tailSlot_valid = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  pred_rdata_hold_data_1_entry_pftAddr = _RAND_32[2:0];
  _RAND_33 = {1{`RANDOM}};
  pred_rdata_hold_data_1_entry_carry = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  pred_rdata_hold_data_1_entry_isCall = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  pred_rdata_hold_data_1_entry_isRet = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  pred_rdata_hold_data_1_entry_isJalr = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  pred_rdata_hold_data_1_entry_last_may_be_rvi_call = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  pred_rdata_hold_data_1_entry_always_taken_0 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  pred_rdata_hold_data_1_entry_always_taken_1 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  pred_rdata_hold_data_1_tag = _RAND_40[19:0];
  _RAND_41 = {1{`RANDOM}};
  pred_rdata_hold_data_2_entry_valid = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  pred_rdata_hold_data_2_entry_brSlots_0_offset = _RAND_42[2:0];
  _RAND_43 = {1{`RANDOM}};
  pred_rdata_hold_data_2_entry_brSlots_0_lower = _RAND_43[11:0];
  _RAND_44 = {1{`RANDOM}};
  pred_rdata_hold_data_2_entry_brSlots_0_tarStat = _RAND_44[1:0];
  _RAND_45 = {1{`RANDOM}};
  pred_rdata_hold_data_2_entry_brSlots_0_sharing = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  pred_rdata_hold_data_2_entry_brSlots_0_valid = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  pred_rdata_hold_data_2_entry_tailSlot_offset = _RAND_47[2:0];
  _RAND_48 = {1{`RANDOM}};
  pred_rdata_hold_data_2_entry_tailSlot_lower = _RAND_48[19:0];
  _RAND_49 = {1{`RANDOM}};
  pred_rdata_hold_data_2_entry_tailSlot_tarStat = _RAND_49[1:0];
  _RAND_50 = {1{`RANDOM}};
  pred_rdata_hold_data_2_entry_tailSlot_sharing = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  pred_rdata_hold_data_2_entry_tailSlot_valid = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  pred_rdata_hold_data_2_entry_pftAddr = _RAND_52[2:0];
  _RAND_53 = {1{`RANDOM}};
  pred_rdata_hold_data_2_entry_carry = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  pred_rdata_hold_data_2_entry_isCall = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  pred_rdata_hold_data_2_entry_isRet = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  pred_rdata_hold_data_2_entry_isJalr = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  pred_rdata_hold_data_2_entry_last_may_be_rvi_call = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  pred_rdata_hold_data_2_entry_always_taken_0 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  pred_rdata_hold_data_2_entry_always_taken_1 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  pred_rdata_hold_data_2_tag = _RAND_60[19:0];
  _RAND_61 = {1{`RANDOM}};
  pred_rdata_hold_data_3_entry_valid = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  pred_rdata_hold_data_3_entry_brSlots_0_offset = _RAND_62[2:0];
  _RAND_63 = {1{`RANDOM}};
  pred_rdata_hold_data_3_entry_brSlots_0_lower = _RAND_63[11:0];
  _RAND_64 = {1{`RANDOM}};
  pred_rdata_hold_data_3_entry_brSlots_0_tarStat = _RAND_64[1:0];
  _RAND_65 = {1{`RANDOM}};
  pred_rdata_hold_data_3_entry_brSlots_0_sharing = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  pred_rdata_hold_data_3_entry_brSlots_0_valid = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  pred_rdata_hold_data_3_entry_tailSlot_offset = _RAND_67[2:0];
  _RAND_68 = {1{`RANDOM}};
  pred_rdata_hold_data_3_entry_tailSlot_lower = _RAND_68[19:0];
  _RAND_69 = {1{`RANDOM}};
  pred_rdata_hold_data_3_entry_tailSlot_tarStat = _RAND_69[1:0];
  _RAND_70 = {1{`RANDOM}};
  pred_rdata_hold_data_3_entry_tailSlot_sharing = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  pred_rdata_hold_data_3_entry_tailSlot_valid = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  pred_rdata_hold_data_3_entry_pftAddr = _RAND_72[2:0];
  _RAND_73 = {1{`RANDOM}};
  pred_rdata_hold_data_3_entry_carry = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  pred_rdata_hold_data_3_entry_isCall = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  pred_rdata_hold_data_3_entry_isRet = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  pred_rdata_hold_data_3_entry_isJalr = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  pred_rdata_hold_data_3_entry_last_may_be_rvi_call = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  pred_rdata_hold_data_3_entry_always_taken_0 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  pred_rdata_hold_data_3_entry_always_taken_1 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  pred_rdata_hold_data_3_tag = _RAND_80[19:0];
  _RAND_81 = {1{`RANDOM}};
  req_tag = _RAND_81[19:0];
  _RAND_82 = {1{`RANDOM}};
  req_idx = _RAND_82[8:0];
  _RAND_83 = {1{`RANDOM}};
  u_req_tag = _RAND_83[19:0];
  _RAND_84 = {1{`RANDOM}};
  u_total_hits_REG = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  u_total_hits_REG_1 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  u_total_hits_REG_2 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  u_total_hits_REG_3 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  state_vec_0 = _RAND_88[2:0];
  _RAND_89 = {1{`RANDOM}};
  state_vec_1 = _RAND_89[2:0];
  _RAND_90 = {1{`RANDOM}};
  state_vec_2 = _RAND_90[2:0];
  _RAND_91 = {1{`RANDOM}};
  state_vec_3 = _RAND_91[2:0];
  _RAND_92 = {1{`RANDOM}};
  state_vec_4 = _RAND_92[2:0];
  _RAND_93 = {1{`RANDOM}};
  state_vec_5 = _RAND_93[2:0];
  _RAND_94 = {1{`RANDOM}};
  state_vec_6 = _RAND_94[2:0];
  _RAND_95 = {1{`RANDOM}};
  state_vec_7 = _RAND_95[2:0];
  _RAND_96 = {1{`RANDOM}};
  state_vec_8 = _RAND_96[2:0];
  _RAND_97 = {1{`RANDOM}};
  state_vec_9 = _RAND_97[2:0];
  _RAND_98 = {1{`RANDOM}};
  state_vec_10 = _RAND_98[2:0];
  _RAND_99 = {1{`RANDOM}};
  state_vec_11 = _RAND_99[2:0];
  _RAND_100 = {1{`RANDOM}};
  state_vec_12 = _RAND_100[2:0];
  _RAND_101 = {1{`RANDOM}};
  state_vec_13 = _RAND_101[2:0];
  _RAND_102 = {1{`RANDOM}};
  state_vec_14 = _RAND_102[2:0];
  _RAND_103 = {1{`RANDOM}};
  state_vec_15 = _RAND_103[2:0];
  _RAND_104 = {1{`RANDOM}};
  state_vec_16 = _RAND_104[2:0];
  _RAND_105 = {1{`RANDOM}};
  state_vec_17 = _RAND_105[2:0];
  _RAND_106 = {1{`RANDOM}};
  state_vec_18 = _RAND_106[2:0];
  _RAND_107 = {1{`RANDOM}};
  state_vec_19 = _RAND_107[2:0];
  _RAND_108 = {1{`RANDOM}};
  state_vec_20 = _RAND_108[2:0];
  _RAND_109 = {1{`RANDOM}};
  state_vec_21 = _RAND_109[2:0];
  _RAND_110 = {1{`RANDOM}};
  state_vec_22 = _RAND_110[2:0];
  _RAND_111 = {1{`RANDOM}};
  state_vec_23 = _RAND_111[2:0];
  _RAND_112 = {1{`RANDOM}};
  state_vec_24 = _RAND_112[2:0];
  _RAND_113 = {1{`RANDOM}};
  state_vec_25 = _RAND_113[2:0];
  _RAND_114 = {1{`RANDOM}};
  state_vec_26 = _RAND_114[2:0];
  _RAND_115 = {1{`RANDOM}};
  state_vec_27 = _RAND_115[2:0];
  _RAND_116 = {1{`RANDOM}};
  state_vec_28 = _RAND_116[2:0];
  _RAND_117 = {1{`RANDOM}};
  state_vec_29 = _RAND_117[2:0];
  _RAND_118 = {1{`RANDOM}};
  state_vec_30 = _RAND_118[2:0];
  _RAND_119 = {1{`RANDOM}};
  state_vec_31 = _RAND_119[2:0];
  _RAND_120 = {1{`RANDOM}};
  state_vec_32 = _RAND_120[2:0];
  _RAND_121 = {1{`RANDOM}};
  state_vec_33 = _RAND_121[2:0];
  _RAND_122 = {1{`RANDOM}};
  state_vec_34 = _RAND_122[2:0];
  _RAND_123 = {1{`RANDOM}};
  state_vec_35 = _RAND_123[2:0];
  _RAND_124 = {1{`RANDOM}};
  state_vec_36 = _RAND_124[2:0];
  _RAND_125 = {1{`RANDOM}};
  state_vec_37 = _RAND_125[2:0];
  _RAND_126 = {1{`RANDOM}};
  state_vec_38 = _RAND_126[2:0];
  _RAND_127 = {1{`RANDOM}};
  state_vec_39 = _RAND_127[2:0];
  _RAND_128 = {1{`RANDOM}};
  state_vec_40 = _RAND_128[2:0];
  _RAND_129 = {1{`RANDOM}};
  state_vec_41 = _RAND_129[2:0];
  _RAND_130 = {1{`RANDOM}};
  state_vec_42 = _RAND_130[2:0];
  _RAND_131 = {1{`RANDOM}};
  state_vec_43 = _RAND_131[2:0];
  _RAND_132 = {1{`RANDOM}};
  state_vec_44 = _RAND_132[2:0];
  _RAND_133 = {1{`RANDOM}};
  state_vec_45 = _RAND_133[2:0];
  _RAND_134 = {1{`RANDOM}};
  state_vec_46 = _RAND_134[2:0];
  _RAND_135 = {1{`RANDOM}};
  state_vec_47 = _RAND_135[2:0];
  _RAND_136 = {1{`RANDOM}};
  state_vec_48 = _RAND_136[2:0];
  _RAND_137 = {1{`RANDOM}};
  state_vec_49 = _RAND_137[2:0];
  _RAND_138 = {1{`RANDOM}};
  state_vec_50 = _RAND_138[2:0];
  _RAND_139 = {1{`RANDOM}};
  state_vec_51 = _RAND_139[2:0];
  _RAND_140 = {1{`RANDOM}};
  state_vec_52 = _RAND_140[2:0];
  _RAND_141 = {1{`RANDOM}};
  state_vec_53 = _RAND_141[2:0];
  _RAND_142 = {1{`RANDOM}};
  state_vec_54 = _RAND_142[2:0];
  _RAND_143 = {1{`RANDOM}};
  state_vec_55 = _RAND_143[2:0];
  _RAND_144 = {1{`RANDOM}};
  state_vec_56 = _RAND_144[2:0];
  _RAND_145 = {1{`RANDOM}};
  state_vec_57 = _RAND_145[2:0];
  _RAND_146 = {1{`RANDOM}};
  state_vec_58 = _RAND_146[2:0];
  _RAND_147 = {1{`RANDOM}};
  state_vec_59 = _RAND_147[2:0];
  _RAND_148 = {1{`RANDOM}};
  state_vec_60 = _RAND_148[2:0];
  _RAND_149 = {1{`RANDOM}};
  state_vec_61 = _RAND_149[2:0];
  _RAND_150 = {1{`RANDOM}};
  state_vec_62 = _RAND_150[2:0];
  _RAND_151 = {1{`RANDOM}};
  state_vec_63 = _RAND_151[2:0];
  _RAND_152 = {1{`RANDOM}};
  state_vec_64 = _RAND_152[2:0];
  _RAND_153 = {1{`RANDOM}};
  state_vec_65 = _RAND_153[2:0];
  _RAND_154 = {1{`RANDOM}};
  state_vec_66 = _RAND_154[2:0];
  _RAND_155 = {1{`RANDOM}};
  state_vec_67 = _RAND_155[2:0];
  _RAND_156 = {1{`RANDOM}};
  state_vec_68 = _RAND_156[2:0];
  _RAND_157 = {1{`RANDOM}};
  state_vec_69 = _RAND_157[2:0];
  _RAND_158 = {1{`RANDOM}};
  state_vec_70 = _RAND_158[2:0];
  _RAND_159 = {1{`RANDOM}};
  state_vec_71 = _RAND_159[2:0];
  _RAND_160 = {1{`RANDOM}};
  state_vec_72 = _RAND_160[2:0];
  _RAND_161 = {1{`RANDOM}};
  state_vec_73 = _RAND_161[2:0];
  _RAND_162 = {1{`RANDOM}};
  state_vec_74 = _RAND_162[2:0];
  _RAND_163 = {1{`RANDOM}};
  state_vec_75 = _RAND_163[2:0];
  _RAND_164 = {1{`RANDOM}};
  state_vec_76 = _RAND_164[2:0];
  _RAND_165 = {1{`RANDOM}};
  state_vec_77 = _RAND_165[2:0];
  _RAND_166 = {1{`RANDOM}};
  state_vec_78 = _RAND_166[2:0];
  _RAND_167 = {1{`RANDOM}};
  state_vec_79 = _RAND_167[2:0];
  _RAND_168 = {1{`RANDOM}};
  state_vec_80 = _RAND_168[2:0];
  _RAND_169 = {1{`RANDOM}};
  state_vec_81 = _RAND_169[2:0];
  _RAND_170 = {1{`RANDOM}};
  state_vec_82 = _RAND_170[2:0];
  _RAND_171 = {1{`RANDOM}};
  state_vec_83 = _RAND_171[2:0];
  _RAND_172 = {1{`RANDOM}};
  state_vec_84 = _RAND_172[2:0];
  _RAND_173 = {1{`RANDOM}};
  state_vec_85 = _RAND_173[2:0];
  _RAND_174 = {1{`RANDOM}};
  state_vec_86 = _RAND_174[2:0];
  _RAND_175 = {1{`RANDOM}};
  state_vec_87 = _RAND_175[2:0];
  _RAND_176 = {1{`RANDOM}};
  state_vec_88 = _RAND_176[2:0];
  _RAND_177 = {1{`RANDOM}};
  state_vec_89 = _RAND_177[2:0];
  _RAND_178 = {1{`RANDOM}};
  state_vec_90 = _RAND_178[2:0];
  _RAND_179 = {1{`RANDOM}};
  state_vec_91 = _RAND_179[2:0];
  _RAND_180 = {1{`RANDOM}};
  state_vec_92 = _RAND_180[2:0];
  _RAND_181 = {1{`RANDOM}};
  state_vec_93 = _RAND_181[2:0];
  _RAND_182 = {1{`RANDOM}};
  state_vec_94 = _RAND_182[2:0];
  _RAND_183 = {1{`RANDOM}};
  state_vec_95 = _RAND_183[2:0];
  _RAND_184 = {1{`RANDOM}};
  state_vec_96 = _RAND_184[2:0];
  _RAND_185 = {1{`RANDOM}};
  state_vec_97 = _RAND_185[2:0];
  _RAND_186 = {1{`RANDOM}};
  state_vec_98 = _RAND_186[2:0];
  _RAND_187 = {1{`RANDOM}};
  state_vec_99 = _RAND_187[2:0];
  _RAND_188 = {1{`RANDOM}};
  state_vec_100 = _RAND_188[2:0];
  _RAND_189 = {1{`RANDOM}};
  state_vec_101 = _RAND_189[2:0];
  _RAND_190 = {1{`RANDOM}};
  state_vec_102 = _RAND_190[2:0];
  _RAND_191 = {1{`RANDOM}};
  state_vec_103 = _RAND_191[2:0];
  _RAND_192 = {1{`RANDOM}};
  state_vec_104 = _RAND_192[2:0];
  _RAND_193 = {1{`RANDOM}};
  state_vec_105 = _RAND_193[2:0];
  _RAND_194 = {1{`RANDOM}};
  state_vec_106 = _RAND_194[2:0];
  _RAND_195 = {1{`RANDOM}};
  state_vec_107 = _RAND_195[2:0];
  _RAND_196 = {1{`RANDOM}};
  state_vec_108 = _RAND_196[2:0];
  _RAND_197 = {1{`RANDOM}};
  state_vec_109 = _RAND_197[2:0];
  _RAND_198 = {1{`RANDOM}};
  state_vec_110 = _RAND_198[2:0];
  _RAND_199 = {1{`RANDOM}};
  state_vec_111 = _RAND_199[2:0];
  _RAND_200 = {1{`RANDOM}};
  state_vec_112 = _RAND_200[2:0];
  _RAND_201 = {1{`RANDOM}};
  state_vec_113 = _RAND_201[2:0];
  _RAND_202 = {1{`RANDOM}};
  state_vec_114 = _RAND_202[2:0];
  _RAND_203 = {1{`RANDOM}};
  state_vec_115 = _RAND_203[2:0];
  _RAND_204 = {1{`RANDOM}};
  state_vec_116 = _RAND_204[2:0];
  _RAND_205 = {1{`RANDOM}};
  state_vec_117 = _RAND_205[2:0];
  _RAND_206 = {1{`RANDOM}};
  state_vec_118 = _RAND_206[2:0];
  _RAND_207 = {1{`RANDOM}};
  state_vec_119 = _RAND_207[2:0];
  _RAND_208 = {1{`RANDOM}};
  state_vec_120 = _RAND_208[2:0];
  _RAND_209 = {1{`RANDOM}};
  state_vec_121 = _RAND_209[2:0];
  _RAND_210 = {1{`RANDOM}};
  state_vec_122 = _RAND_210[2:0];
  _RAND_211 = {1{`RANDOM}};
  state_vec_123 = _RAND_211[2:0];
  _RAND_212 = {1{`RANDOM}};
  state_vec_124 = _RAND_212[2:0];
  _RAND_213 = {1{`RANDOM}};
  state_vec_125 = _RAND_213[2:0];
  _RAND_214 = {1{`RANDOM}};
  state_vec_126 = _RAND_214[2:0];
  _RAND_215 = {1{`RANDOM}};
  state_vec_127 = _RAND_215[2:0];
  _RAND_216 = {1{`RANDOM}};
  state_vec_128 = _RAND_216[2:0];
  _RAND_217 = {1{`RANDOM}};
  state_vec_129 = _RAND_217[2:0];
  _RAND_218 = {1{`RANDOM}};
  state_vec_130 = _RAND_218[2:0];
  _RAND_219 = {1{`RANDOM}};
  state_vec_131 = _RAND_219[2:0];
  _RAND_220 = {1{`RANDOM}};
  state_vec_132 = _RAND_220[2:0];
  _RAND_221 = {1{`RANDOM}};
  state_vec_133 = _RAND_221[2:0];
  _RAND_222 = {1{`RANDOM}};
  state_vec_134 = _RAND_222[2:0];
  _RAND_223 = {1{`RANDOM}};
  state_vec_135 = _RAND_223[2:0];
  _RAND_224 = {1{`RANDOM}};
  state_vec_136 = _RAND_224[2:0];
  _RAND_225 = {1{`RANDOM}};
  state_vec_137 = _RAND_225[2:0];
  _RAND_226 = {1{`RANDOM}};
  state_vec_138 = _RAND_226[2:0];
  _RAND_227 = {1{`RANDOM}};
  state_vec_139 = _RAND_227[2:0];
  _RAND_228 = {1{`RANDOM}};
  state_vec_140 = _RAND_228[2:0];
  _RAND_229 = {1{`RANDOM}};
  state_vec_141 = _RAND_229[2:0];
  _RAND_230 = {1{`RANDOM}};
  state_vec_142 = _RAND_230[2:0];
  _RAND_231 = {1{`RANDOM}};
  state_vec_143 = _RAND_231[2:0];
  _RAND_232 = {1{`RANDOM}};
  state_vec_144 = _RAND_232[2:0];
  _RAND_233 = {1{`RANDOM}};
  state_vec_145 = _RAND_233[2:0];
  _RAND_234 = {1{`RANDOM}};
  state_vec_146 = _RAND_234[2:0];
  _RAND_235 = {1{`RANDOM}};
  state_vec_147 = _RAND_235[2:0];
  _RAND_236 = {1{`RANDOM}};
  state_vec_148 = _RAND_236[2:0];
  _RAND_237 = {1{`RANDOM}};
  state_vec_149 = _RAND_237[2:0];
  _RAND_238 = {1{`RANDOM}};
  state_vec_150 = _RAND_238[2:0];
  _RAND_239 = {1{`RANDOM}};
  state_vec_151 = _RAND_239[2:0];
  _RAND_240 = {1{`RANDOM}};
  state_vec_152 = _RAND_240[2:0];
  _RAND_241 = {1{`RANDOM}};
  state_vec_153 = _RAND_241[2:0];
  _RAND_242 = {1{`RANDOM}};
  state_vec_154 = _RAND_242[2:0];
  _RAND_243 = {1{`RANDOM}};
  state_vec_155 = _RAND_243[2:0];
  _RAND_244 = {1{`RANDOM}};
  state_vec_156 = _RAND_244[2:0];
  _RAND_245 = {1{`RANDOM}};
  state_vec_157 = _RAND_245[2:0];
  _RAND_246 = {1{`RANDOM}};
  state_vec_158 = _RAND_246[2:0];
  _RAND_247 = {1{`RANDOM}};
  state_vec_159 = _RAND_247[2:0];
  _RAND_248 = {1{`RANDOM}};
  state_vec_160 = _RAND_248[2:0];
  _RAND_249 = {1{`RANDOM}};
  state_vec_161 = _RAND_249[2:0];
  _RAND_250 = {1{`RANDOM}};
  state_vec_162 = _RAND_250[2:0];
  _RAND_251 = {1{`RANDOM}};
  state_vec_163 = _RAND_251[2:0];
  _RAND_252 = {1{`RANDOM}};
  state_vec_164 = _RAND_252[2:0];
  _RAND_253 = {1{`RANDOM}};
  state_vec_165 = _RAND_253[2:0];
  _RAND_254 = {1{`RANDOM}};
  state_vec_166 = _RAND_254[2:0];
  _RAND_255 = {1{`RANDOM}};
  state_vec_167 = _RAND_255[2:0];
  _RAND_256 = {1{`RANDOM}};
  state_vec_168 = _RAND_256[2:0];
  _RAND_257 = {1{`RANDOM}};
  state_vec_169 = _RAND_257[2:0];
  _RAND_258 = {1{`RANDOM}};
  state_vec_170 = _RAND_258[2:0];
  _RAND_259 = {1{`RANDOM}};
  state_vec_171 = _RAND_259[2:0];
  _RAND_260 = {1{`RANDOM}};
  state_vec_172 = _RAND_260[2:0];
  _RAND_261 = {1{`RANDOM}};
  state_vec_173 = _RAND_261[2:0];
  _RAND_262 = {1{`RANDOM}};
  state_vec_174 = _RAND_262[2:0];
  _RAND_263 = {1{`RANDOM}};
  state_vec_175 = _RAND_263[2:0];
  _RAND_264 = {1{`RANDOM}};
  state_vec_176 = _RAND_264[2:0];
  _RAND_265 = {1{`RANDOM}};
  state_vec_177 = _RAND_265[2:0];
  _RAND_266 = {1{`RANDOM}};
  state_vec_178 = _RAND_266[2:0];
  _RAND_267 = {1{`RANDOM}};
  state_vec_179 = _RAND_267[2:0];
  _RAND_268 = {1{`RANDOM}};
  state_vec_180 = _RAND_268[2:0];
  _RAND_269 = {1{`RANDOM}};
  state_vec_181 = _RAND_269[2:0];
  _RAND_270 = {1{`RANDOM}};
  state_vec_182 = _RAND_270[2:0];
  _RAND_271 = {1{`RANDOM}};
  state_vec_183 = _RAND_271[2:0];
  _RAND_272 = {1{`RANDOM}};
  state_vec_184 = _RAND_272[2:0];
  _RAND_273 = {1{`RANDOM}};
  state_vec_185 = _RAND_273[2:0];
  _RAND_274 = {1{`RANDOM}};
  state_vec_186 = _RAND_274[2:0];
  _RAND_275 = {1{`RANDOM}};
  state_vec_187 = _RAND_275[2:0];
  _RAND_276 = {1{`RANDOM}};
  state_vec_188 = _RAND_276[2:0];
  _RAND_277 = {1{`RANDOM}};
  state_vec_189 = _RAND_277[2:0];
  _RAND_278 = {1{`RANDOM}};
  state_vec_190 = _RAND_278[2:0];
  _RAND_279 = {1{`RANDOM}};
  state_vec_191 = _RAND_279[2:0];
  _RAND_280 = {1{`RANDOM}};
  state_vec_192 = _RAND_280[2:0];
  _RAND_281 = {1{`RANDOM}};
  state_vec_193 = _RAND_281[2:0];
  _RAND_282 = {1{`RANDOM}};
  state_vec_194 = _RAND_282[2:0];
  _RAND_283 = {1{`RANDOM}};
  state_vec_195 = _RAND_283[2:0];
  _RAND_284 = {1{`RANDOM}};
  state_vec_196 = _RAND_284[2:0];
  _RAND_285 = {1{`RANDOM}};
  state_vec_197 = _RAND_285[2:0];
  _RAND_286 = {1{`RANDOM}};
  state_vec_198 = _RAND_286[2:0];
  _RAND_287 = {1{`RANDOM}};
  state_vec_199 = _RAND_287[2:0];
  _RAND_288 = {1{`RANDOM}};
  state_vec_200 = _RAND_288[2:0];
  _RAND_289 = {1{`RANDOM}};
  state_vec_201 = _RAND_289[2:0];
  _RAND_290 = {1{`RANDOM}};
  state_vec_202 = _RAND_290[2:0];
  _RAND_291 = {1{`RANDOM}};
  state_vec_203 = _RAND_291[2:0];
  _RAND_292 = {1{`RANDOM}};
  state_vec_204 = _RAND_292[2:0];
  _RAND_293 = {1{`RANDOM}};
  state_vec_205 = _RAND_293[2:0];
  _RAND_294 = {1{`RANDOM}};
  state_vec_206 = _RAND_294[2:0];
  _RAND_295 = {1{`RANDOM}};
  state_vec_207 = _RAND_295[2:0];
  _RAND_296 = {1{`RANDOM}};
  state_vec_208 = _RAND_296[2:0];
  _RAND_297 = {1{`RANDOM}};
  state_vec_209 = _RAND_297[2:0];
  _RAND_298 = {1{`RANDOM}};
  state_vec_210 = _RAND_298[2:0];
  _RAND_299 = {1{`RANDOM}};
  state_vec_211 = _RAND_299[2:0];
  _RAND_300 = {1{`RANDOM}};
  state_vec_212 = _RAND_300[2:0];
  _RAND_301 = {1{`RANDOM}};
  state_vec_213 = _RAND_301[2:0];
  _RAND_302 = {1{`RANDOM}};
  state_vec_214 = _RAND_302[2:0];
  _RAND_303 = {1{`RANDOM}};
  state_vec_215 = _RAND_303[2:0];
  _RAND_304 = {1{`RANDOM}};
  state_vec_216 = _RAND_304[2:0];
  _RAND_305 = {1{`RANDOM}};
  state_vec_217 = _RAND_305[2:0];
  _RAND_306 = {1{`RANDOM}};
  state_vec_218 = _RAND_306[2:0];
  _RAND_307 = {1{`RANDOM}};
  state_vec_219 = _RAND_307[2:0];
  _RAND_308 = {1{`RANDOM}};
  state_vec_220 = _RAND_308[2:0];
  _RAND_309 = {1{`RANDOM}};
  state_vec_221 = _RAND_309[2:0];
  _RAND_310 = {1{`RANDOM}};
  state_vec_222 = _RAND_310[2:0];
  _RAND_311 = {1{`RANDOM}};
  state_vec_223 = _RAND_311[2:0];
  _RAND_312 = {1{`RANDOM}};
  state_vec_224 = _RAND_312[2:0];
  _RAND_313 = {1{`RANDOM}};
  state_vec_225 = _RAND_313[2:0];
  _RAND_314 = {1{`RANDOM}};
  state_vec_226 = _RAND_314[2:0];
  _RAND_315 = {1{`RANDOM}};
  state_vec_227 = _RAND_315[2:0];
  _RAND_316 = {1{`RANDOM}};
  state_vec_228 = _RAND_316[2:0];
  _RAND_317 = {1{`RANDOM}};
  state_vec_229 = _RAND_317[2:0];
  _RAND_318 = {1{`RANDOM}};
  state_vec_230 = _RAND_318[2:0];
  _RAND_319 = {1{`RANDOM}};
  state_vec_231 = _RAND_319[2:0];
  _RAND_320 = {1{`RANDOM}};
  state_vec_232 = _RAND_320[2:0];
  _RAND_321 = {1{`RANDOM}};
  state_vec_233 = _RAND_321[2:0];
  _RAND_322 = {1{`RANDOM}};
  state_vec_234 = _RAND_322[2:0];
  _RAND_323 = {1{`RANDOM}};
  state_vec_235 = _RAND_323[2:0];
  _RAND_324 = {1{`RANDOM}};
  state_vec_236 = _RAND_324[2:0];
  _RAND_325 = {1{`RANDOM}};
  state_vec_237 = _RAND_325[2:0];
  _RAND_326 = {1{`RANDOM}};
  state_vec_238 = _RAND_326[2:0];
  _RAND_327 = {1{`RANDOM}};
  state_vec_239 = _RAND_327[2:0];
  _RAND_328 = {1{`RANDOM}};
  state_vec_240 = _RAND_328[2:0];
  _RAND_329 = {1{`RANDOM}};
  state_vec_241 = _RAND_329[2:0];
  _RAND_330 = {1{`RANDOM}};
  state_vec_242 = _RAND_330[2:0];
  _RAND_331 = {1{`RANDOM}};
  state_vec_243 = _RAND_331[2:0];
  _RAND_332 = {1{`RANDOM}};
  state_vec_244 = _RAND_332[2:0];
  _RAND_333 = {1{`RANDOM}};
  state_vec_245 = _RAND_333[2:0];
  _RAND_334 = {1{`RANDOM}};
  state_vec_246 = _RAND_334[2:0];
  _RAND_335 = {1{`RANDOM}};
  state_vec_247 = _RAND_335[2:0];
  _RAND_336 = {1{`RANDOM}};
  state_vec_248 = _RAND_336[2:0];
  _RAND_337 = {1{`RANDOM}};
  state_vec_249 = _RAND_337[2:0];
  _RAND_338 = {1{`RANDOM}};
  state_vec_250 = _RAND_338[2:0];
  _RAND_339 = {1{`RANDOM}};
  state_vec_251 = _RAND_339[2:0];
  _RAND_340 = {1{`RANDOM}};
  state_vec_252 = _RAND_340[2:0];
  _RAND_341 = {1{`RANDOM}};
  state_vec_253 = _RAND_341[2:0];
  _RAND_342 = {1{`RANDOM}};
  state_vec_254 = _RAND_342[2:0];
  _RAND_343 = {1{`RANDOM}};
  state_vec_255 = _RAND_343[2:0];
  _RAND_344 = {1{`RANDOM}};
  state_vec_256 = _RAND_344[2:0];
  _RAND_345 = {1{`RANDOM}};
  state_vec_257 = _RAND_345[2:0];
  _RAND_346 = {1{`RANDOM}};
  state_vec_258 = _RAND_346[2:0];
  _RAND_347 = {1{`RANDOM}};
  state_vec_259 = _RAND_347[2:0];
  _RAND_348 = {1{`RANDOM}};
  state_vec_260 = _RAND_348[2:0];
  _RAND_349 = {1{`RANDOM}};
  state_vec_261 = _RAND_349[2:0];
  _RAND_350 = {1{`RANDOM}};
  state_vec_262 = _RAND_350[2:0];
  _RAND_351 = {1{`RANDOM}};
  state_vec_263 = _RAND_351[2:0];
  _RAND_352 = {1{`RANDOM}};
  state_vec_264 = _RAND_352[2:0];
  _RAND_353 = {1{`RANDOM}};
  state_vec_265 = _RAND_353[2:0];
  _RAND_354 = {1{`RANDOM}};
  state_vec_266 = _RAND_354[2:0];
  _RAND_355 = {1{`RANDOM}};
  state_vec_267 = _RAND_355[2:0];
  _RAND_356 = {1{`RANDOM}};
  state_vec_268 = _RAND_356[2:0];
  _RAND_357 = {1{`RANDOM}};
  state_vec_269 = _RAND_357[2:0];
  _RAND_358 = {1{`RANDOM}};
  state_vec_270 = _RAND_358[2:0];
  _RAND_359 = {1{`RANDOM}};
  state_vec_271 = _RAND_359[2:0];
  _RAND_360 = {1{`RANDOM}};
  state_vec_272 = _RAND_360[2:0];
  _RAND_361 = {1{`RANDOM}};
  state_vec_273 = _RAND_361[2:0];
  _RAND_362 = {1{`RANDOM}};
  state_vec_274 = _RAND_362[2:0];
  _RAND_363 = {1{`RANDOM}};
  state_vec_275 = _RAND_363[2:0];
  _RAND_364 = {1{`RANDOM}};
  state_vec_276 = _RAND_364[2:0];
  _RAND_365 = {1{`RANDOM}};
  state_vec_277 = _RAND_365[2:0];
  _RAND_366 = {1{`RANDOM}};
  state_vec_278 = _RAND_366[2:0];
  _RAND_367 = {1{`RANDOM}};
  state_vec_279 = _RAND_367[2:0];
  _RAND_368 = {1{`RANDOM}};
  state_vec_280 = _RAND_368[2:0];
  _RAND_369 = {1{`RANDOM}};
  state_vec_281 = _RAND_369[2:0];
  _RAND_370 = {1{`RANDOM}};
  state_vec_282 = _RAND_370[2:0];
  _RAND_371 = {1{`RANDOM}};
  state_vec_283 = _RAND_371[2:0];
  _RAND_372 = {1{`RANDOM}};
  state_vec_284 = _RAND_372[2:0];
  _RAND_373 = {1{`RANDOM}};
  state_vec_285 = _RAND_373[2:0];
  _RAND_374 = {1{`RANDOM}};
  state_vec_286 = _RAND_374[2:0];
  _RAND_375 = {1{`RANDOM}};
  state_vec_287 = _RAND_375[2:0];
  _RAND_376 = {1{`RANDOM}};
  state_vec_288 = _RAND_376[2:0];
  _RAND_377 = {1{`RANDOM}};
  state_vec_289 = _RAND_377[2:0];
  _RAND_378 = {1{`RANDOM}};
  state_vec_290 = _RAND_378[2:0];
  _RAND_379 = {1{`RANDOM}};
  state_vec_291 = _RAND_379[2:0];
  _RAND_380 = {1{`RANDOM}};
  state_vec_292 = _RAND_380[2:0];
  _RAND_381 = {1{`RANDOM}};
  state_vec_293 = _RAND_381[2:0];
  _RAND_382 = {1{`RANDOM}};
  state_vec_294 = _RAND_382[2:0];
  _RAND_383 = {1{`RANDOM}};
  state_vec_295 = _RAND_383[2:0];
  _RAND_384 = {1{`RANDOM}};
  state_vec_296 = _RAND_384[2:0];
  _RAND_385 = {1{`RANDOM}};
  state_vec_297 = _RAND_385[2:0];
  _RAND_386 = {1{`RANDOM}};
  state_vec_298 = _RAND_386[2:0];
  _RAND_387 = {1{`RANDOM}};
  state_vec_299 = _RAND_387[2:0];
  _RAND_388 = {1{`RANDOM}};
  state_vec_300 = _RAND_388[2:0];
  _RAND_389 = {1{`RANDOM}};
  state_vec_301 = _RAND_389[2:0];
  _RAND_390 = {1{`RANDOM}};
  state_vec_302 = _RAND_390[2:0];
  _RAND_391 = {1{`RANDOM}};
  state_vec_303 = _RAND_391[2:0];
  _RAND_392 = {1{`RANDOM}};
  state_vec_304 = _RAND_392[2:0];
  _RAND_393 = {1{`RANDOM}};
  state_vec_305 = _RAND_393[2:0];
  _RAND_394 = {1{`RANDOM}};
  state_vec_306 = _RAND_394[2:0];
  _RAND_395 = {1{`RANDOM}};
  state_vec_307 = _RAND_395[2:0];
  _RAND_396 = {1{`RANDOM}};
  state_vec_308 = _RAND_396[2:0];
  _RAND_397 = {1{`RANDOM}};
  state_vec_309 = _RAND_397[2:0];
  _RAND_398 = {1{`RANDOM}};
  state_vec_310 = _RAND_398[2:0];
  _RAND_399 = {1{`RANDOM}};
  state_vec_311 = _RAND_399[2:0];
  _RAND_400 = {1{`RANDOM}};
  state_vec_312 = _RAND_400[2:0];
  _RAND_401 = {1{`RANDOM}};
  state_vec_313 = _RAND_401[2:0];
  _RAND_402 = {1{`RANDOM}};
  state_vec_314 = _RAND_402[2:0];
  _RAND_403 = {1{`RANDOM}};
  state_vec_315 = _RAND_403[2:0];
  _RAND_404 = {1{`RANDOM}};
  state_vec_316 = _RAND_404[2:0];
  _RAND_405 = {1{`RANDOM}};
  state_vec_317 = _RAND_405[2:0];
  _RAND_406 = {1{`RANDOM}};
  state_vec_318 = _RAND_406[2:0];
  _RAND_407 = {1{`RANDOM}};
  state_vec_319 = _RAND_407[2:0];
  _RAND_408 = {1{`RANDOM}};
  state_vec_320 = _RAND_408[2:0];
  _RAND_409 = {1{`RANDOM}};
  state_vec_321 = _RAND_409[2:0];
  _RAND_410 = {1{`RANDOM}};
  state_vec_322 = _RAND_410[2:0];
  _RAND_411 = {1{`RANDOM}};
  state_vec_323 = _RAND_411[2:0];
  _RAND_412 = {1{`RANDOM}};
  state_vec_324 = _RAND_412[2:0];
  _RAND_413 = {1{`RANDOM}};
  state_vec_325 = _RAND_413[2:0];
  _RAND_414 = {1{`RANDOM}};
  state_vec_326 = _RAND_414[2:0];
  _RAND_415 = {1{`RANDOM}};
  state_vec_327 = _RAND_415[2:0];
  _RAND_416 = {1{`RANDOM}};
  state_vec_328 = _RAND_416[2:0];
  _RAND_417 = {1{`RANDOM}};
  state_vec_329 = _RAND_417[2:0];
  _RAND_418 = {1{`RANDOM}};
  state_vec_330 = _RAND_418[2:0];
  _RAND_419 = {1{`RANDOM}};
  state_vec_331 = _RAND_419[2:0];
  _RAND_420 = {1{`RANDOM}};
  state_vec_332 = _RAND_420[2:0];
  _RAND_421 = {1{`RANDOM}};
  state_vec_333 = _RAND_421[2:0];
  _RAND_422 = {1{`RANDOM}};
  state_vec_334 = _RAND_422[2:0];
  _RAND_423 = {1{`RANDOM}};
  state_vec_335 = _RAND_423[2:0];
  _RAND_424 = {1{`RANDOM}};
  state_vec_336 = _RAND_424[2:0];
  _RAND_425 = {1{`RANDOM}};
  state_vec_337 = _RAND_425[2:0];
  _RAND_426 = {1{`RANDOM}};
  state_vec_338 = _RAND_426[2:0];
  _RAND_427 = {1{`RANDOM}};
  state_vec_339 = _RAND_427[2:0];
  _RAND_428 = {1{`RANDOM}};
  state_vec_340 = _RAND_428[2:0];
  _RAND_429 = {1{`RANDOM}};
  state_vec_341 = _RAND_429[2:0];
  _RAND_430 = {1{`RANDOM}};
  state_vec_342 = _RAND_430[2:0];
  _RAND_431 = {1{`RANDOM}};
  state_vec_343 = _RAND_431[2:0];
  _RAND_432 = {1{`RANDOM}};
  state_vec_344 = _RAND_432[2:0];
  _RAND_433 = {1{`RANDOM}};
  state_vec_345 = _RAND_433[2:0];
  _RAND_434 = {1{`RANDOM}};
  state_vec_346 = _RAND_434[2:0];
  _RAND_435 = {1{`RANDOM}};
  state_vec_347 = _RAND_435[2:0];
  _RAND_436 = {1{`RANDOM}};
  state_vec_348 = _RAND_436[2:0];
  _RAND_437 = {1{`RANDOM}};
  state_vec_349 = _RAND_437[2:0];
  _RAND_438 = {1{`RANDOM}};
  state_vec_350 = _RAND_438[2:0];
  _RAND_439 = {1{`RANDOM}};
  state_vec_351 = _RAND_439[2:0];
  _RAND_440 = {1{`RANDOM}};
  state_vec_352 = _RAND_440[2:0];
  _RAND_441 = {1{`RANDOM}};
  state_vec_353 = _RAND_441[2:0];
  _RAND_442 = {1{`RANDOM}};
  state_vec_354 = _RAND_442[2:0];
  _RAND_443 = {1{`RANDOM}};
  state_vec_355 = _RAND_443[2:0];
  _RAND_444 = {1{`RANDOM}};
  state_vec_356 = _RAND_444[2:0];
  _RAND_445 = {1{`RANDOM}};
  state_vec_357 = _RAND_445[2:0];
  _RAND_446 = {1{`RANDOM}};
  state_vec_358 = _RAND_446[2:0];
  _RAND_447 = {1{`RANDOM}};
  state_vec_359 = _RAND_447[2:0];
  _RAND_448 = {1{`RANDOM}};
  state_vec_360 = _RAND_448[2:0];
  _RAND_449 = {1{`RANDOM}};
  state_vec_361 = _RAND_449[2:0];
  _RAND_450 = {1{`RANDOM}};
  state_vec_362 = _RAND_450[2:0];
  _RAND_451 = {1{`RANDOM}};
  state_vec_363 = _RAND_451[2:0];
  _RAND_452 = {1{`RANDOM}};
  state_vec_364 = _RAND_452[2:0];
  _RAND_453 = {1{`RANDOM}};
  state_vec_365 = _RAND_453[2:0];
  _RAND_454 = {1{`RANDOM}};
  state_vec_366 = _RAND_454[2:0];
  _RAND_455 = {1{`RANDOM}};
  state_vec_367 = _RAND_455[2:0];
  _RAND_456 = {1{`RANDOM}};
  state_vec_368 = _RAND_456[2:0];
  _RAND_457 = {1{`RANDOM}};
  state_vec_369 = _RAND_457[2:0];
  _RAND_458 = {1{`RANDOM}};
  state_vec_370 = _RAND_458[2:0];
  _RAND_459 = {1{`RANDOM}};
  state_vec_371 = _RAND_459[2:0];
  _RAND_460 = {1{`RANDOM}};
  state_vec_372 = _RAND_460[2:0];
  _RAND_461 = {1{`RANDOM}};
  state_vec_373 = _RAND_461[2:0];
  _RAND_462 = {1{`RANDOM}};
  state_vec_374 = _RAND_462[2:0];
  _RAND_463 = {1{`RANDOM}};
  state_vec_375 = _RAND_463[2:0];
  _RAND_464 = {1{`RANDOM}};
  state_vec_376 = _RAND_464[2:0];
  _RAND_465 = {1{`RANDOM}};
  state_vec_377 = _RAND_465[2:0];
  _RAND_466 = {1{`RANDOM}};
  state_vec_378 = _RAND_466[2:0];
  _RAND_467 = {1{`RANDOM}};
  state_vec_379 = _RAND_467[2:0];
  _RAND_468 = {1{`RANDOM}};
  state_vec_380 = _RAND_468[2:0];
  _RAND_469 = {1{`RANDOM}};
  state_vec_381 = _RAND_469[2:0];
  _RAND_470 = {1{`RANDOM}};
  state_vec_382 = _RAND_470[2:0];
  _RAND_471 = {1{`RANDOM}};
  state_vec_383 = _RAND_471[2:0];
  _RAND_472 = {1{`RANDOM}};
  state_vec_384 = _RAND_472[2:0];
  _RAND_473 = {1{`RANDOM}};
  state_vec_385 = _RAND_473[2:0];
  _RAND_474 = {1{`RANDOM}};
  state_vec_386 = _RAND_474[2:0];
  _RAND_475 = {1{`RANDOM}};
  state_vec_387 = _RAND_475[2:0];
  _RAND_476 = {1{`RANDOM}};
  state_vec_388 = _RAND_476[2:0];
  _RAND_477 = {1{`RANDOM}};
  state_vec_389 = _RAND_477[2:0];
  _RAND_478 = {1{`RANDOM}};
  state_vec_390 = _RAND_478[2:0];
  _RAND_479 = {1{`RANDOM}};
  state_vec_391 = _RAND_479[2:0];
  _RAND_480 = {1{`RANDOM}};
  state_vec_392 = _RAND_480[2:0];
  _RAND_481 = {1{`RANDOM}};
  state_vec_393 = _RAND_481[2:0];
  _RAND_482 = {1{`RANDOM}};
  state_vec_394 = _RAND_482[2:0];
  _RAND_483 = {1{`RANDOM}};
  state_vec_395 = _RAND_483[2:0];
  _RAND_484 = {1{`RANDOM}};
  state_vec_396 = _RAND_484[2:0];
  _RAND_485 = {1{`RANDOM}};
  state_vec_397 = _RAND_485[2:0];
  _RAND_486 = {1{`RANDOM}};
  state_vec_398 = _RAND_486[2:0];
  _RAND_487 = {1{`RANDOM}};
  state_vec_399 = _RAND_487[2:0];
  _RAND_488 = {1{`RANDOM}};
  state_vec_400 = _RAND_488[2:0];
  _RAND_489 = {1{`RANDOM}};
  state_vec_401 = _RAND_489[2:0];
  _RAND_490 = {1{`RANDOM}};
  state_vec_402 = _RAND_490[2:0];
  _RAND_491 = {1{`RANDOM}};
  state_vec_403 = _RAND_491[2:0];
  _RAND_492 = {1{`RANDOM}};
  state_vec_404 = _RAND_492[2:0];
  _RAND_493 = {1{`RANDOM}};
  state_vec_405 = _RAND_493[2:0];
  _RAND_494 = {1{`RANDOM}};
  state_vec_406 = _RAND_494[2:0];
  _RAND_495 = {1{`RANDOM}};
  state_vec_407 = _RAND_495[2:0];
  _RAND_496 = {1{`RANDOM}};
  state_vec_408 = _RAND_496[2:0];
  _RAND_497 = {1{`RANDOM}};
  state_vec_409 = _RAND_497[2:0];
  _RAND_498 = {1{`RANDOM}};
  state_vec_410 = _RAND_498[2:0];
  _RAND_499 = {1{`RANDOM}};
  state_vec_411 = _RAND_499[2:0];
  _RAND_500 = {1{`RANDOM}};
  state_vec_412 = _RAND_500[2:0];
  _RAND_501 = {1{`RANDOM}};
  state_vec_413 = _RAND_501[2:0];
  _RAND_502 = {1{`RANDOM}};
  state_vec_414 = _RAND_502[2:0];
  _RAND_503 = {1{`RANDOM}};
  state_vec_415 = _RAND_503[2:0];
  _RAND_504 = {1{`RANDOM}};
  state_vec_416 = _RAND_504[2:0];
  _RAND_505 = {1{`RANDOM}};
  state_vec_417 = _RAND_505[2:0];
  _RAND_506 = {1{`RANDOM}};
  state_vec_418 = _RAND_506[2:0];
  _RAND_507 = {1{`RANDOM}};
  state_vec_419 = _RAND_507[2:0];
  _RAND_508 = {1{`RANDOM}};
  state_vec_420 = _RAND_508[2:0];
  _RAND_509 = {1{`RANDOM}};
  state_vec_421 = _RAND_509[2:0];
  _RAND_510 = {1{`RANDOM}};
  state_vec_422 = _RAND_510[2:0];
  _RAND_511 = {1{`RANDOM}};
  state_vec_423 = _RAND_511[2:0];
  _RAND_512 = {1{`RANDOM}};
  state_vec_424 = _RAND_512[2:0];
  _RAND_513 = {1{`RANDOM}};
  state_vec_425 = _RAND_513[2:0];
  _RAND_514 = {1{`RANDOM}};
  state_vec_426 = _RAND_514[2:0];
  _RAND_515 = {1{`RANDOM}};
  state_vec_427 = _RAND_515[2:0];
  _RAND_516 = {1{`RANDOM}};
  state_vec_428 = _RAND_516[2:0];
  _RAND_517 = {1{`RANDOM}};
  state_vec_429 = _RAND_517[2:0];
  _RAND_518 = {1{`RANDOM}};
  state_vec_430 = _RAND_518[2:0];
  _RAND_519 = {1{`RANDOM}};
  state_vec_431 = _RAND_519[2:0];
  _RAND_520 = {1{`RANDOM}};
  state_vec_432 = _RAND_520[2:0];
  _RAND_521 = {1{`RANDOM}};
  state_vec_433 = _RAND_521[2:0];
  _RAND_522 = {1{`RANDOM}};
  state_vec_434 = _RAND_522[2:0];
  _RAND_523 = {1{`RANDOM}};
  state_vec_435 = _RAND_523[2:0];
  _RAND_524 = {1{`RANDOM}};
  state_vec_436 = _RAND_524[2:0];
  _RAND_525 = {1{`RANDOM}};
  state_vec_437 = _RAND_525[2:0];
  _RAND_526 = {1{`RANDOM}};
  state_vec_438 = _RAND_526[2:0];
  _RAND_527 = {1{`RANDOM}};
  state_vec_439 = _RAND_527[2:0];
  _RAND_528 = {1{`RANDOM}};
  state_vec_440 = _RAND_528[2:0];
  _RAND_529 = {1{`RANDOM}};
  state_vec_441 = _RAND_529[2:0];
  _RAND_530 = {1{`RANDOM}};
  state_vec_442 = _RAND_530[2:0];
  _RAND_531 = {1{`RANDOM}};
  state_vec_443 = _RAND_531[2:0];
  _RAND_532 = {1{`RANDOM}};
  state_vec_444 = _RAND_532[2:0];
  _RAND_533 = {1{`RANDOM}};
  state_vec_445 = _RAND_533[2:0];
  _RAND_534 = {1{`RANDOM}};
  state_vec_446 = _RAND_534[2:0];
  _RAND_535 = {1{`RANDOM}};
  state_vec_447 = _RAND_535[2:0];
  _RAND_536 = {1{`RANDOM}};
  state_vec_448 = _RAND_536[2:0];
  _RAND_537 = {1{`RANDOM}};
  state_vec_449 = _RAND_537[2:0];
  _RAND_538 = {1{`RANDOM}};
  state_vec_450 = _RAND_538[2:0];
  _RAND_539 = {1{`RANDOM}};
  state_vec_451 = _RAND_539[2:0];
  _RAND_540 = {1{`RANDOM}};
  state_vec_452 = _RAND_540[2:0];
  _RAND_541 = {1{`RANDOM}};
  state_vec_453 = _RAND_541[2:0];
  _RAND_542 = {1{`RANDOM}};
  state_vec_454 = _RAND_542[2:0];
  _RAND_543 = {1{`RANDOM}};
  state_vec_455 = _RAND_543[2:0];
  _RAND_544 = {1{`RANDOM}};
  state_vec_456 = _RAND_544[2:0];
  _RAND_545 = {1{`RANDOM}};
  state_vec_457 = _RAND_545[2:0];
  _RAND_546 = {1{`RANDOM}};
  state_vec_458 = _RAND_546[2:0];
  _RAND_547 = {1{`RANDOM}};
  state_vec_459 = _RAND_547[2:0];
  _RAND_548 = {1{`RANDOM}};
  state_vec_460 = _RAND_548[2:0];
  _RAND_549 = {1{`RANDOM}};
  state_vec_461 = _RAND_549[2:0];
  _RAND_550 = {1{`RANDOM}};
  state_vec_462 = _RAND_550[2:0];
  _RAND_551 = {1{`RANDOM}};
  state_vec_463 = _RAND_551[2:0];
  _RAND_552 = {1{`RANDOM}};
  state_vec_464 = _RAND_552[2:0];
  _RAND_553 = {1{`RANDOM}};
  state_vec_465 = _RAND_553[2:0];
  _RAND_554 = {1{`RANDOM}};
  state_vec_466 = _RAND_554[2:0];
  _RAND_555 = {1{`RANDOM}};
  state_vec_467 = _RAND_555[2:0];
  _RAND_556 = {1{`RANDOM}};
  state_vec_468 = _RAND_556[2:0];
  _RAND_557 = {1{`RANDOM}};
  state_vec_469 = _RAND_557[2:0];
  _RAND_558 = {1{`RANDOM}};
  state_vec_470 = _RAND_558[2:0];
  _RAND_559 = {1{`RANDOM}};
  state_vec_471 = _RAND_559[2:0];
  _RAND_560 = {1{`RANDOM}};
  state_vec_472 = _RAND_560[2:0];
  _RAND_561 = {1{`RANDOM}};
  state_vec_473 = _RAND_561[2:0];
  _RAND_562 = {1{`RANDOM}};
  state_vec_474 = _RAND_562[2:0];
  _RAND_563 = {1{`RANDOM}};
  state_vec_475 = _RAND_563[2:0];
  _RAND_564 = {1{`RANDOM}};
  state_vec_476 = _RAND_564[2:0];
  _RAND_565 = {1{`RANDOM}};
  state_vec_477 = _RAND_565[2:0];
  _RAND_566 = {1{`RANDOM}};
  state_vec_478 = _RAND_566[2:0];
  _RAND_567 = {1{`RANDOM}};
  state_vec_479 = _RAND_567[2:0];
  _RAND_568 = {1{`RANDOM}};
  state_vec_480 = _RAND_568[2:0];
  _RAND_569 = {1{`RANDOM}};
  state_vec_481 = _RAND_569[2:0];
  _RAND_570 = {1{`RANDOM}};
  state_vec_482 = _RAND_570[2:0];
  _RAND_571 = {1{`RANDOM}};
  state_vec_483 = _RAND_571[2:0];
  _RAND_572 = {1{`RANDOM}};
  state_vec_484 = _RAND_572[2:0];
  _RAND_573 = {1{`RANDOM}};
  state_vec_485 = _RAND_573[2:0];
  _RAND_574 = {1{`RANDOM}};
  state_vec_486 = _RAND_574[2:0];
  _RAND_575 = {1{`RANDOM}};
  state_vec_487 = _RAND_575[2:0];
  _RAND_576 = {1{`RANDOM}};
  state_vec_488 = _RAND_576[2:0];
  _RAND_577 = {1{`RANDOM}};
  state_vec_489 = _RAND_577[2:0];
  _RAND_578 = {1{`RANDOM}};
  state_vec_490 = _RAND_578[2:0];
  _RAND_579 = {1{`RANDOM}};
  state_vec_491 = _RAND_579[2:0];
  _RAND_580 = {1{`RANDOM}};
  state_vec_492 = _RAND_580[2:0];
  _RAND_581 = {1{`RANDOM}};
  state_vec_493 = _RAND_581[2:0];
  _RAND_582 = {1{`RANDOM}};
  state_vec_494 = _RAND_582[2:0];
  _RAND_583 = {1{`RANDOM}};
  state_vec_495 = _RAND_583[2:0];
  _RAND_584 = {1{`RANDOM}};
  state_vec_496 = _RAND_584[2:0];
  _RAND_585 = {1{`RANDOM}};
  state_vec_497 = _RAND_585[2:0];
  _RAND_586 = {1{`RANDOM}};
  state_vec_498 = _RAND_586[2:0];
  _RAND_587 = {1{`RANDOM}};
  state_vec_499 = _RAND_587[2:0];
  _RAND_588 = {1{`RANDOM}};
  state_vec_500 = _RAND_588[2:0];
  _RAND_589 = {1{`RANDOM}};
  state_vec_501 = _RAND_589[2:0];
  _RAND_590 = {1{`RANDOM}};
  state_vec_502 = _RAND_590[2:0];
  _RAND_591 = {1{`RANDOM}};
  state_vec_503 = _RAND_591[2:0];
  _RAND_592 = {1{`RANDOM}};
  state_vec_504 = _RAND_592[2:0];
  _RAND_593 = {1{`RANDOM}};
  state_vec_505 = _RAND_593[2:0];
  _RAND_594 = {1{`RANDOM}};
  state_vec_506 = _RAND_594[2:0];
  _RAND_595 = {1{`RANDOM}};
  state_vec_507 = _RAND_595[2:0];
  _RAND_596 = {1{`RANDOM}};
  state_vec_508 = _RAND_596[2:0];
  _RAND_597 = {1{`RANDOM}};
  state_vec_509 = _RAND_597[2:0];
  _RAND_598 = {1{`RANDOM}};
  state_vec_510 = _RAND_598[2:0];
  _RAND_599 = {1{`RANDOM}};
  state_vec_511 = _RAND_599[2:0];
  _RAND_600 = {1{`RANDOM}};
  allocWriteWay_REG_3 = _RAND_600[0:0];
  _RAND_601 = {1{`RANDOM}};
  allocWriteWay_REG_2 = _RAND_601[0:0];
  _RAND_602 = {1{`RANDOM}};
  allocWriteWay_REG_1 = _RAND_602[0:0];
  _RAND_603 = {1{`RANDOM}};
  allocWriteWay_REG_0 = _RAND_603[0:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    state_vec_0 = 3'h0;
  end
  if (reset) begin
    state_vec_1 = 3'h0;
  end
  if (reset) begin
    state_vec_2 = 3'h0;
  end
  if (reset) begin
    state_vec_3 = 3'h0;
  end
  if (reset) begin
    state_vec_4 = 3'h0;
  end
  if (reset) begin
    state_vec_5 = 3'h0;
  end
  if (reset) begin
    state_vec_6 = 3'h0;
  end
  if (reset) begin
    state_vec_7 = 3'h0;
  end
  if (reset) begin
    state_vec_8 = 3'h0;
  end
  if (reset) begin
    state_vec_9 = 3'h0;
  end
  if (reset) begin
    state_vec_10 = 3'h0;
  end
  if (reset) begin
    state_vec_11 = 3'h0;
  end
  if (reset) begin
    state_vec_12 = 3'h0;
  end
  if (reset) begin
    state_vec_13 = 3'h0;
  end
  if (reset) begin
    state_vec_14 = 3'h0;
  end
  if (reset) begin
    state_vec_15 = 3'h0;
  end
  if (reset) begin
    state_vec_16 = 3'h0;
  end
  if (reset) begin
    state_vec_17 = 3'h0;
  end
  if (reset) begin
    state_vec_18 = 3'h0;
  end
  if (reset) begin
    state_vec_19 = 3'h0;
  end
  if (reset) begin
    state_vec_20 = 3'h0;
  end
  if (reset) begin
    state_vec_21 = 3'h0;
  end
  if (reset) begin
    state_vec_22 = 3'h0;
  end
  if (reset) begin
    state_vec_23 = 3'h0;
  end
  if (reset) begin
    state_vec_24 = 3'h0;
  end
  if (reset) begin
    state_vec_25 = 3'h0;
  end
  if (reset) begin
    state_vec_26 = 3'h0;
  end
  if (reset) begin
    state_vec_27 = 3'h0;
  end
  if (reset) begin
    state_vec_28 = 3'h0;
  end
  if (reset) begin
    state_vec_29 = 3'h0;
  end
  if (reset) begin
    state_vec_30 = 3'h0;
  end
  if (reset) begin
    state_vec_31 = 3'h0;
  end
  if (reset) begin
    state_vec_32 = 3'h0;
  end
  if (reset) begin
    state_vec_33 = 3'h0;
  end
  if (reset) begin
    state_vec_34 = 3'h0;
  end
  if (reset) begin
    state_vec_35 = 3'h0;
  end
  if (reset) begin
    state_vec_36 = 3'h0;
  end
  if (reset) begin
    state_vec_37 = 3'h0;
  end
  if (reset) begin
    state_vec_38 = 3'h0;
  end
  if (reset) begin
    state_vec_39 = 3'h0;
  end
  if (reset) begin
    state_vec_40 = 3'h0;
  end
  if (reset) begin
    state_vec_41 = 3'h0;
  end
  if (reset) begin
    state_vec_42 = 3'h0;
  end
  if (reset) begin
    state_vec_43 = 3'h0;
  end
  if (reset) begin
    state_vec_44 = 3'h0;
  end
  if (reset) begin
    state_vec_45 = 3'h0;
  end
  if (reset) begin
    state_vec_46 = 3'h0;
  end
  if (reset) begin
    state_vec_47 = 3'h0;
  end
  if (reset) begin
    state_vec_48 = 3'h0;
  end
  if (reset) begin
    state_vec_49 = 3'h0;
  end
  if (reset) begin
    state_vec_50 = 3'h0;
  end
  if (reset) begin
    state_vec_51 = 3'h0;
  end
  if (reset) begin
    state_vec_52 = 3'h0;
  end
  if (reset) begin
    state_vec_53 = 3'h0;
  end
  if (reset) begin
    state_vec_54 = 3'h0;
  end
  if (reset) begin
    state_vec_55 = 3'h0;
  end
  if (reset) begin
    state_vec_56 = 3'h0;
  end
  if (reset) begin
    state_vec_57 = 3'h0;
  end
  if (reset) begin
    state_vec_58 = 3'h0;
  end
  if (reset) begin
    state_vec_59 = 3'h0;
  end
  if (reset) begin
    state_vec_60 = 3'h0;
  end
  if (reset) begin
    state_vec_61 = 3'h0;
  end
  if (reset) begin
    state_vec_62 = 3'h0;
  end
  if (reset) begin
    state_vec_63 = 3'h0;
  end
  if (reset) begin
    state_vec_64 = 3'h0;
  end
  if (reset) begin
    state_vec_65 = 3'h0;
  end
  if (reset) begin
    state_vec_66 = 3'h0;
  end
  if (reset) begin
    state_vec_67 = 3'h0;
  end
  if (reset) begin
    state_vec_68 = 3'h0;
  end
  if (reset) begin
    state_vec_69 = 3'h0;
  end
  if (reset) begin
    state_vec_70 = 3'h0;
  end
  if (reset) begin
    state_vec_71 = 3'h0;
  end
  if (reset) begin
    state_vec_72 = 3'h0;
  end
  if (reset) begin
    state_vec_73 = 3'h0;
  end
  if (reset) begin
    state_vec_74 = 3'h0;
  end
  if (reset) begin
    state_vec_75 = 3'h0;
  end
  if (reset) begin
    state_vec_76 = 3'h0;
  end
  if (reset) begin
    state_vec_77 = 3'h0;
  end
  if (reset) begin
    state_vec_78 = 3'h0;
  end
  if (reset) begin
    state_vec_79 = 3'h0;
  end
  if (reset) begin
    state_vec_80 = 3'h0;
  end
  if (reset) begin
    state_vec_81 = 3'h0;
  end
  if (reset) begin
    state_vec_82 = 3'h0;
  end
  if (reset) begin
    state_vec_83 = 3'h0;
  end
  if (reset) begin
    state_vec_84 = 3'h0;
  end
  if (reset) begin
    state_vec_85 = 3'h0;
  end
  if (reset) begin
    state_vec_86 = 3'h0;
  end
  if (reset) begin
    state_vec_87 = 3'h0;
  end
  if (reset) begin
    state_vec_88 = 3'h0;
  end
  if (reset) begin
    state_vec_89 = 3'h0;
  end
  if (reset) begin
    state_vec_90 = 3'h0;
  end
  if (reset) begin
    state_vec_91 = 3'h0;
  end
  if (reset) begin
    state_vec_92 = 3'h0;
  end
  if (reset) begin
    state_vec_93 = 3'h0;
  end
  if (reset) begin
    state_vec_94 = 3'h0;
  end
  if (reset) begin
    state_vec_95 = 3'h0;
  end
  if (reset) begin
    state_vec_96 = 3'h0;
  end
  if (reset) begin
    state_vec_97 = 3'h0;
  end
  if (reset) begin
    state_vec_98 = 3'h0;
  end
  if (reset) begin
    state_vec_99 = 3'h0;
  end
  if (reset) begin
    state_vec_100 = 3'h0;
  end
  if (reset) begin
    state_vec_101 = 3'h0;
  end
  if (reset) begin
    state_vec_102 = 3'h0;
  end
  if (reset) begin
    state_vec_103 = 3'h0;
  end
  if (reset) begin
    state_vec_104 = 3'h0;
  end
  if (reset) begin
    state_vec_105 = 3'h0;
  end
  if (reset) begin
    state_vec_106 = 3'h0;
  end
  if (reset) begin
    state_vec_107 = 3'h0;
  end
  if (reset) begin
    state_vec_108 = 3'h0;
  end
  if (reset) begin
    state_vec_109 = 3'h0;
  end
  if (reset) begin
    state_vec_110 = 3'h0;
  end
  if (reset) begin
    state_vec_111 = 3'h0;
  end
  if (reset) begin
    state_vec_112 = 3'h0;
  end
  if (reset) begin
    state_vec_113 = 3'h0;
  end
  if (reset) begin
    state_vec_114 = 3'h0;
  end
  if (reset) begin
    state_vec_115 = 3'h0;
  end
  if (reset) begin
    state_vec_116 = 3'h0;
  end
  if (reset) begin
    state_vec_117 = 3'h0;
  end
  if (reset) begin
    state_vec_118 = 3'h0;
  end
  if (reset) begin
    state_vec_119 = 3'h0;
  end
  if (reset) begin
    state_vec_120 = 3'h0;
  end
  if (reset) begin
    state_vec_121 = 3'h0;
  end
  if (reset) begin
    state_vec_122 = 3'h0;
  end
  if (reset) begin
    state_vec_123 = 3'h0;
  end
  if (reset) begin
    state_vec_124 = 3'h0;
  end
  if (reset) begin
    state_vec_125 = 3'h0;
  end
  if (reset) begin
    state_vec_126 = 3'h0;
  end
  if (reset) begin
    state_vec_127 = 3'h0;
  end
  if (reset) begin
    state_vec_128 = 3'h0;
  end
  if (reset) begin
    state_vec_129 = 3'h0;
  end
  if (reset) begin
    state_vec_130 = 3'h0;
  end
  if (reset) begin
    state_vec_131 = 3'h0;
  end
  if (reset) begin
    state_vec_132 = 3'h0;
  end
  if (reset) begin
    state_vec_133 = 3'h0;
  end
  if (reset) begin
    state_vec_134 = 3'h0;
  end
  if (reset) begin
    state_vec_135 = 3'h0;
  end
  if (reset) begin
    state_vec_136 = 3'h0;
  end
  if (reset) begin
    state_vec_137 = 3'h0;
  end
  if (reset) begin
    state_vec_138 = 3'h0;
  end
  if (reset) begin
    state_vec_139 = 3'h0;
  end
  if (reset) begin
    state_vec_140 = 3'h0;
  end
  if (reset) begin
    state_vec_141 = 3'h0;
  end
  if (reset) begin
    state_vec_142 = 3'h0;
  end
  if (reset) begin
    state_vec_143 = 3'h0;
  end
  if (reset) begin
    state_vec_144 = 3'h0;
  end
  if (reset) begin
    state_vec_145 = 3'h0;
  end
  if (reset) begin
    state_vec_146 = 3'h0;
  end
  if (reset) begin
    state_vec_147 = 3'h0;
  end
  if (reset) begin
    state_vec_148 = 3'h0;
  end
  if (reset) begin
    state_vec_149 = 3'h0;
  end
  if (reset) begin
    state_vec_150 = 3'h0;
  end
  if (reset) begin
    state_vec_151 = 3'h0;
  end
  if (reset) begin
    state_vec_152 = 3'h0;
  end
  if (reset) begin
    state_vec_153 = 3'h0;
  end
  if (reset) begin
    state_vec_154 = 3'h0;
  end
  if (reset) begin
    state_vec_155 = 3'h0;
  end
  if (reset) begin
    state_vec_156 = 3'h0;
  end
  if (reset) begin
    state_vec_157 = 3'h0;
  end
  if (reset) begin
    state_vec_158 = 3'h0;
  end
  if (reset) begin
    state_vec_159 = 3'h0;
  end
  if (reset) begin
    state_vec_160 = 3'h0;
  end
  if (reset) begin
    state_vec_161 = 3'h0;
  end
  if (reset) begin
    state_vec_162 = 3'h0;
  end
  if (reset) begin
    state_vec_163 = 3'h0;
  end
  if (reset) begin
    state_vec_164 = 3'h0;
  end
  if (reset) begin
    state_vec_165 = 3'h0;
  end
  if (reset) begin
    state_vec_166 = 3'h0;
  end
  if (reset) begin
    state_vec_167 = 3'h0;
  end
  if (reset) begin
    state_vec_168 = 3'h0;
  end
  if (reset) begin
    state_vec_169 = 3'h0;
  end
  if (reset) begin
    state_vec_170 = 3'h0;
  end
  if (reset) begin
    state_vec_171 = 3'h0;
  end
  if (reset) begin
    state_vec_172 = 3'h0;
  end
  if (reset) begin
    state_vec_173 = 3'h0;
  end
  if (reset) begin
    state_vec_174 = 3'h0;
  end
  if (reset) begin
    state_vec_175 = 3'h0;
  end
  if (reset) begin
    state_vec_176 = 3'h0;
  end
  if (reset) begin
    state_vec_177 = 3'h0;
  end
  if (reset) begin
    state_vec_178 = 3'h0;
  end
  if (reset) begin
    state_vec_179 = 3'h0;
  end
  if (reset) begin
    state_vec_180 = 3'h0;
  end
  if (reset) begin
    state_vec_181 = 3'h0;
  end
  if (reset) begin
    state_vec_182 = 3'h0;
  end
  if (reset) begin
    state_vec_183 = 3'h0;
  end
  if (reset) begin
    state_vec_184 = 3'h0;
  end
  if (reset) begin
    state_vec_185 = 3'h0;
  end
  if (reset) begin
    state_vec_186 = 3'h0;
  end
  if (reset) begin
    state_vec_187 = 3'h0;
  end
  if (reset) begin
    state_vec_188 = 3'h0;
  end
  if (reset) begin
    state_vec_189 = 3'h0;
  end
  if (reset) begin
    state_vec_190 = 3'h0;
  end
  if (reset) begin
    state_vec_191 = 3'h0;
  end
  if (reset) begin
    state_vec_192 = 3'h0;
  end
  if (reset) begin
    state_vec_193 = 3'h0;
  end
  if (reset) begin
    state_vec_194 = 3'h0;
  end
  if (reset) begin
    state_vec_195 = 3'h0;
  end
  if (reset) begin
    state_vec_196 = 3'h0;
  end
  if (reset) begin
    state_vec_197 = 3'h0;
  end
  if (reset) begin
    state_vec_198 = 3'h0;
  end
  if (reset) begin
    state_vec_199 = 3'h0;
  end
  if (reset) begin
    state_vec_200 = 3'h0;
  end
  if (reset) begin
    state_vec_201 = 3'h0;
  end
  if (reset) begin
    state_vec_202 = 3'h0;
  end
  if (reset) begin
    state_vec_203 = 3'h0;
  end
  if (reset) begin
    state_vec_204 = 3'h0;
  end
  if (reset) begin
    state_vec_205 = 3'h0;
  end
  if (reset) begin
    state_vec_206 = 3'h0;
  end
  if (reset) begin
    state_vec_207 = 3'h0;
  end
  if (reset) begin
    state_vec_208 = 3'h0;
  end
  if (reset) begin
    state_vec_209 = 3'h0;
  end
  if (reset) begin
    state_vec_210 = 3'h0;
  end
  if (reset) begin
    state_vec_211 = 3'h0;
  end
  if (reset) begin
    state_vec_212 = 3'h0;
  end
  if (reset) begin
    state_vec_213 = 3'h0;
  end
  if (reset) begin
    state_vec_214 = 3'h0;
  end
  if (reset) begin
    state_vec_215 = 3'h0;
  end
  if (reset) begin
    state_vec_216 = 3'h0;
  end
  if (reset) begin
    state_vec_217 = 3'h0;
  end
  if (reset) begin
    state_vec_218 = 3'h0;
  end
  if (reset) begin
    state_vec_219 = 3'h0;
  end
  if (reset) begin
    state_vec_220 = 3'h0;
  end
  if (reset) begin
    state_vec_221 = 3'h0;
  end
  if (reset) begin
    state_vec_222 = 3'h0;
  end
  if (reset) begin
    state_vec_223 = 3'h0;
  end
  if (reset) begin
    state_vec_224 = 3'h0;
  end
  if (reset) begin
    state_vec_225 = 3'h0;
  end
  if (reset) begin
    state_vec_226 = 3'h0;
  end
  if (reset) begin
    state_vec_227 = 3'h0;
  end
  if (reset) begin
    state_vec_228 = 3'h0;
  end
  if (reset) begin
    state_vec_229 = 3'h0;
  end
  if (reset) begin
    state_vec_230 = 3'h0;
  end
  if (reset) begin
    state_vec_231 = 3'h0;
  end
  if (reset) begin
    state_vec_232 = 3'h0;
  end
  if (reset) begin
    state_vec_233 = 3'h0;
  end
  if (reset) begin
    state_vec_234 = 3'h0;
  end
  if (reset) begin
    state_vec_235 = 3'h0;
  end
  if (reset) begin
    state_vec_236 = 3'h0;
  end
  if (reset) begin
    state_vec_237 = 3'h0;
  end
  if (reset) begin
    state_vec_238 = 3'h0;
  end
  if (reset) begin
    state_vec_239 = 3'h0;
  end
  if (reset) begin
    state_vec_240 = 3'h0;
  end
  if (reset) begin
    state_vec_241 = 3'h0;
  end
  if (reset) begin
    state_vec_242 = 3'h0;
  end
  if (reset) begin
    state_vec_243 = 3'h0;
  end
  if (reset) begin
    state_vec_244 = 3'h0;
  end
  if (reset) begin
    state_vec_245 = 3'h0;
  end
  if (reset) begin
    state_vec_246 = 3'h0;
  end
  if (reset) begin
    state_vec_247 = 3'h0;
  end
  if (reset) begin
    state_vec_248 = 3'h0;
  end
  if (reset) begin
    state_vec_249 = 3'h0;
  end
  if (reset) begin
    state_vec_250 = 3'h0;
  end
  if (reset) begin
    state_vec_251 = 3'h0;
  end
  if (reset) begin
    state_vec_252 = 3'h0;
  end
  if (reset) begin
    state_vec_253 = 3'h0;
  end
  if (reset) begin
    state_vec_254 = 3'h0;
  end
  if (reset) begin
    state_vec_255 = 3'h0;
  end
  if (reset) begin
    state_vec_256 = 3'h0;
  end
  if (reset) begin
    state_vec_257 = 3'h0;
  end
  if (reset) begin
    state_vec_258 = 3'h0;
  end
  if (reset) begin
    state_vec_259 = 3'h0;
  end
  if (reset) begin
    state_vec_260 = 3'h0;
  end
  if (reset) begin
    state_vec_261 = 3'h0;
  end
  if (reset) begin
    state_vec_262 = 3'h0;
  end
  if (reset) begin
    state_vec_263 = 3'h0;
  end
  if (reset) begin
    state_vec_264 = 3'h0;
  end
  if (reset) begin
    state_vec_265 = 3'h0;
  end
  if (reset) begin
    state_vec_266 = 3'h0;
  end
  if (reset) begin
    state_vec_267 = 3'h0;
  end
  if (reset) begin
    state_vec_268 = 3'h0;
  end
  if (reset) begin
    state_vec_269 = 3'h0;
  end
  if (reset) begin
    state_vec_270 = 3'h0;
  end
  if (reset) begin
    state_vec_271 = 3'h0;
  end
  if (reset) begin
    state_vec_272 = 3'h0;
  end
  if (reset) begin
    state_vec_273 = 3'h0;
  end
  if (reset) begin
    state_vec_274 = 3'h0;
  end
  if (reset) begin
    state_vec_275 = 3'h0;
  end
  if (reset) begin
    state_vec_276 = 3'h0;
  end
  if (reset) begin
    state_vec_277 = 3'h0;
  end
  if (reset) begin
    state_vec_278 = 3'h0;
  end
  if (reset) begin
    state_vec_279 = 3'h0;
  end
  if (reset) begin
    state_vec_280 = 3'h0;
  end
  if (reset) begin
    state_vec_281 = 3'h0;
  end
  if (reset) begin
    state_vec_282 = 3'h0;
  end
  if (reset) begin
    state_vec_283 = 3'h0;
  end
  if (reset) begin
    state_vec_284 = 3'h0;
  end
  if (reset) begin
    state_vec_285 = 3'h0;
  end
  if (reset) begin
    state_vec_286 = 3'h0;
  end
  if (reset) begin
    state_vec_287 = 3'h0;
  end
  if (reset) begin
    state_vec_288 = 3'h0;
  end
  if (reset) begin
    state_vec_289 = 3'h0;
  end
  if (reset) begin
    state_vec_290 = 3'h0;
  end
  if (reset) begin
    state_vec_291 = 3'h0;
  end
  if (reset) begin
    state_vec_292 = 3'h0;
  end
  if (reset) begin
    state_vec_293 = 3'h0;
  end
  if (reset) begin
    state_vec_294 = 3'h0;
  end
  if (reset) begin
    state_vec_295 = 3'h0;
  end
  if (reset) begin
    state_vec_296 = 3'h0;
  end
  if (reset) begin
    state_vec_297 = 3'h0;
  end
  if (reset) begin
    state_vec_298 = 3'h0;
  end
  if (reset) begin
    state_vec_299 = 3'h0;
  end
  if (reset) begin
    state_vec_300 = 3'h0;
  end
  if (reset) begin
    state_vec_301 = 3'h0;
  end
  if (reset) begin
    state_vec_302 = 3'h0;
  end
  if (reset) begin
    state_vec_303 = 3'h0;
  end
  if (reset) begin
    state_vec_304 = 3'h0;
  end
  if (reset) begin
    state_vec_305 = 3'h0;
  end
  if (reset) begin
    state_vec_306 = 3'h0;
  end
  if (reset) begin
    state_vec_307 = 3'h0;
  end
  if (reset) begin
    state_vec_308 = 3'h0;
  end
  if (reset) begin
    state_vec_309 = 3'h0;
  end
  if (reset) begin
    state_vec_310 = 3'h0;
  end
  if (reset) begin
    state_vec_311 = 3'h0;
  end
  if (reset) begin
    state_vec_312 = 3'h0;
  end
  if (reset) begin
    state_vec_313 = 3'h0;
  end
  if (reset) begin
    state_vec_314 = 3'h0;
  end
  if (reset) begin
    state_vec_315 = 3'h0;
  end
  if (reset) begin
    state_vec_316 = 3'h0;
  end
  if (reset) begin
    state_vec_317 = 3'h0;
  end
  if (reset) begin
    state_vec_318 = 3'h0;
  end
  if (reset) begin
    state_vec_319 = 3'h0;
  end
  if (reset) begin
    state_vec_320 = 3'h0;
  end
  if (reset) begin
    state_vec_321 = 3'h0;
  end
  if (reset) begin
    state_vec_322 = 3'h0;
  end
  if (reset) begin
    state_vec_323 = 3'h0;
  end
  if (reset) begin
    state_vec_324 = 3'h0;
  end
  if (reset) begin
    state_vec_325 = 3'h0;
  end
  if (reset) begin
    state_vec_326 = 3'h0;
  end
  if (reset) begin
    state_vec_327 = 3'h0;
  end
  if (reset) begin
    state_vec_328 = 3'h0;
  end
  if (reset) begin
    state_vec_329 = 3'h0;
  end
  if (reset) begin
    state_vec_330 = 3'h0;
  end
  if (reset) begin
    state_vec_331 = 3'h0;
  end
  if (reset) begin
    state_vec_332 = 3'h0;
  end
  if (reset) begin
    state_vec_333 = 3'h0;
  end
  if (reset) begin
    state_vec_334 = 3'h0;
  end
  if (reset) begin
    state_vec_335 = 3'h0;
  end
  if (reset) begin
    state_vec_336 = 3'h0;
  end
  if (reset) begin
    state_vec_337 = 3'h0;
  end
  if (reset) begin
    state_vec_338 = 3'h0;
  end
  if (reset) begin
    state_vec_339 = 3'h0;
  end
  if (reset) begin
    state_vec_340 = 3'h0;
  end
  if (reset) begin
    state_vec_341 = 3'h0;
  end
  if (reset) begin
    state_vec_342 = 3'h0;
  end
  if (reset) begin
    state_vec_343 = 3'h0;
  end
  if (reset) begin
    state_vec_344 = 3'h0;
  end
  if (reset) begin
    state_vec_345 = 3'h0;
  end
  if (reset) begin
    state_vec_346 = 3'h0;
  end
  if (reset) begin
    state_vec_347 = 3'h0;
  end
  if (reset) begin
    state_vec_348 = 3'h0;
  end
  if (reset) begin
    state_vec_349 = 3'h0;
  end
  if (reset) begin
    state_vec_350 = 3'h0;
  end
  if (reset) begin
    state_vec_351 = 3'h0;
  end
  if (reset) begin
    state_vec_352 = 3'h0;
  end
  if (reset) begin
    state_vec_353 = 3'h0;
  end
  if (reset) begin
    state_vec_354 = 3'h0;
  end
  if (reset) begin
    state_vec_355 = 3'h0;
  end
  if (reset) begin
    state_vec_356 = 3'h0;
  end
  if (reset) begin
    state_vec_357 = 3'h0;
  end
  if (reset) begin
    state_vec_358 = 3'h0;
  end
  if (reset) begin
    state_vec_359 = 3'h0;
  end
  if (reset) begin
    state_vec_360 = 3'h0;
  end
  if (reset) begin
    state_vec_361 = 3'h0;
  end
  if (reset) begin
    state_vec_362 = 3'h0;
  end
  if (reset) begin
    state_vec_363 = 3'h0;
  end
  if (reset) begin
    state_vec_364 = 3'h0;
  end
  if (reset) begin
    state_vec_365 = 3'h0;
  end
  if (reset) begin
    state_vec_366 = 3'h0;
  end
  if (reset) begin
    state_vec_367 = 3'h0;
  end
  if (reset) begin
    state_vec_368 = 3'h0;
  end
  if (reset) begin
    state_vec_369 = 3'h0;
  end
  if (reset) begin
    state_vec_370 = 3'h0;
  end
  if (reset) begin
    state_vec_371 = 3'h0;
  end
  if (reset) begin
    state_vec_372 = 3'h0;
  end
  if (reset) begin
    state_vec_373 = 3'h0;
  end
  if (reset) begin
    state_vec_374 = 3'h0;
  end
  if (reset) begin
    state_vec_375 = 3'h0;
  end
  if (reset) begin
    state_vec_376 = 3'h0;
  end
  if (reset) begin
    state_vec_377 = 3'h0;
  end
  if (reset) begin
    state_vec_378 = 3'h0;
  end
  if (reset) begin
    state_vec_379 = 3'h0;
  end
  if (reset) begin
    state_vec_380 = 3'h0;
  end
  if (reset) begin
    state_vec_381 = 3'h0;
  end
  if (reset) begin
    state_vec_382 = 3'h0;
  end
  if (reset) begin
    state_vec_383 = 3'h0;
  end
  if (reset) begin
    state_vec_384 = 3'h0;
  end
  if (reset) begin
    state_vec_385 = 3'h0;
  end
  if (reset) begin
    state_vec_386 = 3'h0;
  end
  if (reset) begin
    state_vec_387 = 3'h0;
  end
  if (reset) begin
    state_vec_388 = 3'h0;
  end
  if (reset) begin
    state_vec_389 = 3'h0;
  end
  if (reset) begin
    state_vec_390 = 3'h0;
  end
  if (reset) begin
    state_vec_391 = 3'h0;
  end
  if (reset) begin
    state_vec_392 = 3'h0;
  end
  if (reset) begin
    state_vec_393 = 3'h0;
  end
  if (reset) begin
    state_vec_394 = 3'h0;
  end
  if (reset) begin
    state_vec_395 = 3'h0;
  end
  if (reset) begin
    state_vec_396 = 3'h0;
  end
  if (reset) begin
    state_vec_397 = 3'h0;
  end
  if (reset) begin
    state_vec_398 = 3'h0;
  end
  if (reset) begin
    state_vec_399 = 3'h0;
  end
  if (reset) begin
    state_vec_400 = 3'h0;
  end
  if (reset) begin
    state_vec_401 = 3'h0;
  end
  if (reset) begin
    state_vec_402 = 3'h0;
  end
  if (reset) begin
    state_vec_403 = 3'h0;
  end
  if (reset) begin
    state_vec_404 = 3'h0;
  end
  if (reset) begin
    state_vec_405 = 3'h0;
  end
  if (reset) begin
    state_vec_406 = 3'h0;
  end
  if (reset) begin
    state_vec_407 = 3'h0;
  end
  if (reset) begin
    state_vec_408 = 3'h0;
  end
  if (reset) begin
    state_vec_409 = 3'h0;
  end
  if (reset) begin
    state_vec_410 = 3'h0;
  end
  if (reset) begin
    state_vec_411 = 3'h0;
  end
  if (reset) begin
    state_vec_412 = 3'h0;
  end
  if (reset) begin
    state_vec_413 = 3'h0;
  end
  if (reset) begin
    state_vec_414 = 3'h0;
  end
  if (reset) begin
    state_vec_415 = 3'h0;
  end
  if (reset) begin
    state_vec_416 = 3'h0;
  end
  if (reset) begin
    state_vec_417 = 3'h0;
  end
  if (reset) begin
    state_vec_418 = 3'h0;
  end
  if (reset) begin
    state_vec_419 = 3'h0;
  end
  if (reset) begin
    state_vec_420 = 3'h0;
  end
  if (reset) begin
    state_vec_421 = 3'h0;
  end
  if (reset) begin
    state_vec_422 = 3'h0;
  end
  if (reset) begin
    state_vec_423 = 3'h0;
  end
  if (reset) begin
    state_vec_424 = 3'h0;
  end
  if (reset) begin
    state_vec_425 = 3'h0;
  end
  if (reset) begin
    state_vec_426 = 3'h0;
  end
  if (reset) begin
    state_vec_427 = 3'h0;
  end
  if (reset) begin
    state_vec_428 = 3'h0;
  end
  if (reset) begin
    state_vec_429 = 3'h0;
  end
  if (reset) begin
    state_vec_430 = 3'h0;
  end
  if (reset) begin
    state_vec_431 = 3'h0;
  end
  if (reset) begin
    state_vec_432 = 3'h0;
  end
  if (reset) begin
    state_vec_433 = 3'h0;
  end
  if (reset) begin
    state_vec_434 = 3'h0;
  end
  if (reset) begin
    state_vec_435 = 3'h0;
  end
  if (reset) begin
    state_vec_436 = 3'h0;
  end
  if (reset) begin
    state_vec_437 = 3'h0;
  end
  if (reset) begin
    state_vec_438 = 3'h0;
  end
  if (reset) begin
    state_vec_439 = 3'h0;
  end
  if (reset) begin
    state_vec_440 = 3'h0;
  end
  if (reset) begin
    state_vec_441 = 3'h0;
  end
  if (reset) begin
    state_vec_442 = 3'h0;
  end
  if (reset) begin
    state_vec_443 = 3'h0;
  end
  if (reset) begin
    state_vec_444 = 3'h0;
  end
  if (reset) begin
    state_vec_445 = 3'h0;
  end
  if (reset) begin
    state_vec_446 = 3'h0;
  end
  if (reset) begin
    state_vec_447 = 3'h0;
  end
  if (reset) begin
    state_vec_448 = 3'h0;
  end
  if (reset) begin
    state_vec_449 = 3'h0;
  end
  if (reset) begin
    state_vec_450 = 3'h0;
  end
  if (reset) begin
    state_vec_451 = 3'h0;
  end
  if (reset) begin
    state_vec_452 = 3'h0;
  end
  if (reset) begin
    state_vec_453 = 3'h0;
  end
  if (reset) begin
    state_vec_454 = 3'h0;
  end
  if (reset) begin
    state_vec_455 = 3'h0;
  end
  if (reset) begin
    state_vec_456 = 3'h0;
  end
  if (reset) begin
    state_vec_457 = 3'h0;
  end
  if (reset) begin
    state_vec_458 = 3'h0;
  end
  if (reset) begin
    state_vec_459 = 3'h0;
  end
  if (reset) begin
    state_vec_460 = 3'h0;
  end
  if (reset) begin
    state_vec_461 = 3'h0;
  end
  if (reset) begin
    state_vec_462 = 3'h0;
  end
  if (reset) begin
    state_vec_463 = 3'h0;
  end
  if (reset) begin
    state_vec_464 = 3'h0;
  end
  if (reset) begin
    state_vec_465 = 3'h0;
  end
  if (reset) begin
    state_vec_466 = 3'h0;
  end
  if (reset) begin
    state_vec_467 = 3'h0;
  end
  if (reset) begin
    state_vec_468 = 3'h0;
  end
  if (reset) begin
    state_vec_469 = 3'h0;
  end
  if (reset) begin
    state_vec_470 = 3'h0;
  end
  if (reset) begin
    state_vec_471 = 3'h0;
  end
  if (reset) begin
    state_vec_472 = 3'h0;
  end
  if (reset) begin
    state_vec_473 = 3'h0;
  end
  if (reset) begin
    state_vec_474 = 3'h0;
  end
  if (reset) begin
    state_vec_475 = 3'h0;
  end
  if (reset) begin
    state_vec_476 = 3'h0;
  end
  if (reset) begin
    state_vec_477 = 3'h0;
  end
  if (reset) begin
    state_vec_478 = 3'h0;
  end
  if (reset) begin
    state_vec_479 = 3'h0;
  end
  if (reset) begin
    state_vec_480 = 3'h0;
  end
  if (reset) begin
    state_vec_481 = 3'h0;
  end
  if (reset) begin
    state_vec_482 = 3'h0;
  end
  if (reset) begin
    state_vec_483 = 3'h0;
  end
  if (reset) begin
    state_vec_484 = 3'h0;
  end
  if (reset) begin
    state_vec_485 = 3'h0;
  end
  if (reset) begin
    state_vec_486 = 3'h0;
  end
  if (reset) begin
    state_vec_487 = 3'h0;
  end
  if (reset) begin
    state_vec_488 = 3'h0;
  end
  if (reset) begin
    state_vec_489 = 3'h0;
  end
  if (reset) begin
    state_vec_490 = 3'h0;
  end
  if (reset) begin
    state_vec_491 = 3'h0;
  end
  if (reset) begin
    state_vec_492 = 3'h0;
  end
  if (reset) begin
    state_vec_493 = 3'h0;
  end
  if (reset) begin
    state_vec_494 = 3'h0;
  end
  if (reset) begin
    state_vec_495 = 3'h0;
  end
  if (reset) begin
    state_vec_496 = 3'h0;
  end
  if (reset) begin
    state_vec_497 = 3'h0;
  end
  if (reset) begin
    state_vec_498 = 3'h0;
  end
  if (reset) begin
    state_vec_499 = 3'h0;
  end
  if (reset) begin
    state_vec_500 = 3'h0;
  end
  if (reset) begin
    state_vec_501 = 3'h0;
  end
  if (reset) begin
    state_vec_502 = 3'h0;
  end
  if (reset) begin
    state_vec_503 = 3'h0;
  end
  if (reset) begin
    state_vec_504 = 3'h0;
  end
  if (reset) begin
    state_vec_505 = 3'h0;
  end
  if (reset) begin
    state_vec_506 = 3'h0;
  end
  if (reset) begin
    state_vec_507 = 3'h0;
  end
  if (reset) begin
    state_vec_508 = 3'h0;
  end
  if (reset) begin
    state_vec_509 = 3'h0;
  end
  if (reset) begin
    state_vec_510 = 3'h0;
  end
  if (reset) begin
    state_vec_511 = 3'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule

