module LFST(
  input        clock,
  input        reset,
  input        io_redirect_valid,
  input        io_redirect_bits_robIdx_flag,
  input  [4:0] io_redirect_bits_robIdx_value,
  input        io_redirect_bits_level,
  input        io_dispatch_req_0_valid,
  input        io_dispatch_req_0_bits_isstore,
  input  [4:0] io_dispatch_req_0_bits_ssid,
  input        io_dispatch_req_0_bits_robIdx_flag,
  input  [4:0] io_dispatch_req_0_bits_robIdx_value,
  input        io_dispatch_req_1_valid,
  input        io_dispatch_req_1_bits_isstore,
  input  [4:0] io_dispatch_req_1_bits_ssid,
  input        io_dispatch_req_1_bits_robIdx_flag,
  input  [4:0] io_dispatch_req_1_bits_robIdx_value,
  output       io_dispatch_resp_0_bits_shouldWait,
  output       io_dispatch_resp_0_bits_robIdx_flag,
  output [4:0] io_dispatch_resp_0_bits_robIdx_value,
  output       io_dispatch_resp_1_bits_shouldWait,
  output       io_dispatch_resp_1_bits_robIdx_flag,
  output [4:0] io_dispatch_resp_1_bits_robIdx_value,
  input        io_storeIssue_0_valid,
  input        io_storeIssue_0_bits_uop_cf_storeSetHit,
  input  [4:0] io_storeIssue_0_bits_uop_cf_ssid,
  input  [4:0] io_storeIssue_0_bits_uop_robIdx_value,
  input        io_storeIssue_1_valid,
  input        io_storeIssue_1_bits_uop_cf_storeSetHit,
  input  [4:0] io_storeIssue_1_bits_uop_cf_ssid,
  input  [4:0] io_storeIssue_1_bits_uop_robIdx_value,
  input        io_csrCtrl_lvpred_disable,
  input        io_csrCtrl_no_spec_load,
  input        io_csrCtrl_storeset_wait_store
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
`endif // RANDOMIZE_REG_INIT
  reg  validVec_0_0; // @[StoreSet.scala 491:25]
  reg  validVec_0_1; // @[StoreSet.scala 491:25]
  reg  validVec_0_2; // @[StoreSet.scala 491:25]
  reg  validVec_0_3; // @[StoreSet.scala 491:25]
  reg  validVec_1_0; // @[StoreSet.scala 491:25]
  reg  validVec_1_1; // @[StoreSet.scala 491:25]
  reg  validVec_1_2; // @[StoreSet.scala 491:25]
  reg  validVec_1_3; // @[StoreSet.scala 491:25]
  reg  validVec_2_0; // @[StoreSet.scala 491:25]
  reg  validVec_2_1; // @[StoreSet.scala 491:25]
  reg  validVec_2_2; // @[StoreSet.scala 491:25]
  reg  validVec_2_3; // @[StoreSet.scala 491:25]
  reg  validVec_3_0; // @[StoreSet.scala 491:25]
  reg  validVec_3_1; // @[StoreSet.scala 491:25]
  reg  validVec_3_2; // @[StoreSet.scala 491:25]
  reg  validVec_3_3; // @[StoreSet.scala 491:25]
  reg  validVec_4_0; // @[StoreSet.scala 491:25]
  reg  validVec_4_1; // @[StoreSet.scala 491:25]
  reg  validVec_4_2; // @[StoreSet.scala 491:25]
  reg  validVec_4_3; // @[StoreSet.scala 491:25]
  reg  validVec_5_0; // @[StoreSet.scala 491:25]
  reg  validVec_5_1; // @[StoreSet.scala 491:25]
  reg  validVec_5_2; // @[StoreSet.scala 491:25]
  reg  validVec_5_3; // @[StoreSet.scala 491:25]
  reg  validVec_6_0; // @[StoreSet.scala 491:25]
  reg  validVec_6_1; // @[StoreSet.scala 491:25]
  reg  validVec_6_2; // @[StoreSet.scala 491:25]
  reg  validVec_6_3; // @[StoreSet.scala 491:25]
  reg  validVec_7_0; // @[StoreSet.scala 491:25]
  reg  validVec_7_1; // @[StoreSet.scala 491:25]
  reg  validVec_7_2; // @[StoreSet.scala 491:25]
  reg  validVec_7_3; // @[StoreSet.scala 491:25]
  reg  validVec_8_0; // @[StoreSet.scala 491:25]
  reg  validVec_8_1; // @[StoreSet.scala 491:25]
  reg  validVec_8_2; // @[StoreSet.scala 491:25]
  reg  validVec_8_3; // @[StoreSet.scala 491:25]
  reg  validVec_9_0; // @[StoreSet.scala 491:25]
  reg  validVec_9_1; // @[StoreSet.scala 491:25]
  reg  validVec_9_2; // @[StoreSet.scala 491:25]
  reg  validVec_9_3; // @[StoreSet.scala 491:25]
  reg  validVec_10_0; // @[StoreSet.scala 491:25]
  reg  validVec_10_1; // @[StoreSet.scala 491:25]
  reg  validVec_10_2; // @[StoreSet.scala 491:25]
  reg  validVec_10_3; // @[StoreSet.scala 491:25]
  reg  validVec_11_0; // @[StoreSet.scala 491:25]
  reg  validVec_11_1; // @[StoreSet.scala 491:25]
  reg  validVec_11_2; // @[StoreSet.scala 491:25]
  reg  validVec_11_3; // @[StoreSet.scala 491:25]
  reg  validVec_12_0; // @[StoreSet.scala 491:25]
  reg  validVec_12_1; // @[StoreSet.scala 491:25]
  reg  validVec_12_2; // @[StoreSet.scala 491:25]
  reg  validVec_12_3; // @[StoreSet.scala 491:25]
  reg  validVec_13_0; // @[StoreSet.scala 491:25]
  reg  validVec_13_1; // @[StoreSet.scala 491:25]
  reg  validVec_13_2; // @[StoreSet.scala 491:25]
  reg  validVec_13_3; // @[StoreSet.scala 491:25]
  reg  validVec_14_0; // @[StoreSet.scala 491:25]
  reg  validVec_14_1; // @[StoreSet.scala 491:25]
  reg  validVec_14_2; // @[StoreSet.scala 491:25]
  reg  validVec_14_3; // @[StoreSet.scala 491:25]
  reg  validVec_15_0; // @[StoreSet.scala 491:25]
  reg  validVec_15_1; // @[StoreSet.scala 491:25]
  reg  validVec_15_2; // @[StoreSet.scala 491:25]
  reg  validVec_15_3; // @[StoreSet.scala 491:25]
  reg  validVec_16_0; // @[StoreSet.scala 491:25]
  reg  validVec_16_1; // @[StoreSet.scala 491:25]
  reg  validVec_16_2; // @[StoreSet.scala 491:25]
  reg  validVec_16_3; // @[StoreSet.scala 491:25]
  reg  validVec_17_0; // @[StoreSet.scala 491:25]
  reg  validVec_17_1; // @[StoreSet.scala 491:25]
  reg  validVec_17_2; // @[StoreSet.scala 491:25]
  reg  validVec_17_3; // @[StoreSet.scala 491:25]
  reg  validVec_18_0; // @[StoreSet.scala 491:25]
  reg  validVec_18_1; // @[StoreSet.scala 491:25]
  reg  validVec_18_2; // @[StoreSet.scala 491:25]
  reg  validVec_18_3; // @[StoreSet.scala 491:25]
  reg  validVec_19_0; // @[StoreSet.scala 491:25]
  reg  validVec_19_1; // @[StoreSet.scala 491:25]
  reg  validVec_19_2; // @[StoreSet.scala 491:25]
  reg  validVec_19_3; // @[StoreSet.scala 491:25]
  reg  validVec_20_0; // @[StoreSet.scala 491:25]
  reg  validVec_20_1; // @[StoreSet.scala 491:25]
  reg  validVec_20_2; // @[StoreSet.scala 491:25]
  reg  validVec_20_3; // @[StoreSet.scala 491:25]
  reg  validVec_21_0; // @[StoreSet.scala 491:25]
  reg  validVec_21_1; // @[StoreSet.scala 491:25]
  reg  validVec_21_2; // @[StoreSet.scala 491:25]
  reg  validVec_21_3; // @[StoreSet.scala 491:25]
  reg  validVec_22_0; // @[StoreSet.scala 491:25]
  reg  validVec_22_1; // @[StoreSet.scala 491:25]
  reg  validVec_22_2; // @[StoreSet.scala 491:25]
  reg  validVec_22_3; // @[StoreSet.scala 491:25]
  reg  validVec_23_0; // @[StoreSet.scala 491:25]
  reg  validVec_23_1; // @[StoreSet.scala 491:25]
  reg  validVec_23_2; // @[StoreSet.scala 491:25]
  reg  validVec_23_3; // @[StoreSet.scala 491:25]
  reg  validVec_24_0; // @[StoreSet.scala 491:25]
  reg  validVec_24_1; // @[StoreSet.scala 491:25]
  reg  validVec_24_2; // @[StoreSet.scala 491:25]
  reg  validVec_24_3; // @[StoreSet.scala 491:25]
  reg  validVec_25_0; // @[StoreSet.scala 491:25]
  reg  validVec_25_1; // @[StoreSet.scala 491:25]
  reg  validVec_25_2; // @[StoreSet.scala 491:25]
  reg  validVec_25_3; // @[StoreSet.scala 491:25]
  reg  validVec_26_0; // @[StoreSet.scala 491:25]
  reg  validVec_26_1; // @[StoreSet.scala 491:25]
  reg  validVec_26_2; // @[StoreSet.scala 491:25]
  reg  validVec_26_3; // @[StoreSet.scala 491:25]
  reg  validVec_27_0; // @[StoreSet.scala 491:25]
  reg  validVec_27_1; // @[StoreSet.scala 491:25]
  reg  validVec_27_2; // @[StoreSet.scala 491:25]
  reg  validVec_27_3; // @[StoreSet.scala 491:25]
  reg  validVec_28_0; // @[StoreSet.scala 491:25]
  reg  validVec_28_1; // @[StoreSet.scala 491:25]
  reg  validVec_28_2; // @[StoreSet.scala 491:25]
  reg  validVec_28_3; // @[StoreSet.scala 491:25]
  reg  validVec_29_0; // @[StoreSet.scala 491:25]
  reg  validVec_29_1; // @[StoreSet.scala 491:25]
  reg  validVec_29_2; // @[StoreSet.scala 491:25]
  reg  validVec_29_3; // @[StoreSet.scala 491:25]
  reg  validVec_30_0; // @[StoreSet.scala 491:25]
  reg  validVec_30_1; // @[StoreSet.scala 491:25]
  reg  validVec_30_2; // @[StoreSet.scala 491:25]
  reg  validVec_30_3; // @[StoreSet.scala 491:25]
  reg  validVec_31_0; // @[StoreSet.scala 491:25]
  reg  validVec_31_1; // @[StoreSet.scala 491:25]
  reg  validVec_31_2; // @[StoreSet.scala 491:25]
  reg  validVec_31_3; // @[StoreSet.scala 491:25]
  reg  robIdxVec_0_0_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_0_0_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_0_1_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_0_1_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_0_2_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_0_2_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_0_3_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_0_3_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_1_0_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_1_0_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_1_1_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_1_1_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_1_2_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_1_2_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_1_3_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_1_3_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_2_0_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_2_0_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_2_1_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_2_1_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_2_2_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_2_2_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_2_3_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_2_3_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_3_0_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_3_0_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_3_1_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_3_1_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_3_2_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_3_2_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_3_3_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_3_3_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_4_0_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_4_0_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_4_1_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_4_1_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_4_2_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_4_2_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_4_3_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_4_3_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_5_0_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_5_0_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_5_1_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_5_1_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_5_2_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_5_2_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_5_3_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_5_3_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_6_0_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_6_0_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_6_1_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_6_1_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_6_2_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_6_2_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_6_3_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_6_3_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_7_0_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_7_0_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_7_1_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_7_1_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_7_2_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_7_2_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_7_3_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_7_3_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_8_0_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_8_0_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_8_1_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_8_1_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_8_2_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_8_2_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_8_3_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_8_3_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_9_0_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_9_0_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_9_1_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_9_1_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_9_2_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_9_2_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_9_3_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_9_3_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_10_0_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_10_0_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_10_1_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_10_1_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_10_2_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_10_2_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_10_3_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_10_3_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_11_0_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_11_0_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_11_1_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_11_1_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_11_2_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_11_2_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_11_3_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_11_3_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_12_0_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_12_0_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_12_1_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_12_1_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_12_2_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_12_2_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_12_3_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_12_3_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_13_0_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_13_0_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_13_1_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_13_1_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_13_2_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_13_2_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_13_3_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_13_3_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_14_0_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_14_0_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_14_1_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_14_1_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_14_2_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_14_2_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_14_3_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_14_3_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_15_0_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_15_0_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_15_1_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_15_1_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_15_2_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_15_2_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_15_3_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_15_3_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_16_0_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_16_0_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_16_1_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_16_1_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_16_2_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_16_2_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_16_3_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_16_3_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_17_0_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_17_0_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_17_1_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_17_1_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_17_2_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_17_2_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_17_3_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_17_3_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_18_0_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_18_0_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_18_1_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_18_1_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_18_2_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_18_2_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_18_3_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_18_3_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_19_0_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_19_0_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_19_1_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_19_1_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_19_2_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_19_2_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_19_3_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_19_3_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_20_0_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_20_0_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_20_1_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_20_1_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_20_2_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_20_2_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_20_3_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_20_3_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_21_0_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_21_0_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_21_1_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_21_1_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_21_2_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_21_2_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_21_3_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_21_3_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_22_0_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_22_0_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_22_1_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_22_1_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_22_2_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_22_2_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_22_3_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_22_3_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_23_0_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_23_0_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_23_1_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_23_1_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_23_2_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_23_2_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_23_3_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_23_3_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_24_0_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_24_0_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_24_1_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_24_1_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_24_2_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_24_2_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_24_3_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_24_3_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_25_0_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_25_0_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_25_1_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_25_1_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_25_2_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_25_2_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_25_3_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_25_3_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_26_0_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_26_0_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_26_1_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_26_1_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_26_2_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_26_2_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_26_3_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_26_3_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_27_0_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_27_0_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_27_1_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_27_1_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_27_2_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_27_2_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_27_3_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_27_3_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_28_0_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_28_0_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_28_1_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_28_1_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_28_2_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_28_2_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_28_3_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_28_3_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_29_0_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_29_0_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_29_1_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_29_1_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_29_2_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_29_2_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_29_3_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_29_3_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_30_0_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_30_0_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_30_1_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_30_1_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_30_2_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_30_2_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_30_3_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_30_3_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_31_0_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_31_0_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_31_1_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_31_1_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_31_2_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_31_2_value; // @[StoreSet.scala 492:22]
  reg  robIdxVec_31_3_flag; // @[StoreSet.scala 492:22]
  reg [4:0] robIdxVec_31_3_value; // @[StoreSet.scala 492:22]
  reg [1:0] allocPtr_0; // @[StoreSet.scala 493:25]
  reg [1:0] allocPtr_1; // @[StoreSet.scala 493:25]
  reg [1:0] allocPtr_2; // @[StoreSet.scala 493:25]
  reg [1:0] allocPtr_3; // @[StoreSet.scala 493:25]
  reg [1:0] allocPtr_4; // @[StoreSet.scala 493:25]
  reg [1:0] allocPtr_5; // @[StoreSet.scala 493:25]
  reg [1:0] allocPtr_6; // @[StoreSet.scala 493:25]
  reg [1:0] allocPtr_7; // @[StoreSet.scala 493:25]
  reg [1:0] allocPtr_8; // @[StoreSet.scala 493:25]
  reg [1:0] allocPtr_9; // @[StoreSet.scala 493:25]
  reg [1:0] allocPtr_10; // @[StoreSet.scala 493:25]
  reg [1:0] allocPtr_11; // @[StoreSet.scala 493:25]
  reg [1:0] allocPtr_12; // @[StoreSet.scala 493:25]
  reg [1:0] allocPtr_13; // @[StoreSet.scala 493:25]
  reg [1:0] allocPtr_14; // @[StoreSet.scala 493:25]
  reg [1:0] allocPtr_15; // @[StoreSet.scala 493:25]
  reg [1:0] allocPtr_16; // @[StoreSet.scala 493:25]
  reg [1:0] allocPtr_17; // @[StoreSet.scala 493:25]
  reg [1:0] allocPtr_18; // @[StoreSet.scala 493:25]
  reg [1:0] allocPtr_19; // @[StoreSet.scala 493:25]
  reg [1:0] allocPtr_20; // @[StoreSet.scala 493:25]
  reg [1:0] allocPtr_21; // @[StoreSet.scala 493:25]
  reg [1:0] allocPtr_22; // @[StoreSet.scala 493:25]
  reg [1:0] allocPtr_23; // @[StoreSet.scala 493:25]
  reg [1:0] allocPtr_24; // @[StoreSet.scala 493:25]
  reg [1:0] allocPtr_25; // @[StoreSet.scala 493:25]
  reg [1:0] allocPtr_26; // @[StoreSet.scala 493:25]
  reg [1:0] allocPtr_27; // @[StoreSet.scala 493:25]
  reg [1:0] allocPtr_28; // @[StoreSet.scala 493:25]
  reg [1:0] allocPtr_29; // @[StoreSet.scala 493:25]
  reg [1:0] allocPtr_30; // @[StoreSet.scala 493:25]
  reg [1:0] allocPtr_31; // @[StoreSet.scala 493:25]
  wire [3:0] _valid_0_T = {validVec_0_3,validVec_0_2,validVec_0_1,validVec_0_0}; // @[StoreSet.scala 496:29]
  wire  valid_0 = |_valid_0_T; // @[StoreSet.scala 496:36]
  wire [3:0] _valid_1_T = {validVec_1_3,validVec_1_2,validVec_1_1,validVec_1_0}; // @[StoreSet.scala 496:29]
  wire  valid_1 = |_valid_1_T; // @[StoreSet.scala 496:36]
  wire [3:0] _valid_2_T = {validVec_2_3,validVec_2_2,validVec_2_1,validVec_2_0}; // @[StoreSet.scala 496:29]
  wire  valid_2 = |_valid_2_T; // @[StoreSet.scala 496:36]
  wire [3:0] _valid_3_T = {validVec_3_3,validVec_3_2,validVec_3_1,validVec_3_0}; // @[StoreSet.scala 496:29]
  wire  valid_3 = |_valid_3_T; // @[StoreSet.scala 496:36]
  wire [3:0] _valid_4_T = {validVec_4_3,validVec_4_2,validVec_4_1,validVec_4_0}; // @[StoreSet.scala 496:29]
  wire  valid_4 = |_valid_4_T; // @[StoreSet.scala 496:36]
  wire [3:0] _valid_5_T = {validVec_5_3,validVec_5_2,validVec_5_1,validVec_5_0}; // @[StoreSet.scala 496:29]
  wire  valid_5 = |_valid_5_T; // @[StoreSet.scala 496:36]
  wire [3:0] _valid_6_T = {validVec_6_3,validVec_6_2,validVec_6_1,validVec_6_0}; // @[StoreSet.scala 496:29]
  wire  valid_6 = |_valid_6_T; // @[StoreSet.scala 496:36]
  wire [3:0] _valid_7_T = {validVec_7_3,validVec_7_2,validVec_7_1,validVec_7_0}; // @[StoreSet.scala 496:29]
  wire  valid_7 = |_valid_7_T; // @[StoreSet.scala 496:36]
  wire [3:0] _valid_8_T = {validVec_8_3,validVec_8_2,validVec_8_1,validVec_8_0}; // @[StoreSet.scala 496:29]
  wire  valid_8 = |_valid_8_T; // @[StoreSet.scala 496:36]
  wire [3:0] _valid_9_T = {validVec_9_3,validVec_9_2,validVec_9_1,validVec_9_0}; // @[StoreSet.scala 496:29]
  wire  valid_9 = |_valid_9_T; // @[StoreSet.scala 496:36]
  wire [3:0] _valid_10_T = {validVec_10_3,validVec_10_2,validVec_10_1,validVec_10_0}; // @[StoreSet.scala 496:29]
  wire  valid_10 = |_valid_10_T; // @[StoreSet.scala 496:36]
  wire [3:0] _valid_11_T = {validVec_11_3,validVec_11_2,validVec_11_1,validVec_11_0}; // @[StoreSet.scala 496:29]
  wire  valid_11 = |_valid_11_T; // @[StoreSet.scala 496:36]
  wire [3:0] _valid_12_T = {validVec_12_3,validVec_12_2,validVec_12_1,validVec_12_0}; // @[StoreSet.scala 496:29]
  wire  valid_12 = |_valid_12_T; // @[StoreSet.scala 496:36]
  wire [3:0] _valid_13_T = {validVec_13_3,validVec_13_2,validVec_13_1,validVec_13_0}; // @[StoreSet.scala 496:29]
  wire  valid_13 = |_valid_13_T; // @[StoreSet.scala 496:36]
  wire [3:0] _valid_14_T = {validVec_14_3,validVec_14_2,validVec_14_1,validVec_14_0}; // @[StoreSet.scala 496:29]
  wire  valid_14 = |_valid_14_T; // @[StoreSet.scala 496:36]
  wire [3:0] _valid_15_T = {validVec_15_3,validVec_15_2,validVec_15_1,validVec_15_0}; // @[StoreSet.scala 496:29]
  wire  valid_15 = |_valid_15_T; // @[StoreSet.scala 496:36]
  wire [3:0] _valid_16_T = {validVec_16_3,validVec_16_2,validVec_16_1,validVec_16_0}; // @[StoreSet.scala 496:29]
  wire  valid_16 = |_valid_16_T; // @[StoreSet.scala 496:36]
  wire [3:0] _valid_17_T = {validVec_17_3,validVec_17_2,validVec_17_1,validVec_17_0}; // @[StoreSet.scala 496:29]
  wire  valid_17 = |_valid_17_T; // @[StoreSet.scala 496:36]
  wire [3:0] _valid_18_T = {validVec_18_3,validVec_18_2,validVec_18_1,validVec_18_0}; // @[StoreSet.scala 496:29]
  wire  valid_18 = |_valid_18_T; // @[StoreSet.scala 496:36]
  wire [3:0] _valid_19_T = {validVec_19_3,validVec_19_2,validVec_19_1,validVec_19_0}; // @[StoreSet.scala 496:29]
  wire  valid_19 = |_valid_19_T; // @[StoreSet.scala 496:36]
  wire [3:0] _valid_20_T = {validVec_20_3,validVec_20_2,validVec_20_1,validVec_20_0}; // @[StoreSet.scala 496:29]
  wire  valid_20 = |_valid_20_T; // @[StoreSet.scala 496:36]
  wire [3:0] _valid_21_T = {validVec_21_3,validVec_21_2,validVec_21_1,validVec_21_0}; // @[StoreSet.scala 496:29]
  wire  valid_21 = |_valid_21_T; // @[StoreSet.scala 496:36]
  wire [3:0] _valid_22_T = {validVec_22_3,validVec_22_2,validVec_22_1,validVec_22_0}; // @[StoreSet.scala 496:29]
  wire  valid_22 = |_valid_22_T; // @[StoreSet.scala 496:36]
  wire [3:0] _valid_23_T = {validVec_23_3,validVec_23_2,validVec_23_1,validVec_23_0}; // @[StoreSet.scala 496:29]
  wire  valid_23 = |_valid_23_T; // @[StoreSet.scala 496:36]
  wire [3:0] _valid_24_T = {validVec_24_3,validVec_24_2,validVec_24_1,validVec_24_0}; // @[StoreSet.scala 496:29]
  wire  valid_24 = |_valid_24_T; // @[StoreSet.scala 496:36]
  wire [3:0] _valid_25_T = {validVec_25_3,validVec_25_2,validVec_25_1,validVec_25_0}; // @[StoreSet.scala 496:29]
  wire  valid_25 = |_valid_25_T; // @[StoreSet.scala 496:36]
  wire [3:0] _valid_26_T = {validVec_26_3,validVec_26_2,validVec_26_1,validVec_26_0}; // @[StoreSet.scala 496:29]
  wire  valid_26 = |_valid_26_T; // @[StoreSet.scala 496:36]
  wire [3:0] _valid_27_T = {validVec_27_3,validVec_27_2,validVec_27_1,validVec_27_0}; // @[StoreSet.scala 496:29]
  wire  valid_27 = |_valid_27_T; // @[StoreSet.scala 496:36]
  wire [3:0] _valid_28_T = {validVec_28_3,validVec_28_2,validVec_28_1,validVec_28_0}; // @[StoreSet.scala 496:29]
  wire  valid_28 = |_valid_28_T; // @[StoreSet.scala 496:36]
  wire [3:0] _valid_29_T = {validVec_29_3,validVec_29_2,validVec_29_1,validVec_29_0}; // @[StoreSet.scala 496:29]
  wire  valid_29 = |_valid_29_T; // @[StoreSet.scala 496:36]
  wire [3:0] _valid_30_T = {validVec_30_3,validVec_30_2,validVec_30_1,validVec_30_0}; // @[StoreSet.scala 496:29]
  wire  valid_30 = |_valid_30_T; // @[StoreSet.scala 496:36]
  wire [3:0] _valid_31_T = {validVec_31_3,validVec_31_2,validVec_31_1,validVec_31_0}; // @[StoreSet.scala 496:29]
  wire  valid_31 = |_valid_31_T; // @[StoreSet.scala 496:36]
  wire  _GEN_1 = 5'h1 == io_dispatch_req_0_bits_ssid ? valid_1 : valid_0; // @[StoreSet.scala 516:{46,46}]
  wire  _GEN_2 = 5'h2 == io_dispatch_req_0_bits_ssid ? valid_2 : _GEN_1; // @[StoreSet.scala 516:{46,46}]
  wire  _GEN_3 = 5'h3 == io_dispatch_req_0_bits_ssid ? valid_3 : _GEN_2; // @[StoreSet.scala 516:{46,46}]
  wire  _GEN_4 = 5'h4 == io_dispatch_req_0_bits_ssid ? valid_4 : _GEN_3; // @[StoreSet.scala 516:{46,46}]
  wire  _GEN_5 = 5'h5 == io_dispatch_req_0_bits_ssid ? valid_5 : _GEN_4; // @[StoreSet.scala 516:{46,46}]
  wire  _GEN_6 = 5'h6 == io_dispatch_req_0_bits_ssid ? valid_6 : _GEN_5; // @[StoreSet.scala 516:{46,46}]
  wire  _GEN_7 = 5'h7 == io_dispatch_req_0_bits_ssid ? valid_7 : _GEN_6; // @[StoreSet.scala 516:{46,46}]
  wire  _GEN_8 = 5'h8 == io_dispatch_req_0_bits_ssid ? valid_8 : _GEN_7; // @[StoreSet.scala 516:{46,46}]
  wire  _GEN_9 = 5'h9 == io_dispatch_req_0_bits_ssid ? valid_9 : _GEN_8; // @[StoreSet.scala 516:{46,46}]
  wire  _GEN_10 = 5'ha == io_dispatch_req_0_bits_ssid ? valid_10 : _GEN_9; // @[StoreSet.scala 516:{46,46}]
  wire  _GEN_11 = 5'hb == io_dispatch_req_0_bits_ssid ? valid_11 : _GEN_10; // @[StoreSet.scala 516:{46,46}]
  wire  _GEN_12 = 5'hc == io_dispatch_req_0_bits_ssid ? valid_12 : _GEN_11; // @[StoreSet.scala 516:{46,46}]
  wire  _GEN_13 = 5'hd == io_dispatch_req_0_bits_ssid ? valid_13 : _GEN_12; // @[StoreSet.scala 516:{46,46}]
  wire  _GEN_14 = 5'he == io_dispatch_req_0_bits_ssid ? valid_14 : _GEN_13; // @[StoreSet.scala 516:{46,46}]
  wire  _GEN_15 = 5'hf == io_dispatch_req_0_bits_ssid ? valid_15 : _GEN_14; // @[StoreSet.scala 516:{46,46}]
  wire  _GEN_16 = 5'h10 == io_dispatch_req_0_bits_ssid ? valid_16 : _GEN_15; // @[StoreSet.scala 516:{46,46}]
  wire  _GEN_17 = 5'h11 == io_dispatch_req_0_bits_ssid ? valid_17 : _GEN_16; // @[StoreSet.scala 516:{46,46}]
  wire  _GEN_18 = 5'h12 == io_dispatch_req_0_bits_ssid ? valid_18 : _GEN_17; // @[StoreSet.scala 516:{46,46}]
  wire  _GEN_19 = 5'h13 == io_dispatch_req_0_bits_ssid ? valid_19 : _GEN_18; // @[StoreSet.scala 516:{46,46}]
  wire  _GEN_20 = 5'h14 == io_dispatch_req_0_bits_ssid ? valid_20 : _GEN_19; // @[StoreSet.scala 516:{46,46}]
  wire  _GEN_21 = 5'h15 == io_dispatch_req_0_bits_ssid ? valid_21 : _GEN_20; // @[StoreSet.scala 516:{46,46}]
  wire  _GEN_22 = 5'h16 == io_dispatch_req_0_bits_ssid ? valid_22 : _GEN_21; // @[StoreSet.scala 516:{46,46}]
  wire  _GEN_23 = 5'h17 == io_dispatch_req_0_bits_ssid ? valid_23 : _GEN_22; // @[StoreSet.scala 516:{46,46}]
  wire  _GEN_24 = 5'h18 == io_dispatch_req_0_bits_ssid ? valid_24 : _GEN_23; // @[StoreSet.scala 516:{46,46}]
  wire  _GEN_25 = 5'h19 == io_dispatch_req_0_bits_ssid ? valid_25 : _GEN_24; // @[StoreSet.scala 516:{46,46}]
  wire  _GEN_26 = 5'h1a == io_dispatch_req_0_bits_ssid ? valid_26 : _GEN_25; // @[StoreSet.scala 516:{46,46}]
  wire  _GEN_27 = 5'h1b == io_dispatch_req_0_bits_ssid ? valid_27 : _GEN_26; // @[StoreSet.scala 516:{46,46}]
  wire  _GEN_28 = 5'h1c == io_dispatch_req_0_bits_ssid ? valid_28 : _GEN_27; // @[StoreSet.scala 516:{46,46}]
  wire  _GEN_29 = 5'h1d == io_dispatch_req_0_bits_ssid ? valid_29 : _GEN_28; // @[StoreSet.scala 516:{46,46}]
  wire  _GEN_30 = 5'h1e == io_dispatch_req_0_bits_ssid ? valid_30 : _GEN_29; // @[StoreSet.scala 516:{46,46}]
  wire  _GEN_31 = 5'h1f == io_dispatch_req_0_bits_ssid ? valid_31 : _GEN_30; // @[StoreSet.scala 516:{46,46}]
  wire  _io_dispatch_resp_0_bits_shouldWait_T_1 = _GEN_31 & io_dispatch_req_0_valid; // @[StoreSet.scala 516:70]
  wire  _io_dispatch_resp_0_bits_shouldWait_T_3 = ~io_dispatch_req_0_bits_isstore | io_csrCtrl_storeset_wait_store; // @[StoreSet.scala 518:43]
  wire  _io_dispatch_resp_0_bits_shouldWait_T_4 = _io_dispatch_resp_0_bits_shouldWait_T_1 &
    _io_dispatch_resp_0_bits_shouldWait_T_3; // @[StoreSet.scala 517:34]
  wire [1:0] _GEN_33 = 5'h1 == io_dispatch_req_0_bits_ssid ? allocPtr_1 : allocPtr_0; // @[StoreSet.scala 520:{118,118}]
  wire [1:0] _GEN_34 = 5'h2 == io_dispatch_req_0_bits_ssid ? allocPtr_2 : _GEN_33; // @[StoreSet.scala 520:{118,118}]
  wire [1:0] _GEN_35 = 5'h3 == io_dispatch_req_0_bits_ssid ? allocPtr_3 : _GEN_34; // @[StoreSet.scala 520:{118,118}]
  wire [1:0] _GEN_36 = 5'h4 == io_dispatch_req_0_bits_ssid ? allocPtr_4 : _GEN_35; // @[StoreSet.scala 520:{118,118}]
  wire [1:0] _GEN_37 = 5'h5 == io_dispatch_req_0_bits_ssid ? allocPtr_5 : _GEN_36; // @[StoreSet.scala 520:{118,118}]
  wire [1:0] _GEN_38 = 5'h6 == io_dispatch_req_0_bits_ssid ? allocPtr_6 : _GEN_37; // @[StoreSet.scala 520:{118,118}]
  wire [1:0] _GEN_39 = 5'h7 == io_dispatch_req_0_bits_ssid ? allocPtr_7 : _GEN_38; // @[StoreSet.scala 520:{118,118}]
  wire [1:0] _GEN_40 = 5'h8 == io_dispatch_req_0_bits_ssid ? allocPtr_8 : _GEN_39; // @[StoreSet.scala 520:{118,118}]
  wire [1:0] _GEN_41 = 5'h9 == io_dispatch_req_0_bits_ssid ? allocPtr_9 : _GEN_40; // @[StoreSet.scala 520:{118,118}]
  wire [1:0] _GEN_42 = 5'ha == io_dispatch_req_0_bits_ssid ? allocPtr_10 : _GEN_41; // @[StoreSet.scala 520:{118,118}]
  wire [1:0] _GEN_43 = 5'hb == io_dispatch_req_0_bits_ssid ? allocPtr_11 : _GEN_42; // @[StoreSet.scala 520:{118,118}]
  wire [1:0] _GEN_44 = 5'hc == io_dispatch_req_0_bits_ssid ? allocPtr_12 : _GEN_43; // @[StoreSet.scala 520:{118,118}]
  wire [1:0] _GEN_45 = 5'hd == io_dispatch_req_0_bits_ssid ? allocPtr_13 : _GEN_44; // @[StoreSet.scala 520:{118,118}]
  wire [1:0] _GEN_46 = 5'he == io_dispatch_req_0_bits_ssid ? allocPtr_14 : _GEN_45; // @[StoreSet.scala 520:{118,118}]
  wire [1:0] _GEN_47 = 5'hf == io_dispatch_req_0_bits_ssid ? allocPtr_15 : _GEN_46; // @[StoreSet.scala 520:{118,118}]
  wire [1:0] _GEN_48 = 5'h10 == io_dispatch_req_0_bits_ssid ? allocPtr_16 : _GEN_47; // @[StoreSet.scala 520:{118,118}]
  wire [1:0] _GEN_49 = 5'h11 == io_dispatch_req_0_bits_ssid ? allocPtr_17 : _GEN_48; // @[StoreSet.scala 520:{118,118}]
  wire [1:0] _GEN_50 = 5'h12 == io_dispatch_req_0_bits_ssid ? allocPtr_18 : _GEN_49; // @[StoreSet.scala 520:{118,118}]
  wire [1:0] _GEN_51 = 5'h13 == io_dispatch_req_0_bits_ssid ? allocPtr_19 : _GEN_50; // @[StoreSet.scala 520:{118,118}]
  wire [1:0] _GEN_52 = 5'h14 == io_dispatch_req_0_bits_ssid ? allocPtr_20 : _GEN_51; // @[StoreSet.scala 520:{118,118}]
  wire [1:0] _GEN_53 = 5'h15 == io_dispatch_req_0_bits_ssid ? allocPtr_21 : _GEN_52; // @[StoreSet.scala 520:{118,118}]
  wire [1:0] _GEN_54 = 5'h16 == io_dispatch_req_0_bits_ssid ? allocPtr_22 : _GEN_53; // @[StoreSet.scala 520:{118,118}]
  wire [1:0] _GEN_55 = 5'h17 == io_dispatch_req_0_bits_ssid ? allocPtr_23 : _GEN_54; // @[StoreSet.scala 520:{118,118}]
  wire [1:0] _GEN_56 = 5'h18 == io_dispatch_req_0_bits_ssid ? allocPtr_24 : _GEN_55; // @[StoreSet.scala 520:{118,118}]
  wire [1:0] _GEN_57 = 5'h19 == io_dispatch_req_0_bits_ssid ? allocPtr_25 : _GEN_56; // @[StoreSet.scala 520:{118,118}]
  wire [1:0] _GEN_58 = 5'h1a == io_dispatch_req_0_bits_ssid ? allocPtr_26 : _GEN_57; // @[StoreSet.scala 520:{118,118}]
  wire [1:0] _GEN_59 = 5'h1b == io_dispatch_req_0_bits_ssid ? allocPtr_27 : _GEN_58; // @[StoreSet.scala 520:{118,118}]
  wire [1:0] _GEN_60 = 5'h1c == io_dispatch_req_0_bits_ssid ? allocPtr_28 : _GEN_59; // @[StoreSet.scala 520:{118,118}]
  wire [1:0] _GEN_61 = 5'h1d == io_dispatch_req_0_bits_ssid ? allocPtr_29 : _GEN_60; // @[StoreSet.scala 520:{118,118}]
  wire [1:0] _GEN_62 = 5'h1e == io_dispatch_req_0_bits_ssid ? allocPtr_30 : _GEN_61; // @[StoreSet.scala 520:{118,118}]
  wire [1:0] _GEN_63 = 5'h1f == io_dispatch_req_0_bits_ssid ? allocPtr_31 : _GEN_62; // @[StoreSet.scala 520:{118,118}]
  wire [1:0] _io_dispatch_resp_0_bits_robIdx_T_1 = _GEN_63 - 2'h1; // @[StoreSet.scala 520:118]
  wire  _GEN_3874 = 5'h0 == io_dispatch_req_0_bits_ssid; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_65 = 5'h0 == io_dispatch_req_0_bits_ssid & 2'h1 == _io_dispatch_resp_0_bits_robIdx_T_1 ? robIdxVec_0_1_flag
     : robIdxVec_0_0_flag; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_66 = 5'h0 == io_dispatch_req_0_bits_ssid & 2'h2 == _io_dispatch_resp_0_bits_robIdx_T_1 ? robIdxVec_0_2_flag
     : _GEN_65; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_67 = 5'h0 == io_dispatch_req_0_bits_ssid & 2'h3 == _io_dispatch_resp_0_bits_robIdx_T_1 ? robIdxVec_0_3_flag
     : _GEN_66; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_3880 = 5'h1 == io_dispatch_req_0_bits_ssid; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_68 = 5'h1 == io_dispatch_req_0_bits_ssid & 2'h0 == _io_dispatch_resp_0_bits_robIdx_T_1 ? robIdxVec_1_0_flag
     : _GEN_67; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_69 = 5'h1 == io_dispatch_req_0_bits_ssid & 2'h1 == _io_dispatch_resp_0_bits_robIdx_T_1 ? robIdxVec_1_1_flag
     : _GEN_68; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_70 = 5'h1 == io_dispatch_req_0_bits_ssid & 2'h2 == _io_dispatch_resp_0_bits_robIdx_T_1 ? robIdxVec_1_2_flag
     : _GEN_69; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_71 = 5'h1 == io_dispatch_req_0_bits_ssid & 2'h3 == _io_dispatch_resp_0_bits_robIdx_T_1 ? robIdxVec_1_3_flag
     : _GEN_70; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_3888 = 5'h2 == io_dispatch_req_0_bits_ssid; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_72 = 5'h2 == io_dispatch_req_0_bits_ssid & 2'h0 == _io_dispatch_resp_0_bits_robIdx_T_1 ? robIdxVec_2_0_flag
     : _GEN_71; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_73 = 5'h2 == io_dispatch_req_0_bits_ssid & 2'h1 == _io_dispatch_resp_0_bits_robIdx_T_1 ? robIdxVec_2_1_flag
     : _GEN_72; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_74 = 5'h2 == io_dispatch_req_0_bits_ssid & 2'h2 == _io_dispatch_resp_0_bits_robIdx_T_1 ? robIdxVec_2_2_flag
     : _GEN_73; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_75 = 5'h2 == io_dispatch_req_0_bits_ssid & 2'h3 == _io_dispatch_resp_0_bits_robIdx_T_1 ? robIdxVec_2_3_flag
     : _GEN_74; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_3896 = 5'h3 == io_dispatch_req_0_bits_ssid; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_76 = 5'h3 == io_dispatch_req_0_bits_ssid & 2'h0 == _io_dispatch_resp_0_bits_robIdx_T_1 ? robIdxVec_3_0_flag
     : _GEN_75; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_77 = 5'h3 == io_dispatch_req_0_bits_ssid & 2'h1 == _io_dispatch_resp_0_bits_robIdx_T_1 ? robIdxVec_3_1_flag
     : _GEN_76; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_78 = 5'h3 == io_dispatch_req_0_bits_ssid & 2'h2 == _io_dispatch_resp_0_bits_robIdx_T_1 ? robIdxVec_3_2_flag
     : _GEN_77; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_79 = 5'h3 == io_dispatch_req_0_bits_ssid & 2'h3 == _io_dispatch_resp_0_bits_robIdx_T_1 ? robIdxVec_3_3_flag
     : _GEN_78; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_3904 = 5'h4 == io_dispatch_req_0_bits_ssid; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_80 = 5'h4 == io_dispatch_req_0_bits_ssid & 2'h0 == _io_dispatch_resp_0_bits_robIdx_T_1 ? robIdxVec_4_0_flag
     : _GEN_79; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_81 = 5'h4 == io_dispatch_req_0_bits_ssid & 2'h1 == _io_dispatch_resp_0_bits_robIdx_T_1 ? robIdxVec_4_1_flag
     : _GEN_80; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_82 = 5'h4 == io_dispatch_req_0_bits_ssid & 2'h2 == _io_dispatch_resp_0_bits_robIdx_T_1 ? robIdxVec_4_2_flag
     : _GEN_81; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_83 = 5'h4 == io_dispatch_req_0_bits_ssid & 2'h3 == _io_dispatch_resp_0_bits_robIdx_T_1 ? robIdxVec_4_3_flag
     : _GEN_82; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_3912 = 5'h5 == io_dispatch_req_0_bits_ssid; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_84 = 5'h5 == io_dispatch_req_0_bits_ssid & 2'h0 == _io_dispatch_resp_0_bits_robIdx_T_1 ? robIdxVec_5_0_flag
     : _GEN_83; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_85 = 5'h5 == io_dispatch_req_0_bits_ssid & 2'h1 == _io_dispatch_resp_0_bits_robIdx_T_1 ? robIdxVec_5_1_flag
     : _GEN_84; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_86 = 5'h5 == io_dispatch_req_0_bits_ssid & 2'h2 == _io_dispatch_resp_0_bits_robIdx_T_1 ? robIdxVec_5_2_flag
     : _GEN_85; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_87 = 5'h5 == io_dispatch_req_0_bits_ssid & 2'h3 == _io_dispatch_resp_0_bits_robIdx_T_1 ? robIdxVec_5_3_flag
     : _GEN_86; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_3920 = 5'h6 == io_dispatch_req_0_bits_ssid; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_88 = 5'h6 == io_dispatch_req_0_bits_ssid & 2'h0 == _io_dispatch_resp_0_bits_robIdx_T_1 ? robIdxVec_6_0_flag
     : _GEN_87; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_89 = 5'h6 == io_dispatch_req_0_bits_ssid & 2'h1 == _io_dispatch_resp_0_bits_robIdx_T_1 ? robIdxVec_6_1_flag
     : _GEN_88; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_90 = 5'h6 == io_dispatch_req_0_bits_ssid & 2'h2 == _io_dispatch_resp_0_bits_robIdx_T_1 ? robIdxVec_6_2_flag
     : _GEN_89; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_91 = 5'h6 == io_dispatch_req_0_bits_ssid & 2'h3 == _io_dispatch_resp_0_bits_robIdx_T_1 ? robIdxVec_6_3_flag
     : _GEN_90; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_3928 = 5'h7 == io_dispatch_req_0_bits_ssid; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_92 = 5'h7 == io_dispatch_req_0_bits_ssid & 2'h0 == _io_dispatch_resp_0_bits_robIdx_T_1 ? robIdxVec_7_0_flag
     : _GEN_91; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_93 = 5'h7 == io_dispatch_req_0_bits_ssid & 2'h1 == _io_dispatch_resp_0_bits_robIdx_T_1 ? robIdxVec_7_1_flag
     : _GEN_92; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_94 = 5'h7 == io_dispatch_req_0_bits_ssid & 2'h2 == _io_dispatch_resp_0_bits_robIdx_T_1 ? robIdxVec_7_2_flag
     : _GEN_93; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_95 = 5'h7 == io_dispatch_req_0_bits_ssid & 2'h3 == _io_dispatch_resp_0_bits_robIdx_T_1 ? robIdxVec_7_3_flag
     : _GEN_94; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_3936 = 5'h8 == io_dispatch_req_0_bits_ssid; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_96 = 5'h8 == io_dispatch_req_0_bits_ssid & 2'h0 == _io_dispatch_resp_0_bits_robIdx_T_1 ? robIdxVec_8_0_flag
     : _GEN_95; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_97 = 5'h8 == io_dispatch_req_0_bits_ssid & 2'h1 == _io_dispatch_resp_0_bits_robIdx_T_1 ? robIdxVec_8_1_flag
     : _GEN_96; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_98 = 5'h8 == io_dispatch_req_0_bits_ssid & 2'h2 == _io_dispatch_resp_0_bits_robIdx_T_1 ? robIdxVec_8_2_flag
     : _GEN_97; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_99 = 5'h8 == io_dispatch_req_0_bits_ssid & 2'h3 == _io_dispatch_resp_0_bits_robIdx_T_1 ? robIdxVec_8_3_flag
     : _GEN_98; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_3944 = 5'h9 == io_dispatch_req_0_bits_ssid; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_100 = 5'h9 == io_dispatch_req_0_bits_ssid & 2'h0 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_9_0_flag : _GEN_99; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_101 = 5'h9 == io_dispatch_req_0_bits_ssid & 2'h1 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_9_1_flag : _GEN_100; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_102 = 5'h9 == io_dispatch_req_0_bits_ssid & 2'h2 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_9_2_flag : _GEN_101; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_103 = 5'h9 == io_dispatch_req_0_bits_ssid & 2'h3 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_9_3_flag : _GEN_102; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_3952 = 5'ha == io_dispatch_req_0_bits_ssid; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_104 = 5'ha == io_dispatch_req_0_bits_ssid & 2'h0 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_10_0_flag : _GEN_103; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_105 = 5'ha == io_dispatch_req_0_bits_ssid & 2'h1 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_10_1_flag : _GEN_104; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_106 = 5'ha == io_dispatch_req_0_bits_ssid & 2'h2 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_10_2_flag : _GEN_105; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_107 = 5'ha == io_dispatch_req_0_bits_ssid & 2'h3 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_10_3_flag : _GEN_106; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_3960 = 5'hb == io_dispatch_req_0_bits_ssid; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_108 = 5'hb == io_dispatch_req_0_bits_ssid & 2'h0 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_11_0_flag : _GEN_107; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_109 = 5'hb == io_dispatch_req_0_bits_ssid & 2'h1 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_11_1_flag : _GEN_108; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_110 = 5'hb == io_dispatch_req_0_bits_ssid & 2'h2 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_11_2_flag : _GEN_109; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_111 = 5'hb == io_dispatch_req_0_bits_ssid & 2'h3 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_11_3_flag : _GEN_110; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_3968 = 5'hc == io_dispatch_req_0_bits_ssid; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_112 = 5'hc == io_dispatch_req_0_bits_ssid & 2'h0 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_12_0_flag : _GEN_111; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_113 = 5'hc == io_dispatch_req_0_bits_ssid & 2'h1 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_12_1_flag : _GEN_112; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_114 = 5'hc == io_dispatch_req_0_bits_ssid & 2'h2 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_12_2_flag : _GEN_113; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_115 = 5'hc == io_dispatch_req_0_bits_ssid & 2'h3 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_12_3_flag : _GEN_114; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_3976 = 5'hd == io_dispatch_req_0_bits_ssid; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_116 = 5'hd == io_dispatch_req_0_bits_ssid & 2'h0 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_13_0_flag : _GEN_115; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_117 = 5'hd == io_dispatch_req_0_bits_ssid & 2'h1 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_13_1_flag : _GEN_116; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_118 = 5'hd == io_dispatch_req_0_bits_ssid & 2'h2 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_13_2_flag : _GEN_117; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_119 = 5'hd == io_dispatch_req_0_bits_ssid & 2'h3 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_13_3_flag : _GEN_118; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_3984 = 5'he == io_dispatch_req_0_bits_ssid; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_120 = 5'he == io_dispatch_req_0_bits_ssid & 2'h0 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_14_0_flag : _GEN_119; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_121 = 5'he == io_dispatch_req_0_bits_ssid & 2'h1 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_14_1_flag : _GEN_120; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_122 = 5'he == io_dispatch_req_0_bits_ssid & 2'h2 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_14_2_flag : _GEN_121; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_123 = 5'he == io_dispatch_req_0_bits_ssid & 2'h3 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_14_3_flag : _GEN_122; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_3992 = 5'hf == io_dispatch_req_0_bits_ssid; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_124 = 5'hf == io_dispatch_req_0_bits_ssid & 2'h0 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_15_0_flag : _GEN_123; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_125 = 5'hf == io_dispatch_req_0_bits_ssid & 2'h1 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_15_1_flag : _GEN_124; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_126 = 5'hf == io_dispatch_req_0_bits_ssid & 2'h2 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_15_2_flag : _GEN_125; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_127 = 5'hf == io_dispatch_req_0_bits_ssid & 2'h3 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_15_3_flag : _GEN_126; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_4000 = 5'h10 == io_dispatch_req_0_bits_ssid; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_128 = 5'h10 == io_dispatch_req_0_bits_ssid & 2'h0 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_16_0_flag : _GEN_127; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_129 = 5'h10 == io_dispatch_req_0_bits_ssid & 2'h1 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_16_1_flag : _GEN_128; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_130 = 5'h10 == io_dispatch_req_0_bits_ssid & 2'h2 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_16_2_flag : _GEN_129; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_131 = 5'h10 == io_dispatch_req_0_bits_ssid & 2'h3 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_16_3_flag : _GEN_130; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_4008 = 5'h11 == io_dispatch_req_0_bits_ssid; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_132 = 5'h11 == io_dispatch_req_0_bits_ssid & 2'h0 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_17_0_flag : _GEN_131; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_133 = 5'h11 == io_dispatch_req_0_bits_ssid & 2'h1 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_17_1_flag : _GEN_132; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_134 = 5'h11 == io_dispatch_req_0_bits_ssid & 2'h2 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_17_2_flag : _GEN_133; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_135 = 5'h11 == io_dispatch_req_0_bits_ssid & 2'h3 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_17_3_flag : _GEN_134; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_4016 = 5'h12 == io_dispatch_req_0_bits_ssid; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_136 = 5'h12 == io_dispatch_req_0_bits_ssid & 2'h0 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_18_0_flag : _GEN_135; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_137 = 5'h12 == io_dispatch_req_0_bits_ssid & 2'h1 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_18_1_flag : _GEN_136; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_138 = 5'h12 == io_dispatch_req_0_bits_ssid & 2'h2 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_18_2_flag : _GEN_137; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_139 = 5'h12 == io_dispatch_req_0_bits_ssid & 2'h3 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_18_3_flag : _GEN_138; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_4024 = 5'h13 == io_dispatch_req_0_bits_ssid; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_140 = 5'h13 == io_dispatch_req_0_bits_ssid & 2'h0 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_19_0_flag : _GEN_139; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_141 = 5'h13 == io_dispatch_req_0_bits_ssid & 2'h1 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_19_1_flag : _GEN_140; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_142 = 5'h13 == io_dispatch_req_0_bits_ssid & 2'h2 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_19_2_flag : _GEN_141; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_143 = 5'h13 == io_dispatch_req_0_bits_ssid & 2'h3 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_19_3_flag : _GEN_142; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_4032 = 5'h14 == io_dispatch_req_0_bits_ssid; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_144 = 5'h14 == io_dispatch_req_0_bits_ssid & 2'h0 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_20_0_flag : _GEN_143; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_145 = 5'h14 == io_dispatch_req_0_bits_ssid & 2'h1 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_20_1_flag : _GEN_144; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_146 = 5'h14 == io_dispatch_req_0_bits_ssid & 2'h2 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_20_2_flag : _GEN_145; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_147 = 5'h14 == io_dispatch_req_0_bits_ssid & 2'h3 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_20_3_flag : _GEN_146; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_4040 = 5'h15 == io_dispatch_req_0_bits_ssid; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_148 = 5'h15 == io_dispatch_req_0_bits_ssid & 2'h0 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_21_0_flag : _GEN_147; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_149 = 5'h15 == io_dispatch_req_0_bits_ssid & 2'h1 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_21_1_flag : _GEN_148; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_150 = 5'h15 == io_dispatch_req_0_bits_ssid & 2'h2 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_21_2_flag : _GEN_149; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_151 = 5'h15 == io_dispatch_req_0_bits_ssid & 2'h3 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_21_3_flag : _GEN_150; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_4048 = 5'h16 == io_dispatch_req_0_bits_ssid; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_152 = 5'h16 == io_dispatch_req_0_bits_ssid & 2'h0 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_22_0_flag : _GEN_151; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_153 = 5'h16 == io_dispatch_req_0_bits_ssid & 2'h1 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_22_1_flag : _GEN_152; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_154 = 5'h16 == io_dispatch_req_0_bits_ssid & 2'h2 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_22_2_flag : _GEN_153; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_155 = 5'h16 == io_dispatch_req_0_bits_ssid & 2'h3 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_22_3_flag : _GEN_154; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_4056 = 5'h17 == io_dispatch_req_0_bits_ssid; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_156 = 5'h17 == io_dispatch_req_0_bits_ssid & 2'h0 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_23_0_flag : _GEN_155; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_157 = 5'h17 == io_dispatch_req_0_bits_ssid & 2'h1 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_23_1_flag : _GEN_156; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_158 = 5'h17 == io_dispatch_req_0_bits_ssid & 2'h2 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_23_2_flag : _GEN_157; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_159 = 5'h17 == io_dispatch_req_0_bits_ssid & 2'h3 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_23_3_flag : _GEN_158; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_4064 = 5'h18 == io_dispatch_req_0_bits_ssid; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_160 = 5'h18 == io_dispatch_req_0_bits_ssid & 2'h0 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_24_0_flag : _GEN_159; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_161 = 5'h18 == io_dispatch_req_0_bits_ssid & 2'h1 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_24_1_flag : _GEN_160; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_162 = 5'h18 == io_dispatch_req_0_bits_ssid & 2'h2 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_24_2_flag : _GEN_161; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_163 = 5'h18 == io_dispatch_req_0_bits_ssid & 2'h3 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_24_3_flag : _GEN_162; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_4072 = 5'h19 == io_dispatch_req_0_bits_ssid; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_164 = 5'h19 == io_dispatch_req_0_bits_ssid & 2'h0 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_25_0_flag : _GEN_163; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_165 = 5'h19 == io_dispatch_req_0_bits_ssid & 2'h1 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_25_1_flag : _GEN_164; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_166 = 5'h19 == io_dispatch_req_0_bits_ssid & 2'h2 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_25_2_flag : _GEN_165; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_167 = 5'h19 == io_dispatch_req_0_bits_ssid & 2'h3 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_25_3_flag : _GEN_166; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_4080 = 5'h1a == io_dispatch_req_0_bits_ssid; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_168 = 5'h1a == io_dispatch_req_0_bits_ssid & 2'h0 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_26_0_flag : _GEN_167; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_169 = 5'h1a == io_dispatch_req_0_bits_ssid & 2'h1 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_26_1_flag : _GEN_168; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_170 = 5'h1a == io_dispatch_req_0_bits_ssid & 2'h2 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_26_2_flag : _GEN_169; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_171 = 5'h1a == io_dispatch_req_0_bits_ssid & 2'h3 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_26_3_flag : _GEN_170; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_4088 = 5'h1b == io_dispatch_req_0_bits_ssid; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_172 = 5'h1b == io_dispatch_req_0_bits_ssid & 2'h0 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_27_0_flag : _GEN_171; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_173 = 5'h1b == io_dispatch_req_0_bits_ssid & 2'h1 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_27_1_flag : _GEN_172; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_174 = 5'h1b == io_dispatch_req_0_bits_ssid & 2'h2 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_27_2_flag : _GEN_173; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_175 = 5'h1b == io_dispatch_req_0_bits_ssid & 2'h3 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_27_3_flag : _GEN_174; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_4096 = 5'h1c == io_dispatch_req_0_bits_ssid; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_176 = 5'h1c == io_dispatch_req_0_bits_ssid & 2'h0 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_28_0_flag : _GEN_175; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_177 = 5'h1c == io_dispatch_req_0_bits_ssid & 2'h1 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_28_1_flag : _GEN_176; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_178 = 5'h1c == io_dispatch_req_0_bits_ssid & 2'h2 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_28_2_flag : _GEN_177; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_179 = 5'h1c == io_dispatch_req_0_bits_ssid & 2'h3 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_28_3_flag : _GEN_178; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_4104 = 5'h1d == io_dispatch_req_0_bits_ssid; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_180 = 5'h1d == io_dispatch_req_0_bits_ssid & 2'h0 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_29_0_flag : _GEN_179; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_181 = 5'h1d == io_dispatch_req_0_bits_ssid & 2'h1 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_29_1_flag : _GEN_180; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_182 = 5'h1d == io_dispatch_req_0_bits_ssid & 2'h2 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_29_2_flag : _GEN_181; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_183 = 5'h1d == io_dispatch_req_0_bits_ssid & 2'h3 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_29_3_flag : _GEN_182; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_4112 = 5'h1e == io_dispatch_req_0_bits_ssid; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_184 = 5'h1e == io_dispatch_req_0_bits_ssid & 2'h0 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_30_0_flag : _GEN_183; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_185 = 5'h1e == io_dispatch_req_0_bits_ssid & 2'h1 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_30_1_flag : _GEN_184; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_186 = 5'h1e == io_dispatch_req_0_bits_ssid & 2'h2 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_30_2_flag : _GEN_185; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_187 = 5'h1e == io_dispatch_req_0_bits_ssid & 2'h3 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_30_3_flag : _GEN_186; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_4120 = 5'h1f == io_dispatch_req_0_bits_ssid; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_188 = 5'h1f == io_dispatch_req_0_bits_ssid & 2'h0 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_31_0_flag : _GEN_187; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_189 = 5'h1f == io_dispatch_req_0_bits_ssid & 2'h1 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_31_1_flag : _GEN_188; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_190 = 5'h1f == io_dispatch_req_0_bits_ssid & 2'h2 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_31_2_flag : _GEN_189; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_193 = 5'h0 == io_dispatch_req_0_bits_ssid & 2'h1 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_0_1_value : robIdxVec_0_0_value; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_194 = 5'h0 == io_dispatch_req_0_bits_ssid & 2'h2 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_0_2_value : _GEN_193; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_195 = 5'h0 == io_dispatch_req_0_bits_ssid & 2'h3 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_0_3_value : _GEN_194; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_196 = 5'h1 == io_dispatch_req_0_bits_ssid & 2'h0 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_1_0_value : _GEN_195; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_197 = 5'h1 == io_dispatch_req_0_bits_ssid & 2'h1 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_1_1_value : _GEN_196; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_198 = 5'h1 == io_dispatch_req_0_bits_ssid & 2'h2 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_1_2_value : _GEN_197; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_199 = 5'h1 == io_dispatch_req_0_bits_ssid & 2'h3 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_1_3_value : _GEN_198; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_200 = 5'h2 == io_dispatch_req_0_bits_ssid & 2'h0 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_2_0_value : _GEN_199; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_201 = 5'h2 == io_dispatch_req_0_bits_ssid & 2'h1 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_2_1_value : _GEN_200; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_202 = 5'h2 == io_dispatch_req_0_bits_ssid & 2'h2 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_2_2_value : _GEN_201; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_203 = 5'h2 == io_dispatch_req_0_bits_ssid & 2'h3 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_2_3_value : _GEN_202; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_204 = 5'h3 == io_dispatch_req_0_bits_ssid & 2'h0 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_3_0_value : _GEN_203; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_205 = 5'h3 == io_dispatch_req_0_bits_ssid & 2'h1 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_3_1_value : _GEN_204; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_206 = 5'h3 == io_dispatch_req_0_bits_ssid & 2'h2 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_3_2_value : _GEN_205; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_207 = 5'h3 == io_dispatch_req_0_bits_ssid & 2'h3 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_3_3_value : _GEN_206; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_208 = 5'h4 == io_dispatch_req_0_bits_ssid & 2'h0 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_4_0_value : _GEN_207; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_209 = 5'h4 == io_dispatch_req_0_bits_ssid & 2'h1 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_4_1_value : _GEN_208; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_210 = 5'h4 == io_dispatch_req_0_bits_ssid & 2'h2 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_4_2_value : _GEN_209; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_211 = 5'h4 == io_dispatch_req_0_bits_ssid & 2'h3 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_4_3_value : _GEN_210; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_212 = 5'h5 == io_dispatch_req_0_bits_ssid & 2'h0 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_5_0_value : _GEN_211; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_213 = 5'h5 == io_dispatch_req_0_bits_ssid & 2'h1 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_5_1_value : _GEN_212; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_214 = 5'h5 == io_dispatch_req_0_bits_ssid & 2'h2 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_5_2_value : _GEN_213; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_215 = 5'h5 == io_dispatch_req_0_bits_ssid & 2'h3 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_5_3_value : _GEN_214; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_216 = 5'h6 == io_dispatch_req_0_bits_ssid & 2'h0 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_6_0_value : _GEN_215; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_217 = 5'h6 == io_dispatch_req_0_bits_ssid & 2'h1 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_6_1_value : _GEN_216; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_218 = 5'h6 == io_dispatch_req_0_bits_ssid & 2'h2 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_6_2_value : _GEN_217; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_219 = 5'h6 == io_dispatch_req_0_bits_ssid & 2'h3 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_6_3_value : _GEN_218; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_220 = 5'h7 == io_dispatch_req_0_bits_ssid & 2'h0 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_7_0_value : _GEN_219; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_221 = 5'h7 == io_dispatch_req_0_bits_ssid & 2'h1 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_7_1_value : _GEN_220; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_222 = 5'h7 == io_dispatch_req_0_bits_ssid & 2'h2 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_7_2_value : _GEN_221; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_223 = 5'h7 == io_dispatch_req_0_bits_ssid & 2'h3 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_7_3_value : _GEN_222; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_224 = 5'h8 == io_dispatch_req_0_bits_ssid & 2'h0 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_8_0_value : _GEN_223; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_225 = 5'h8 == io_dispatch_req_0_bits_ssid & 2'h1 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_8_1_value : _GEN_224; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_226 = 5'h8 == io_dispatch_req_0_bits_ssid & 2'h2 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_8_2_value : _GEN_225; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_227 = 5'h8 == io_dispatch_req_0_bits_ssid & 2'h3 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_8_3_value : _GEN_226; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_228 = 5'h9 == io_dispatch_req_0_bits_ssid & 2'h0 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_9_0_value : _GEN_227; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_229 = 5'h9 == io_dispatch_req_0_bits_ssid & 2'h1 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_9_1_value : _GEN_228; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_230 = 5'h9 == io_dispatch_req_0_bits_ssid & 2'h2 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_9_2_value : _GEN_229; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_231 = 5'h9 == io_dispatch_req_0_bits_ssid & 2'h3 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_9_3_value : _GEN_230; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_232 = 5'ha == io_dispatch_req_0_bits_ssid & 2'h0 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_10_0_value : _GEN_231; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_233 = 5'ha == io_dispatch_req_0_bits_ssid & 2'h1 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_10_1_value : _GEN_232; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_234 = 5'ha == io_dispatch_req_0_bits_ssid & 2'h2 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_10_2_value : _GEN_233; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_235 = 5'ha == io_dispatch_req_0_bits_ssid & 2'h3 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_10_3_value : _GEN_234; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_236 = 5'hb == io_dispatch_req_0_bits_ssid & 2'h0 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_11_0_value : _GEN_235; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_237 = 5'hb == io_dispatch_req_0_bits_ssid & 2'h1 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_11_1_value : _GEN_236; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_238 = 5'hb == io_dispatch_req_0_bits_ssid & 2'h2 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_11_2_value : _GEN_237; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_239 = 5'hb == io_dispatch_req_0_bits_ssid & 2'h3 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_11_3_value : _GEN_238; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_240 = 5'hc == io_dispatch_req_0_bits_ssid & 2'h0 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_12_0_value : _GEN_239; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_241 = 5'hc == io_dispatch_req_0_bits_ssid & 2'h1 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_12_1_value : _GEN_240; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_242 = 5'hc == io_dispatch_req_0_bits_ssid & 2'h2 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_12_2_value : _GEN_241; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_243 = 5'hc == io_dispatch_req_0_bits_ssid & 2'h3 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_12_3_value : _GEN_242; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_244 = 5'hd == io_dispatch_req_0_bits_ssid & 2'h0 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_13_0_value : _GEN_243; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_245 = 5'hd == io_dispatch_req_0_bits_ssid & 2'h1 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_13_1_value : _GEN_244; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_246 = 5'hd == io_dispatch_req_0_bits_ssid & 2'h2 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_13_2_value : _GEN_245; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_247 = 5'hd == io_dispatch_req_0_bits_ssid & 2'h3 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_13_3_value : _GEN_246; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_248 = 5'he == io_dispatch_req_0_bits_ssid & 2'h0 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_14_0_value : _GEN_247; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_249 = 5'he == io_dispatch_req_0_bits_ssid & 2'h1 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_14_1_value : _GEN_248; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_250 = 5'he == io_dispatch_req_0_bits_ssid & 2'h2 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_14_2_value : _GEN_249; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_251 = 5'he == io_dispatch_req_0_bits_ssid & 2'h3 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_14_3_value : _GEN_250; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_252 = 5'hf == io_dispatch_req_0_bits_ssid & 2'h0 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_15_0_value : _GEN_251; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_253 = 5'hf == io_dispatch_req_0_bits_ssid & 2'h1 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_15_1_value : _GEN_252; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_254 = 5'hf == io_dispatch_req_0_bits_ssid & 2'h2 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_15_2_value : _GEN_253; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_255 = 5'hf == io_dispatch_req_0_bits_ssid & 2'h3 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_15_3_value : _GEN_254; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_256 = 5'h10 == io_dispatch_req_0_bits_ssid & 2'h0 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_16_0_value : _GEN_255; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_257 = 5'h10 == io_dispatch_req_0_bits_ssid & 2'h1 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_16_1_value : _GEN_256; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_258 = 5'h10 == io_dispatch_req_0_bits_ssid & 2'h2 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_16_2_value : _GEN_257; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_259 = 5'h10 == io_dispatch_req_0_bits_ssid & 2'h3 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_16_3_value : _GEN_258; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_260 = 5'h11 == io_dispatch_req_0_bits_ssid & 2'h0 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_17_0_value : _GEN_259; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_261 = 5'h11 == io_dispatch_req_0_bits_ssid & 2'h1 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_17_1_value : _GEN_260; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_262 = 5'h11 == io_dispatch_req_0_bits_ssid & 2'h2 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_17_2_value : _GEN_261; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_263 = 5'h11 == io_dispatch_req_0_bits_ssid & 2'h3 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_17_3_value : _GEN_262; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_264 = 5'h12 == io_dispatch_req_0_bits_ssid & 2'h0 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_18_0_value : _GEN_263; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_265 = 5'h12 == io_dispatch_req_0_bits_ssid & 2'h1 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_18_1_value : _GEN_264; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_266 = 5'h12 == io_dispatch_req_0_bits_ssid & 2'h2 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_18_2_value : _GEN_265; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_267 = 5'h12 == io_dispatch_req_0_bits_ssid & 2'h3 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_18_3_value : _GEN_266; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_268 = 5'h13 == io_dispatch_req_0_bits_ssid & 2'h0 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_19_0_value : _GEN_267; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_269 = 5'h13 == io_dispatch_req_0_bits_ssid & 2'h1 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_19_1_value : _GEN_268; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_270 = 5'h13 == io_dispatch_req_0_bits_ssid & 2'h2 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_19_2_value : _GEN_269; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_271 = 5'h13 == io_dispatch_req_0_bits_ssid & 2'h3 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_19_3_value : _GEN_270; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_272 = 5'h14 == io_dispatch_req_0_bits_ssid & 2'h0 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_20_0_value : _GEN_271; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_273 = 5'h14 == io_dispatch_req_0_bits_ssid & 2'h1 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_20_1_value : _GEN_272; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_274 = 5'h14 == io_dispatch_req_0_bits_ssid & 2'h2 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_20_2_value : _GEN_273; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_275 = 5'h14 == io_dispatch_req_0_bits_ssid & 2'h3 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_20_3_value : _GEN_274; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_276 = 5'h15 == io_dispatch_req_0_bits_ssid & 2'h0 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_21_0_value : _GEN_275; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_277 = 5'h15 == io_dispatch_req_0_bits_ssid & 2'h1 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_21_1_value : _GEN_276; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_278 = 5'h15 == io_dispatch_req_0_bits_ssid & 2'h2 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_21_2_value : _GEN_277; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_279 = 5'h15 == io_dispatch_req_0_bits_ssid & 2'h3 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_21_3_value : _GEN_278; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_280 = 5'h16 == io_dispatch_req_0_bits_ssid & 2'h0 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_22_0_value : _GEN_279; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_281 = 5'h16 == io_dispatch_req_0_bits_ssid & 2'h1 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_22_1_value : _GEN_280; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_282 = 5'h16 == io_dispatch_req_0_bits_ssid & 2'h2 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_22_2_value : _GEN_281; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_283 = 5'h16 == io_dispatch_req_0_bits_ssid & 2'h3 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_22_3_value : _GEN_282; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_284 = 5'h17 == io_dispatch_req_0_bits_ssid & 2'h0 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_23_0_value : _GEN_283; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_285 = 5'h17 == io_dispatch_req_0_bits_ssid & 2'h1 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_23_1_value : _GEN_284; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_286 = 5'h17 == io_dispatch_req_0_bits_ssid & 2'h2 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_23_2_value : _GEN_285; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_287 = 5'h17 == io_dispatch_req_0_bits_ssid & 2'h3 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_23_3_value : _GEN_286; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_288 = 5'h18 == io_dispatch_req_0_bits_ssid & 2'h0 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_24_0_value : _GEN_287; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_289 = 5'h18 == io_dispatch_req_0_bits_ssid & 2'h1 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_24_1_value : _GEN_288; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_290 = 5'h18 == io_dispatch_req_0_bits_ssid & 2'h2 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_24_2_value : _GEN_289; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_291 = 5'h18 == io_dispatch_req_0_bits_ssid & 2'h3 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_24_3_value : _GEN_290; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_292 = 5'h19 == io_dispatch_req_0_bits_ssid & 2'h0 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_25_0_value : _GEN_291; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_293 = 5'h19 == io_dispatch_req_0_bits_ssid & 2'h1 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_25_1_value : _GEN_292; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_294 = 5'h19 == io_dispatch_req_0_bits_ssid & 2'h2 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_25_2_value : _GEN_293; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_295 = 5'h19 == io_dispatch_req_0_bits_ssid & 2'h3 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_25_3_value : _GEN_294; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_296 = 5'h1a == io_dispatch_req_0_bits_ssid & 2'h0 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_26_0_value : _GEN_295; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_297 = 5'h1a == io_dispatch_req_0_bits_ssid & 2'h1 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_26_1_value : _GEN_296; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_298 = 5'h1a == io_dispatch_req_0_bits_ssid & 2'h2 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_26_2_value : _GEN_297; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_299 = 5'h1a == io_dispatch_req_0_bits_ssid & 2'h3 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_26_3_value : _GEN_298; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_300 = 5'h1b == io_dispatch_req_0_bits_ssid & 2'h0 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_27_0_value : _GEN_299; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_301 = 5'h1b == io_dispatch_req_0_bits_ssid & 2'h1 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_27_1_value : _GEN_300; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_302 = 5'h1b == io_dispatch_req_0_bits_ssid & 2'h2 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_27_2_value : _GEN_301; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_303 = 5'h1b == io_dispatch_req_0_bits_ssid & 2'h3 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_27_3_value : _GEN_302; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_304 = 5'h1c == io_dispatch_req_0_bits_ssid & 2'h0 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_28_0_value : _GEN_303; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_305 = 5'h1c == io_dispatch_req_0_bits_ssid & 2'h1 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_28_1_value : _GEN_304; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_306 = 5'h1c == io_dispatch_req_0_bits_ssid & 2'h2 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_28_2_value : _GEN_305; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_307 = 5'h1c == io_dispatch_req_0_bits_ssid & 2'h3 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_28_3_value : _GEN_306; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_308 = 5'h1d == io_dispatch_req_0_bits_ssid & 2'h0 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_29_0_value : _GEN_307; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_309 = 5'h1d == io_dispatch_req_0_bits_ssid & 2'h1 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_29_1_value : _GEN_308; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_310 = 5'h1d == io_dispatch_req_0_bits_ssid & 2'h2 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_29_2_value : _GEN_309; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_311 = 5'h1d == io_dispatch_req_0_bits_ssid & 2'h3 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_29_3_value : _GEN_310; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_312 = 5'h1e == io_dispatch_req_0_bits_ssid & 2'h0 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_30_0_value : _GEN_311; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_313 = 5'h1e == io_dispatch_req_0_bits_ssid & 2'h1 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_30_1_value : _GEN_312; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_314 = 5'h1e == io_dispatch_req_0_bits_ssid & 2'h2 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_30_2_value : _GEN_313; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_315 = 5'h1e == io_dispatch_req_0_bits_ssid & 2'h3 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_30_3_value : _GEN_314; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_316 = 5'h1f == io_dispatch_req_0_bits_ssid & 2'h0 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_31_0_value : _GEN_315; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_317 = 5'h1f == io_dispatch_req_0_bits_ssid & 2'h1 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_31_1_value : _GEN_316; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_318 = 5'h1f == io_dispatch_req_0_bits_ssid & 2'h2 == _io_dispatch_resp_0_bits_robIdx_T_1 ?
    robIdxVec_31_2_value : _GEN_317; // @[StoreSet.scala 520:{37,37}]
  wire  _hitInDispatchBundleVec_T = io_dispatch_req_0_valid & io_dispatch_req_0_bits_isstore; // @[StoreSet.scala 506:34]
  wire  _hitInDispatchBundleVec_T_1 = io_dispatch_req_0_bits_ssid == io_dispatch_req_1_bits_ssid; // @[StoreSet.scala 508:38]
  wire  hitInDispatchBundleVec_1_0 = _hitInDispatchBundleVec_T & _hitInDispatchBundleVec_T_1; // @[StoreSet.scala 507:41]
  wire  hitInDispatchBundle_1 = |hitInDispatchBundleVec_1_0; // @[StoreSet.scala 513:61]
  wire  _GEN_321 = 5'h1 == io_dispatch_req_1_bits_ssid ? valid_1 : valid_0; // @[StoreSet.scala 516:{46,46}]
  wire  _GEN_322 = 5'h2 == io_dispatch_req_1_bits_ssid ? valid_2 : _GEN_321; // @[StoreSet.scala 516:{46,46}]
  wire  _GEN_323 = 5'h3 == io_dispatch_req_1_bits_ssid ? valid_3 : _GEN_322; // @[StoreSet.scala 516:{46,46}]
  wire  _GEN_324 = 5'h4 == io_dispatch_req_1_bits_ssid ? valid_4 : _GEN_323; // @[StoreSet.scala 516:{46,46}]
  wire  _GEN_325 = 5'h5 == io_dispatch_req_1_bits_ssid ? valid_5 : _GEN_324; // @[StoreSet.scala 516:{46,46}]
  wire  _GEN_326 = 5'h6 == io_dispatch_req_1_bits_ssid ? valid_6 : _GEN_325; // @[StoreSet.scala 516:{46,46}]
  wire  _GEN_327 = 5'h7 == io_dispatch_req_1_bits_ssid ? valid_7 : _GEN_326; // @[StoreSet.scala 516:{46,46}]
  wire  _GEN_328 = 5'h8 == io_dispatch_req_1_bits_ssid ? valid_8 : _GEN_327; // @[StoreSet.scala 516:{46,46}]
  wire  _GEN_329 = 5'h9 == io_dispatch_req_1_bits_ssid ? valid_9 : _GEN_328; // @[StoreSet.scala 516:{46,46}]
  wire  _GEN_330 = 5'ha == io_dispatch_req_1_bits_ssid ? valid_10 : _GEN_329; // @[StoreSet.scala 516:{46,46}]
  wire  _GEN_331 = 5'hb == io_dispatch_req_1_bits_ssid ? valid_11 : _GEN_330; // @[StoreSet.scala 516:{46,46}]
  wire  _GEN_332 = 5'hc == io_dispatch_req_1_bits_ssid ? valid_12 : _GEN_331; // @[StoreSet.scala 516:{46,46}]
  wire  _GEN_333 = 5'hd == io_dispatch_req_1_bits_ssid ? valid_13 : _GEN_332; // @[StoreSet.scala 516:{46,46}]
  wire  _GEN_334 = 5'he == io_dispatch_req_1_bits_ssid ? valid_14 : _GEN_333; // @[StoreSet.scala 516:{46,46}]
  wire  _GEN_335 = 5'hf == io_dispatch_req_1_bits_ssid ? valid_15 : _GEN_334; // @[StoreSet.scala 516:{46,46}]
  wire  _GEN_336 = 5'h10 == io_dispatch_req_1_bits_ssid ? valid_16 : _GEN_335; // @[StoreSet.scala 516:{46,46}]
  wire  _GEN_337 = 5'h11 == io_dispatch_req_1_bits_ssid ? valid_17 : _GEN_336; // @[StoreSet.scala 516:{46,46}]
  wire  _GEN_338 = 5'h12 == io_dispatch_req_1_bits_ssid ? valid_18 : _GEN_337; // @[StoreSet.scala 516:{46,46}]
  wire  _GEN_339 = 5'h13 == io_dispatch_req_1_bits_ssid ? valid_19 : _GEN_338; // @[StoreSet.scala 516:{46,46}]
  wire  _GEN_340 = 5'h14 == io_dispatch_req_1_bits_ssid ? valid_20 : _GEN_339; // @[StoreSet.scala 516:{46,46}]
  wire  _GEN_341 = 5'h15 == io_dispatch_req_1_bits_ssid ? valid_21 : _GEN_340; // @[StoreSet.scala 516:{46,46}]
  wire  _GEN_342 = 5'h16 == io_dispatch_req_1_bits_ssid ? valid_22 : _GEN_341; // @[StoreSet.scala 516:{46,46}]
  wire  _GEN_343 = 5'h17 == io_dispatch_req_1_bits_ssid ? valid_23 : _GEN_342; // @[StoreSet.scala 516:{46,46}]
  wire  _GEN_344 = 5'h18 == io_dispatch_req_1_bits_ssid ? valid_24 : _GEN_343; // @[StoreSet.scala 516:{46,46}]
  wire  _GEN_345 = 5'h19 == io_dispatch_req_1_bits_ssid ? valid_25 : _GEN_344; // @[StoreSet.scala 516:{46,46}]
  wire  _GEN_346 = 5'h1a == io_dispatch_req_1_bits_ssid ? valid_26 : _GEN_345; // @[StoreSet.scala 516:{46,46}]
  wire  _GEN_347 = 5'h1b == io_dispatch_req_1_bits_ssid ? valid_27 : _GEN_346; // @[StoreSet.scala 516:{46,46}]
  wire  _GEN_348 = 5'h1c == io_dispatch_req_1_bits_ssid ? valid_28 : _GEN_347; // @[StoreSet.scala 516:{46,46}]
  wire  _GEN_349 = 5'h1d == io_dispatch_req_1_bits_ssid ? valid_29 : _GEN_348; // @[StoreSet.scala 516:{46,46}]
  wire  _GEN_350 = 5'h1e == io_dispatch_req_1_bits_ssid ? valid_30 : _GEN_349; // @[StoreSet.scala 516:{46,46}]
  wire  _GEN_351 = 5'h1f == io_dispatch_req_1_bits_ssid ? valid_31 : _GEN_350; // @[StoreSet.scala 516:{46,46}]
  wire  _io_dispatch_resp_1_bits_shouldWait_T_1 = (_GEN_351 | hitInDispatchBundle_1) & io_dispatch_req_1_valid; // @[StoreSet.scala 516:70]
  wire  _io_dispatch_resp_1_bits_shouldWait_T_3 = ~io_dispatch_req_1_bits_isstore | io_csrCtrl_storeset_wait_store; // @[StoreSet.scala 518:43]
  wire  _io_dispatch_resp_1_bits_shouldWait_T_4 = _io_dispatch_resp_1_bits_shouldWait_T_1 &
    _io_dispatch_resp_1_bits_shouldWait_T_3; // @[StoreSet.scala 517:34]
  wire [1:0] _GEN_353 = 5'h1 == io_dispatch_req_1_bits_ssid ? allocPtr_1 : allocPtr_0; // @[StoreSet.scala 520:{118,118}]
  wire [1:0] _GEN_354 = 5'h2 == io_dispatch_req_1_bits_ssid ? allocPtr_2 : _GEN_353; // @[StoreSet.scala 520:{118,118}]
  wire [1:0] _GEN_355 = 5'h3 == io_dispatch_req_1_bits_ssid ? allocPtr_3 : _GEN_354; // @[StoreSet.scala 520:{118,118}]
  wire [1:0] _GEN_356 = 5'h4 == io_dispatch_req_1_bits_ssid ? allocPtr_4 : _GEN_355; // @[StoreSet.scala 520:{118,118}]
  wire [1:0] _GEN_357 = 5'h5 == io_dispatch_req_1_bits_ssid ? allocPtr_5 : _GEN_356; // @[StoreSet.scala 520:{118,118}]
  wire [1:0] _GEN_358 = 5'h6 == io_dispatch_req_1_bits_ssid ? allocPtr_6 : _GEN_357; // @[StoreSet.scala 520:{118,118}]
  wire [1:0] _GEN_359 = 5'h7 == io_dispatch_req_1_bits_ssid ? allocPtr_7 : _GEN_358; // @[StoreSet.scala 520:{118,118}]
  wire [1:0] _GEN_360 = 5'h8 == io_dispatch_req_1_bits_ssid ? allocPtr_8 : _GEN_359; // @[StoreSet.scala 520:{118,118}]
  wire [1:0] _GEN_361 = 5'h9 == io_dispatch_req_1_bits_ssid ? allocPtr_9 : _GEN_360; // @[StoreSet.scala 520:{118,118}]
  wire [1:0] _GEN_362 = 5'ha == io_dispatch_req_1_bits_ssid ? allocPtr_10 : _GEN_361; // @[StoreSet.scala 520:{118,118}]
  wire [1:0] _GEN_363 = 5'hb == io_dispatch_req_1_bits_ssid ? allocPtr_11 : _GEN_362; // @[StoreSet.scala 520:{118,118}]
  wire [1:0] _GEN_364 = 5'hc == io_dispatch_req_1_bits_ssid ? allocPtr_12 : _GEN_363; // @[StoreSet.scala 520:{118,118}]
  wire [1:0] _GEN_365 = 5'hd == io_dispatch_req_1_bits_ssid ? allocPtr_13 : _GEN_364; // @[StoreSet.scala 520:{118,118}]
  wire [1:0] _GEN_366 = 5'he == io_dispatch_req_1_bits_ssid ? allocPtr_14 : _GEN_365; // @[StoreSet.scala 520:{118,118}]
  wire [1:0] _GEN_367 = 5'hf == io_dispatch_req_1_bits_ssid ? allocPtr_15 : _GEN_366; // @[StoreSet.scala 520:{118,118}]
  wire [1:0] _GEN_368 = 5'h10 == io_dispatch_req_1_bits_ssid ? allocPtr_16 : _GEN_367; // @[StoreSet.scala 520:{118,118}]
  wire [1:0] _GEN_369 = 5'h11 == io_dispatch_req_1_bits_ssid ? allocPtr_17 : _GEN_368; // @[StoreSet.scala 520:{118,118}]
  wire [1:0] _GEN_370 = 5'h12 == io_dispatch_req_1_bits_ssid ? allocPtr_18 : _GEN_369; // @[StoreSet.scala 520:{118,118}]
  wire [1:0] _GEN_371 = 5'h13 == io_dispatch_req_1_bits_ssid ? allocPtr_19 : _GEN_370; // @[StoreSet.scala 520:{118,118}]
  wire [1:0] _GEN_372 = 5'h14 == io_dispatch_req_1_bits_ssid ? allocPtr_20 : _GEN_371; // @[StoreSet.scala 520:{118,118}]
  wire [1:0] _GEN_373 = 5'h15 == io_dispatch_req_1_bits_ssid ? allocPtr_21 : _GEN_372; // @[StoreSet.scala 520:{118,118}]
  wire [1:0] _GEN_374 = 5'h16 == io_dispatch_req_1_bits_ssid ? allocPtr_22 : _GEN_373; // @[StoreSet.scala 520:{118,118}]
  wire [1:0] _GEN_375 = 5'h17 == io_dispatch_req_1_bits_ssid ? allocPtr_23 : _GEN_374; // @[StoreSet.scala 520:{118,118}]
  wire [1:0] _GEN_376 = 5'h18 == io_dispatch_req_1_bits_ssid ? allocPtr_24 : _GEN_375; // @[StoreSet.scala 520:{118,118}]
  wire [1:0] _GEN_377 = 5'h19 == io_dispatch_req_1_bits_ssid ? allocPtr_25 : _GEN_376; // @[StoreSet.scala 520:{118,118}]
  wire [1:0] _GEN_378 = 5'h1a == io_dispatch_req_1_bits_ssid ? allocPtr_26 : _GEN_377; // @[StoreSet.scala 520:{118,118}]
  wire [1:0] _GEN_379 = 5'h1b == io_dispatch_req_1_bits_ssid ? allocPtr_27 : _GEN_378; // @[StoreSet.scala 520:{118,118}]
  wire [1:0] _GEN_380 = 5'h1c == io_dispatch_req_1_bits_ssid ? allocPtr_28 : _GEN_379; // @[StoreSet.scala 520:{118,118}]
  wire [1:0] _GEN_381 = 5'h1d == io_dispatch_req_1_bits_ssid ? allocPtr_29 : _GEN_380; // @[StoreSet.scala 520:{118,118}]
  wire [1:0] _GEN_382 = 5'h1e == io_dispatch_req_1_bits_ssid ? allocPtr_30 : _GEN_381; // @[StoreSet.scala 520:{118,118}]
  wire [1:0] _GEN_383 = 5'h1f == io_dispatch_req_1_bits_ssid ? allocPtr_31 : _GEN_382; // @[StoreSet.scala 520:{118,118}]
  wire [1:0] _io_dispatch_resp_1_bits_robIdx_T_1 = _GEN_383 - 2'h1; // @[StoreSet.scala 520:118]
  wire  _GEN_4382 = 5'h0 == io_dispatch_req_1_bits_ssid; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_385 = 5'h0 == io_dispatch_req_1_bits_ssid & 2'h1 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_0_1_flag : robIdxVec_0_0_flag; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_386 = 5'h0 == io_dispatch_req_1_bits_ssid & 2'h2 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_0_2_flag : _GEN_385; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_387 = 5'h0 == io_dispatch_req_1_bits_ssid & 2'h3 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_0_3_flag : _GEN_386; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_4388 = 5'h1 == io_dispatch_req_1_bits_ssid; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_388 = 5'h1 == io_dispatch_req_1_bits_ssid & 2'h0 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_1_0_flag : _GEN_387; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_389 = 5'h1 == io_dispatch_req_1_bits_ssid & 2'h1 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_1_1_flag : _GEN_388; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_390 = 5'h1 == io_dispatch_req_1_bits_ssid & 2'h2 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_1_2_flag : _GEN_389; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_391 = 5'h1 == io_dispatch_req_1_bits_ssid & 2'h3 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_1_3_flag : _GEN_390; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_4396 = 5'h2 == io_dispatch_req_1_bits_ssid; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_392 = 5'h2 == io_dispatch_req_1_bits_ssid & 2'h0 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_2_0_flag : _GEN_391; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_393 = 5'h2 == io_dispatch_req_1_bits_ssid & 2'h1 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_2_1_flag : _GEN_392; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_394 = 5'h2 == io_dispatch_req_1_bits_ssid & 2'h2 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_2_2_flag : _GEN_393; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_395 = 5'h2 == io_dispatch_req_1_bits_ssid & 2'h3 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_2_3_flag : _GEN_394; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_4404 = 5'h3 == io_dispatch_req_1_bits_ssid; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_396 = 5'h3 == io_dispatch_req_1_bits_ssid & 2'h0 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_3_0_flag : _GEN_395; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_397 = 5'h3 == io_dispatch_req_1_bits_ssid & 2'h1 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_3_1_flag : _GEN_396; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_398 = 5'h3 == io_dispatch_req_1_bits_ssid & 2'h2 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_3_2_flag : _GEN_397; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_399 = 5'h3 == io_dispatch_req_1_bits_ssid & 2'h3 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_3_3_flag : _GEN_398; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_4412 = 5'h4 == io_dispatch_req_1_bits_ssid; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_400 = 5'h4 == io_dispatch_req_1_bits_ssid & 2'h0 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_4_0_flag : _GEN_399; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_401 = 5'h4 == io_dispatch_req_1_bits_ssid & 2'h1 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_4_1_flag : _GEN_400; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_402 = 5'h4 == io_dispatch_req_1_bits_ssid & 2'h2 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_4_2_flag : _GEN_401; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_403 = 5'h4 == io_dispatch_req_1_bits_ssid & 2'h3 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_4_3_flag : _GEN_402; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_4420 = 5'h5 == io_dispatch_req_1_bits_ssid; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_404 = 5'h5 == io_dispatch_req_1_bits_ssid & 2'h0 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_5_0_flag : _GEN_403; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_405 = 5'h5 == io_dispatch_req_1_bits_ssid & 2'h1 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_5_1_flag : _GEN_404; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_406 = 5'h5 == io_dispatch_req_1_bits_ssid & 2'h2 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_5_2_flag : _GEN_405; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_407 = 5'h5 == io_dispatch_req_1_bits_ssid & 2'h3 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_5_3_flag : _GEN_406; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_4428 = 5'h6 == io_dispatch_req_1_bits_ssid; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_408 = 5'h6 == io_dispatch_req_1_bits_ssid & 2'h0 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_6_0_flag : _GEN_407; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_409 = 5'h6 == io_dispatch_req_1_bits_ssid & 2'h1 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_6_1_flag : _GEN_408; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_410 = 5'h6 == io_dispatch_req_1_bits_ssid & 2'h2 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_6_2_flag : _GEN_409; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_411 = 5'h6 == io_dispatch_req_1_bits_ssid & 2'h3 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_6_3_flag : _GEN_410; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_4436 = 5'h7 == io_dispatch_req_1_bits_ssid; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_412 = 5'h7 == io_dispatch_req_1_bits_ssid & 2'h0 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_7_0_flag : _GEN_411; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_413 = 5'h7 == io_dispatch_req_1_bits_ssid & 2'h1 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_7_1_flag : _GEN_412; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_414 = 5'h7 == io_dispatch_req_1_bits_ssid & 2'h2 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_7_2_flag : _GEN_413; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_415 = 5'h7 == io_dispatch_req_1_bits_ssid & 2'h3 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_7_3_flag : _GEN_414; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_4444 = 5'h8 == io_dispatch_req_1_bits_ssid; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_416 = 5'h8 == io_dispatch_req_1_bits_ssid & 2'h0 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_8_0_flag : _GEN_415; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_417 = 5'h8 == io_dispatch_req_1_bits_ssid & 2'h1 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_8_1_flag : _GEN_416; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_418 = 5'h8 == io_dispatch_req_1_bits_ssid & 2'h2 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_8_2_flag : _GEN_417; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_419 = 5'h8 == io_dispatch_req_1_bits_ssid & 2'h3 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_8_3_flag : _GEN_418; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_4452 = 5'h9 == io_dispatch_req_1_bits_ssid; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_420 = 5'h9 == io_dispatch_req_1_bits_ssid & 2'h0 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_9_0_flag : _GEN_419; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_421 = 5'h9 == io_dispatch_req_1_bits_ssid & 2'h1 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_9_1_flag : _GEN_420; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_422 = 5'h9 == io_dispatch_req_1_bits_ssid & 2'h2 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_9_2_flag : _GEN_421; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_423 = 5'h9 == io_dispatch_req_1_bits_ssid & 2'h3 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_9_3_flag : _GEN_422; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_4460 = 5'ha == io_dispatch_req_1_bits_ssid; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_424 = 5'ha == io_dispatch_req_1_bits_ssid & 2'h0 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_10_0_flag : _GEN_423; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_425 = 5'ha == io_dispatch_req_1_bits_ssid & 2'h1 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_10_1_flag : _GEN_424; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_426 = 5'ha == io_dispatch_req_1_bits_ssid & 2'h2 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_10_2_flag : _GEN_425; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_427 = 5'ha == io_dispatch_req_1_bits_ssid & 2'h3 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_10_3_flag : _GEN_426; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_4468 = 5'hb == io_dispatch_req_1_bits_ssid; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_428 = 5'hb == io_dispatch_req_1_bits_ssid & 2'h0 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_11_0_flag : _GEN_427; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_429 = 5'hb == io_dispatch_req_1_bits_ssid & 2'h1 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_11_1_flag : _GEN_428; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_430 = 5'hb == io_dispatch_req_1_bits_ssid & 2'h2 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_11_2_flag : _GEN_429; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_431 = 5'hb == io_dispatch_req_1_bits_ssid & 2'h3 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_11_3_flag : _GEN_430; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_4476 = 5'hc == io_dispatch_req_1_bits_ssid; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_432 = 5'hc == io_dispatch_req_1_bits_ssid & 2'h0 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_12_0_flag : _GEN_431; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_433 = 5'hc == io_dispatch_req_1_bits_ssid & 2'h1 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_12_1_flag : _GEN_432; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_434 = 5'hc == io_dispatch_req_1_bits_ssid & 2'h2 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_12_2_flag : _GEN_433; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_435 = 5'hc == io_dispatch_req_1_bits_ssid & 2'h3 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_12_3_flag : _GEN_434; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_4484 = 5'hd == io_dispatch_req_1_bits_ssid; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_436 = 5'hd == io_dispatch_req_1_bits_ssid & 2'h0 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_13_0_flag : _GEN_435; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_437 = 5'hd == io_dispatch_req_1_bits_ssid & 2'h1 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_13_1_flag : _GEN_436; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_438 = 5'hd == io_dispatch_req_1_bits_ssid & 2'h2 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_13_2_flag : _GEN_437; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_439 = 5'hd == io_dispatch_req_1_bits_ssid & 2'h3 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_13_3_flag : _GEN_438; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_4492 = 5'he == io_dispatch_req_1_bits_ssid; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_440 = 5'he == io_dispatch_req_1_bits_ssid & 2'h0 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_14_0_flag : _GEN_439; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_441 = 5'he == io_dispatch_req_1_bits_ssid & 2'h1 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_14_1_flag : _GEN_440; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_442 = 5'he == io_dispatch_req_1_bits_ssid & 2'h2 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_14_2_flag : _GEN_441; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_443 = 5'he == io_dispatch_req_1_bits_ssid & 2'h3 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_14_3_flag : _GEN_442; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_4500 = 5'hf == io_dispatch_req_1_bits_ssid; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_444 = 5'hf == io_dispatch_req_1_bits_ssid & 2'h0 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_15_0_flag : _GEN_443; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_445 = 5'hf == io_dispatch_req_1_bits_ssid & 2'h1 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_15_1_flag : _GEN_444; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_446 = 5'hf == io_dispatch_req_1_bits_ssid & 2'h2 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_15_2_flag : _GEN_445; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_447 = 5'hf == io_dispatch_req_1_bits_ssid & 2'h3 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_15_3_flag : _GEN_446; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_4508 = 5'h10 == io_dispatch_req_1_bits_ssid; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_448 = 5'h10 == io_dispatch_req_1_bits_ssid & 2'h0 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_16_0_flag : _GEN_447; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_449 = 5'h10 == io_dispatch_req_1_bits_ssid & 2'h1 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_16_1_flag : _GEN_448; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_450 = 5'h10 == io_dispatch_req_1_bits_ssid & 2'h2 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_16_2_flag : _GEN_449; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_451 = 5'h10 == io_dispatch_req_1_bits_ssid & 2'h3 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_16_3_flag : _GEN_450; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_4516 = 5'h11 == io_dispatch_req_1_bits_ssid; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_452 = 5'h11 == io_dispatch_req_1_bits_ssid & 2'h0 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_17_0_flag : _GEN_451; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_453 = 5'h11 == io_dispatch_req_1_bits_ssid & 2'h1 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_17_1_flag : _GEN_452; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_454 = 5'h11 == io_dispatch_req_1_bits_ssid & 2'h2 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_17_2_flag : _GEN_453; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_455 = 5'h11 == io_dispatch_req_1_bits_ssid & 2'h3 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_17_3_flag : _GEN_454; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_4524 = 5'h12 == io_dispatch_req_1_bits_ssid; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_456 = 5'h12 == io_dispatch_req_1_bits_ssid & 2'h0 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_18_0_flag : _GEN_455; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_457 = 5'h12 == io_dispatch_req_1_bits_ssid & 2'h1 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_18_1_flag : _GEN_456; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_458 = 5'h12 == io_dispatch_req_1_bits_ssid & 2'h2 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_18_2_flag : _GEN_457; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_459 = 5'h12 == io_dispatch_req_1_bits_ssid & 2'h3 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_18_3_flag : _GEN_458; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_4532 = 5'h13 == io_dispatch_req_1_bits_ssid; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_460 = 5'h13 == io_dispatch_req_1_bits_ssid & 2'h0 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_19_0_flag : _GEN_459; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_461 = 5'h13 == io_dispatch_req_1_bits_ssid & 2'h1 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_19_1_flag : _GEN_460; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_462 = 5'h13 == io_dispatch_req_1_bits_ssid & 2'h2 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_19_2_flag : _GEN_461; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_463 = 5'h13 == io_dispatch_req_1_bits_ssid & 2'h3 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_19_3_flag : _GEN_462; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_4540 = 5'h14 == io_dispatch_req_1_bits_ssid; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_464 = 5'h14 == io_dispatch_req_1_bits_ssid & 2'h0 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_20_0_flag : _GEN_463; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_465 = 5'h14 == io_dispatch_req_1_bits_ssid & 2'h1 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_20_1_flag : _GEN_464; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_466 = 5'h14 == io_dispatch_req_1_bits_ssid & 2'h2 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_20_2_flag : _GEN_465; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_467 = 5'h14 == io_dispatch_req_1_bits_ssid & 2'h3 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_20_3_flag : _GEN_466; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_4548 = 5'h15 == io_dispatch_req_1_bits_ssid; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_468 = 5'h15 == io_dispatch_req_1_bits_ssid & 2'h0 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_21_0_flag : _GEN_467; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_469 = 5'h15 == io_dispatch_req_1_bits_ssid & 2'h1 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_21_1_flag : _GEN_468; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_470 = 5'h15 == io_dispatch_req_1_bits_ssid & 2'h2 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_21_2_flag : _GEN_469; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_471 = 5'h15 == io_dispatch_req_1_bits_ssid & 2'h3 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_21_3_flag : _GEN_470; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_4556 = 5'h16 == io_dispatch_req_1_bits_ssid; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_472 = 5'h16 == io_dispatch_req_1_bits_ssid & 2'h0 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_22_0_flag : _GEN_471; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_473 = 5'h16 == io_dispatch_req_1_bits_ssid & 2'h1 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_22_1_flag : _GEN_472; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_474 = 5'h16 == io_dispatch_req_1_bits_ssid & 2'h2 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_22_2_flag : _GEN_473; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_475 = 5'h16 == io_dispatch_req_1_bits_ssid & 2'h3 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_22_3_flag : _GEN_474; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_4564 = 5'h17 == io_dispatch_req_1_bits_ssid; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_476 = 5'h17 == io_dispatch_req_1_bits_ssid & 2'h0 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_23_0_flag : _GEN_475; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_477 = 5'h17 == io_dispatch_req_1_bits_ssid & 2'h1 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_23_1_flag : _GEN_476; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_478 = 5'h17 == io_dispatch_req_1_bits_ssid & 2'h2 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_23_2_flag : _GEN_477; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_479 = 5'h17 == io_dispatch_req_1_bits_ssid & 2'h3 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_23_3_flag : _GEN_478; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_4572 = 5'h18 == io_dispatch_req_1_bits_ssid; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_480 = 5'h18 == io_dispatch_req_1_bits_ssid & 2'h0 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_24_0_flag : _GEN_479; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_481 = 5'h18 == io_dispatch_req_1_bits_ssid & 2'h1 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_24_1_flag : _GEN_480; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_482 = 5'h18 == io_dispatch_req_1_bits_ssid & 2'h2 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_24_2_flag : _GEN_481; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_483 = 5'h18 == io_dispatch_req_1_bits_ssid & 2'h3 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_24_3_flag : _GEN_482; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_4580 = 5'h19 == io_dispatch_req_1_bits_ssid; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_484 = 5'h19 == io_dispatch_req_1_bits_ssid & 2'h0 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_25_0_flag : _GEN_483; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_485 = 5'h19 == io_dispatch_req_1_bits_ssid & 2'h1 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_25_1_flag : _GEN_484; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_486 = 5'h19 == io_dispatch_req_1_bits_ssid & 2'h2 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_25_2_flag : _GEN_485; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_487 = 5'h19 == io_dispatch_req_1_bits_ssid & 2'h3 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_25_3_flag : _GEN_486; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_4588 = 5'h1a == io_dispatch_req_1_bits_ssid; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_488 = 5'h1a == io_dispatch_req_1_bits_ssid & 2'h0 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_26_0_flag : _GEN_487; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_489 = 5'h1a == io_dispatch_req_1_bits_ssid & 2'h1 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_26_1_flag : _GEN_488; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_490 = 5'h1a == io_dispatch_req_1_bits_ssid & 2'h2 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_26_2_flag : _GEN_489; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_491 = 5'h1a == io_dispatch_req_1_bits_ssid & 2'h3 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_26_3_flag : _GEN_490; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_4596 = 5'h1b == io_dispatch_req_1_bits_ssid; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_492 = 5'h1b == io_dispatch_req_1_bits_ssid & 2'h0 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_27_0_flag : _GEN_491; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_493 = 5'h1b == io_dispatch_req_1_bits_ssid & 2'h1 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_27_1_flag : _GEN_492; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_494 = 5'h1b == io_dispatch_req_1_bits_ssid & 2'h2 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_27_2_flag : _GEN_493; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_495 = 5'h1b == io_dispatch_req_1_bits_ssid & 2'h3 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_27_3_flag : _GEN_494; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_4604 = 5'h1c == io_dispatch_req_1_bits_ssid; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_496 = 5'h1c == io_dispatch_req_1_bits_ssid & 2'h0 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_28_0_flag : _GEN_495; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_497 = 5'h1c == io_dispatch_req_1_bits_ssid & 2'h1 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_28_1_flag : _GEN_496; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_498 = 5'h1c == io_dispatch_req_1_bits_ssid & 2'h2 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_28_2_flag : _GEN_497; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_499 = 5'h1c == io_dispatch_req_1_bits_ssid & 2'h3 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_28_3_flag : _GEN_498; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_4612 = 5'h1d == io_dispatch_req_1_bits_ssid; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_500 = 5'h1d == io_dispatch_req_1_bits_ssid & 2'h0 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_29_0_flag : _GEN_499; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_501 = 5'h1d == io_dispatch_req_1_bits_ssid & 2'h1 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_29_1_flag : _GEN_500; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_502 = 5'h1d == io_dispatch_req_1_bits_ssid & 2'h2 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_29_2_flag : _GEN_501; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_503 = 5'h1d == io_dispatch_req_1_bits_ssid & 2'h3 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_29_3_flag : _GEN_502; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_4620 = 5'h1e == io_dispatch_req_1_bits_ssid; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_504 = 5'h1e == io_dispatch_req_1_bits_ssid & 2'h0 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_30_0_flag : _GEN_503; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_505 = 5'h1e == io_dispatch_req_1_bits_ssid & 2'h1 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_30_1_flag : _GEN_504; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_506 = 5'h1e == io_dispatch_req_1_bits_ssid & 2'h2 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_30_2_flag : _GEN_505; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_507 = 5'h1e == io_dispatch_req_1_bits_ssid & 2'h3 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_30_3_flag : _GEN_506; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_4628 = 5'h1f == io_dispatch_req_1_bits_ssid; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_508 = 5'h1f == io_dispatch_req_1_bits_ssid & 2'h0 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_31_0_flag : _GEN_507; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_509 = 5'h1f == io_dispatch_req_1_bits_ssid & 2'h1 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_31_1_flag : _GEN_508; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_510 = 5'h1f == io_dispatch_req_1_bits_ssid & 2'h2 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_31_2_flag : _GEN_509; // @[StoreSet.scala 520:{37,37}]
  wire  _GEN_511 = 5'h1f == io_dispatch_req_1_bits_ssid & 2'h3 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_31_3_flag : _GEN_510; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_513 = 5'h0 == io_dispatch_req_1_bits_ssid & 2'h1 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_0_1_value : robIdxVec_0_0_value; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_514 = 5'h0 == io_dispatch_req_1_bits_ssid & 2'h2 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_0_2_value : _GEN_513; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_515 = 5'h0 == io_dispatch_req_1_bits_ssid & 2'h3 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_0_3_value : _GEN_514; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_516 = 5'h1 == io_dispatch_req_1_bits_ssid & 2'h0 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_1_0_value : _GEN_515; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_517 = 5'h1 == io_dispatch_req_1_bits_ssid & 2'h1 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_1_1_value : _GEN_516; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_518 = 5'h1 == io_dispatch_req_1_bits_ssid & 2'h2 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_1_2_value : _GEN_517; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_519 = 5'h1 == io_dispatch_req_1_bits_ssid & 2'h3 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_1_3_value : _GEN_518; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_520 = 5'h2 == io_dispatch_req_1_bits_ssid & 2'h0 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_2_0_value : _GEN_519; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_521 = 5'h2 == io_dispatch_req_1_bits_ssid & 2'h1 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_2_1_value : _GEN_520; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_522 = 5'h2 == io_dispatch_req_1_bits_ssid & 2'h2 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_2_2_value : _GEN_521; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_523 = 5'h2 == io_dispatch_req_1_bits_ssid & 2'h3 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_2_3_value : _GEN_522; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_524 = 5'h3 == io_dispatch_req_1_bits_ssid & 2'h0 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_3_0_value : _GEN_523; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_525 = 5'h3 == io_dispatch_req_1_bits_ssid & 2'h1 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_3_1_value : _GEN_524; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_526 = 5'h3 == io_dispatch_req_1_bits_ssid & 2'h2 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_3_2_value : _GEN_525; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_527 = 5'h3 == io_dispatch_req_1_bits_ssid & 2'h3 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_3_3_value : _GEN_526; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_528 = 5'h4 == io_dispatch_req_1_bits_ssid & 2'h0 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_4_0_value : _GEN_527; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_529 = 5'h4 == io_dispatch_req_1_bits_ssid & 2'h1 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_4_1_value : _GEN_528; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_530 = 5'h4 == io_dispatch_req_1_bits_ssid & 2'h2 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_4_2_value : _GEN_529; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_531 = 5'h4 == io_dispatch_req_1_bits_ssid & 2'h3 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_4_3_value : _GEN_530; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_532 = 5'h5 == io_dispatch_req_1_bits_ssid & 2'h0 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_5_0_value : _GEN_531; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_533 = 5'h5 == io_dispatch_req_1_bits_ssid & 2'h1 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_5_1_value : _GEN_532; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_534 = 5'h5 == io_dispatch_req_1_bits_ssid & 2'h2 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_5_2_value : _GEN_533; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_535 = 5'h5 == io_dispatch_req_1_bits_ssid & 2'h3 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_5_3_value : _GEN_534; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_536 = 5'h6 == io_dispatch_req_1_bits_ssid & 2'h0 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_6_0_value : _GEN_535; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_537 = 5'h6 == io_dispatch_req_1_bits_ssid & 2'h1 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_6_1_value : _GEN_536; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_538 = 5'h6 == io_dispatch_req_1_bits_ssid & 2'h2 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_6_2_value : _GEN_537; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_539 = 5'h6 == io_dispatch_req_1_bits_ssid & 2'h3 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_6_3_value : _GEN_538; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_540 = 5'h7 == io_dispatch_req_1_bits_ssid & 2'h0 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_7_0_value : _GEN_539; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_541 = 5'h7 == io_dispatch_req_1_bits_ssid & 2'h1 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_7_1_value : _GEN_540; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_542 = 5'h7 == io_dispatch_req_1_bits_ssid & 2'h2 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_7_2_value : _GEN_541; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_543 = 5'h7 == io_dispatch_req_1_bits_ssid & 2'h3 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_7_3_value : _GEN_542; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_544 = 5'h8 == io_dispatch_req_1_bits_ssid & 2'h0 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_8_0_value : _GEN_543; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_545 = 5'h8 == io_dispatch_req_1_bits_ssid & 2'h1 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_8_1_value : _GEN_544; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_546 = 5'h8 == io_dispatch_req_1_bits_ssid & 2'h2 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_8_2_value : _GEN_545; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_547 = 5'h8 == io_dispatch_req_1_bits_ssid & 2'h3 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_8_3_value : _GEN_546; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_548 = 5'h9 == io_dispatch_req_1_bits_ssid & 2'h0 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_9_0_value : _GEN_547; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_549 = 5'h9 == io_dispatch_req_1_bits_ssid & 2'h1 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_9_1_value : _GEN_548; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_550 = 5'h9 == io_dispatch_req_1_bits_ssid & 2'h2 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_9_2_value : _GEN_549; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_551 = 5'h9 == io_dispatch_req_1_bits_ssid & 2'h3 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_9_3_value : _GEN_550; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_552 = 5'ha == io_dispatch_req_1_bits_ssid & 2'h0 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_10_0_value : _GEN_551; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_553 = 5'ha == io_dispatch_req_1_bits_ssid & 2'h1 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_10_1_value : _GEN_552; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_554 = 5'ha == io_dispatch_req_1_bits_ssid & 2'h2 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_10_2_value : _GEN_553; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_555 = 5'ha == io_dispatch_req_1_bits_ssid & 2'h3 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_10_3_value : _GEN_554; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_556 = 5'hb == io_dispatch_req_1_bits_ssid & 2'h0 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_11_0_value : _GEN_555; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_557 = 5'hb == io_dispatch_req_1_bits_ssid & 2'h1 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_11_1_value : _GEN_556; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_558 = 5'hb == io_dispatch_req_1_bits_ssid & 2'h2 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_11_2_value : _GEN_557; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_559 = 5'hb == io_dispatch_req_1_bits_ssid & 2'h3 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_11_3_value : _GEN_558; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_560 = 5'hc == io_dispatch_req_1_bits_ssid & 2'h0 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_12_0_value : _GEN_559; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_561 = 5'hc == io_dispatch_req_1_bits_ssid & 2'h1 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_12_1_value : _GEN_560; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_562 = 5'hc == io_dispatch_req_1_bits_ssid & 2'h2 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_12_2_value : _GEN_561; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_563 = 5'hc == io_dispatch_req_1_bits_ssid & 2'h3 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_12_3_value : _GEN_562; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_564 = 5'hd == io_dispatch_req_1_bits_ssid & 2'h0 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_13_0_value : _GEN_563; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_565 = 5'hd == io_dispatch_req_1_bits_ssid & 2'h1 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_13_1_value : _GEN_564; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_566 = 5'hd == io_dispatch_req_1_bits_ssid & 2'h2 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_13_2_value : _GEN_565; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_567 = 5'hd == io_dispatch_req_1_bits_ssid & 2'h3 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_13_3_value : _GEN_566; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_568 = 5'he == io_dispatch_req_1_bits_ssid & 2'h0 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_14_0_value : _GEN_567; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_569 = 5'he == io_dispatch_req_1_bits_ssid & 2'h1 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_14_1_value : _GEN_568; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_570 = 5'he == io_dispatch_req_1_bits_ssid & 2'h2 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_14_2_value : _GEN_569; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_571 = 5'he == io_dispatch_req_1_bits_ssid & 2'h3 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_14_3_value : _GEN_570; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_572 = 5'hf == io_dispatch_req_1_bits_ssid & 2'h0 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_15_0_value : _GEN_571; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_573 = 5'hf == io_dispatch_req_1_bits_ssid & 2'h1 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_15_1_value : _GEN_572; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_574 = 5'hf == io_dispatch_req_1_bits_ssid & 2'h2 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_15_2_value : _GEN_573; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_575 = 5'hf == io_dispatch_req_1_bits_ssid & 2'h3 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_15_3_value : _GEN_574; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_576 = 5'h10 == io_dispatch_req_1_bits_ssid & 2'h0 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_16_0_value : _GEN_575; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_577 = 5'h10 == io_dispatch_req_1_bits_ssid & 2'h1 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_16_1_value : _GEN_576; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_578 = 5'h10 == io_dispatch_req_1_bits_ssid & 2'h2 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_16_2_value : _GEN_577; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_579 = 5'h10 == io_dispatch_req_1_bits_ssid & 2'h3 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_16_3_value : _GEN_578; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_580 = 5'h11 == io_dispatch_req_1_bits_ssid & 2'h0 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_17_0_value : _GEN_579; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_581 = 5'h11 == io_dispatch_req_1_bits_ssid & 2'h1 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_17_1_value : _GEN_580; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_582 = 5'h11 == io_dispatch_req_1_bits_ssid & 2'h2 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_17_2_value : _GEN_581; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_583 = 5'h11 == io_dispatch_req_1_bits_ssid & 2'h3 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_17_3_value : _GEN_582; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_584 = 5'h12 == io_dispatch_req_1_bits_ssid & 2'h0 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_18_0_value : _GEN_583; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_585 = 5'h12 == io_dispatch_req_1_bits_ssid & 2'h1 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_18_1_value : _GEN_584; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_586 = 5'h12 == io_dispatch_req_1_bits_ssid & 2'h2 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_18_2_value : _GEN_585; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_587 = 5'h12 == io_dispatch_req_1_bits_ssid & 2'h3 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_18_3_value : _GEN_586; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_588 = 5'h13 == io_dispatch_req_1_bits_ssid & 2'h0 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_19_0_value : _GEN_587; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_589 = 5'h13 == io_dispatch_req_1_bits_ssid & 2'h1 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_19_1_value : _GEN_588; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_590 = 5'h13 == io_dispatch_req_1_bits_ssid & 2'h2 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_19_2_value : _GEN_589; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_591 = 5'h13 == io_dispatch_req_1_bits_ssid & 2'h3 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_19_3_value : _GEN_590; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_592 = 5'h14 == io_dispatch_req_1_bits_ssid & 2'h0 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_20_0_value : _GEN_591; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_593 = 5'h14 == io_dispatch_req_1_bits_ssid & 2'h1 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_20_1_value : _GEN_592; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_594 = 5'h14 == io_dispatch_req_1_bits_ssid & 2'h2 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_20_2_value : _GEN_593; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_595 = 5'h14 == io_dispatch_req_1_bits_ssid & 2'h3 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_20_3_value : _GEN_594; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_596 = 5'h15 == io_dispatch_req_1_bits_ssid & 2'h0 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_21_0_value : _GEN_595; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_597 = 5'h15 == io_dispatch_req_1_bits_ssid & 2'h1 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_21_1_value : _GEN_596; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_598 = 5'h15 == io_dispatch_req_1_bits_ssid & 2'h2 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_21_2_value : _GEN_597; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_599 = 5'h15 == io_dispatch_req_1_bits_ssid & 2'h3 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_21_3_value : _GEN_598; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_600 = 5'h16 == io_dispatch_req_1_bits_ssid & 2'h0 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_22_0_value : _GEN_599; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_601 = 5'h16 == io_dispatch_req_1_bits_ssid & 2'h1 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_22_1_value : _GEN_600; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_602 = 5'h16 == io_dispatch_req_1_bits_ssid & 2'h2 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_22_2_value : _GEN_601; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_603 = 5'h16 == io_dispatch_req_1_bits_ssid & 2'h3 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_22_3_value : _GEN_602; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_604 = 5'h17 == io_dispatch_req_1_bits_ssid & 2'h0 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_23_0_value : _GEN_603; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_605 = 5'h17 == io_dispatch_req_1_bits_ssid & 2'h1 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_23_1_value : _GEN_604; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_606 = 5'h17 == io_dispatch_req_1_bits_ssid & 2'h2 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_23_2_value : _GEN_605; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_607 = 5'h17 == io_dispatch_req_1_bits_ssid & 2'h3 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_23_3_value : _GEN_606; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_608 = 5'h18 == io_dispatch_req_1_bits_ssid & 2'h0 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_24_0_value : _GEN_607; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_609 = 5'h18 == io_dispatch_req_1_bits_ssid & 2'h1 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_24_1_value : _GEN_608; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_610 = 5'h18 == io_dispatch_req_1_bits_ssid & 2'h2 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_24_2_value : _GEN_609; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_611 = 5'h18 == io_dispatch_req_1_bits_ssid & 2'h3 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_24_3_value : _GEN_610; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_612 = 5'h19 == io_dispatch_req_1_bits_ssid & 2'h0 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_25_0_value : _GEN_611; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_613 = 5'h19 == io_dispatch_req_1_bits_ssid & 2'h1 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_25_1_value : _GEN_612; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_614 = 5'h19 == io_dispatch_req_1_bits_ssid & 2'h2 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_25_2_value : _GEN_613; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_615 = 5'h19 == io_dispatch_req_1_bits_ssid & 2'h3 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_25_3_value : _GEN_614; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_616 = 5'h1a == io_dispatch_req_1_bits_ssid & 2'h0 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_26_0_value : _GEN_615; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_617 = 5'h1a == io_dispatch_req_1_bits_ssid & 2'h1 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_26_1_value : _GEN_616; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_618 = 5'h1a == io_dispatch_req_1_bits_ssid & 2'h2 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_26_2_value : _GEN_617; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_619 = 5'h1a == io_dispatch_req_1_bits_ssid & 2'h3 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_26_3_value : _GEN_618; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_620 = 5'h1b == io_dispatch_req_1_bits_ssid & 2'h0 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_27_0_value : _GEN_619; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_621 = 5'h1b == io_dispatch_req_1_bits_ssid & 2'h1 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_27_1_value : _GEN_620; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_622 = 5'h1b == io_dispatch_req_1_bits_ssid & 2'h2 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_27_2_value : _GEN_621; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_623 = 5'h1b == io_dispatch_req_1_bits_ssid & 2'h3 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_27_3_value : _GEN_622; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_624 = 5'h1c == io_dispatch_req_1_bits_ssid & 2'h0 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_28_0_value : _GEN_623; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_625 = 5'h1c == io_dispatch_req_1_bits_ssid & 2'h1 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_28_1_value : _GEN_624; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_626 = 5'h1c == io_dispatch_req_1_bits_ssid & 2'h2 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_28_2_value : _GEN_625; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_627 = 5'h1c == io_dispatch_req_1_bits_ssid & 2'h3 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_28_3_value : _GEN_626; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_628 = 5'h1d == io_dispatch_req_1_bits_ssid & 2'h0 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_29_0_value : _GEN_627; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_629 = 5'h1d == io_dispatch_req_1_bits_ssid & 2'h1 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_29_1_value : _GEN_628; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_630 = 5'h1d == io_dispatch_req_1_bits_ssid & 2'h2 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_29_2_value : _GEN_629; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_631 = 5'h1d == io_dispatch_req_1_bits_ssid & 2'h3 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_29_3_value : _GEN_630; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_632 = 5'h1e == io_dispatch_req_1_bits_ssid & 2'h0 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_30_0_value : _GEN_631; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_633 = 5'h1e == io_dispatch_req_1_bits_ssid & 2'h1 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_30_1_value : _GEN_632; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_634 = 5'h1e == io_dispatch_req_1_bits_ssid & 2'h2 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_30_2_value : _GEN_633; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_635 = 5'h1e == io_dispatch_req_1_bits_ssid & 2'h3 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_30_3_value : _GEN_634; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_636 = 5'h1f == io_dispatch_req_1_bits_ssid & 2'h0 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_31_0_value : _GEN_635; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_637 = 5'h1f == io_dispatch_req_1_bits_ssid & 2'h1 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_31_1_value : _GEN_636; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_638 = 5'h1f == io_dispatch_req_1_bits_ssid & 2'h2 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_31_2_value : _GEN_637; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_639 = 5'h1f == io_dispatch_req_1_bits_ssid & 2'h3 == _io_dispatch_resp_1_bits_robIdx_T_1 ?
    robIdxVec_31_3_value : _GEN_638; // @[StoreSet.scala 520:{37,37}]
  wire [4:0] _GEN_643 = 5'h1 == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_1_0_value : robIdxVec_0_0_value; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_644 = 5'h2 == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_2_0_value : _GEN_643; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_645 = 5'h3 == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_3_0_value : _GEN_644; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_646 = 5'h4 == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_4_0_value : _GEN_645; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_647 = 5'h5 == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_5_0_value : _GEN_646; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_648 = 5'h6 == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_6_0_value : _GEN_647; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_649 = 5'h7 == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_7_0_value : _GEN_648; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_650 = 5'h8 == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_8_0_value : _GEN_649; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_651 = 5'h9 == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_9_0_value : _GEN_650; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_652 = 5'ha == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_10_0_value : _GEN_651; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_653 = 5'hb == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_11_0_value : _GEN_652; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_654 = 5'hc == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_12_0_value : _GEN_653; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_655 = 5'hd == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_13_0_value : _GEN_654; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_656 = 5'he == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_14_0_value : _GEN_655; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_657 = 5'hf == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_15_0_value : _GEN_656; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_658 = 5'h10 == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_16_0_value : _GEN_657; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_659 = 5'h11 == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_17_0_value : _GEN_658; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_660 = 5'h12 == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_18_0_value : _GEN_659; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_661 = 5'h13 == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_19_0_value : _GEN_660; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_662 = 5'h14 == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_20_0_value : _GEN_661; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_663 = 5'h15 == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_21_0_value : _GEN_662; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_664 = 5'h16 == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_22_0_value : _GEN_663; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_665 = 5'h17 == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_23_0_value : _GEN_664; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_666 = 5'h18 == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_24_0_value : _GEN_665; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_667 = 5'h19 == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_25_0_value : _GEN_666; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_668 = 5'h1a == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_26_0_value : _GEN_667; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_669 = 5'h1b == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_27_0_value : _GEN_668; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_670 = 5'h1c == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_28_0_value : _GEN_669; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_671 = 5'h1d == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_29_0_value : _GEN_670; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_672 = 5'h1e == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_30_0_value : _GEN_671; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_673 = 5'h1f == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_31_0_value : _GEN_672; // @[StoreSet.scala 534:{121,121}]
  wire  _GEN_674 = 5'h0 == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_0_0; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_675 = 5'h1 == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_1_0; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_676 = 5'h2 == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_2_0; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_677 = 5'h3 == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_3_0; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_678 = 5'h4 == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_4_0; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_679 = 5'h5 == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_5_0; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_680 = 5'h6 == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_6_0; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_681 = 5'h7 == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_7_0; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_682 = 5'h8 == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_8_0; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_683 = 5'h9 == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_9_0; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_684 = 5'ha == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_10_0; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_685 = 5'hb == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_11_0; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_686 = 5'hc == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_12_0; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_687 = 5'hd == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_13_0; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_688 = 5'he == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_14_0; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_689 = 5'hf == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_15_0; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_690 = 5'h10 == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_16_0; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_691 = 5'h11 == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_17_0; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_692 = 5'h12 == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_18_0; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_693 = 5'h13 == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_19_0; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_694 = 5'h14 == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_20_0; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_695 = 5'h15 == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_21_0; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_696 = 5'h16 == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_22_0; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_697 = 5'h17 == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_23_0; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_698 = 5'h18 == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_24_0; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_699 = 5'h19 == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_25_0; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_700 = 5'h1a == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_26_0; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_701 = 5'h1b == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_27_0; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_702 = 5'h1c == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_28_0; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_703 = 5'h1d == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_29_0; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_704 = 5'h1e == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_30_0; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_705 = 5'h1f == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_31_0; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_706 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_673 ? _GEN_674 : validVec_0_0; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_707 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_673 ? _GEN_675 : validVec_1_0; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_708 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_673 ? _GEN_676 : validVec_2_0; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_709 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_673 ? _GEN_677 : validVec_3_0; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_710 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_673 ? _GEN_678 : validVec_4_0; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_711 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_673 ? _GEN_679 : validVec_5_0; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_712 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_673 ? _GEN_680 : validVec_6_0; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_713 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_673 ? _GEN_681 : validVec_7_0; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_714 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_673 ? _GEN_682 : validVec_8_0; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_715 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_673 ? _GEN_683 : validVec_9_0; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_716 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_673 ? _GEN_684 : validVec_10_0; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_717 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_673 ? _GEN_685 : validVec_11_0; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_718 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_673 ? _GEN_686 : validVec_12_0; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_719 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_673 ? _GEN_687 : validVec_13_0; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_720 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_673 ? _GEN_688 : validVec_14_0; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_721 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_673 ? _GEN_689 : validVec_15_0; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_722 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_673 ? _GEN_690 : validVec_16_0; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_723 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_673 ? _GEN_691 : validVec_17_0; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_724 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_673 ? _GEN_692 : validVec_18_0; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_725 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_673 ? _GEN_693 : validVec_19_0; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_726 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_673 ? _GEN_694 : validVec_20_0; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_727 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_673 ? _GEN_695 : validVec_21_0; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_728 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_673 ? _GEN_696 : validVec_22_0; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_729 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_673 ? _GEN_697 : validVec_23_0; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_730 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_673 ? _GEN_698 : validVec_24_0; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_731 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_673 ? _GEN_699 : validVec_25_0; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_732 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_673 ? _GEN_700 : validVec_26_0; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_733 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_673 ? _GEN_701 : validVec_27_0; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_734 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_673 ? _GEN_702 : validVec_28_0; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_735 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_673 ? _GEN_703 : validVec_29_0; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_736 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_673 ? _GEN_704 : validVec_30_0; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_737 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_673 ? _GEN_705 : validVec_31_0; // @[StoreSet.scala 534:179 491:25]
  wire [4:0] _GEN_739 = 5'h1 == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_1_1_value : robIdxVec_0_1_value; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_740 = 5'h2 == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_2_1_value : _GEN_739; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_741 = 5'h3 == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_3_1_value : _GEN_740; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_742 = 5'h4 == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_4_1_value : _GEN_741; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_743 = 5'h5 == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_5_1_value : _GEN_742; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_744 = 5'h6 == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_6_1_value : _GEN_743; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_745 = 5'h7 == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_7_1_value : _GEN_744; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_746 = 5'h8 == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_8_1_value : _GEN_745; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_747 = 5'h9 == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_9_1_value : _GEN_746; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_748 = 5'ha == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_10_1_value : _GEN_747; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_749 = 5'hb == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_11_1_value : _GEN_748; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_750 = 5'hc == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_12_1_value : _GEN_749; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_751 = 5'hd == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_13_1_value : _GEN_750; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_752 = 5'he == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_14_1_value : _GEN_751; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_753 = 5'hf == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_15_1_value : _GEN_752; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_754 = 5'h10 == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_16_1_value : _GEN_753; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_755 = 5'h11 == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_17_1_value : _GEN_754; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_756 = 5'h12 == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_18_1_value : _GEN_755; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_757 = 5'h13 == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_19_1_value : _GEN_756; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_758 = 5'h14 == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_20_1_value : _GEN_757; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_759 = 5'h15 == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_21_1_value : _GEN_758; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_760 = 5'h16 == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_22_1_value : _GEN_759; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_761 = 5'h17 == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_23_1_value : _GEN_760; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_762 = 5'h18 == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_24_1_value : _GEN_761; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_763 = 5'h19 == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_25_1_value : _GEN_762; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_764 = 5'h1a == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_26_1_value : _GEN_763; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_765 = 5'h1b == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_27_1_value : _GEN_764; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_766 = 5'h1c == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_28_1_value : _GEN_765; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_767 = 5'h1d == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_29_1_value : _GEN_766; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_768 = 5'h1e == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_30_1_value : _GEN_767; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_769 = 5'h1f == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_31_1_value : _GEN_768; // @[StoreSet.scala 534:{121,121}]
  wire  _GEN_770 = 5'h0 == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_0_1; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_771 = 5'h1 == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_1_1; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_772 = 5'h2 == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_2_1; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_773 = 5'h3 == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_3_1; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_774 = 5'h4 == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_4_1; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_775 = 5'h5 == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_5_1; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_776 = 5'h6 == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_6_1; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_777 = 5'h7 == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_7_1; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_778 = 5'h8 == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_8_1; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_779 = 5'h9 == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_9_1; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_780 = 5'ha == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_10_1; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_781 = 5'hb == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_11_1; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_782 = 5'hc == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_12_1; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_783 = 5'hd == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_13_1; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_784 = 5'he == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_14_1; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_785 = 5'hf == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_15_1; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_786 = 5'h10 == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_16_1; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_787 = 5'h11 == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_17_1; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_788 = 5'h12 == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_18_1; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_789 = 5'h13 == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_19_1; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_790 = 5'h14 == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_20_1; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_791 = 5'h15 == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_21_1; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_792 = 5'h16 == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_22_1; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_793 = 5'h17 == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_23_1; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_794 = 5'h18 == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_24_1; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_795 = 5'h19 == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_25_1; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_796 = 5'h1a == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_26_1; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_797 = 5'h1b == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_27_1; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_798 = 5'h1c == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_28_1; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_799 = 5'h1d == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_29_1; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_800 = 5'h1e == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_30_1; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_801 = 5'h1f == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_31_1; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_802 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_769 ? _GEN_770 : validVec_0_1; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_803 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_769 ? _GEN_771 : validVec_1_1; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_804 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_769 ? _GEN_772 : validVec_2_1; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_805 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_769 ? _GEN_773 : validVec_3_1; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_806 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_769 ? _GEN_774 : validVec_4_1; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_807 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_769 ? _GEN_775 : validVec_5_1; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_808 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_769 ? _GEN_776 : validVec_6_1; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_809 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_769 ? _GEN_777 : validVec_7_1; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_810 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_769 ? _GEN_778 : validVec_8_1; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_811 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_769 ? _GEN_779 : validVec_9_1; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_812 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_769 ? _GEN_780 : validVec_10_1; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_813 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_769 ? _GEN_781 : validVec_11_1; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_814 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_769 ? _GEN_782 : validVec_12_1; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_815 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_769 ? _GEN_783 : validVec_13_1; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_816 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_769 ? _GEN_784 : validVec_14_1; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_817 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_769 ? _GEN_785 : validVec_15_1; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_818 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_769 ? _GEN_786 : validVec_16_1; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_819 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_769 ? _GEN_787 : validVec_17_1; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_820 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_769 ? _GEN_788 : validVec_18_1; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_821 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_769 ? _GEN_789 : validVec_19_1; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_822 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_769 ? _GEN_790 : validVec_20_1; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_823 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_769 ? _GEN_791 : validVec_21_1; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_824 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_769 ? _GEN_792 : validVec_22_1; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_825 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_769 ? _GEN_793 : validVec_23_1; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_826 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_769 ? _GEN_794 : validVec_24_1; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_827 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_769 ? _GEN_795 : validVec_25_1; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_828 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_769 ? _GEN_796 : validVec_26_1; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_829 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_769 ? _GEN_797 : validVec_27_1; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_830 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_769 ? _GEN_798 : validVec_28_1; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_831 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_769 ? _GEN_799 : validVec_29_1; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_832 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_769 ? _GEN_800 : validVec_30_1; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_833 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_769 ? _GEN_801 : validVec_31_1; // @[StoreSet.scala 534:179 491:25]
  wire [4:0] _GEN_835 = 5'h1 == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_1_2_value : robIdxVec_0_2_value; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_836 = 5'h2 == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_2_2_value : _GEN_835; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_837 = 5'h3 == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_3_2_value : _GEN_836; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_838 = 5'h4 == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_4_2_value : _GEN_837; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_839 = 5'h5 == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_5_2_value : _GEN_838; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_840 = 5'h6 == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_6_2_value : _GEN_839; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_841 = 5'h7 == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_7_2_value : _GEN_840; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_842 = 5'h8 == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_8_2_value : _GEN_841; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_843 = 5'h9 == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_9_2_value : _GEN_842; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_844 = 5'ha == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_10_2_value : _GEN_843; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_845 = 5'hb == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_11_2_value : _GEN_844; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_846 = 5'hc == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_12_2_value : _GEN_845; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_847 = 5'hd == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_13_2_value : _GEN_846; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_848 = 5'he == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_14_2_value : _GEN_847; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_849 = 5'hf == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_15_2_value : _GEN_848; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_850 = 5'h10 == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_16_2_value : _GEN_849; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_851 = 5'h11 == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_17_2_value : _GEN_850; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_852 = 5'h12 == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_18_2_value : _GEN_851; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_853 = 5'h13 == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_19_2_value : _GEN_852; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_854 = 5'h14 == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_20_2_value : _GEN_853; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_855 = 5'h15 == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_21_2_value : _GEN_854; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_856 = 5'h16 == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_22_2_value : _GEN_855; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_857 = 5'h17 == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_23_2_value : _GEN_856; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_858 = 5'h18 == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_24_2_value : _GEN_857; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_859 = 5'h19 == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_25_2_value : _GEN_858; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_860 = 5'h1a == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_26_2_value : _GEN_859; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_861 = 5'h1b == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_27_2_value : _GEN_860; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_862 = 5'h1c == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_28_2_value : _GEN_861; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_863 = 5'h1d == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_29_2_value : _GEN_862; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_864 = 5'h1e == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_30_2_value : _GEN_863; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_865 = 5'h1f == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_31_2_value : _GEN_864; // @[StoreSet.scala 534:{121,121}]
  wire  _GEN_866 = 5'h0 == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_0_2; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_867 = 5'h1 == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_1_2; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_868 = 5'h2 == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_2_2; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_869 = 5'h3 == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_3_2; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_870 = 5'h4 == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_4_2; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_871 = 5'h5 == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_5_2; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_872 = 5'h6 == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_6_2; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_873 = 5'h7 == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_7_2; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_874 = 5'h8 == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_8_2; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_875 = 5'h9 == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_9_2; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_876 = 5'ha == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_10_2; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_877 = 5'hb == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_11_2; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_878 = 5'hc == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_12_2; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_879 = 5'hd == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_13_2; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_880 = 5'he == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_14_2; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_881 = 5'hf == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_15_2; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_882 = 5'h10 == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_16_2; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_883 = 5'h11 == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_17_2; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_884 = 5'h12 == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_18_2; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_885 = 5'h13 == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_19_2; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_886 = 5'h14 == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_20_2; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_887 = 5'h15 == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_21_2; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_888 = 5'h16 == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_22_2; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_889 = 5'h17 == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_23_2; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_890 = 5'h18 == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_24_2; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_891 = 5'h19 == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_25_2; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_892 = 5'h1a == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_26_2; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_893 = 5'h1b == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_27_2; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_894 = 5'h1c == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_28_2; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_895 = 5'h1d == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_29_2; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_896 = 5'h1e == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_30_2; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_897 = 5'h1f == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_31_2; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_898 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_865 ? _GEN_866 : validVec_0_2; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_899 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_865 ? _GEN_867 : validVec_1_2; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_900 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_865 ? _GEN_868 : validVec_2_2; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_901 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_865 ? _GEN_869 : validVec_3_2; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_902 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_865 ? _GEN_870 : validVec_4_2; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_903 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_865 ? _GEN_871 : validVec_5_2; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_904 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_865 ? _GEN_872 : validVec_6_2; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_905 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_865 ? _GEN_873 : validVec_7_2; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_906 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_865 ? _GEN_874 : validVec_8_2; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_907 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_865 ? _GEN_875 : validVec_9_2; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_908 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_865 ? _GEN_876 : validVec_10_2; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_909 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_865 ? _GEN_877 : validVec_11_2; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_910 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_865 ? _GEN_878 : validVec_12_2; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_911 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_865 ? _GEN_879 : validVec_13_2; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_912 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_865 ? _GEN_880 : validVec_14_2; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_913 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_865 ? _GEN_881 : validVec_15_2; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_914 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_865 ? _GEN_882 : validVec_16_2; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_915 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_865 ? _GEN_883 : validVec_17_2; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_916 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_865 ? _GEN_884 : validVec_18_2; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_917 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_865 ? _GEN_885 : validVec_19_2; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_918 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_865 ? _GEN_886 : validVec_20_2; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_919 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_865 ? _GEN_887 : validVec_21_2; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_920 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_865 ? _GEN_888 : validVec_22_2; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_921 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_865 ? _GEN_889 : validVec_23_2; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_922 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_865 ? _GEN_890 : validVec_24_2; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_923 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_865 ? _GEN_891 : validVec_25_2; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_924 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_865 ? _GEN_892 : validVec_26_2; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_925 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_865 ? _GEN_893 : validVec_27_2; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_926 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_865 ? _GEN_894 : validVec_28_2; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_927 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_865 ? _GEN_895 : validVec_29_2; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_928 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_865 ? _GEN_896 : validVec_30_2; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_929 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_865 ? _GEN_897 : validVec_31_2; // @[StoreSet.scala 534:179 491:25]
  wire [4:0] _GEN_931 = 5'h1 == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_1_3_value : robIdxVec_0_3_value; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_932 = 5'h2 == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_2_3_value : _GEN_931; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_933 = 5'h3 == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_3_3_value : _GEN_932; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_934 = 5'h4 == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_4_3_value : _GEN_933; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_935 = 5'h5 == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_5_3_value : _GEN_934; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_936 = 5'h6 == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_6_3_value : _GEN_935; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_937 = 5'h7 == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_7_3_value : _GEN_936; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_938 = 5'h8 == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_8_3_value : _GEN_937; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_939 = 5'h9 == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_9_3_value : _GEN_938; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_940 = 5'ha == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_10_3_value : _GEN_939; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_941 = 5'hb == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_11_3_value : _GEN_940; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_942 = 5'hc == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_12_3_value : _GEN_941; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_943 = 5'hd == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_13_3_value : _GEN_942; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_944 = 5'he == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_14_3_value : _GEN_943; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_945 = 5'hf == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_15_3_value : _GEN_944; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_946 = 5'h10 == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_16_3_value : _GEN_945; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_947 = 5'h11 == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_17_3_value : _GEN_946; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_948 = 5'h12 == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_18_3_value : _GEN_947; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_949 = 5'h13 == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_19_3_value : _GEN_948; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_950 = 5'h14 == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_20_3_value : _GEN_949; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_951 = 5'h15 == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_21_3_value : _GEN_950; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_952 = 5'h16 == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_22_3_value : _GEN_951; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_953 = 5'h17 == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_23_3_value : _GEN_952; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_954 = 5'h18 == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_24_3_value : _GEN_953; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_955 = 5'h19 == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_25_3_value : _GEN_954; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_956 = 5'h1a == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_26_3_value : _GEN_955; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_957 = 5'h1b == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_27_3_value : _GEN_956; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_958 = 5'h1c == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_28_3_value : _GEN_957; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_959 = 5'h1d == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_29_3_value : _GEN_958; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_960 = 5'h1e == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_30_3_value : _GEN_959; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_961 = 5'h1f == io_storeIssue_0_bits_uop_cf_ssid ? robIdxVec_31_3_value : _GEN_960; // @[StoreSet.scala 534:{121,121}]
  wire  _GEN_962 = 5'h0 == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_0_3; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_963 = 5'h1 == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_1_3; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_964 = 5'h2 == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_2_3; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_965 = 5'h3 == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_3_3; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_966 = 5'h4 == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_4_3; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_967 = 5'h5 == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_5_3; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_968 = 5'h6 == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_6_3; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_969 = 5'h7 == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_7_3; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_970 = 5'h8 == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_8_3; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_971 = 5'h9 == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_9_3; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_972 = 5'ha == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_10_3; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_973 = 5'hb == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_11_3; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_974 = 5'hc == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_12_3; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_975 = 5'hd == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_13_3; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_976 = 5'he == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_14_3; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_977 = 5'hf == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_15_3; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_978 = 5'h10 == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_16_3; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_979 = 5'h11 == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_17_3; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_980 = 5'h12 == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_18_3; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_981 = 5'h13 == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_19_3; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_982 = 5'h14 == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_20_3; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_983 = 5'h15 == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_21_3; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_984 = 5'h16 == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_22_3; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_985 = 5'h17 == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_23_3; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_986 = 5'h18 == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_24_3; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_987 = 5'h19 == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_25_3; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_988 = 5'h1a == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_26_3; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_989 = 5'h1b == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_27_3; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_990 = 5'h1c == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_28_3; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_991 = 5'h1d == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_29_3; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_992 = 5'h1e == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_30_3; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_993 = 5'h1f == io_storeIssue_0_bits_uop_cf_ssid ? 1'h0 : validVec_31_3; // @[StoreSet.scala 491:25 535:{56,56}]
  wire  _GEN_994 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_961 ? _GEN_962 : validVec_0_3; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_995 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_961 ? _GEN_963 : validVec_1_3; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_996 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_961 ? _GEN_964 : validVec_2_3; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_997 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_961 ? _GEN_965 : validVec_3_3; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_998 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_961 ? _GEN_966 : validVec_4_3; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_999 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_961 ? _GEN_967 : validVec_5_3; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_1000 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_961 ? _GEN_968 : validVec_6_3; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_1001 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_961 ? _GEN_969 : validVec_7_3; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_1002 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_961 ? _GEN_970 : validVec_8_3; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_1003 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_961 ? _GEN_971 : validVec_9_3; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_1004 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_961 ? _GEN_972 : validVec_10_3; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_1005 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_961 ? _GEN_973 : validVec_11_3; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_1006 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_961 ? _GEN_974 : validVec_12_3; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_1007 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_961 ? _GEN_975 : validVec_13_3; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_1008 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_961 ? _GEN_976 : validVec_14_3; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_1009 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_961 ? _GEN_977 : validVec_15_3; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_1010 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_961 ? _GEN_978 : validVec_16_3; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_1011 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_961 ? _GEN_979 : validVec_17_3; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_1012 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_961 ? _GEN_980 : validVec_18_3; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_1013 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_961 ? _GEN_981 : validVec_19_3; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_1014 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_961 ? _GEN_982 : validVec_20_3; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_1015 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_961 ? _GEN_983 : validVec_21_3; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_1016 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_961 ? _GEN_984 : validVec_22_3; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_1017 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_961 ? _GEN_985 : validVec_23_3; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_1018 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_961 ? _GEN_986 : validVec_24_3; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_1019 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_961 ? _GEN_987 : validVec_25_3; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_1020 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_961 ? _GEN_988 : validVec_26_3; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_1021 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_961 ? _GEN_989 : validVec_27_3; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_1022 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_961 ? _GEN_990 : validVec_28_3; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_1023 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_961 ? _GEN_991 : validVec_29_3; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_1024 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_961 ? _GEN_992 : validVec_30_3; // @[StoreSet.scala 534:179 491:25]
  wire  _GEN_1025 = io_storeIssue_0_valid & io_storeIssue_0_bits_uop_cf_storeSetHit &
    io_storeIssue_0_bits_uop_robIdx_value == _GEN_961 ? _GEN_993 : validVec_31_3; // @[StoreSet.scala 534:179 491:25]
  wire [4:0] _GEN_1027 = 5'h1 == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_1_0_value : robIdxVec_0_0_value; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1028 = 5'h2 == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_2_0_value : _GEN_1027; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1029 = 5'h3 == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_3_0_value : _GEN_1028; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1030 = 5'h4 == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_4_0_value : _GEN_1029; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1031 = 5'h5 == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_5_0_value : _GEN_1030; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1032 = 5'h6 == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_6_0_value : _GEN_1031; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1033 = 5'h7 == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_7_0_value : _GEN_1032; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1034 = 5'h8 == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_8_0_value : _GEN_1033; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1035 = 5'h9 == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_9_0_value : _GEN_1034; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1036 = 5'ha == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_10_0_value : _GEN_1035; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1037 = 5'hb == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_11_0_value : _GEN_1036; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1038 = 5'hc == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_12_0_value : _GEN_1037; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1039 = 5'hd == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_13_0_value : _GEN_1038; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1040 = 5'he == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_14_0_value : _GEN_1039; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1041 = 5'hf == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_15_0_value : _GEN_1040; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1042 = 5'h10 == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_16_0_value : _GEN_1041; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1043 = 5'h11 == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_17_0_value : _GEN_1042; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1044 = 5'h12 == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_18_0_value : _GEN_1043; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1045 = 5'h13 == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_19_0_value : _GEN_1044; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1046 = 5'h14 == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_20_0_value : _GEN_1045; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1047 = 5'h15 == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_21_0_value : _GEN_1046; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1048 = 5'h16 == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_22_0_value : _GEN_1047; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1049 = 5'h17 == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_23_0_value : _GEN_1048; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1050 = 5'h18 == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_24_0_value : _GEN_1049; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1051 = 5'h19 == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_25_0_value : _GEN_1050; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1052 = 5'h1a == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_26_0_value : _GEN_1051; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1053 = 5'h1b == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_27_0_value : _GEN_1052; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1054 = 5'h1c == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_28_0_value : _GEN_1053; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1055 = 5'h1d == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_29_0_value : _GEN_1054; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1056 = 5'h1e == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_30_0_value : _GEN_1055; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1057 = 5'h1f == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_31_0_value : _GEN_1056; // @[StoreSet.scala 534:{121,121}]
  wire  _GEN_1058 = 5'h0 == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_706; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1059 = 5'h1 == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_707; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1060 = 5'h2 == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_708; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1061 = 5'h3 == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_709; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1062 = 5'h4 == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_710; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1063 = 5'h5 == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_711; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1064 = 5'h6 == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_712; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1065 = 5'h7 == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_713; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1066 = 5'h8 == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_714; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1067 = 5'h9 == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_715; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1068 = 5'ha == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_716; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1069 = 5'hb == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_717; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1070 = 5'hc == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_718; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1071 = 5'hd == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_719; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1072 = 5'he == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_720; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1073 = 5'hf == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_721; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1074 = 5'h10 == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_722; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1075 = 5'h11 == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_723; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1076 = 5'h12 == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_724; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1077 = 5'h13 == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_725; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1078 = 5'h14 == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_726; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1079 = 5'h15 == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_727; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1080 = 5'h16 == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_728; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1081 = 5'h17 == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_729; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1082 = 5'h18 == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_730; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1083 = 5'h19 == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_731; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1084 = 5'h1a == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_732; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1085 = 5'h1b == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_733; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1086 = 5'h1c == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_734; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1087 = 5'h1d == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_735; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1088 = 5'h1e == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_736; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1089 = 5'h1f == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_737; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1090 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1057 ? _GEN_1058 : _GEN_706; // @[StoreSet.scala 534:179]
  wire  _GEN_1091 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1057 ? _GEN_1059 : _GEN_707; // @[StoreSet.scala 534:179]
  wire  _GEN_1092 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1057 ? _GEN_1060 : _GEN_708; // @[StoreSet.scala 534:179]
  wire  _GEN_1093 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1057 ? _GEN_1061 : _GEN_709; // @[StoreSet.scala 534:179]
  wire  _GEN_1094 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1057 ? _GEN_1062 : _GEN_710; // @[StoreSet.scala 534:179]
  wire  _GEN_1095 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1057 ? _GEN_1063 : _GEN_711; // @[StoreSet.scala 534:179]
  wire  _GEN_1096 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1057 ? _GEN_1064 : _GEN_712; // @[StoreSet.scala 534:179]
  wire  _GEN_1097 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1057 ? _GEN_1065 : _GEN_713; // @[StoreSet.scala 534:179]
  wire  _GEN_1098 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1057 ? _GEN_1066 : _GEN_714; // @[StoreSet.scala 534:179]
  wire  _GEN_1099 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1057 ? _GEN_1067 : _GEN_715; // @[StoreSet.scala 534:179]
  wire  _GEN_1100 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1057 ? _GEN_1068 : _GEN_716; // @[StoreSet.scala 534:179]
  wire  _GEN_1101 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1057 ? _GEN_1069 : _GEN_717; // @[StoreSet.scala 534:179]
  wire  _GEN_1102 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1057 ? _GEN_1070 : _GEN_718; // @[StoreSet.scala 534:179]
  wire  _GEN_1103 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1057 ? _GEN_1071 : _GEN_719; // @[StoreSet.scala 534:179]
  wire  _GEN_1104 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1057 ? _GEN_1072 : _GEN_720; // @[StoreSet.scala 534:179]
  wire  _GEN_1105 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1057 ? _GEN_1073 : _GEN_721; // @[StoreSet.scala 534:179]
  wire  _GEN_1106 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1057 ? _GEN_1074 : _GEN_722; // @[StoreSet.scala 534:179]
  wire  _GEN_1107 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1057 ? _GEN_1075 : _GEN_723; // @[StoreSet.scala 534:179]
  wire  _GEN_1108 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1057 ? _GEN_1076 : _GEN_724; // @[StoreSet.scala 534:179]
  wire  _GEN_1109 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1057 ? _GEN_1077 : _GEN_725; // @[StoreSet.scala 534:179]
  wire  _GEN_1110 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1057 ? _GEN_1078 : _GEN_726; // @[StoreSet.scala 534:179]
  wire  _GEN_1111 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1057 ? _GEN_1079 : _GEN_727; // @[StoreSet.scala 534:179]
  wire  _GEN_1112 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1057 ? _GEN_1080 : _GEN_728; // @[StoreSet.scala 534:179]
  wire  _GEN_1113 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1057 ? _GEN_1081 : _GEN_729; // @[StoreSet.scala 534:179]
  wire  _GEN_1114 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1057 ? _GEN_1082 : _GEN_730; // @[StoreSet.scala 534:179]
  wire  _GEN_1115 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1057 ? _GEN_1083 : _GEN_731; // @[StoreSet.scala 534:179]
  wire  _GEN_1116 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1057 ? _GEN_1084 : _GEN_732; // @[StoreSet.scala 534:179]
  wire  _GEN_1117 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1057 ? _GEN_1085 : _GEN_733; // @[StoreSet.scala 534:179]
  wire  _GEN_1118 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1057 ? _GEN_1086 : _GEN_734; // @[StoreSet.scala 534:179]
  wire  _GEN_1119 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1057 ? _GEN_1087 : _GEN_735; // @[StoreSet.scala 534:179]
  wire  _GEN_1120 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1057 ? _GEN_1088 : _GEN_736; // @[StoreSet.scala 534:179]
  wire  _GEN_1121 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1057 ? _GEN_1089 : _GEN_737; // @[StoreSet.scala 534:179]
  wire [4:0] _GEN_1123 = 5'h1 == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_1_1_value : robIdxVec_0_1_value; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1124 = 5'h2 == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_2_1_value : _GEN_1123; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1125 = 5'h3 == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_3_1_value : _GEN_1124; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1126 = 5'h4 == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_4_1_value : _GEN_1125; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1127 = 5'h5 == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_5_1_value : _GEN_1126; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1128 = 5'h6 == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_6_1_value : _GEN_1127; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1129 = 5'h7 == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_7_1_value : _GEN_1128; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1130 = 5'h8 == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_8_1_value : _GEN_1129; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1131 = 5'h9 == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_9_1_value : _GEN_1130; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1132 = 5'ha == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_10_1_value : _GEN_1131; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1133 = 5'hb == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_11_1_value : _GEN_1132; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1134 = 5'hc == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_12_1_value : _GEN_1133; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1135 = 5'hd == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_13_1_value : _GEN_1134; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1136 = 5'he == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_14_1_value : _GEN_1135; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1137 = 5'hf == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_15_1_value : _GEN_1136; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1138 = 5'h10 == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_16_1_value : _GEN_1137; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1139 = 5'h11 == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_17_1_value : _GEN_1138; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1140 = 5'h12 == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_18_1_value : _GEN_1139; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1141 = 5'h13 == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_19_1_value : _GEN_1140; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1142 = 5'h14 == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_20_1_value : _GEN_1141; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1143 = 5'h15 == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_21_1_value : _GEN_1142; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1144 = 5'h16 == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_22_1_value : _GEN_1143; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1145 = 5'h17 == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_23_1_value : _GEN_1144; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1146 = 5'h18 == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_24_1_value : _GEN_1145; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1147 = 5'h19 == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_25_1_value : _GEN_1146; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1148 = 5'h1a == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_26_1_value : _GEN_1147; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1149 = 5'h1b == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_27_1_value : _GEN_1148; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1150 = 5'h1c == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_28_1_value : _GEN_1149; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1151 = 5'h1d == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_29_1_value : _GEN_1150; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1152 = 5'h1e == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_30_1_value : _GEN_1151; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1153 = 5'h1f == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_31_1_value : _GEN_1152; // @[StoreSet.scala 534:{121,121}]
  wire  _GEN_1154 = 5'h0 == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_802; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1155 = 5'h1 == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_803; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1156 = 5'h2 == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_804; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1157 = 5'h3 == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_805; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1158 = 5'h4 == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_806; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1159 = 5'h5 == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_807; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1160 = 5'h6 == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_808; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1161 = 5'h7 == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_809; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1162 = 5'h8 == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_810; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1163 = 5'h9 == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_811; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1164 = 5'ha == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_812; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1165 = 5'hb == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_813; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1166 = 5'hc == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_814; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1167 = 5'hd == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_815; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1168 = 5'he == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_816; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1169 = 5'hf == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_817; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1170 = 5'h10 == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_818; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1171 = 5'h11 == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_819; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1172 = 5'h12 == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_820; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1173 = 5'h13 == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_821; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1174 = 5'h14 == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_822; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1175 = 5'h15 == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_823; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1176 = 5'h16 == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_824; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1177 = 5'h17 == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_825; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1178 = 5'h18 == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_826; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1179 = 5'h19 == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_827; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1180 = 5'h1a == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_828; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1181 = 5'h1b == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_829; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1182 = 5'h1c == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_830; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1183 = 5'h1d == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_831; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1184 = 5'h1e == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_832; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1185 = 5'h1f == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_833; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1186 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1153 ? _GEN_1154 : _GEN_802; // @[StoreSet.scala 534:179]
  wire  _GEN_1187 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1153 ? _GEN_1155 : _GEN_803; // @[StoreSet.scala 534:179]
  wire  _GEN_1188 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1153 ? _GEN_1156 : _GEN_804; // @[StoreSet.scala 534:179]
  wire  _GEN_1189 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1153 ? _GEN_1157 : _GEN_805; // @[StoreSet.scala 534:179]
  wire  _GEN_1190 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1153 ? _GEN_1158 : _GEN_806; // @[StoreSet.scala 534:179]
  wire  _GEN_1191 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1153 ? _GEN_1159 : _GEN_807; // @[StoreSet.scala 534:179]
  wire  _GEN_1192 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1153 ? _GEN_1160 : _GEN_808; // @[StoreSet.scala 534:179]
  wire  _GEN_1193 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1153 ? _GEN_1161 : _GEN_809; // @[StoreSet.scala 534:179]
  wire  _GEN_1194 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1153 ? _GEN_1162 : _GEN_810; // @[StoreSet.scala 534:179]
  wire  _GEN_1195 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1153 ? _GEN_1163 : _GEN_811; // @[StoreSet.scala 534:179]
  wire  _GEN_1196 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1153 ? _GEN_1164 : _GEN_812; // @[StoreSet.scala 534:179]
  wire  _GEN_1197 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1153 ? _GEN_1165 : _GEN_813; // @[StoreSet.scala 534:179]
  wire  _GEN_1198 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1153 ? _GEN_1166 : _GEN_814; // @[StoreSet.scala 534:179]
  wire  _GEN_1199 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1153 ? _GEN_1167 : _GEN_815; // @[StoreSet.scala 534:179]
  wire  _GEN_1200 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1153 ? _GEN_1168 : _GEN_816; // @[StoreSet.scala 534:179]
  wire  _GEN_1201 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1153 ? _GEN_1169 : _GEN_817; // @[StoreSet.scala 534:179]
  wire  _GEN_1202 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1153 ? _GEN_1170 : _GEN_818; // @[StoreSet.scala 534:179]
  wire  _GEN_1203 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1153 ? _GEN_1171 : _GEN_819; // @[StoreSet.scala 534:179]
  wire  _GEN_1204 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1153 ? _GEN_1172 : _GEN_820; // @[StoreSet.scala 534:179]
  wire  _GEN_1205 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1153 ? _GEN_1173 : _GEN_821; // @[StoreSet.scala 534:179]
  wire  _GEN_1206 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1153 ? _GEN_1174 : _GEN_822; // @[StoreSet.scala 534:179]
  wire  _GEN_1207 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1153 ? _GEN_1175 : _GEN_823; // @[StoreSet.scala 534:179]
  wire  _GEN_1208 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1153 ? _GEN_1176 : _GEN_824; // @[StoreSet.scala 534:179]
  wire  _GEN_1209 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1153 ? _GEN_1177 : _GEN_825; // @[StoreSet.scala 534:179]
  wire  _GEN_1210 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1153 ? _GEN_1178 : _GEN_826; // @[StoreSet.scala 534:179]
  wire  _GEN_1211 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1153 ? _GEN_1179 : _GEN_827; // @[StoreSet.scala 534:179]
  wire  _GEN_1212 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1153 ? _GEN_1180 : _GEN_828; // @[StoreSet.scala 534:179]
  wire  _GEN_1213 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1153 ? _GEN_1181 : _GEN_829; // @[StoreSet.scala 534:179]
  wire  _GEN_1214 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1153 ? _GEN_1182 : _GEN_830; // @[StoreSet.scala 534:179]
  wire  _GEN_1215 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1153 ? _GEN_1183 : _GEN_831; // @[StoreSet.scala 534:179]
  wire  _GEN_1216 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1153 ? _GEN_1184 : _GEN_832; // @[StoreSet.scala 534:179]
  wire  _GEN_1217 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1153 ? _GEN_1185 : _GEN_833; // @[StoreSet.scala 534:179]
  wire [4:0] _GEN_1219 = 5'h1 == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_1_2_value : robIdxVec_0_2_value; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1220 = 5'h2 == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_2_2_value : _GEN_1219; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1221 = 5'h3 == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_3_2_value : _GEN_1220; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1222 = 5'h4 == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_4_2_value : _GEN_1221; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1223 = 5'h5 == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_5_2_value : _GEN_1222; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1224 = 5'h6 == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_6_2_value : _GEN_1223; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1225 = 5'h7 == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_7_2_value : _GEN_1224; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1226 = 5'h8 == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_8_2_value : _GEN_1225; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1227 = 5'h9 == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_9_2_value : _GEN_1226; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1228 = 5'ha == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_10_2_value : _GEN_1227; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1229 = 5'hb == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_11_2_value : _GEN_1228; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1230 = 5'hc == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_12_2_value : _GEN_1229; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1231 = 5'hd == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_13_2_value : _GEN_1230; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1232 = 5'he == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_14_2_value : _GEN_1231; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1233 = 5'hf == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_15_2_value : _GEN_1232; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1234 = 5'h10 == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_16_2_value : _GEN_1233; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1235 = 5'h11 == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_17_2_value : _GEN_1234; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1236 = 5'h12 == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_18_2_value : _GEN_1235; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1237 = 5'h13 == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_19_2_value : _GEN_1236; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1238 = 5'h14 == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_20_2_value : _GEN_1237; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1239 = 5'h15 == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_21_2_value : _GEN_1238; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1240 = 5'h16 == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_22_2_value : _GEN_1239; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1241 = 5'h17 == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_23_2_value : _GEN_1240; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1242 = 5'h18 == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_24_2_value : _GEN_1241; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1243 = 5'h19 == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_25_2_value : _GEN_1242; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1244 = 5'h1a == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_26_2_value : _GEN_1243; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1245 = 5'h1b == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_27_2_value : _GEN_1244; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1246 = 5'h1c == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_28_2_value : _GEN_1245; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1247 = 5'h1d == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_29_2_value : _GEN_1246; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1248 = 5'h1e == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_30_2_value : _GEN_1247; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1249 = 5'h1f == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_31_2_value : _GEN_1248; // @[StoreSet.scala 534:{121,121}]
  wire  _GEN_1250 = 5'h0 == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_898; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1251 = 5'h1 == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_899; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1252 = 5'h2 == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_900; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1253 = 5'h3 == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_901; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1254 = 5'h4 == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_902; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1255 = 5'h5 == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_903; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1256 = 5'h6 == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_904; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1257 = 5'h7 == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_905; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1258 = 5'h8 == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_906; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1259 = 5'h9 == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_907; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1260 = 5'ha == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_908; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1261 = 5'hb == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_909; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1262 = 5'hc == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_910; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1263 = 5'hd == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_911; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1264 = 5'he == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_912; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1265 = 5'hf == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_913; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1266 = 5'h10 == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_914; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1267 = 5'h11 == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_915; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1268 = 5'h12 == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_916; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1269 = 5'h13 == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_917; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1270 = 5'h14 == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_918; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1271 = 5'h15 == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_919; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1272 = 5'h16 == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_920; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1273 = 5'h17 == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_921; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1274 = 5'h18 == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_922; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1275 = 5'h19 == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_923; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1276 = 5'h1a == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_924; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1277 = 5'h1b == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_925; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1278 = 5'h1c == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_926; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1279 = 5'h1d == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_927; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1280 = 5'h1e == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_928; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1281 = 5'h1f == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_929; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1282 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1249 ? _GEN_1250 : _GEN_898; // @[StoreSet.scala 534:179]
  wire  _GEN_1283 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1249 ? _GEN_1251 : _GEN_899; // @[StoreSet.scala 534:179]
  wire  _GEN_1284 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1249 ? _GEN_1252 : _GEN_900; // @[StoreSet.scala 534:179]
  wire  _GEN_1285 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1249 ? _GEN_1253 : _GEN_901; // @[StoreSet.scala 534:179]
  wire  _GEN_1286 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1249 ? _GEN_1254 : _GEN_902; // @[StoreSet.scala 534:179]
  wire  _GEN_1287 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1249 ? _GEN_1255 : _GEN_903; // @[StoreSet.scala 534:179]
  wire  _GEN_1288 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1249 ? _GEN_1256 : _GEN_904; // @[StoreSet.scala 534:179]
  wire  _GEN_1289 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1249 ? _GEN_1257 : _GEN_905; // @[StoreSet.scala 534:179]
  wire  _GEN_1290 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1249 ? _GEN_1258 : _GEN_906; // @[StoreSet.scala 534:179]
  wire  _GEN_1291 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1249 ? _GEN_1259 : _GEN_907; // @[StoreSet.scala 534:179]
  wire  _GEN_1292 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1249 ? _GEN_1260 : _GEN_908; // @[StoreSet.scala 534:179]
  wire  _GEN_1293 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1249 ? _GEN_1261 : _GEN_909; // @[StoreSet.scala 534:179]
  wire  _GEN_1294 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1249 ? _GEN_1262 : _GEN_910; // @[StoreSet.scala 534:179]
  wire  _GEN_1295 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1249 ? _GEN_1263 : _GEN_911; // @[StoreSet.scala 534:179]
  wire  _GEN_1296 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1249 ? _GEN_1264 : _GEN_912; // @[StoreSet.scala 534:179]
  wire  _GEN_1297 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1249 ? _GEN_1265 : _GEN_913; // @[StoreSet.scala 534:179]
  wire  _GEN_1298 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1249 ? _GEN_1266 : _GEN_914; // @[StoreSet.scala 534:179]
  wire  _GEN_1299 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1249 ? _GEN_1267 : _GEN_915; // @[StoreSet.scala 534:179]
  wire  _GEN_1300 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1249 ? _GEN_1268 : _GEN_916; // @[StoreSet.scala 534:179]
  wire  _GEN_1301 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1249 ? _GEN_1269 : _GEN_917; // @[StoreSet.scala 534:179]
  wire  _GEN_1302 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1249 ? _GEN_1270 : _GEN_918; // @[StoreSet.scala 534:179]
  wire  _GEN_1303 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1249 ? _GEN_1271 : _GEN_919; // @[StoreSet.scala 534:179]
  wire  _GEN_1304 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1249 ? _GEN_1272 : _GEN_920; // @[StoreSet.scala 534:179]
  wire  _GEN_1305 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1249 ? _GEN_1273 : _GEN_921; // @[StoreSet.scala 534:179]
  wire  _GEN_1306 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1249 ? _GEN_1274 : _GEN_922; // @[StoreSet.scala 534:179]
  wire  _GEN_1307 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1249 ? _GEN_1275 : _GEN_923; // @[StoreSet.scala 534:179]
  wire  _GEN_1308 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1249 ? _GEN_1276 : _GEN_924; // @[StoreSet.scala 534:179]
  wire  _GEN_1309 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1249 ? _GEN_1277 : _GEN_925; // @[StoreSet.scala 534:179]
  wire  _GEN_1310 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1249 ? _GEN_1278 : _GEN_926; // @[StoreSet.scala 534:179]
  wire  _GEN_1311 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1249 ? _GEN_1279 : _GEN_927; // @[StoreSet.scala 534:179]
  wire  _GEN_1312 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1249 ? _GEN_1280 : _GEN_928; // @[StoreSet.scala 534:179]
  wire  _GEN_1313 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1249 ? _GEN_1281 : _GEN_929; // @[StoreSet.scala 534:179]
  wire [4:0] _GEN_1315 = 5'h1 == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_1_3_value : robIdxVec_0_3_value; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1316 = 5'h2 == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_2_3_value : _GEN_1315; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1317 = 5'h3 == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_3_3_value : _GEN_1316; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1318 = 5'h4 == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_4_3_value : _GEN_1317; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1319 = 5'h5 == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_5_3_value : _GEN_1318; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1320 = 5'h6 == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_6_3_value : _GEN_1319; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1321 = 5'h7 == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_7_3_value : _GEN_1320; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1322 = 5'h8 == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_8_3_value : _GEN_1321; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1323 = 5'h9 == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_9_3_value : _GEN_1322; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1324 = 5'ha == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_10_3_value : _GEN_1323; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1325 = 5'hb == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_11_3_value : _GEN_1324; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1326 = 5'hc == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_12_3_value : _GEN_1325; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1327 = 5'hd == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_13_3_value : _GEN_1326; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1328 = 5'he == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_14_3_value : _GEN_1327; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1329 = 5'hf == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_15_3_value : _GEN_1328; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1330 = 5'h10 == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_16_3_value : _GEN_1329; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1331 = 5'h11 == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_17_3_value : _GEN_1330; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1332 = 5'h12 == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_18_3_value : _GEN_1331; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1333 = 5'h13 == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_19_3_value : _GEN_1332; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1334 = 5'h14 == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_20_3_value : _GEN_1333; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1335 = 5'h15 == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_21_3_value : _GEN_1334; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1336 = 5'h16 == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_22_3_value : _GEN_1335; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1337 = 5'h17 == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_23_3_value : _GEN_1336; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1338 = 5'h18 == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_24_3_value : _GEN_1337; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1339 = 5'h19 == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_25_3_value : _GEN_1338; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1340 = 5'h1a == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_26_3_value : _GEN_1339; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1341 = 5'h1b == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_27_3_value : _GEN_1340; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1342 = 5'h1c == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_28_3_value : _GEN_1341; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1343 = 5'h1d == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_29_3_value : _GEN_1342; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1344 = 5'h1e == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_30_3_value : _GEN_1343; // @[StoreSet.scala 534:{121,121}]
  wire [4:0] _GEN_1345 = 5'h1f == io_storeIssue_1_bits_uop_cf_ssid ? robIdxVec_31_3_value : _GEN_1344; // @[StoreSet.scala 534:{121,121}]
  wire  _GEN_1346 = 5'h0 == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_994; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1347 = 5'h1 == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_995; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1348 = 5'h2 == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_996; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1349 = 5'h3 == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_997; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1350 = 5'h4 == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_998; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1351 = 5'h5 == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_999; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1352 = 5'h6 == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_1000; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1353 = 5'h7 == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_1001; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1354 = 5'h8 == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_1002; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1355 = 5'h9 == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_1003; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1356 = 5'ha == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_1004; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1357 = 5'hb == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_1005; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1358 = 5'hc == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_1006; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1359 = 5'hd == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_1007; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1360 = 5'he == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_1008; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1361 = 5'hf == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_1009; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1362 = 5'h10 == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_1010; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1363 = 5'h11 == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_1011; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1364 = 5'h12 == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_1012; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1365 = 5'h13 == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_1013; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1366 = 5'h14 == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_1014; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1367 = 5'h15 == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_1015; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1368 = 5'h16 == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_1016; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1369 = 5'h17 == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_1017; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1370 = 5'h18 == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_1018; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1371 = 5'h19 == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_1019; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1372 = 5'h1a == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_1020; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1373 = 5'h1b == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_1021; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1374 = 5'h1c == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_1022; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1375 = 5'h1d == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_1023; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1376 = 5'h1e == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_1024; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1377 = 5'h1f == io_storeIssue_1_bits_uop_cf_ssid ? 1'h0 : _GEN_1025; // @[StoreSet.scala 535:{56,56}]
  wire  _GEN_1378 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1345 ? _GEN_1346 : _GEN_994; // @[StoreSet.scala 534:179]
  wire  _GEN_1379 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1345 ? _GEN_1347 : _GEN_995; // @[StoreSet.scala 534:179]
  wire  _GEN_1380 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1345 ? _GEN_1348 : _GEN_996; // @[StoreSet.scala 534:179]
  wire  _GEN_1381 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1345 ? _GEN_1349 : _GEN_997; // @[StoreSet.scala 534:179]
  wire  _GEN_1382 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1345 ? _GEN_1350 : _GEN_998; // @[StoreSet.scala 534:179]
  wire  _GEN_1383 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1345 ? _GEN_1351 : _GEN_999; // @[StoreSet.scala 534:179]
  wire  _GEN_1384 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1345 ? _GEN_1352 : _GEN_1000; // @[StoreSet.scala 534:179]
  wire  _GEN_1385 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1345 ? _GEN_1353 : _GEN_1001; // @[StoreSet.scala 534:179]
  wire  _GEN_1386 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1345 ? _GEN_1354 : _GEN_1002; // @[StoreSet.scala 534:179]
  wire  _GEN_1387 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1345 ? _GEN_1355 : _GEN_1003; // @[StoreSet.scala 534:179]
  wire  _GEN_1388 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1345 ? _GEN_1356 : _GEN_1004; // @[StoreSet.scala 534:179]
  wire  _GEN_1389 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1345 ? _GEN_1357 : _GEN_1005; // @[StoreSet.scala 534:179]
  wire  _GEN_1390 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1345 ? _GEN_1358 : _GEN_1006; // @[StoreSet.scala 534:179]
  wire  _GEN_1391 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1345 ? _GEN_1359 : _GEN_1007; // @[StoreSet.scala 534:179]
  wire  _GEN_1392 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1345 ? _GEN_1360 : _GEN_1008; // @[StoreSet.scala 534:179]
  wire  _GEN_1393 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1345 ? _GEN_1361 : _GEN_1009; // @[StoreSet.scala 534:179]
  wire  _GEN_1394 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1345 ? _GEN_1362 : _GEN_1010; // @[StoreSet.scala 534:179]
  wire  _GEN_1395 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1345 ? _GEN_1363 : _GEN_1011; // @[StoreSet.scala 534:179]
  wire  _GEN_1396 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1345 ? _GEN_1364 : _GEN_1012; // @[StoreSet.scala 534:179]
  wire  _GEN_1397 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1345 ? _GEN_1365 : _GEN_1013; // @[StoreSet.scala 534:179]
  wire  _GEN_1398 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1345 ? _GEN_1366 : _GEN_1014; // @[StoreSet.scala 534:179]
  wire  _GEN_1399 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1345 ? _GEN_1367 : _GEN_1015; // @[StoreSet.scala 534:179]
  wire  _GEN_1400 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1345 ? _GEN_1368 : _GEN_1016; // @[StoreSet.scala 534:179]
  wire  _GEN_1401 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1345 ? _GEN_1369 : _GEN_1017; // @[StoreSet.scala 534:179]
  wire  _GEN_1402 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1345 ? _GEN_1370 : _GEN_1018; // @[StoreSet.scala 534:179]
  wire  _GEN_1403 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1345 ? _GEN_1371 : _GEN_1019; // @[StoreSet.scala 534:179]
  wire  _GEN_1404 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1345 ? _GEN_1372 : _GEN_1020; // @[StoreSet.scala 534:179]
  wire  _GEN_1405 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1345 ? _GEN_1373 : _GEN_1021; // @[StoreSet.scala 534:179]
  wire  _GEN_1406 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1345 ? _GEN_1374 : _GEN_1022; // @[StoreSet.scala 534:179]
  wire  _GEN_1407 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1345 ? _GEN_1375 : _GEN_1023; // @[StoreSet.scala 534:179]
  wire  _GEN_1408 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1345 ? _GEN_1376 : _GEN_1024; // @[StoreSet.scala 534:179]
  wire  _GEN_1409 = io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit &
    io_storeIssue_1_bits_uop_robIdx_value == _GEN_1345 ? _GEN_1377 : _GEN_1025; // @[StoreSet.scala 534:179]
  wire [1:0] _allocPtr_T_1 = _GEN_63 + 2'h1; // @[StoreSet.scala 545:42]
  wire [1:0] _GEN_1410 = 5'h0 == io_dispatch_req_0_bits_ssid ? _allocPtr_T_1 : allocPtr_0; // @[StoreSet.scala 545:{23,23} 493:25]
  wire [1:0] _GEN_1411 = 5'h1 == io_dispatch_req_0_bits_ssid ? _allocPtr_T_1 : allocPtr_1; // @[StoreSet.scala 545:{23,23} 493:25]
  wire [1:0] _GEN_1412 = 5'h2 == io_dispatch_req_0_bits_ssid ? _allocPtr_T_1 : allocPtr_2; // @[StoreSet.scala 545:{23,23} 493:25]
  wire [1:0] _GEN_1413 = 5'h3 == io_dispatch_req_0_bits_ssid ? _allocPtr_T_1 : allocPtr_3; // @[StoreSet.scala 545:{23,23} 493:25]
  wire [1:0] _GEN_1414 = 5'h4 == io_dispatch_req_0_bits_ssid ? _allocPtr_T_1 : allocPtr_4; // @[StoreSet.scala 545:{23,23} 493:25]
  wire [1:0] _GEN_1415 = 5'h5 == io_dispatch_req_0_bits_ssid ? _allocPtr_T_1 : allocPtr_5; // @[StoreSet.scala 545:{23,23} 493:25]
  wire [1:0] _GEN_1416 = 5'h6 == io_dispatch_req_0_bits_ssid ? _allocPtr_T_1 : allocPtr_6; // @[StoreSet.scala 545:{23,23} 493:25]
  wire [1:0] _GEN_1417 = 5'h7 == io_dispatch_req_0_bits_ssid ? _allocPtr_T_1 : allocPtr_7; // @[StoreSet.scala 545:{23,23} 493:25]
  wire [1:0] _GEN_1418 = 5'h8 == io_dispatch_req_0_bits_ssid ? _allocPtr_T_1 : allocPtr_8; // @[StoreSet.scala 545:{23,23} 493:25]
  wire [1:0] _GEN_1419 = 5'h9 == io_dispatch_req_0_bits_ssid ? _allocPtr_T_1 : allocPtr_9; // @[StoreSet.scala 545:{23,23} 493:25]
  wire [1:0] _GEN_1420 = 5'ha == io_dispatch_req_0_bits_ssid ? _allocPtr_T_1 : allocPtr_10; // @[StoreSet.scala 545:{23,23} 493:25]
  wire [1:0] _GEN_1421 = 5'hb == io_dispatch_req_0_bits_ssid ? _allocPtr_T_1 : allocPtr_11; // @[StoreSet.scala 545:{23,23} 493:25]
  wire [1:0] _GEN_1422 = 5'hc == io_dispatch_req_0_bits_ssid ? _allocPtr_T_1 : allocPtr_12; // @[StoreSet.scala 545:{23,23} 493:25]
  wire [1:0] _GEN_1423 = 5'hd == io_dispatch_req_0_bits_ssid ? _allocPtr_T_1 : allocPtr_13; // @[StoreSet.scala 545:{23,23} 493:25]
  wire [1:0] _GEN_1424 = 5'he == io_dispatch_req_0_bits_ssid ? _allocPtr_T_1 : allocPtr_14; // @[StoreSet.scala 545:{23,23} 493:25]
  wire [1:0] _GEN_1425 = 5'hf == io_dispatch_req_0_bits_ssid ? _allocPtr_T_1 : allocPtr_15; // @[StoreSet.scala 545:{23,23} 493:25]
  wire [1:0] _GEN_1426 = 5'h10 == io_dispatch_req_0_bits_ssid ? _allocPtr_T_1 : allocPtr_16; // @[StoreSet.scala 545:{23,23} 493:25]
  wire [1:0] _GEN_1427 = 5'h11 == io_dispatch_req_0_bits_ssid ? _allocPtr_T_1 : allocPtr_17; // @[StoreSet.scala 545:{23,23} 493:25]
  wire [1:0] _GEN_1428 = 5'h12 == io_dispatch_req_0_bits_ssid ? _allocPtr_T_1 : allocPtr_18; // @[StoreSet.scala 545:{23,23} 493:25]
  wire [1:0] _GEN_1429 = 5'h13 == io_dispatch_req_0_bits_ssid ? _allocPtr_T_1 : allocPtr_19; // @[StoreSet.scala 545:{23,23} 493:25]
  wire [1:0] _GEN_1430 = 5'h14 == io_dispatch_req_0_bits_ssid ? _allocPtr_T_1 : allocPtr_20; // @[StoreSet.scala 545:{23,23} 493:25]
  wire [1:0] _GEN_1431 = 5'h15 == io_dispatch_req_0_bits_ssid ? _allocPtr_T_1 : allocPtr_21; // @[StoreSet.scala 545:{23,23} 493:25]
  wire [1:0] _GEN_1432 = 5'h16 == io_dispatch_req_0_bits_ssid ? _allocPtr_T_1 : allocPtr_22; // @[StoreSet.scala 545:{23,23} 493:25]
  wire [1:0] _GEN_1433 = 5'h17 == io_dispatch_req_0_bits_ssid ? _allocPtr_T_1 : allocPtr_23; // @[StoreSet.scala 545:{23,23} 493:25]
  wire [1:0] _GEN_1434 = 5'h18 == io_dispatch_req_0_bits_ssid ? _allocPtr_T_1 : allocPtr_24; // @[StoreSet.scala 545:{23,23} 493:25]
  wire [1:0] _GEN_1435 = 5'h19 == io_dispatch_req_0_bits_ssid ? _allocPtr_T_1 : allocPtr_25; // @[StoreSet.scala 545:{23,23} 493:25]
  wire [1:0] _GEN_1436 = 5'h1a == io_dispatch_req_0_bits_ssid ? _allocPtr_T_1 : allocPtr_26; // @[StoreSet.scala 545:{23,23} 493:25]
  wire [1:0] _GEN_1437 = 5'h1b == io_dispatch_req_0_bits_ssid ? _allocPtr_T_1 : allocPtr_27; // @[StoreSet.scala 545:{23,23} 493:25]
  wire [1:0] _GEN_1438 = 5'h1c == io_dispatch_req_0_bits_ssid ? _allocPtr_T_1 : allocPtr_28; // @[StoreSet.scala 545:{23,23} 493:25]
  wire [1:0] _GEN_1439 = 5'h1d == io_dispatch_req_0_bits_ssid ? _allocPtr_T_1 : allocPtr_29; // @[StoreSet.scala 545:{23,23} 493:25]
  wire [1:0] _GEN_1440 = 5'h1e == io_dispatch_req_0_bits_ssid ? _allocPtr_T_1 : allocPtr_30; // @[StoreSet.scala 545:{23,23} 493:25]
  wire [1:0] _GEN_1441 = 5'h1f == io_dispatch_req_0_bits_ssid ? _allocPtr_T_1 : allocPtr_31; // @[StoreSet.scala 545:{23,23} 493:25]
  wire  _GEN_4891 = 2'h0 == _GEN_63; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1442 = _GEN_3874 & 2'h0 == _GEN_63 | _GEN_1090; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_4894 = 2'h1 == _GEN_63; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1443 = _GEN_3874 & 2'h1 == _GEN_63 | _GEN_1186; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_4897 = 2'h2 == _GEN_63; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1444 = _GEN_3874 & 2'h2 == _GEN_63 | _GEN_1282; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_4900 = 2'h3 == _GEN_63; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1445 = _GEN_3874 & 2'h3 == _GEN_63 | _GEN_1378; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1446 = _GEN_3880 & 2'h0 == _GEN_63 | _GEN_1091; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1447 = _GEN_3880 & 2'h1 == _GEN_63 | _GEN_1187; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1448 = _GEN_3880 & 2'h2 == _GEN_63 | _GEN_1283; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1449 = _GEN_3880 & 2'h3 == _GEN_63 | _GEN_1379; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1450 = _GEN_3888 & 2'h0 == _GEN_63 | _GEN_1092; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1451 = _GEN_3888 & 2'h1 == _GEN_63 | _GEN_1188; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1452 = _GEN_3888 & 2'h2 == _GEN_63 | _GEN_1284; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1453 = _GEN_3888 & 2'h3 == _GEN_63 | _GEN_1380; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1454 = _GEN_3896 & 2'h0 == _GEN_63 | _GEN_1093; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1455 = _GEN_3896 & 2'h1 == _GEN_63 | _GEN_1189; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1456 = _GEN_3896 & 2'h2 == _GEN_63 | _GEN_1285; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1457 = _GEN_3896 & 2'h3 == _GEN_63 | _GEN_1381; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1458 = _GEN_3904 & 2'h0 == _GEN_63 | _GEN_1094; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1459 = _GEN_3904 & 2'h1 == _GEN_63 | _GEN_1190; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1460 = _GEN_3904 & 2'h2 == _GEN_63 | _GEN_1286; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1461 = _GEN_3904 & 2'h3 == _GEN_63 | _GEN_1382; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1462 = _GEN_3912 & 2'h0 == _GEN_63 | _GEN_1095; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1463 = _GEN_3912 & 2'h1 == _GEN_63 | _GEN_1191; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1464 = _GEN_3912 & 2'h2 == _GEN_63 | _GEN_1287; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1465 = _GEN_3912 & 2'h3 == _GEN_63 | _GEN_1383; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1466 = _GEN_3920 & 2'h0 == _GEN_63 | _GEN_1096; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1467 = _GEN_3920 & 2'h1 == _GEN_63 | _GEN_1192; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1468 = _GEN_3920 & 2'h2 == _GEN_63 | _GEN_1288; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1469 = _GEN_3920 & 2'h3 == _GEN_63 | _GEN_1384; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1470 = _GEN_3928 & 2'h0 == _GEN_63 | _GEN_1097; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1471 = _GEN_3928 & 2'h1 == _GEN_63 | _GEN_1193; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1472 = _GEN_3928 & 2'h2 == _GEN_63 | _GEN_1289; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1473 = _GEN_3928 & 2'h3 == _GEN_63 | _GEN_1385; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1474 = _GEN_3936 & 2'h0 == _GEN_63 | _GEN_1098; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1475 = _GEN_3936 & 2'h1 == _GEN_63 | _GEN_1194; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1476 = _GEN_3936 & 2'h2 == _GEN_63 | _GEN_1290; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1477 = _GEN_3936 & 2'h3 == _GEN_63 | _GEN_1386; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1478 = _GEN_3944 & 2'h0 == _GEN_63 | _GEN_1099; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1479 = _GEN_3944 & 2'h1 == _GEN_63 | _GEN_1195; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1480 = _GEN_3944 & 2'h2 == _GEN_63 | _GEN_1291; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1481 = _GEN_3944 & 2'h3 == _GEN_63 | _GEN_1387; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1482 = _GEN_3952 & 2'h0 == _GEN_63 | _GEN_1100; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1483 = _GEN_3952 & 2'h1 == _GEN_63 | _GEN_1196; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1484 = _GEN_3952 & 2'h2 == _GEN_63 | _GEN_1292; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1485 = _GEN_3952 & 2'h3 == _GEN_63 | _GEN_1388; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1486 = _GEN_3960 & 2'h0 == _GEN_63 | _GEN_1101; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1487 = _GEN_3960 & 2'h1 == _GEN_63 | _GEN_1197; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1488 = _GEN_3960 & 2'h2 == _GEN_63 | _GEN_1293; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1489 = _GEN_3960 & 2'h3 == _GEN_63 | _GEN_1389; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1490 = _GEN_3968 & 2'h0 == _GEN_63 | _GEN_1102; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1491 = _GEN_3968 & 2'h1 == _GEN_63 | _GEN_1198; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1492 = _GEN_3968 & 2'h2 == _GEN_63 | _GEN_1294; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1493 = _GEN_3968 & 2'h3 == _GEN_63 | _GEN_1390; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1494 = _GEN_3976 & 2'h0 == _GEN_63 | _GEN_1103; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1495 = _GEN_3976 & 2'h1 == _GEN_63 | _GEN_1199; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1496 = _GEN_3976 & 2'h2 == _GEN_63 | _GEN_1295; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1497 = _GEN_3976 & 2'h3 == _GEN_63 | _GEN_1391; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1498 = _GEN_3984 & 2'h0 == _GEN_63 | _GEN_1104; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1499 = _GEN_3984 & 2'h1 == _GEN_63 | _GEN_1200; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1500 = _GEN_3984 & 2'h2 == _GEN_63 | _GEN_1296; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1501 = _GEN_3984 & 2'h3 == _GEN_63 | _GEN_1392; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1502 = _GEN_3992 & 2'h0 == _GEN_63 | _GEN_1105; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1503 = _GEN_3992 & 2'h1 == _GEN_63 | _GEN_1201; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1504 = _GEN_3992 & 2'h2 == _GEN_63 | _GEN_1297; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1505 = _GEN_3992 & 2'h3 == _GEN_63 | _GEN_1393; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1506 = _GEN_4000 & 2'h0 == _GEN_63 | _GEN_1106; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1507 = _GEN_4000 & 2'h1 == _GEN_63 | _GEN_1202; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1508 = _GEN_4000 & 2'h2 == _GEN_63 | _GEN_1298; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1509 = _GEN_4000 & 2'h3 == _GEN_63 | _GEN_1394; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1510 = _GEN_4008 & 2'h0 == _GEN_63 | _GEN_1107; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1511 = _GEN_4008 & 2'h1 == _GEN_63 | _GEN_1203; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1512 = _GEN_4008 & 2'h2 == _GEN_63 | _GEN_1299; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1513 = _GEN_4008 & 2'h3 == _GEN_63 | _GEN_1395; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1514 = _GEN_4016 & 2'h0 == _GEN_63 | _GEN_1108; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1515 = _GEN_4016 & 2'h1 == _GEN_63 | _GEN_1204; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1516 = _GEN_4016 & 2'h2 == _GEN_63 | _GEN_1300; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1517 = _GEN_4016 & 2'h3 == _GEN_63 | _GEN_1396; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1518 = _GEN_4024 & 2'h0 == _GEN_63 | _GEN_1109; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1519 = _GEN_4024 & 2'h1 == _GEN_63 | _GEN_1205; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1520 = _GEN_4024 & 2'h2 == _GEN_63 | _GEN_1301; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1521 = _GEN_4024 & 2'h3 == _GEN_63 | _GEN_1397; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1522 = _GEN_4032 & 2'h0 == _GEN_63 | _GEN_1110; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1523 = _GEN_4032 & 2'h1 == _GEN_63 | _GEN_1206; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1524 = _GEN_4032 & 2'h2 == _GEN_63 | _GEN_1302; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1525 = _GEN_4032 & 2'h3 == _GEN_63 | _GEN_1398; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1526 = _GEN_4040 & 2'h0 == _GEN_63 | _GEN_1111; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1527 = _GEN_4040 & 2'h1 == _GEN_63 | _GEN_1207; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1528 = _GEN_4040 & 2'h2 == _GEN_63 | _GEN_1303; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1529 = _GEN_4040 & 2'h3 == _GEN_63 | _GEN_1399; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1530 = _GEN_4048 & 2'h0 == _GEN_63 | _GEN_1112; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1531 = _GEN_4048 & 2'h1 == _GEN_63 | _GEN_1208; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1532 = _GEN_4048 & 2'h2 == _GEN_63 | _GEN_1304; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1533 = _GEN_4048 & 2'h3 == _GEN_63 | _GEN_1400; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1534 = _GEN_4056 & 2'h0 == _GEN_63 | _GEN_1113; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1535 = _GEN_4056 & 2'h1 == _GEN_63 | _GEN_1209; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1536 = _GEN_4056 & 2'h2 == _GEN_63 | _GEN_1305; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1537 = _GEN_4056 & 2'h3 == _GEN_63 | _GEN_1401; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1538 = _GEN_4064 & 2'h0 == _GEN_63 | _GEN_1114; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1539 = _GEN_4064 & 2'h1 == _GEN_63 | _GEN_1210; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1540 = _GEN_4064 & 2'h2 == _GEN_63 | _GEN_1306; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1541 = _GEN_4064 & 2'h3 == _GEN_63 | _GEN_1402; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1542 = _GEN_4072 & 2'h0 == _GEN_63 | _GEN_1115; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1543 = _GEN_4072 & 2'h1 == _GEN_63 | _GEN_1211; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1544 = _GEN_4072 & 2'h2 == _GEN_63 | _GEN_1307; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1545 = _GEN_4072 & 2'h3 == _GEN_63 | _GEN_1403; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1546 = _GEN_4080 & 2'h0 == _GEN_63 | _GEN_1116; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1547 = _GEN_4080 & 2'h1 == _GEN_63 | _GEN_1212; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1548 = _GEN_4080 & 2'h2 == _GEN_63 | _GEN_1308; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1549 = _GEN_4080 & 2'h3 == _GEN_63 | _GEN_1404; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1550 = _GEN_4088 & 2'h0 == _GEN_63 | _GEN_1117; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1551 = _GEN_4088 & 2'h1 == _GEN_63 | _GEN_1213; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1552 = _GEN_4088 & 2'h2 == _GEN_63 | _GEN_1309; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1553 = _GEN_4088 & 2'h3 == _GEN_63 | _GEN_1405; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1554 = _GEN_4096 & 2'h0 == _GEN_63 | _GEN_1118; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1555 = _GEN_4096 & 2'h1 == _GEN_63 | _GEN_1214; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1556 = _GEN_4096 & 2'h2 == _GEN_63 | _GEN_1310; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1557 = _GEN_4096 & 2'h3 == _GEN_63 | _GEN_1406; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1558 = _GEN_4104 & 2'h0 == _GEN_63 | _GEN_1119; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1559 = _GEN_4104 & 2'h1 == _GEN_63 | _GEN_1215; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1560 = _GEN_4104 & 2'h2 == _GEN_63 | _GEN_1311; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1561 = _GEN_4104 & 2'h3 == _GEN_63 | _GEN_1407; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1562 = _GEN_4112 & 2'h0 == _GEN_63 | _GEN_1120; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1563 = _GEN_4112 & 2'h1 == _GEN_63 | _GEN_1216; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1564 = _GEN_4112 & 2'h2 == _GEN_63 | _GEN_1312; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1565 = _GEN_4112 & 2'h3 == _GEN_63 | _GEN_1408; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1566 = _GEN_4120 & 2'h0 == _GEN_63 | _GEN_1121; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1567 = _GEN_4120 & 2'h1 == _GEN_63 | _GEN_1217; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1568 = _GEN_4120 & 2'h2 == _GEN_63 | _GEN_1313; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1569 = _GEN_4120 & 2'h3 == _GEN_63 | _GEN_1409; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_1570 = _GEN_3874 & _GEN_4891 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_0_0_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1571 = _GEN_3874 & _GEN_4894 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_0_1_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1572 = _GEN_3874 & _GEN_4897 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_0_2_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1573 = _GEN_3874 & _GEN_4900 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_0_3_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1574 = _GEN_3880 & _GEN_4891 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_1_0_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1575 = _GEN_3880 & _GEN_4894 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_1_1_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1576 = _GEN_3880 & _GEN_4897 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_1_2_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1577 = _GEN_3880 & _GEN_4900 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_1_3_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1578 = _GEN_3888 & _GEN_4891 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_2_0_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1579 = _GEN_3888 & _GEN_4894 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_2_1_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1580 = _GEN_3888 & _GEN_4897 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_2_2_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1581 = _GEN_3888 & _GEN_4900 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_2_3_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1582 = _GEN_3896 & _GEN_4891 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_3_0_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1583 = _GEN_3896 & _GEN_4894 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_3_1_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1584 = _GEN_3896 & _GEN_4897 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_3_2_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1585 = _GEN_3896 & _GEN_4900 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_3_3_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1586 = _GEN_3904 & _GEN_4891 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_4_0_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1587 = _GEN_3904 & _GEN_4894 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_4_1_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1588 = _GEN_3904 & _GEN_4897 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_4_2_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1589 = _GEN_3904 & _GEN_4900 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_4_3_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1590 = _GEN_3912 & _GEN_4891 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_5_0_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1591 = _GEN_3912 & _GEN_4894 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_5_1_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1592 = _GEN_3912 & _GEN_4897 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_5_2_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1593 = _GEN_3912 & _GEN_4900 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_5_3_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1594 = _GEN_3920 & _GEN_4891 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_6_0_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1595 = _GEN_3920 & _GEN_4894 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_6_1_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1596 = _GEN_3920 & _GEN_4897 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_6_2_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1597 = _GEN_3920 & _GEN_4900 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_6_3_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1598 = _GEN_3928 & _GEN_4891 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_7_0_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1599 = _GEN_3928 & _GEN_4894 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_7_1_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1600 = _GEN_3928 & _GEN_4897 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_7_2_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1601 = _GEN_3928 & _GEN_4900 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_7_3_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1602 = _GEN_3936 & _GEN_4891 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_8_0_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1603 = _GEN_3936 & _GEN_4894 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_8_1_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1604 = _GEN_3936 & _GEN_4897 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_8_2_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1605 = _GEN_3936 & _GEN_4900 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_8_3_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1606 = _GEN_3944 & _GEN_4891 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_9_0_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1607 = _GEN_3944 & _GEN_4894 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_9_1_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1608 = _GEN_3944 & _GEN_4897 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_9_2_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1609 = _GEN_3944 & _GEN_4900 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_9_3_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1610 = _GEN_3952 & _GEN_4891 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_10_0_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1611 = _GEN_3952 & _GEN_4894 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_10_1_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1612 = _GEN_3952 & _GEN_4897 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_10_2_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1613 = _GEN_3952 & _GEN_4900 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_10_3_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1614 = _GEN_3960 & _GEN_4891 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_11_0_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1615 = _GEN_3960 & _GEN_4894 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_11_1_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1616 = _GEN_3960 & _GEN_4897 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_11_2_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1617 = _GEN_3960 & _GEN_4900 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_11_3_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1618 = _GEN_3968 & _GEN_4891 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_12_0_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1619 = _GEN_3968 & _GEN_4894 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_12_1_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1620 = _GEN_3968 & _GEN_4897 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_12_2_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1621 = _GEN_3968 & _GEN_4900 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_12_3_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1622 = _GEN_3976 & _GEN_4891 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_13_0_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1623 = _GEN_3976 & _GEN_4894 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_13_1_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1624 = _GEN_3976 & _GEN_4897 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_13_2_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1625 = _GEN_3976 & _GEN_4900 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_13_3_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1626 = _GEN_3984 & _GEN_4891 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_14_0_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1627 = _GEN_3984 & _GEN_4894 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_14_1_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1628 = _GEN_3984 & _GEN_4897 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_14_2_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1629 = _GEN_3984 & _GEN_4900 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_14_3_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1630 = _GEN_3992 & _GEN_4891 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_15_0_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1631 = _GEN_3992 & _GEN_4894 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_15_1_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1632 = _GEN_3992 & _GEN_4897 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_15_2_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1633 = _GEN_3992 & _GEN_4900 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_15_3_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1634 = _GEN_4000 & _GEN_4891 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_16_0_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1635 = _GEN_4000 & _GEN_4894 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_16_1_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1636 = _GEN_4000 & _GEN_4897 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_16_2_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1637 = _GEN_4000 & _GEN_4900 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_16_3_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1638 = _GEN_4008 & _GEN_4891 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_17_0_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1639 = _GEN_4008 & _GEN_4894 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_17_1_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1640 = _GEN_4008 & _GEN_4897 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_17_2_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1641 = _GEN_4008 & _GEN_4900 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_17_3_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1642 = _GEN_4016 & _GEN_4891 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_18_0_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1643 = _GEN_4016 & _GEN_4894 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_18_1_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1644 = _GEN_4016 & _GEN_4897 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_18_2_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1645 = _GEN_4016 & _GEN_4900 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_18_3_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1646 = _GEN_4024 & _GEN_4891 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_19_0_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1647 = _GEN_4024 & _GEN_4894 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_19_1_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1648 = _GEN_4024 & _GEN_4897 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_19_2_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1649 = _GEN_4024 & _GEN_4900 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_19_3_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1650 = _GEN_4032 & _GEN_4891 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_20_0_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1651 = _GEN_4032 & _GEN_4894 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_20_1_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1652 = _GEN_4032 & _GEN_4897 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_20_2_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1653 = _GEN_4032 & _GEN_4900 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_20_3_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1654 = _GEN_4040 & _GEN_4891 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_21_0_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1655 = _GEN_4040 & _GEN_4894 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_21_1_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1656 = _GEN_4040 & _GEN_4897 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_21_2_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1657 = _GEN_4040 & _GEN_4900 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_21_3_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1658 = _GEN_4048 & _GEN_4891 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_22_0_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1659 = _GEN_4048 & _GEN_4894 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_22_1_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1660 = _GEN_4048 & _GEN_4897 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_22_2_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1661 = _GEN_4048 & _GEN_4900 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_22_3_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1662 = _GEN_4056 & _GEN_4891 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_23_0_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1663 = _GEN_4056 & _GEN_4894 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_23_1_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1664 = _GEN_4056 & _GEN_4897 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_23_2_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1665 = _GEN_4056 & _GEN_4900 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_23_3_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1666 = _GEN_4064 & _GEN_4891 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_24_0_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1667 = _GEN_4064 & _GEN_4894 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_24_1_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1668 = _GEN_4064 & _GEN_4897 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_24_2_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1669 = _GEN_4064 & _GEN_4900 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_24_3_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1670 = _GEN_4072 & _GEN_4891 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_25_0_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1671 = _GEN_4072 & _GEN_4894 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_25_1_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1672 = _GEN_4072 & _GEN_4897 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_25_2_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1673 = _GEN_4072 & _GEN_4900 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_25_3_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1674 = _GEN_4080 & _GEN_4891 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_26_0_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1675 = _GEN_4080 & _GEN_4894 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_26_1_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1676 = _GEN_4080 & _GEN_4897 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_26_2_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1677 = _GEN_4080 & _GEN_4900 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_26_3_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1678 = _GEN_4088 & _GEN_4891 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_27_0_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1679 = _GEN_4088 & _GEN_4894 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_27_1_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1680 = _GEN_4088 & _GEN_4897 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_27_2_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1681 = _GEN_4088 & _GEN_4900 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_27_3_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1682 = _GEN_4096 & _GEN_4891 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_28_0_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1683 = _GEN_4096 & _GEN_4894 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_28_1_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1684 = _GEN_4096 & _GEN_4897 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_28_2_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1685 = _GEN_4096 & _GEN_4900 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_28_3_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1686 = _GEN_4104 & _GEN_4891 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_29_0_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1687 = _GEN_4104 & _GEN_4894 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_29_1_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1688 = _GEN_4104 & _GEN_4897 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_29_2_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1689 = _GEN_4104 & _GEN_4900 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_29_3_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1690 = _GEN_4112 & _GEN_4891 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_30_0_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1691 = _GEN_4112 & _GEN_4894 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_30_1_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1692 = _GEN_4112 & _GEN_4897 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_30_2_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1693 = _GEN_4112 & _GEN_4900 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_30_3_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1694 = _GEN_4120 & _GEN_4891 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_31_0_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1695 = _GEN_4120 & _GEN_4894 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_31_1_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1696 = _GEN_4120 & _GEN_4897 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_31_2_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire  _GEN_1697 = _GEN_4120 & _GEN_4900 ? io_dispatch_req_0_bits_robIdx_flag : robIdxVec_31_3_flag; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1698 = _GEN_3874 & _GEN_4891 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_0_0_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1699 = _GEN_3874 & _GEN_4894 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_0_1_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1700 = _GEN_3874 & _GEN_4897 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_0_2_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1701 = _GEN_3874 & _GEN_4900 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_0_3_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1702 = _GEN_3880 & _GEN_4891 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_1_0_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1703 = _GEN_3880 & _GEN_4894 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_1_1_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1704 = _GEN_3880 & _GEN_4897 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_1_2_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1705 = _GEN_3880 & _GEN_4900 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_1_3_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1706 = _GEN_3888 & _GEN_4891 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_2_0_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1707 = _GEN_3888 & _GEN_4894 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_2_1_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1708 = _GEN_3888 & _GEN_4897 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_2_2_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1709 = _GEN_3888 & _GEN_4900 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_2_3_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1710 = _GEN_3896 & _GEN_4891 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_3_0_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1711 = _GEN_3896 & _GEN_4894 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_3_1_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1712 = _GEN_3896 & _GEN_4897 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_3_2_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1713 = _GEN_3896 & _GEN_4900 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_3_3_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1714 = _GEN_3904 & _GEN_4891 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_4_0_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1715 = _GEN_3904 & _GEN_4894 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_4_1_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1716 = _GEN_3904 & _GEN_4897 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_4_2_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1717 = _GEN_3904 & _GEN_4900 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_4_3_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1718 = _GEN_3912 & _GEN_4891 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_5_0_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1719 = _GEN_3912 & _GEN_4894 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_5_1_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1720 = _GEN_3912 & _GEN_4897 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_5_2_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1721 = _GEN_3912 & _GEN_4900 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_5_3_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1722 = _GEN_3920 & _GEN_4891 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_6_0_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1723 = _GEN_3920 & _GEN_4894 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_6_1_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1724 = _GEN_3920 & _GEN_4897 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_6_2_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1725 = _GEN_3920 & _GEN_4900 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_6_3_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1726 = _GEN_3928 & _GEN_4891 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_7_0_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1727 = _GEN_3928 & _GEN_4894 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_7_1_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1728 = _GEN_3928 & _GEN_4897 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_7_2_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1729 = _GEN_3928 & _GEN_4900 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_7_3_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1730 = _GEN_3936 & _GEN_4891 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_8_0_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1731 = _GEN_3936 & _GEN_4894 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_8_1_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1732 = _GEN_3936 & _GEN_4897 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_8_2_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1733 = _GEN_3936 & _GEN_4900 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_8_3_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1734 = _GEN_3944 & _GEN_4891 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_9_0_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1735 = _GEN_3944 & _GEN_4894 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_9_1_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1736 = _GEN_3944 & _GEN_4897 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_9_2_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1737 = _GEN_3944 & _GEN_4900 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_9_3_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1738 = _GEN_3952 & _GEN_4891 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_10_0_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1739 = _GEN_3952 & _GEN_4894 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_10_1_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1740 = _GEN_3952 & _GEN_4897 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_10_2_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1741 = _GEN_3952 & _GEN_4900 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_10_3_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1742 = _GEN_3960 & _GEN_4891 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_11_0_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1743 = _GEN_3960 & _GEN_4894 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_11_1_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1744 = _GEN_3960 & _GEN_4897 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_11_2_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1745 = _GEN_3960 & _GEN_4900 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_11_3_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1746 = _GEN_3968 & _GEN_4891 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_12_0_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1747 = _GEN_3968 & _GEN_4894 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_12_1_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1748 = _GEN_3968 & _GEN_4897 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_12_2_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1749 = _GEN_3968 & _GEN_4900 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_12_3_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1750 = _GEN_3976 & _GEN_4891 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_13_0_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1751 = _GEN_3976 & _GEN_4894 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_13_1_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1752 = _GEN_3976 & _GEN_4897 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_13_2_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1753 = _GEN_3976 & _GEN_4900 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_13_3_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1754 = _GEN_3984 & _GEN_4891 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_14_0_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1755 = _GEN_3984 & _GEN_4894 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_14_1_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1756 = _GEN_3984 & _GEN_4897 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_14_2_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1757 = _GEN_3984 & _GEN_4900 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_14_3_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1758 = _GEN_3992 & _GEN_4891 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_15_0_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1759 = _GEN_3992 & _GEN_4894 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_15_1_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1760 = _GEN_3992 & _GEN_4897 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_15_2_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1761 = _GEN_3992 & _GEN_4900 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_15_3_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1762 = _GEN_4000 & _GEN_4891 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_16_0_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1763 = _GEN_4000 & _GEN_4894 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_16_1_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1764 = _GEN_4000 & _GEN_4897 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_16_2_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1765 = _GEN_4000 & _GEN_4900 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_16_3_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1766 = _GEN_4008 & _GEN_4891 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_17_0_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1767 = _GEN_4008 & _GEN_4894 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_17_1_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1768 = _GEN_4008 & _GEN_4897 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_17_2_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1769 = _GEN_4008 & _GEN_4900 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_17_3_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1770 = _GEN_4016 & _GEN_4891 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_18_0_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1771 = _GEN_4016 & _GEN_4894 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_18_1_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1772 = _GEN_4016 & _GEN_4897 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_18_2_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1773 = _GEN_4016 & _GEN_4900 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_18_3_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1774 = _GEN_4024 & _GEN_4891 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_19_0_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1775 = _GEN_4024 & _GEN_4894 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_19_1_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1776 = _GEN_4024 & _GEN_4897 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_19_2_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1777 = _GEN_4024 & _GEN_4900 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_19_3_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1778 = _GEN_4032 & _GEN_4891 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_20_0_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1779 = _GEN_4032 & _GEN_4894 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_20_1_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1780 = _GEN_4032 & _GEN_4897 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_20_2_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1781 = _GEN_4032 & _GEN_4900 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_20_3_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1782 = _GEN_4040 & _GEN_4891 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_21_0_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1783 = _GEN_4040 & _GEN_4894 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_21_1_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1784 = _GEN_4040 & _GEN_4897 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_21_2_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1785 = _GEN_4040 & _GEN_4900 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_21_3_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1786 = _GEN_4048 & _GEN_4891 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_22_0_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1787 = _GEN_4048 & _GEN_4894 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_22_1_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1788 = _GEN_4048 & _GEN_4897 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_22_2_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1789 = _GEN_4048 & _GEN_4900 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_22_3_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1790 = _GEN_4056 & _GEN_4891 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_23_0_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1791 = _GEN_4056 & _GEN_4894 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_23_1_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1792 = _GEN_4056 & _GEN_4897 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_23_2_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1793 = _GEN_4056 & _GEN_4900 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_23_3_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1794 = _GEN_4064 & _GEN_4891 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_24_0_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1795 = _GEN_4064 & _GEN_4894 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_24_1_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1796 = _GEN_4064 & _GEN_4897 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_24_2_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1797 = _GEN_4064 & _GEN_4900 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_24_3_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1798 = _GEN_4072 & _GEN_4891 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_25_0_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1799 = _GEN_4072 & _GEN_4894 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_25_1_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1800 = _GEN_4072 & _GEN_4897 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_25_2_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1801 = _GEN_4072 & _GEN_4900 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_25_3_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1802 = _GEN_4080 & _GEN_4891 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_26_0_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1803 = _GEN_4080 & _GEN_4894 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_26_1_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1804 = _GEN_4080 & _GEN_4897 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_26_2_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1805 = _GEN_4080 & _GEN_4900 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_26_3_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1806 = _GEN_4088 & _GEN_4891 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_27_0_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1807 = _GEN_4088 & _GEN_4894 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_27_1_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1808 = _GEN_4088 & _GEN_4897 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_27_2_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1809 = _GEN_4088 & _GEN_4900 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_27_3_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1810 = _GEN_4096 & _GEN_4891 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_28_0_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1811 = _GEN_4096 & _GEN_4894 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_28_1_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1812 = _GEN_4096 & _GEN_4897 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_28_2_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1813 = _GEN_4096 & _GEN_4900 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_28_3_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1814 = _GEN_4104 & _GEN_4891 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_29_0_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1815 = _GEN_4104 & _GEN_4894 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_29_1_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1816 = _GEN_4104 & _GEN_4897 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_29_2_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1817 = _GEN_4104 & _GEN_4900 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_29_3_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1818 = _GEN_4112 & _GEN_4891 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_30_0_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1819 = _GEN_4112 & _GEN_4894 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_30_1_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1820 = _GEN_4112 & _GEN_4897 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_30_2_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1821 = _GEN_4112 & _GEN_4900 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_30_3_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1822 = _GEN_4120 & _GEN_4891 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_31_0_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1823 = _GEN_4120 & _GEN_4894 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_31_1_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1824 = _GEN_4120 & _GEN_4897 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_31_2_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [4:0] _GEN_1825 = _GEN_4120 & _GEN_4900 ? io_dispatch_req_0_bits_robIdx_value : robIdxVec_31_3_value; // @[StoreSet.scala 492:22 547:{30,30}]
  wire [1:0] _GEN_1826 = _hitInDispatchBundleVec_T ? _GEN_1410 : allocPtr_0; // @[StoreSet.scala 493:25 542:70]
  wire [1:0] _GEN_1827 = _hitInDispatchBundleVec_T ? _GEN_1411 : allocPtr_1; // @[StoreSet.scala 493:25 542:70]
  wire [1:0] _GEN_1828 = _hitInDispatchBundleVec_T ? _GEN_1412 : allocPtr_2; // @[StoreSet.scala 493:25 542:70]
  wire [1:0] _GEN_1829 = _hitInDispatchBundleVec_T ? _GEN_1413 : allocPtr_3; // @[StoreSet.scala 493:25 542:70]
  wire [1:0] _GEN_1830 = _hitInDispatchBundleVec_T ? _GEN_1414 : allocPtr_4; // @[StoreSet.scala 493:25 542:70]
  wire [1:0] _GEN_1831 = _hitInDispatchBundleVec_T ? _GEN_1415 : allocPtr_5; // @[StoreSet.scala 493:25 542:70]
  wire [1:0] _GEN_1832 = _hitInDispatchBundleVec_T ? _GEN_1416 : allocPtr_6; // @[StoreSet.scala 493:25 542:70]
  wire [1:0] _GEN_1833 = _hitInDispatchBundleVec_T ? _GEN_1417 : allocPtr_7; // @[StoreSet.scala 493:25 542:70]
  wire [1:0] _GEN_1834 = _hitInDispatchBundleVec_T ? _GEN_1418 : allocPtr_8; // @[StoreSet.scala 493:25 542:70]
  wire [1:0] _GEN_1835 = _hitInDispatchBundleVec_T ? _GEN_1419 : allocPtr_9; // @[StoreSet.scala 493:25 542:70]
  wire [1:0] _GEN_1836 = _hitInDispatchBundleVec_T ? _GEN_1420 : allocPtr_10; // @[StoreSet.scala 493:25 542:70]
  wire [1:0] _GEN_1837 = _hitInDispatchBundleVec_T ? _GEN_1421 : allocPtr_11; // @[StoreSet.scala 493:25 542:70]
  wire [1:0] _GEN_1838 = _hitInDispatchBundleVec_T ? _GEN_1422 : allocPtr_12; // @[StoreSet.scala 493:25 542:70]
  wire [1:0] _GEN_1839 = _hitInDispatchBundleVec_T ? _GEN_1423 : allocPtr_13; // @[StoreSet.scala 493:25 542:70]
  wire [1:0] _GEN_1840 = _hitInDispatchBundleVec_T ? _GEN_1424 : allocPtr_14; // @[StoreSet.scala 493:25 542:70]
  wire [1:0] _GEN_1841 = _hitInDispatchBundleVec_T ? _GEN_1425 : allocPtr_15; // @[StoreSet.scala 493:25 542:70]
  wire [1:0] _GEN_1842 = _hitInDispatchBundleVec_T ? _GEN_1426 : allocPtr_16; // @[StoreSet.scala 493:25 542:70]
  wire [1:0] _GEN_1843 = _hitInDispatchBundleVec_T ? _GEN_1427 : allocPtr_17; // @[StoreSet.scala 493:25 542:70]
  wire [1:0] _GEN_1844 = _hitInDispatchBundleVec_T ? _GEN_1428 : allocPtr_18; // @[StoreSet.scala 493:25 542:70]
  wire [1:0] _GEN_1845 = _hitInDispatchBundleVec_T ? _GEN_1429 : allocPtr_19; // @[StoreSet.scala 493:25 542:70]
  wire [1:0] _GEN_1846 = _hitInDispatchBundleVec_T ? _GEN_1430 : allocPtr_20; // @[StoreSet.scala 493:25 542:70]
  wire [1:0] _GEN_1847 = _hitInDispatchBundleVec_T ? _GEN_1431 : allocPtr_21; // @[StoreSet.scala 493:25 542:70]
  wire [1:0] _GEN_1848 = _hitInDispatchBundleVec_T ? _GEN_1432 : allocPtr_22; // @[StoreSet.scala 493:25 542:70]
  wire [1:0] _GEN_1849 = _hitInDispatchBundleVec_T ? _GEN_1433 : allocPtr_23; // @[StoreSet.scala 493:25 542:70]
  wire [1:0] _GEN_1850 = _hitInDispatchBundleVec_T ? _GEN_1434 : allocPtr_24; // @[StoreSet.scala 493:25 542:70]
  wire [1:0] _GEN_1851 = _hitInDispatchBundleVec_T ? _GEN_1435 : allocPtr_25; // @[StoreSet.scala 493:25 542:70]
  wire [1:0] _GEN_1852 = _hitInDispatchBundleVec_T ? _GEN_1436 : allocPtr_26; // @[StoreSet.scala 493:25 542:70]
  wire [1:0] _GEN_1853 = _hitInDispatchBundleVec_T ? _GEN_1437 : allocPtr_27; // @[StoreSet.scala 493:25 542:70]
  wire [1:0] _GEN_1854 = _hitInDispatchBundleVec_T ? _GEN_1438 : allocPtr_28; // @[StoreSet.scala 493:25 542:70]
  wire [1:0] _GEN_1855 = _hitInDispatchBundleVec_T ? _GEN_1439 : allocPtr_29; // @[StoreSet.scala 493:25 542:70]
  wire [1:0] _GEN_1856 = _hitInDispatchBundleVec_T ? _GEN_1440 : allocPtr_30; // @[StoreSet.scala 493:25 542:70]
  wire [1:0] _GEN_1857 = _hitInDispatchBundleVec_T ? _GEN_1441 : allocPtr_31; // @[StoreSet.scala 493:25 542:70]
  wire  _GEN_1858 = _hitInDispatchBundleVec_T ? _GEN_1442 : _GEN_1090; // @[StoreSet.scala 542:70]
  wire  _GEN_1859 = _hitInDispatchBundleVec_T ? _GEN_1443 : _GEN_1186; // @[StoreSet.scala 542:70]
  wire  _GEN_1860 = _hitInDispatchBundleVec_T ? _GEN_1444 : _GEN_1282; // @[StoreSet.scala 542:70]
  wire  _GEN_1861 = _hitInDispatchBundleVec_T ? _GEN_1445 : _GEN_1378; // @[StoreSet.scala 542:70]
  wire  _GEN_1862 = _hitInDispatchBundleVec_T ? _GEN_1446 : _GEN_1091; // @[StoreSet.scala 542:70]
  wire  _GEN_1863 = _hitInDispatchBundleVec_T ? _GEN_1447 : _GEN_1187; // @[StoreSet.scala 542:70]
  wire  _GEN_1864 = _hitInDispatchBundleVec_T ? _GEN_1448 : _GEN_1283; // @[StoreSet.scala 542:70]
  wire  _GEN_1865 = _hitInDispatchBundleVec_T ? _GEN_1449 : _GEN_1379; // @[StoreSet.scala 542:70]
  wire  _GEN_1866 = _hitInDispatchBundleVec_T ? _GEN_1450 : _GEN_1092; // @[StoreSet.scala 542:70]
  wire  _GEN_1867 = _hitInDispatchBundleVec_T ? _GEN_1451 : _GEN_1188; // @[StoreSet.scala 542:70]
  wire  _GEN_1868 = _hitInDispatchBundleVec_T ? _GEN_1452 : _GEN_1284; // @[StoreSet.scala 542:70]
  wire  _GEN_1869 = _hitInDispatchBundleVec_T ? _GEN_1453 : _GEN_1380; // @[StoreSet.scala 542:70]
  wire  _GEN_1870 = _hitInDispatchBundleVec_T ? _GEN_1454 : _GEN_1093; // @[StoreSet.scala 542:70]
  wire  _GEN_1871 = _hitInDispatchBundleVec_T ? _GEN_1455 : _GEN_1189; // @[StoreSet.scala 542:70]
  wire  _GEN_1872 = _hitInDispatchBundleVec_T ? _GEN_1456 : _GEN_1285; // @[StoreSet.scala 542:70]
  wire  _GEN_1873 = _hitInDispatchBundleVec_T ? _GEN_1457 : _GEN_1381; // @[StoreSet.scala 542:70]
  wire  _GEN_1874 = _hitInDispatchBundleVec_T ? _GEN_1458 : _GEN_1094; // @[StoreSet.scala 542:70]
  wire  _GEN_1875 = _hitInDispatchBundleVec_T ? _GEN_1459 : _GEN_1190; // @[StoreSet.scala 542:70]
  wire  _GEN_1876 = _hitInDispatchBundleVec_T ? _GEN_1460 : _GEN_1286; // @[StoreSet.scala 542:70]
  wire  _GEN_1877 = _hitInDispatchBundleVec_T ? _GEN_1461 : _GEN_1382; // @[StoreSet.scala 542:70]
  wire  _GEN_1878 = _hitInDispatchBundleVec_T ? _GEN_1462 : _GEN_1095; // @[StoreSet.scala 542:70]
  wire  _GEN_1879 = _hitInDispatchBundleVec_T ? _GEN_1463 : _GEN_1191; // @[StoreSet.scala 542:70]
  wire  _GEN_1880 = _hitInDispatchBundleVec_T ? _GEN_1464 : _GEN_1287; // @[StoreSet.scala 542:70]
  wire  _GEN_1881 = _hitInDispatchBundleVec_T ? _GEN_1465 : _GEN_1383; // @[StoreSet.scala 542:70]
  wire  _GEN_1882 = _hitInDispatchBundleVec_T ? _GEN_1466 : _GEN_1096; // @[StoreSet.scala 542:70]
  wire  _GEN_1883 = _hitInDispatchBundleVec_T ? _GEN_1467 : _GEN_1192; // @[StoreSet.scala 542:70]
  wire  _GEN_1884 = _hitInDispatchBundleVec_T ? _GEN_1468 : _GEN_1288; // @[StoreSet.scala 542:70]
  wire  _GEN_1885 = _hitInDispatchBundleVec_T ? _GEN_1469 : _GEN_1384; // @[StoreSet.scala 542:70]
  wire  _GEN_1886 = _hitInDispatchBundleVec_T ? _GEN_1470 : _GEN_1097; // @[StoreSet.scala 542:70]
  wire  _GEN_1887 = _hitInDispatchBundleVec_T ? _GEN_1471 : _GEN_1193; // @[StoreSet.scala 542:70]
  wire  _GEN_1888 = _hitInDispatchBundleVec_T ? _GEN_1472 : _GEN_1289; // @[StoreSet.scala 542:70]
  wire  _GEN_1889 = _hitInDispatchBundleVec_T ? _GEN_1473 : _GEN_1385; // @[StoreSet.scala 542:70]
  wire  _GEN_1890 = _hitInDispatchBundleVec_T ? _GEN_1474 : _GEN_1098; // @[StoreSet.scala 542:70]
  wire  _GEN_1891 = _hitInDispatchBundleVec_T ? _GEN_1475 : _GEN_1194; // @[StoreSet.scala 542:70]
  wire  _GEN_1892 = _hitInDispatchBundleVec_T ? _GEN_1476 : _GEN_1290; // @[StoreSet.scala 542:70]
  wire  _GEN_1893 = _hitInDispatchBundleVec_T ? _GEN_1477 : _GEN_1386; // @[StoreSet.scala 542:70]
  wire  _GEN_1894 = _hitInDispatchBundleVec_T ? _GEN_1478 : _GEN_1099; // @[StoreSet.scala 542:70]
  wire  _GEN_1895 = _hitInDispatchBundleVec_T ? _GEN_1479 : _GEN_1195; // @[StoreSet.scala 542:70]
  wire  _GEN_1896 = _hitInDispatchBundleVec_T ? _GEN_1480 : _GEN_1291; // @[StoreSet.scala 542:70]
  wire  _GEN_1897 = _hitInDispatchBundleVec_T ? _GEN_1481 : _GEN_1387; // @[StoreSet.scala 542:70]
  wire  _GEN_1898 = _hitInDispatchBundleVec_T ? _GEN_1482 : _GEN_1100; // @[StoreSet.scala 542:70]
  wire  _GEN_1899 = _hitInDispatchBundleVec_T ? _GEN_1483 : _GEN_1196; // @[StoreSet.scala 542:70]
  wire  _GEN_1900 = _hitInDispatchBundleVec_T ? _GEN_1484 : _GEN_1292; // @[StoreSet.scala 542:70]
  wire  _GEN_1901 = _hitInDispatchBundleVec_T ? _GEN_1485 : _GEN_1388; // @[StoreSet.scala 542:70]
  wire  _GEN_1902 = _hitInDispatchBundleVec_T ? _GEN_1486 : _GEN_1101; // @[StoreSet.scala 542:70]
  wire  _GEN_1903 = _hitInDispatchBundleVec_T ? _GEN_1487 : _GEN_1197; // @[StoreSet.scala 542:70]
  wire  _GEN_1904 = _hitInDispatchBundleVec_T ? _GEN_1488 : _GEN_1293; // @[StoreSet.scala 542:70]
  wire  _GEN_1905 = _hitInDispatchBundleVec_T ? _GEN_1489 : _GEN_1389; // @[StoreSet.scala 542:70]
  wire  _GEN_1906 = _hitInDispatchBundleVec_T ? _GEN_1490 : _GEN_1102; // @[StoreSet.scala 542:70]
  wire  _GEN_1907 = _hitInDispatchBundleVec_T ? _GEN_1491 : _GEN_1198; // @[StoreSet.scala 542:70]
  wire  _GEN_1908 = _hitInDispatchBundleVec_T ? _GEN_1492 : _GEN_1294; // @[StoreSet.scala 542:70]
  wire  _GEN_1909 = _hitInDispatchBundleVec_T ? _GEN_1493 : _GEN_1390; // @[StoreSet.scala 542:70]
  wire  _GEN_1910 = _hitInDispatchBundleVec_T ? _GEN_1494 : _GEN_1103; // @[StoreSet.scala 542:70]
  wire  _GEN_1911 = _hitInDispatchBundleVec_T ? _GEN_1495 : _GEN_1199; // @[StoreSet.scala 542:70]
  wire  _GEN_1912 = _hitInDispatchBundleVec_T ? _GEN_1496 : _GEN_1295; // @[StoreSet.scala 542:70]
  wire  _GEN_1913 = _hitInDispatchBundleVec_T ? _GEN_1497 : _GEN_1391; // @[StoreSet.scala 542:70]
  wire  _GEN_1914 = _hitInDispatchBundleVec_T ? _GEN_1498 : _GEN_1104; // @[StoreSet.scala 542:70]
  wire  _GEN_1915 = _hitInDispatchBundleVec_T ? _GEN_1499 : _GEN_1200; // @[StoreSet.scala 542:70]
  wire  _GEN_1916 = _hitInDispatchBundleVec_T ? _GEN_1500 : _GEN_1296; // @[StoreSet.scala 542:70]
  wire  _GEN_1917 = _hitInDispatchBundleVec_T ? _GEN_1501 : _GEN_1392; // @[StoreSet.scala 542:70]
  wire  _GEN_1918 = _hitInDispatchBundleVec_T ? _GEN_1502 : _GEN_1105; // @[StoreSet.scala 542:70]
  wire  _GEN_1919 = _hitInDispatchBundleVec_T ? _GEN_1503 : _GEN_1201; // @[StoreSet.scala 542:70]
  wire  _GEN_1920 = _hitInDispatchBundleVec_T ? _GEN_1504 : _GEN_1297; // @[StoreSet.scala 542:70]
  wire  _GEN_1921 = _hitInDispatchBundleVec_T ? _GEN_1505 : _GEN_1393; // @[StoreSet.scala 542:70]
  wire  _GEN_1922 = _hitInDispatchBundleVec_T ? _GEN_1506 : _GEN_1106; // @[StoreSet.scala 542:70]
  wire  _GEN_1923 = _hitInDispatchBundleVec_T ? _GEN_1507 : _GEN_1202; // @[StoreSet.scala 542:70]
  wire  _GEN_1924 = _hitInDispatchBundleVec_T ? _GEN_1508 : _GEN_1298; // @[StoreSet.scala 542:70]
  wire  _GEN_1925 = _hitInDispatchBundleVec_T ? _GEN_1509 : _GEN_1394; // @[StoreSet.scala 542:70]
  wire  _GEN_1926 = _hitInDispatchBundleVec_T ? _GEN_1510 : _GEN_1107; // @[StoreSet.scala 542:70]
  wire  _GEN_1927 = _hitInDispatchBundleVec_T ? _GEN_1511 : _GEN_1203; // @[StoreSet.scala 542:70]
  wire  _GEN_1928 = _hitInDispatchBundleVec_T ? _GEN_1512 : _GEN_1299; // @[StoreSet.scala 542:70]
  wire  _GEN_1929 = _hitInDispatchBundleVec_T ? _GEN_1513 : _GEN_1395; // @[StoreSet.scala 542:70]
  wire  _GEN_1930 = _hitInDispatchBundleVec_T ? _GEN_1514 : _GEN_1108; // @[StoreSet.scala 542:70]
  wire  _GEN_1931 = _hitInDispatchBundleVec_T ? _GEN_1515 : _GEN_1204; // @[StoreSet.scala 542:70]
  wire  _GEN_1932 = _hitInDispatchBundleVec_T ? _GEN_1516 : _GEN_1300; // @[StoreSet.scala 542:70]
  wire  _GEN_1933 = _hitInDispatchBundleVec_T ? _GEN_1517 : _GEN_1396; // @[StoreSet.scala 542:70]
  wire  _GEN_1934 = _hitInDispatchBundleVec_T ? _GEN_1518 : _GEN_1109; // @[StoreSet.scala 542:70]
  wire  _GEN_1935 = _hitInDispatchBundleVec_T ? _GEN_1519 : _GEN_1205; // @[StoreSet.scala 542:70]
  wire  _GEN_1936 = _hitInDispatchBundleVec_T ? _GEN_1520 : _GEN_1301; // @[StoreSet.scala 542:70]
  wire  _GEN_1937 = _hitInDispatchBundleVec_T ? _GEN_1521 : _GEN_1397; // @[StoreSet.scala 542:70]
  wire  _GEN_1938 = _hitInDispatchBundleVec_T ? _GEN_1522 : _GEN_1110; // @[StoreSet.scala 542:70]
  wire  _GEN_1939 = _hitInDispatchBundleVec_T ? _GEN_1523 : _GEN_1206; // @[StoreSet.scala 542:70]
  wire  _GEN_1940 = _hitInDispatchBundleVec_T ? _GEN_1524 : _GEN_1302; // @[StoreSet.scala 542:70]
  wire  _GEN_1941 = _hitInDispatchBundleVec_T ? _GEN_1525 : _GEN_1398; // @[StoreSet.scala 542:70]
  wire  _GEN_1942 = _hitInDispatchBundleVec_T ? _GEN_1526 : _GEN_1111; // @[StoreSet.scala 542:70]
  wire  _GEN_1943 = _hitInDispatchBundleVec_T ? _GEN_1527 : _GEN_1207; // @[StoreSet.scala 542:70]
  wire  _GEN_1944 = _hitInDispatchBundleVec_T ? _GEN_1528 : _GEN_1303; // @[StoreSet.scala 542:70]
  wire  _GEN_1945 = _hitInDispatchBundleVec_T ? _GEN_1529 : _GEN_1399; // @[StoreSet.scala 542:70]
  wire  _GEN_1946 = _hitInDispatchBundleVec_T ? _GEN_1530 : _GEN_1112; // @[StoreSet.scala 542:70]
  wire  _GEN_1947 = _hitInDispatchBundleVec_T ? _GEN_1531 : _GEN_1208; // @[StoreSet.scala 542:70]
  wire  _GEN_1948 = _hitInDispatchBundleVec_T ? _GEN_1532 : _GEN_1304; // @[StoreSet.scala 542:70]
  wire  _GEN_1949 = _hitInDispatchBundleVec_T ? _GEN_1533 : _GEN_1400; // @[StoreSet.scala 542:70]
  wire  _GEN_1950 = _hitInDispatchBundleVec_T ? _GEN_1534 : _GEN_1113; // @[StoreSet.scala 542:70]
  wire  _GEN_1951 = _hitInDispatchBundleVec_T ? _GEN_1535 : _GEN_1209; // @[StoreSet.scala 542:70]
  wire  _GEN_1952 = _hitInDispatchBundleVec_T ? _GEN_1536 : _GEN_1305; // @[StoreSet.scala 542:70]
  wire  _GEN_1953 = _hitInDispatchBundleVec_T ? _GEN_1537 : _GEN_1401; // @[StoreSet.scala 542:70]
  wire  _GEN_1954 = _hitInDispatchBundleVec_T ? _GEN_1538 : _GEN_1114; // @[StoreSet.scala 542:70]
  wire  _GEN_1955 = _hitInDispatchBundleVec_T ? _GEN_1539 : _GEN_1210; // @[StoreSet.scala 542:70]
  wire  _GEN_1956 = _hitInDispatchBundleVec_T ? _GEN_1540 : _GEN_1306; // @[StoreSet.scala 542:70]
  wire  _GEN_1957 = _hitInDispatchBundleVec_T ? _GEN_1541 : _GEN_1402; // @[StoreSet.scala 542:70]
  wire  _GEN_1958 = _hitInDispatchBundleVec_T ? _GEN_1542 : _GEN_1115; // @[StoreSet.scala 542:70]
  wire  _GEN_1959 = _hitInDispatchBundleVec_T ? _GEN_1543 : _GEN_1211; // @[StoreSet.scala 542:70]
  wire  _GEN_1960 = _hitInDispatchBundleVec_T ? _GEN_1544 : _GEN_1307; // @[StoreSet.scala 542:70]
  wire  _GEN_1961 = _hitInDispatchBundleVec_T ? _GEN_1545 : _GEN_1403; // @[StoreSet.scala 542:70]
  wire  _GEN_1962 = _hitInDispatchBundleVec_T ? _GEN_1546 : _GEN_1116; // @[StoreSet.scala 542:70]
  wire  _GEN_1963 = _hitInDispatchBundleVec_T ? _GEN_1547 : _GEN_1212; // @[StoreSet.scala 542:70]
  wire  _GEN_1964 = _hitInDispatchBundleVec_T ? _GEN_1548 : _GEN_1308; // @[StoreSet.scala 542:70]
  wire  _GEN_1965 = _hitInDispatchBundleVec_T ? _GEN_1549 : _GEN_1404; // @[StoreSet.scala 542:70]
  wire  _GEN_1966 = _hitInDispatchBundleVec_T ? _GEN_1550 : _GEN_1117; // @[StoreSet.scala 542:70]
  wire  _GEN_1967 = _hitInDispatchBundleVec_T ? _GEN_1551 : _GEN_1213; // @[StoreSet.scala 542:70]
  wire  _GEN_1968 = _hitInDispatchBundleVec_T ? _GEN_1552 : _GEN_1309; // @[StoreSet.scala 542:70]
  wire  _GEN_1969 = _hitInDispatchBundleVec_T ? _GEN_1553 : _GEN_1405; // @[StoreSet.scala 542:70]
  wire  _GEN_1970 = _hitInDispatchBundleVec_T ? _GEN_1554 : _GEN_1118; // @[StoreSet.scala 542:70]
  wire  _GEN_1971 = _hitInDispatchBundleVec_T ? _GEN_1555 : _GEN_1214; // @[StoreSet.scala 542:70]
  wire  _GEN_1972 = _hitInDispatchBundleVec_T ? _GEN_1556 : _GEN_1310; // @[StoreSet.scala 542:70]
  wire  _GEN_1973 = _hitInDispatchBundleVec_T ? _GEN_1557 : _GEN_1406; // @[StoreSet.scala 542:70]
  wire  _GEN_1974 = _hitInDispatchBundleVec_T ? _GEN_1558 : _GEN_1119; // @[StoreSet.scala 542:70]
  wire  _GEN_1975 = _hitInDispatchBundleVec_T ? _GEN_1559 : _GEN_1215; // @[StoreSet.scala 542:70]
  wire  _GEN_1976 = _hitInDispatchBundleVec_T ? _GEN_1560 : _GEN_1311; // @[StoreSet.scala 542:70]
  wire  _GEN_1977 = _hitInDispatchBundleVec_T ? _GEN_1561 : _GEN_1407; // @[StoreSet.scala 542:70]
  wire  _GEN_1978 = _hitInDispatchBundleVec_T ? _GEN_1562 : _GEN_1120; // @[StoreSet.scala 542:70]
  wire  _GEN_1979 = _hitInDispatchBundleVec_T ? _GEN_1563 : _GEN_1216; // @[StoreSet.scala 542:70]
  wire  _GEN_1980 = _hitInDispatchBundleVec_T ? _GEN_1564 : _GEN_1312; // @[StoreSet.scala 542:70]
  wire  _GEN_1981 = _hitInDispatchBundleVec_T ? _GEN_1565 : _GEN_1408; // @[StoreSet.scala 542:70]
  wire  _GEN_1982 = _hitInDispatchBundleVec_T ? _GEN_1566 : _GEN_1121; // @[StoreSet.scala 542:70]
  wire  _GEN_1983 = _hitInDispatchBundleVec_T ? _GEN_1567 : _GEN_1217; // @[StoreSet.scala 542:70]
  wire  _GEN_1984 = _hitInDispatchBundleVec_T ? _GEN_1568 : _GEN_1313; // @[StoreSet.scala 542:70]
  wire  _GEN_1985 = _hitInDispatchBundleVec_T ? _GEN_1569 : _GEN_1409; // @[StoreSet.scala 542:70]
  wire  _GEN_1986 = _hitInDispatchBundleVec_T ? _GEN_1570 : robIdxVec_0_0_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_1987 = _hitInDispatchBundleVec_T ? _GEN_1571 : robIdxVec_0_1_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_1988 = _hitInDispatchBundleVec_T ? _GEN_1572 : robIdxVec_0_2_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_1989 = _hitInDispatchBundleVec_T ? _GEN_1573 : robIdxVec_0_3_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_1990 = _hitInDispatchBundleVec_T ? _GEN_1574 : robIdxVec_1_0_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_1991 = _hitInDispatchBundleVec_T ? _GEN_1575 : robIdxVec_1_1_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_1992 = _hitInDispatchBundleVec_T ? _GEN_1576 : robIdxVec_1_2_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_1993 = _hitInDispatchBundleVec_T ? _GEN_1577 : robIdxVec_1_3_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_1994 = _hitInDispatchBundleVec_T ? _GEN_1578 : robIdxVec_2_0_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_1995 = _hitInDispatchBundleVec_T ? _GEN_1579 : robIdxVec_2_1_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_1996 = _hitInDispatchBundleVec_T ? _GEN_1580 : robIdxVec_2_2_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_1997 = _hitInDispatchBundleVec_T ? _GEN_1581 : robIdxVec_2_3_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_1998 = _hitInDispatchBundleVec_T ? _GEN_1582 : robIdxVec_3_0_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_1999 = _hitInDispatchBundleVec_T ? _GEN_1583 : robIdxVec_3_1_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2000 = _hitInDispatchBundleVec_T ? _GEN_1584 : robIdxVec_3_2_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2001 = _hitInDispatchBundleVec_T ? _GEN_1585 : robIdxVec_3_3_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2002 = _hitInDispatchBundleVec_T ? _GEN_1586 : robIdxVec_4_0_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2003 = _hitInDispatchBundleVec_T ? _GEN_1587 : robIdxVec_4_1_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2004 = _hitInDispatchBundleVec_T ? _GEN_1588 : robIdxVec_4_2_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2005 = _hitInDispatchBundleVec_T ? _GEN_1589 : robIdxVec_4_3_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2006 = _hitInDispatchBundleVec_T ? _GEN_1590 : robIdxVec_5_0_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2007 = _hitInDispatchBundleVec_T ? _GEN_1591 : robIdxVec_5_1_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2008 = _hitInDispatchBundleVec_T ? _GEN_1592 : robIdxVec_5_2_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2009 = _hitInDispatchBundleVec_T ? _GEN_1593 : robIdxVec_5_3_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2010 = _hitInDispatchBundleVec_T ? _GEN_1594 : robIdxVec_6_0_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2011 = _hitInDispatchBundleVec_T ? _GEN_1595 : robIdxVec_6_1_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2012 = _hitInDispatchBundleVec_T ? _GEN_1596 : robIdxVec_6_2_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2013 = _hitInDispatchBundleVec_T ? _GEN_1597 : robIdxVec_6_3_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2014 = _hitInDispatchBundleVec_T ? _GEN_1598 : robIdxVec_7_0_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2015 = _hitInDispatchBundleVec_T ? _GEN_1599 : robIdxVec_7_1_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2016 = _hitInDispatchBundleVec_T ? _GEN_1600 : robIdxVec_7_2_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2017 = _hitInDispatchBundleVec_T ? _GEN_1601 : robIdxVec_7_3_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2018 = _hitInDispatchBundleVec_T ? _GEN_1602 : robIdxVec_8_0_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2019 = _hitInDispatchBundleVec_T ? _GEN_1603 : robIdxVec_8_1_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2020 = _hitInDispatchBundleVec_T ? _GEN_1604 : robIdxVec_8_2_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2021 = _hitInDispatchBundleVec_T ? _GEN_1605 : robIdxVec_8_3_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2022 = _hitInDispatchBundleVec_T ? _GEN_1606 : robIdxVec_9_0_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2023 = _hitInDispatchBundleVec_T ? _GEN_1607 : robIdxVec_9_1_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2024 = _hitInDispatchBundleVec_T ? _GEN_1608 : robIdxVec_9_2_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2025 = _hitInDispatchBundleVec_T ? _GEN_1609 : robIdxVec_9_3_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2026 = _hitInDispatchBundleVec_T ? _GEN_1610 : robIdxVec_10_0_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2027 = _hitInDispatchBundleVec_T ? _GEN_1611 : robIdxVec_10_1_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2028 = _hitInDispatchBundleVec_T ? _GEN_1612 : robIdxVec_10_2_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2029 = _hitInDispatchBundleVec_T ? _GEN_1613 : robIdxVec_10_3_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2030 = _hitInDispatchBundleVec_T ? _GEN_1614 : robIdxVec_11_0_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2031 = _hitInDispatchBundleVec_T ? _GEN_1615 : robIdxVec_11_1_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2032 = _hitInDispatchBundleVec_T ? _GEN_1616 : robIdxVec_11_2_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2033 = _hitInDispatchBundleVec_T ? _GEN_1617 : robIdxVec_11_3_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2034 = _hitInDispatchBundleVec_T ? _GEN_1618 : robIdxVec_12_0_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2035 = _hitInDispatchBundleVec_T ? _GEN_1619 : robIdxVec_12_1_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2036 = _hitInDispatchBundleVec_T ? _GEN_1620 : robIdxVec_12_2_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2037 = _hitInDispatchBundleVec_T ? _GEN_1621 : robIdxVec_12_3_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2038 = _hitInDispatchBundleVec_T ? _GEN_1622 : robIdxVec_13_0_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2039 = _hitInDispatchBundleVec_T ? _GEN_1623 : robIdxVec_13_1_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2040 = _hitInDispatchBundleVec_T ? _GEN_1624 : robIdxVec_13_2_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2041 = _hitInDispatchBundleVec_T ? _GEN_1625 : robIdxVec_13_3_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2042 = _hitInDispatchBundleVec_T ? _GEN_1626 : robIdxVec_14_0_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2043 = _hitInDispatchBundleVec_T ? _GEN_1627 : robIdxVec_14_1_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2044 = _hitInDispatchBundleVec_T ? _GEN_1628 : robIdxVec_14_2_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2045 = _hitInDispatchBundleVec_T ? _GEN_1629 : robIdxVec_14_3_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2046 = _hitInDispatchBundleVec_T ? _GEN_1630 : robIdxVec_15_0_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2047 = _hitInDispatchBundleVec_T ? _GEN_1631 : robIdxVec_15_1_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2048 = _hitInDispatchBundleVec_T ? _GEN_1632 : robIdxVec_15_2_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2049 = _hitInDispatchBundleVec_T ? _GEN_1633 : robIdxVec_15_3_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2050 = _hitInDispatchBundleVec_T ? _GEN_1634 : robIdxVec_16_0_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2051 = _hitInDispatchBundleVec_T ? _GEN_1635 : robIdxVec_16_1_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2052 = _hitInDispatchBundleVec_T ? _GEN_1636 : robIdxVec_16_2_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2053 = _hitInDispatchBundleVec_T ? _GEN_1637 : robIdxVec_16_3_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2054 = _hitInDispatchBundleVec_T ? _GEN_1638 : robIdxVec_17_0_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2055 = _hitInDispatchBundleVec_T ? _GEN_1639 : robIdxVec_17_1_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2056 = _hitInDispatchBundleVec_T ? _GEN_1640 : robIdxVec_17_2_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2057 = _hitInDispatchBundleVec_T ? _GEN_1641 : robIdxVec_17_3_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2058 = _hitInDispatchBundleVec_T ? _GEN_1642 : robIdxVec_18_0_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2059 = _hitInDispatchBundleVec_T ? _GEN_1643 : robIdxVec_18_1_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2060 = _hitInDispatchBundleVec_T ? _GEN_1644 : robIdxVec_18_2_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2061 = _hitInDispatchBundleVec_T ? _GEN_1645 : robIdxVec_18_3_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2062 = _hitInDispatchBundleVec_T ? _GEN_1646 : robIdxVec_19_0_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2063 = _hitInDispatchBundleVec_T ? _GEN_1647 : robIdxVec_19_1_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2064 = _hitInDispatchBundleVec_T ? _GEN_1648 : robIdxVec_19_2_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2065 = _hitInDispatchBundleVec_T ? _GEN_1649 : robIdxVec_19_3_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2066 = _hitInDispatchBundleVec_T ? _GEN_1650 : robIdxVec_20_0_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2067 = _hitInDispatchBundleVec_T ? _GEN_1651 : robIdxVec_20_1_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2068 = _hitInDispatchBundleVec_T ? _GEN_1652 : robIdxVec_20_2_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2069 = _hitInDispatchBundleVec_T ? _GEN_1653 : robIdxVec_20_3_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2070 = _hitInDispatchBundleVec_T ? _GEN_1654 : robIdxVec_21_0_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2071 = _hitInDispatchBundleVec_T ? _GEN_1655 : robIdxVec_21_1_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2072 = _hitInDispatchBundleVec_T ? _GEN_1656 : robIdxVec_21_2_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2073 = _hitInDispatchBundleVec_T ? _GEN_1657 : robIdxVec_21_3_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2074 = _hitInDispatchBundleVec_T ? _GEN_1658 : robIdxVec_22_0_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2075 = _hitInDispatchBundleVec_T ? _GEN_1659 : robIdxVec_22_1_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2076 = _hitInDispatchBundleVec_T ? _GEN_1660 : robIdxVec_22_2_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2077 = _hitInDispatchBundleVec_T ? _GEN_1661 : robIdxVec_22_3_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2078 = _hitInDispatchBundleVec_T ? _GEN_1662 : robIdxVec_23_0_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2079 = _hitInDispatchBundleVec_T ? _GEN_1663 : robIdxVec_23_1_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2080 = _hitInDispatchBundleVec_T ? _GEN_1664 : robIdxVec_23_2_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2081 = _hitInDispatchBundleVec_T ? _GEN_1665 : robIdxVec_23_3_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2082 = _hitInDispatchBundleVec_T ? _GEN_1666 : robIdxVec_24_0_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2083 = _hitInDispatchBundleVec_T ? _GEN_1667 : robIdxVec_24_1_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2084 = _hitInDispatchBundleVec_T ? _GEN_1668 : robIdxVec_24_2_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2085 = _hitInDispatchBundleVec_T ? _GEN_1669 : robIdxVec_24_3_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2086 = _hitInDispatchBundleVec_T ? _GEN_1670 : robIdxVec_25_0_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2087 = _hitInDispatchBundleVec_T ? _GEN_1671 : robIdxVec_25_1_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2088 = _hitInDispatchBundleVec_T ? _GEN_1672 : robIdxVec_25_2_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2089 = _hitInDispatchBundleVec_T ? _GEN_1673 : robIdxVec_25_3_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2090 = _hitInDispatchBundleVec_T ? _GEN_1674 : robIdxVec_26_0_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2091 = _hitInDispatchBundleVec_T ? _GEN_1675 : robIdxVec_26_1_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2092 = _hitInDispatchBundleVec_T ? _GEN_1676 : robIdxVec_26_2_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2093 = _hitInDispatchBundleVec_T ? _GEN_1677 : robIdxVec_26_3_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2094 = _hitInDispatchBundleVec_T ? _GEN_1678 : robIdxVec_27_0_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2095 = _hitInDispatchBundleVec_T ? _GEN_1679 : robIdxVec_27_1_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2096 = _hitInDispatchBundleVec_T ? _GEN_1680 : robIdxVec_27_2_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2097 = _hitInDispatchBundleVec_T ? _GEN_1681 : robIdxVec_27_3_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2098 = _hitInDispatchBundleVec_T ? _GEN_1682 : robIdxVec_28_0_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2099 = _hitInDispatchBundleVec_T ? _GEN_1683 : robIdxVec_28_1_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2100 = _hitInDispatchBundleVec_T ? _GEN_1684 : robIdxVec_28_2_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2101 = _hitInDispatchBundleVec_T ? _GEN_1685 : robIdxVec_28_3_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2102 = _hitInDispatchBundleVec_T ? _GEN_1686 : robIdxVec_29_0_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2103 = _hitInDispatchBundleVec_T ? _GEN_1687 : robIdxVec_29_1_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2104 = _hitInDispatchBundleVec_T ? _GEN_1688 : robIdxVec_29_2_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2105 = _hitInDispatchBundleVec_T ? _GEN_1689 : robIdxVec_29_3_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2106 = _hitInDispatchBundleVec_T ? _GEN_1690 : robIdxVec_30_0_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2107 = _hitInDispatchBundleVec_T ? _GEN_1691 : robIdxVec_30_1_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2108 = _hitInDispatchBundleVec_T ? _GEN_1692 : robIdxVec_30_2_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2109 = _hitInDispatchBundleVec_T ? _GEN_1693 : robIdxVec_30_3_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2110 = _hitInDispatchBundleVec_T ? _GEN_1694 : robIdxVec_31_0_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2111 = _hitInDispatchBundleVec_T ? _GEN_1695 : robIdxVec_31_1_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2112 = _hitInDispatchBundleVec_T ? _GEN_1696 : robIdxVec_31_2_flag; // @[StoreSet.scala 492:22 542:70]
  wire  _GEN_2113 = _hitInDispatchBundleVec_T ? _GEN_1697 : robIdxVec_31_3_flag; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2114 = _hitInDispatchBundleVec_T ? _GEN_1698 : robIdxVec_0_0_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2115 = _hitInDispatchBundleVec_T ? _GEN_1699 : robIdxVec_0_1_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2116 = _hitInDispatchBundleVec_T ? _GEN_1700 : robIdxVec_0_2_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2117 = _hitInDispatchBundleVec_T ? _GEN_1701 : robIdxVec_0_3_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2118 = _hitInDispatchBundleVec_T ? _GEN_1702 : robIdxVec_1_0_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2119 = _hitInDispatchBundleVec_T ? _GEN_1703 : robIdxVec_1_1_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2120 = _hitInDispatchBundleVec_T ? _GEN_1704 : robIdxVec_1_2_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2121 = _hitInDispatchBundleVec_T ? _GEN_1705 : robIdxVec_1_3_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2122 = _hitInDispatchBundleVec_T ? _GEN_1706 : robIdxVec_2_0_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2123 = _hitInDispatchBundleVec_T ? _GEN_1707 : robIdxVec_2_1_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2124 = _hitInDispatchBundleVec_T ? _GEN_1708 : robIdxVec_2_2_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2125 = _hitInDispatchBundleVec_T ? _GEN_1709 : robIdxVec_2_3_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2126 = _hitInDispatchBundleVec_T ? _GEN_1710 : robIdxVec_3_0_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2127 = _hitInDispatchBundleVec_T ? _GEN_1711 : robIdxVec_3_1_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2128 = _hitInDispatchBundleVec_T ? _GEN_1712 : robIdxVec_3_2_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2129 = _hitInDispatchBundleVec_T ? _GEN_1713 : robIdxVec_3_3_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2130 = _hitInDispatchBundleVec_T ? _GEN_1714 : robIdxVec_4_0_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2131 = _hitInDispatchBundleVec_T ? _GEN_1715 : robIdxVec_4_1_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2132 = _hitInDispatchBundleVec_T ? _GEN_1716 : robIdxVec_4_2_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2133 = _hitInDispatchBundleVec_T ? _GEN_1717 : robIdxVec_4_3_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2134 = _hitInDispatchBundleVec_T ? _GEN_1718 : robIdxVec_5_0_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2135 = _hitInDispatchBundleVec_T ? _GEN_1719 : robIdxVec_5_1_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2136 = _hitInDispatchBundleVec_T ? _GEN_1720 : robIdxVec_5_2_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2137 = _hitInDispatchBundleVec_T ? _GEN_1721 : robIdxVec_5_3_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2138 = _hitInDispatchBundleVec_T ? _GEN_1722 : robIdxVec_6_0_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2139 = _hitInDispatchBundleVec_T ? _GEN_1723 : robIdxVec_6_1_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2140 = _hitInDispatchBundleVec_T ? _GEN_1724 : robIdxVec_6_2_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2141 = _hitInDispatchBundleVec_T ? _GEN_1725 : robIdxVec_6_3_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2142 = _hitInDispatchBundleVec_T ? _GEN_1726 : robIdxVec_7_0_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2143 = _hitInDispatchBundleVec_T ? _GEN_1727 : robIdxVec_7_1_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2144 = _hitInDispatchBundleVec_T ? _GEN_1728 : robIdxVec_7_2_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2145 = _hitInDispatchBundleVec_T ? _GEN_1729 : robIdxVec_7_3_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2146 = _hitInDispatchBundleVec_T ? _GEN_1730 : robIdxVec_8_0_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2147 = _hitInDispatchBundleVec_T ? _GEN_1731 : robIdxVec_8_1_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2148 = _hitInDispatchBundleVec_T ? _GEN_1732 : robIdxVec_8_2_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2149 = _hitInDispatchBundleVec_T ? _GEN_1733 : robIdxVec_8_3_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2150 = _hitInDispatchBundleVec_T ? _GEN_1734 : robIdxVec_9_0_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2151 = _hitInDispatchBundleVec_T ? _GEN_1735 : robIdxVec_9_1_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2152 = _hitInDispatchBundleVec_T ? _GEN_1736 : robIdxVec_9_2_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2153 = _hitInDispatchBundleVec_T ? _GEN_1737 : robIdxVec_9_3_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2154 = _hitInDispatchBundleVec_T ? _GEN_1738 : robIdxVec_10_0_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2155 = _hitInDispatchBundleVec_T ? _GEN_1739 : robIdxVec_10_1_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2156 = _hitInDispatchBundleVec_T ? _GEN_1740 : robIdxVec_10_2_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2157 = _hitInDispatchBundleVec_T ? _GEN_1741 : robIdxVec_10_3_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2158 = _hitInDispatchBundleVec_T ? _GEN_1742 : robIdxVec_11_0_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2159 = _hitInDispatchBundleVec_T ? _GEN_1743 : robIdxVec_11_1_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2160 = _hitInDispatchBundleVec_T ? _GEN_1744 : robIdxVec_11_2_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2161 = _hitInDispatchBundleVec_T ? _GEN_1745 : robIdxVec_11_3_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2162 = _hitInDispatchBundleVec_T ? _GEN_1746 : robIdxVec_12_0_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2163 = _hitInDispatchBundleVec_T ? _GEN_1747 : robIdxVec_12_1_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2164 = _hitInDispatchBundleVec_T ? _GEN_1748 : robIdxVec_12_2_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2165 = _hitInDispatchBundleVec_T ? _GEN_1749 : robIdxVec_12_3_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2166 = _hitInDispatchBundleVec_T ? _GEN_1750 : robIdxVec_13_0_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2167 = _hitInDispatchBundleVec_T ? _GEN_1751 : robIdxVec_13_1_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2168 = _hitInDispatchBundleVec_T ? _GEN_1752 : robIdxVec_13_2_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2169 = _hitInDispatchBundleVec_T ? _GEN_1753 : robIdxVec_13_3_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2170 = _hitInDispatchBundleVec_T ? _GEN_1754 : robIdxVec_14_0_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2171 = _hitInDispatchBundleVec_T ? _GEN_1755 : robIdxVec_14_1_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2172 = _hitInDispatchBundleVec_T ? _GEN_1756 : robIdxVec_14_2_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2173 = _hitInDispatchBundleVec_T ? _GEN_1757 : robIdxVec_14_3_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2174 = _hitInDispatchBundleVec_T ? _GEN_1758 : robIdxVec_15_0_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2175 = _hitInDispatchBundleVec_T ? _GEN_1759 : robIdxVec_15_1_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2176 = _hitInDispatchBundleVec_T ? _GEN_1760 : robIdxVec_15_2_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2177 = _hitInDispatchBundleVec_T ? _GEN_1761 : robIdxVec_15_3_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2178 = _hitInDispatchBundleVec_T ? _GEN_1762 : robIdxVec_16_0_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2179 = _hitInDispatchBundleVec_T ? _GEN_1763 : robIdxVec_16_1_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2180 = _hitInDispatchBundleVec_T ? _GEN_1764 : robIdxVec_16_2_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2181 = _hitInDispatchBundleVec_T ? _GEN_1765 : robIdxVec_16_3_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2182 = _hitInDispatchBundleVec_T ? _GEN_1766 : robIdxVec_17_0_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2183 = _hitInDispatchBundleVec_T ? _GEN_1767 : robIdxVec_17_1_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2184 = _hitInDispatchBundleVec_T ? _GEN_1768 : robIdxVec_17_2_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2185 = _hitInDispatchBundleVec_T ? _GEN_1769 : robIdxVec_17_3_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2186 = _hitInDispatchBundleVec_T ? _GEN_1770 : robIdxVec_18_0_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2187 = _hitInDispatchBundleVec_T ? _GEN_1771 : robIdxVec_18_1_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2188 = _hitInDispatchBundleVec_T ? _GEN_1772 : robIdxVec_18_2_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2189 = _hitInDispatchBundleVec_T ? _GEN_1773 : robIdxVec_18_3_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2190 = _hitInDispatchBundleVec_T ? _GEN_1774 : robIdxVec_19_0_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2191 = _hitInDispatchBundleVec_T ? _GEN_1775 : robIdxVec_19_1_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2192 = _hitInDispatchBundleVec_T ? _GEN_1776 : robIdxVec_19_2_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2193 = _hitInDispatchBundleVec_T ? _GEN_1777 : robIdxVec_19_3_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2194 = _hitInDispatchBundleVec_T ? _GEN_1778 : robIdxVec_20_0_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2195 = _hitInDispatchBundleVec_T ? _GEN_1779 : robIdxVec_20_1_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2196 = _hitInDispatchBundleVec_T ? _GEN_1780 : robIdxVec_20_2_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2197 = _hitInDispatchBundleVec_T ? _GEN_1781 : robIdxVec_20_3_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2198 = _hitInDispatchBundleVec_T ? _GEN_1782 : robIdxVec_21_0_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2199 = _hitInDispatchBundleVec_T ? _GEN_1783 : robIdxVec_21_1_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2200 = _hitInDispatchBundleVec_T ? _GEN_1784 : robIdxVec_21_2_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2201 = _hitInDispatchBundleVec_T ? _GEN_1785 : robIdxVec_21_3_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2202 = _hitInDispatchBundleVec_T ? _GEN_1786 : robIdxVec_22_0_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2203 = _hitInDispatchBundleVec_T ? _GEN_1787 : robIdxVec_22_1_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2204 = _hitInDispatchBundleVec_T ? _GEN_1788 : robIdxVec_22_2_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2205 = _hitInDispatchBundleVec_T ? _GEN_1789 : robIdxVec_22_3_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2206 = _hitInDispatchBundleVec_T ? _GEN_1790 : robIdxVec_23_0_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2207 = _hitInDispatchBundleVec_T ? _GEN_1791 : robIdxVec_23_1_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2208 = _hitInDispatchBundleVec_T ? _GEN_1792 : robIdxVec_23_2_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2209 = _hitInDispatchBundleVec_T ? _GEN_1793 : robIdxVec_23_3_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2210 = _hitInDispatchBundleVec_T ? _GEN_1794 : robIdxVec_24_0_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2211 = _hitInDispatchBundleVec_T ? _GEN_1795 : robIdxVec_24_1_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2212 = _hitInDispatchBundleVec_T ? _GEN_1796 : robIdxVec_24_2_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2213 = _hitInDispatchBundleVec_T ? _GEN_1797 : robIdxVec_24_3_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2214 = _hitInDispatchBundleVec_T ? _GEN_1798 : robIdxVec_25_0_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2215 = _hitInDispatchBundleVec_T ? _GEN_1799 : robIdxVec_25_1_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2216 = _hitInDispatchBundleVec_T ? _GEN_1800 : robIdxVec_25_2_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2217 = _hitInDispatchBundleVec_T ? _GEN_1801 : robIdxVec_25_3_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2218 = _hitInDispatchBundleVec_T ? _GEN_1802 : robIdxVec_26_0_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2219 = _hitInDispatchBundleVec_T ? _GEN_1803 : robIdxVec_26_1_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2220 = _hitInDispatchBundleVec_T ? _GEN_1804 : robIdxVec_26_2_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2221 = _hitInDispatchBundleVec_T ? _GEN_1805 : robIdxVec_26_3_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2222 = _hitInDispatchBundleVec_T ? _GEN_1806 : robIdxVec_27_0_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2223 = _hitInDispatchBundleVec_T ? _GEN_1807 : robIdxVec_27_1_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2224 = _hitInDispatchBundleVec_T ? _GEN_1808 : robIdxVec_27_2_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2225 = _hitInDispatchBundleVec_T ? _GEN_1809 : robIdxVec_27_3_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2226 = _hitInDispatchBundleVec_T ? _GEN_1810 : robIdxVec_28_0_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2227 = _hitInDispatchBundleVec_T ? _GEN_1811 : robIdxVec_28_1_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2228 = _hitInDispatchBundleVec_T ? _GEN_1812 : robIdxVec_28_2_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2229 = _hitInDispatchBundleVec_T ? _GEN_1813 : robIdxVec_28_3_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2230 = _hitInDispatchBundleVec_T ? _GEN_1814 : robIdxVec_29_0_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2231 = _hitInDispatchBundleVec_T ? _GEN_1815 : robIdxVec_29_1_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2232 = _hitInDispatchBundleVec_T ? _GEN_1816 : robIdxVec_29_2_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2233 = _hitInDispatchBundleVec_T ? _GEN_1817 : robIdxVec_29_3_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2234 = _hitInDispatchBundleVec_T ? _GEN_1818 : robIdxVec_30_0_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2235 = _hitInDispatchBundleVec_T ? _GEN_1819 : robIdxVec_30_1_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2236 = _hitInDispatchBundleVec_T ? _GEN_1820 : robIdxVec_30_2_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2237 = _hitInDispatchBundleVec_T ? _GEN_1821 : robIdxVec_30_3_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2238 = _hitInDispatchBundleVec_T ? _GEN_1822 : robIdxVec_31_0_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2239 = _hitInDispatchBundleVec_T ? _GEN_1823 : robIdxVec_31_1_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2240 = _hitInDispatchBundleVec_T ? _GEN_1824 : robIdxVec_31_2_value; // @[StoreSet.scala 492:22 542:70]
  wire [4:0] _GEN_2241 = _hitInDispatchBundleVec_T ? _GEN_1825 : robIdxVec_31_3_value; // @[StoreSet.scala 492:22 542:70]
  wire [1:0] _allocPtr_T_3 = _GEN_383 + 2'h1; // @[StoreSet.scala 545:42]
  wire [1:0] _GEN_2242 = 5'h0 == io_dispatch_req_1_bits_ssid ? _allocPtr_T_3 : _GEN_1826; // @[StoreSet.scala 545:{23,23}]
  wire [1:0] _GEN_2243 = 5'h1 == io_dispatch_req_1_bits_ssid ? _allocPtr_T_3 : _GEN_1827; // @[StoreSet.scala 545:{23,23}]
  wire [1:0] _GEN_2244 = 5'h2 == io_dispatch_req_1_bits_ssid ? _allocPtr_T_3 : _GEN_1828; // @[StoreSet.scala 545:{23,23}]
  wire [1:0] _GEN_2245 = 5'h3 == io_dispatch_req_1_bits_ssid ? _allocPtr_T_3 : _GEN_1829; // @[StoreSet.scala 545:{23,23}]
  wire [1:0] _GEN_2246 = 5'h4 == io_dispatch_req_1_bits_ssid ? _allocPtr_T_3 : _GEN_1830; // @[StoreSet.scala 545:{23,23}]
  wire [1:0] _GEN_2247 = 5'h5 == io_dispatch_req_1_bits_ssid ? _allocPtr_T_3 : _GEN_1831; // @[StoreSet.scala 545:{23,23}]
  wire [1:0] _GEN_2248 = 5'h6 == io_dispatch_req_1_bits_ssid ? _allocPtr_T_3 : _GEN_1832; // @[StoreSet.scala 545:{23,23}]
  wire [1:0] _GEN_2249 = 5'h7 == io_dispatch_req_1_bits_ssid ? _allocPtr_T_3 : _GEN_1833; // @[StoreSet.scala 545:{23,23}]
  wire [1:0] _GEN_2250 = 5'h8 == io_dispatch_req_1_bits_ssid ? _allocPtr_T_3 : _GEN_1834; // @[StoreSet.scala 545:{23,23}]
  wire [1:0] _GEN_2251 = 5'h9 == io_dispatch_req_1_bits_ssid ? _allocPtr_T_3 : _GEN_1835; // @[StoreSet.scala 545:{23,23}]
  wire [1:0] _GEN_2252 = 5'ha == io_dispatch_req_1_bits_ssid ? _allocPtr_T_3 : _GEN_1836; // @[StoreSet.scala 545:{23,23}]
  wire [1:0] _GEN_2253 = 5'hb == io_dispatch_req_1_bits_ssid ? _allocPtr_T_3 : _GEN_1837; // @[StoreSet.scala 545:{23,23}]
  wire [1:0] _GEN_2254 = 5'hc == io_dispatch_req_1_bits_ssid ? _allocPtr_T_3 : _GEN_1838; // @[StoreSet.scala 545:{23,23}]
  wire [1:0] _GEN_2255 = 5'hd == io_dispatch_req_1_bits_ssid ? _allocPtr_T_3 : _GEN_1839; // @[StoreSet.scala 545:{23,23}]
  wire [1:0] _GEN_2256 = 5'he == io_dispatch_req_1_bits_ssid ? _allocPtr_T_3 : _GEN_1840; // @[StoreSet.scala 545:{23,23}]
  wire [1:0] _GEN_2257 = 5'hf == io_dispatch_req_1_bits_ssid ? _allocPtr_T_3 : _GEN_1841; // @[StoreSet.scala 545:{23,23}]
  wire [1:0] _GEN_2258 = 5'h10 == io_dispatch_req_1_bits_ssid ? _allocPtr_T_3 : _GEN_1842; // @[StoreSet.scala 545:{23,23}]
  wire [1:0] _GEN_2259 = 5'h11 == io_dispatch_req_1_bits_ssid ? _allocPtr_T_3 : _GEN_1843; // @[StoreSet.scala 545:{23,23}]
  wire [1:0] _GEN_2260 = 5'h12 == io_dispatch_req_1_bits_ssid ? _allocPtr_T_3 : _GEN_1844; // @[StoreSet.scala 545:{23,23}]
  wire [1:0] _GEN_2261 = 5'h13 == io_dispatch_req_1_bits_ssid ? _allocPtr_T_3 : _GEN_1845; // @[StoreSet.scala 545:{23,23}]
  wire [1:0] _GEN_2262 = 5'h14 == io_dispatch_req_1_bits_ssid ? _allocPtr_T_3 : _GEN_1846; // @[StoreSet.scala 545:{23,23}]
  wire [1:0] _GEN_2263 = 5'h15 == io_dispatch_req_1_bits_ssid ? _allocPtr_T_3 : _GEN_1847; // @[StoreSet.scala 545:{23,23}]
  wire [1:0] _GEN_2264 = 5'h16 == io_dispatch_req_1_bits_ssid ? _allocPtr_T_3 : _GEN_1848; // @[StoreSet.scala 545:{23,23}]
  wire [1:0] _GEN_2265 = 5'h17 == io_dispatch_req_1_bits_ssid ? _allocPtr_T_3 : _GEN_1849; // @[StoreSet.scala 545:{23,23}]
  wire [1:0] _GEN_2266 = 5'h18 == io_dispatch_req_1_bits_ssid ? _allocPtr_T_3 : _GEN_1850; // @[StoreSet.scala 545:{23,23}]
  wire [1:0] _GEN_2267 = 5'h19 == io_dispatch_req_1_bits_ssid ? _allocPtr_T_3 : _GEN_1851; // @[StoreSet.scala 545:{23,23}]
  wire [1:0] _GEN_2268 = 5'h1a == io_dispatch_req_1_bits_ssid ? _allocPtr_T_3 : _GEN_1852; // @[StoreSet.scala 545:{23,23}]
  wire [1:0] _GEN_2269 = 5'h1b == io_dispatch_req_1_bits_ssid ? _allocPtr_T_3 : _GEN_1853; // @[StoreSet.scala 545:{23,23}]
  wire [1:0] _GEN_2270 = 5'h1c == io_dispatch_req_1_bits_ssid ? _allocPtr_T_3 : _GEN_1854; // @[StoreSet.scala 545:{23,23}]
  wire [1:0] _GEN_2271 = 5'h1d == io_dispatch_req_1_bits_ssid ? _allocPtr_T_3 : _GEN_1855; // @[StoreSet.scala 545:{23,23}]
  wire [1:0] _GEN_2272 = 5'h1e == io_dispatch_req_1_bits_ssid ? _allocPtr_T_3 : _GEN_1856; // @[StoreSet.scala 545:{23,23}]
  wire [1:0] _GEN_2273 = 5'h1f == io_dispatch_req_1_bits_ssid ? _allocPtr_T_3 : _GEN_1857; // @[StoreSet.scala 545:{23,23}]
  wire  _GEN_5787 = 2'h0 == _GEN_383; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2274 = _GEN_4382 & 2'h0 == _GEN_383 | _GEN_1858; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_5790 = 2'h1 == _GEN_383; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2275 = _GEN_4382 & 2'h1 == _GEN_383 | _GEN_1859; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_5793 = 2'h2 == _GEN_383; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2276 = _GEN_4382 & 2'h2 == _GEN_383 | _GEN_1860; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_5796 = 2'h3 == _GEN_383; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2277 = _GEN_4382 & 2'h3 == _GEN_383 | _GEN_1861; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2278 = _GEN_4388 & 2'h0 == _GEN_383 | _GEN_1862; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2279 = _GEN_4388 & 2'h1 == _GEN_383 | _GEN_1863; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2280 = _GEN_4388 & 2'h2 == _GEN_383 | _GEN_1864; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2281 = _GEN_4388 & 2'h3 == _GEN_383 | _GEN_1865; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2282 = _GEN_4396 & 2'h0 == _GEN_383 | _GEN_1866; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2283 = _GEN_4396 & 2'h1 == _GEN_383 | _GEN_1867; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2284 = _GEN_4396 & 2'h2 == _GEN_383 | _GEN_1868; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2285 = _GEN_4396 & 2'h3 == _GEN_383 | _GEN_1869; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2286 = _GEN_4404 & 2'h0 == _GEN_383 | _GEN_1870; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2287 = _GEN_4404 & 2'h1 == _GEN_383 | _GEN_1871; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2288 = _GEN_4404 & 2'h2 == _GEN_383 | _GEN_1872; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2289 = _GEN_4404 & 2'h3 == _GEN_383 | _GEN_1873; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2290 = _GEN_4412 & 2'h0 == _GEN_383 | _GEN_1874; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2291 = _GEN_4412 & 2'h1 == _GEN_383 | _GEN_1875; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2292 = _GEN_4412 & 2'h2 == _GEN_383 | _GEN_1876; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2293 = _GEN_4412 & 2'h3 == _GEN_383 | _GEN_1877; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2294 = _GEN_4420 & 2'h0 == _GEN_383 | _GEN_1878; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2295 = _GEN_4420 & 2'h1 == _GEN_383 | _GEN_1879; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2296 = _GEN_4420 & 2'h2 == _GEN_383 | _GEN_1880; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2297 = _GEN_4420 & 2'h3 == _GEN_383 | _GEN_1881; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2298 = _GEN_4428 & 2'h0 == _GEN_383 | _GEN_1882; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2299 = _GEN_4428 & 2'h1 == _GEN_383 | _GEN_1883; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2300 = _GEN_4428 & 2'h2 == _GEN_383 | _GEN_1884; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2301 = _GEN_4428 & 2'h3 == _GEN_383 | _GEN_1885; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2302 = _GEN_4436 & 2'h0 == _GEN_383 | _GEN_1886; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2303 = _GEN_4436 & 2'h1 == _GEN_383 | _GEN_1887; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2304 = _GEN_4436 & 2'h2 == _GEN_383 | _GEN_1888; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2305 = _GEN_4436 & 2'h3 == _GEN_383 | _GEN_1889; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2306 = _GEN_4444 & 2'h0 == _GEN_383 | _GEN_1890; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2307 = _GEN_4444 & 2'h1 == _GEN_383 | _GEN_1891; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2308 = _GEN_4444 & 2'h2 == _GEN_383 | _GEN_1892; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2309 = _GEN_4444 & 2'h3 == _GEN_383 | _GEN_1893; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2310 = _GEN_4452 & 2'h0 == _GEN_383 | _GEN_1894; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2311 = _GEN_4452 & 2'h1 == _GEN_383 | _GEN_1895; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2312 = _GEN_4452 & 2'h2 == _GEN_383 | _GEN_1896; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2313 = _GEN_4452 & 2'h3 == _GEN_383 | _GEN_1897; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2314 = _GEN_4460 & 2'h0 == _GEN_383 | _GEN_1898; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2315 = _GEN_4460 & 2'h1 == _GEN_383 | _GEN_1899; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2316 = _GEN_4460 & 2'h2 == _GEN_383 | _GEN_1900; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2317 = _GEN_4460 & 2'h3 == _GEN_383 | _GEN_1901; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2318 = _GEN_4468 & 2'h0 == _GEN_383 | _GEN_1902; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2319 = _GEN_4468 & 2'h1 == _GEN_383 | _GEN_1903; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2320 = _GEN_4468 & 2'h2 == _GEN_383 | _GEN_1904; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2321 = _GEN_4468 & 2'h3 == _GEN_383 | _GEN_1905; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2322 = _GEN_4476 & 2'h0 == _GEN_383 | _GEN_1906; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2323 = _GEN_4476 & 2'h1 == _GEN_383 | _GEN_1907; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2324 = _GEN_4476 & 2'h2 == _GEN_383 | _GEN_1908; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2325 = _GEN_4476 & 2'h3 == _GEN_383 | _GEN_1909; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2326 = _GEN_4484 & 2'h0 == _GEN_383 | _GEN_1910; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2327 = _GEN_4484 & 2'h1 == _GEN_383 | _GEN_1911; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2328 = _GEN_4484 & 2'h2 == _GEN_383 | _GEN_1912; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2329 = _GEN_4484 & 2'h3 == _GEN_383 | _GEN_1913; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2330 = _GEN_4492 & 2'h0 == _GEN_383 | _GEN_1914; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2331 = _GEN_4492 & 2'h1 == _GEN_383 | _GEN_1915; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2332 = _GEN_4492 & 2'h2 == _GEN_383 | _GEN_1916; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2333 = _GEN_4492 & 2'h3 == _GEN_383 | _GEN_1917; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2334 = _GEN_4500 & 2'h0 == _GEN_383 | _GEN_1918; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2335 = _GEN_4500 & 2'h1 == _GEN_383 | _GEN_1919; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2336 = _GEN_4500 & 2'h2 == _GEN_383 | _GEN_1920; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2337 = _GEN_4500 & 2'h3 == _GEN_383 | _GEN_1921; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2338 = _GEN_4508 & 2'h0 == _GEN_383 | _GEN_1922; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2339 = _GEN_4508 & 2'h1 == _GEN_383 | _GEN_1923; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2340 = _GEN_4508 & 2'h2 == _GEN_383 | _GEN_1924; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2341 = _GEN_4508 & 2'h3 == _GEN_383 | _GEN_1925; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2342 = _GEN_4516 & 2'h0 == _GEN_383 | _GEN_1926; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2343 = _GEN_4516 & 2'h1 == _GEN_383 | _GEN_1927; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2344 = _GEN_4516 & 2'h2 == _GEN_383 | _GEN_1928; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2345 = _GEN_4516 & 2'h3 == _GEN_383 | _GEN_1929; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2346 = _GEN_4524 & 2'h0 == _GEN_383 | _GEN_1930; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2347 = _GEN_4524 & 2'h1 == _GEN_383 | _GEN_1931; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2348 = _GEN_4524 & 2'h2 == _GEN_383 | _GEN_1932; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2349 = _GEN_4524 & 2'h3 == _GEN_383 | _GEN_1933; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2350 = _GEN_4532 & 2'h0 == _GEN_383 | _GEN_1934; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2351 = _GEN_4532 & 2'h1 == _GEN_383 | _GEN_1935; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2352 = _GEN_4532 & 2'h2 == _GEN_383 | _GEN_1936; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2353 = _GEN_4532 & 2'h3 == _GEN_383 | _GEN_1937; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2354 = _GEN_4540 & 2'h0 == _GEN_383 | _GEN_1938; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2355 = _GEN_4540 & 2'h1 == _GEN_383 | _GEN_1939; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2356 = _GEN_4540 & 2'h2 == _GEN_383 | _GEN_1940; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2357 = _GEN_4540 & 2'h3 == _GEN_383 | _GEN_1941; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2358 = _GEN_4548 & 2'h0 == _GEN_383 | _GEN_1942; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2359 = _GEN_4548 & 2'h1 == _GEN_383 | _GEN_1943; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2360 = _GEN_4548 & 2'h2 == _GEN_383 | _GEN_1944; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2361 = _GEN_4548 & 2'h3 == _GEN_383 | _GEN_1945; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2362 = _GEN_4556 & 2'h0 == _GEN_383 | _GEN_1946; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2363 = _GEN_4556 & 2'h1 == _GEN_383 | _GEN_1947; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2364 = _GEN_4556 & 2'h2 == _GEN_383 | _GEN_1948; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2365 = _GEN_4556 & 2'h3 == _GEN_383 | _GEN_1949; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2366 = _GEN_4564 & 2'h0 == _GEN_383 | _GEN_1950; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2367 = _GEN_4564 & 2'h1 == _GEN_383 | _GEN_1951; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2368 = _GEN_4564 & 2'h2 == _GEN_383 | _GEN_1952; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2369 = _GEN_4564 & 2'h3 == _GEN_383 | _GEN_1953; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2370 = _GEN_4572 & 2'h0 == _GEN_383 | _GEN_1954; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2371 = _GEN_4572 & 2'h1 == _GEN_383 | _GEN_1955; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2372 = _GEN_4572 & 2'h2 == _GEN_383 | _GEN_1956; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2373 = _GEN_4572 & 2'h3 == _GEN_383 | _GEN_1957; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2374 = _GEN_4580 & 2'h0 == _GEN_383 | _GEN_1958; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2375 = _GEN_4580 & 2'h1 == _GEN_383 | _GEN_1959; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2376 = _GEN_4580 & 2'h2 == _GEN_383 | _GEN_1960; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2377 = _GEN_4580 & 2'h3 == _GEN_383 | _GEN_1961; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2378 = _GEN_4588 & 2'h0 == _GEN_383 | _GEN_1962; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2379 = _GEN_4588 & 2'h1 == _GEN_383 | _GEN_1963; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2380 = _GEN_4588 & 2'h2 == _GEN_383 | _GEN_1964; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2381 = _GEN_4588 & 2'h3 == _GEN_383 | _GEN_1965; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2382 = _GEN_4596 & 2'h0 == _GEN_383 | _GEN_1966; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2383 = _GEN_4596 & 2'h1 == _GEN_383 | _GEN_1967; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2384 = _GEN_4596 & 2'h2 == _GEN_383 | _GEN_1968; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2385 = _GEN_4596 & 2'h3 == _GEN_383 | _GEN_1969; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2386 = _GEN_4604 & 2'h0 == _GEN_383 | _GEN_1970; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2387 = _GEN_4604 & 2'h1 == _GEN_383 | _GEN_1971; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2388 = _GEN_4604 & 2'h2 == _GEN_383 | _GEN_1972; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2389 = _GEN_4604 & 2'h3 == _GEN_383 | _GEN_1973; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2390 = _GEN_4612 & 2'h0 == _GEN_383 | _GEN_1974; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2391 = _GEN_4612 & 2'h1 == _GEN_383 | _GEN_1975; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2392 = _GEN_4612 & 2'h2 == _GEN_383 | _GEN_1976; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2393 = _GEN_4612 & 2'h3 == _GEN_383 | _GEN_1977; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2394 = _GEN_4620 & 2'h0 == _GEN_383 | _GEN_1978; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2395 = _GEN_4620 & 2'h1 == _GEN_383 | _GEN_1979; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2396 = _GEN_4620 & 2'h2 == _GEN_383 | _GEN_1980; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2397 = _GEN_4620 & 2'h3 == _GEN_383 | _GEN_1981; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2398 = _GEN_4628 & 2'h0 == _GEN_383 | _GEN_1982; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2399 = _GEN_4628 & 2'h1 == _GEN_383 | _GEN_1983; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2400 = _GEN_4628 & 2'h2 == _GEN_383 | _GEN_1984; // @[StoreSet.scala 546:{29,29}]
  wire  _GEN_2401 = _GEN_4628 & 2'h3 == _GEN_383 | _GEN_1985; // @[StoreSet.scala 546:{29,29}]
  wire [1:0] _GEN_2658 = io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore ? _GEN_2242 : _GEN_1826; // @[StoreSet.scala 542:70]
  wire [1:0] _GEN_2659 = io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore ? _GEN_2243 : _GEN_1827; // @[StoreSet.scala 542:70]
  wire [1:0] _GEN_2660 = io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore ? _GEN_2244 : _GEN_1828; // @[StoreSet.scala 542:70]
  wire [1:0] _GEN_2661 = io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore ? _GEN_2245 : _GEN_1829; // @[StoreSet.scala 542:70]
  wire [1:0] _GEN_2662 = io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore ? _GEN_2246 : _GEN_1830; // @[StoreSet.scala 542:70]
  wire [1:0] _GEN_2663 = io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore ? _GEN_2247 : _GEN_1831; // @[StoreSet.scala 542:70]
  wire [1:0] _GEN_2664 = io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore ? _GEN_2248 : _GEN_1832; // @[StoreSet.scala 542:70]
  wire [1:0] _GEN_2665 = io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore ? _GEN_2249 : _GEN_1833; // @[StoreSet.scala 542:70]
  wire [1:0] _GEN_2666 = io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore ? _GEN_2250 : _GEN_1834; // @[StoreSet.scala 542:70]
  wire [1:0] _GEN_2667 = io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore ? _GEN_2251 : _GEN_1835; // @[StoreSet.scala 542:70]
  wire [1:0] _GEN_2668 = io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore ? _GEN_2252 : _GEN_1836; // @[StoreSet.scala 542:70]
  wire [1:0] _GEN_2669 = io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore ? _GEN_2253 : _GEN_1837; // @[StoreSet.scala 542:70]
  wire [1:0] _GEN_2670 = io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore ? _GEN_2254 : _GEN_1838; // @[StoreSet.scala 542:70]
  wire [1:0] _GEN_2671 = io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore ? _GEN_2255 : _GEN_1839; // @[StoreSet.scala 542:70]
  wire [1:0] _GEN_2672 = io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore ? _GEN_2256 : _GEN_1840; // @[StoreSet.scala 542:70]
  wire [1:0] _GEN_2673 = io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore ? _GEN_2257 : _GEN_1841; // @[StoreSet.scala 542:70]
  wire [1:0] _GEN_2674 = io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore ? _GEN_2258 : _GEN_1842; // @[StoreSet.scala 542:70]
  wire [1:0] _GEN_2675 = io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore ? _GEN_2259 : _GEN_1843; // @[StoreSet.scala 542:70]
  wire [1:0] _GEN_2676 = io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore ? _GEN_2260 : _GEN_1844; // @[StoreSet.scala 542:70]
  wire [1:0] _GEN_2677 = io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore ? _GEN_2261 : _GEN_1845; // @[StoreSet.scala 542:70]
  wire [1:0] _GEN_2678 = io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore ? _GEN_2262 : _GEN_1846; // @[StoreSet.scala 542:70]
  wire [1:0] _GEN_2679 = io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore ? _GEN_2263 : _GEN_1847; // @[StoreSet.scala 542:70]
  wire [1:0] _GEN_2680 = io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore ? _GEN_2264 : _GEN_1848; // @[StoreSet.scala 542:70]
  wire [1:0] _GEN_2681 = io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore ? _GEN_2265 : _GEN_1849; // @[StoreSet.scala 542:70]
  wire [1:0] _GEN_2682 = io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore ? _GEN_2266 : _GEN_1850; // @[StoreSet.scala 542:70]
  wire [1:0] _GEN_2683 = io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore ? _GEN_2267 : _GEN_1851; // @[StoreSet.scala 542:70]
  wire [1:0] _GEN_2684 = io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore ? _GEN_2268 : _GEN_1852; // @[StoreSet.scala 542:70]
  wire [1:0] _GEN_2685 = io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore ? _GEN_2269 : _GEN_1853; // @[StoreSet.scala 542:70]
  wire [1:0] _GEN_2686 = io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore ? _GEN_2270 : _GEN_1854; // @[StoreSet.scala 542:70]
  wire [1:0] _GEN_2687 = io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore ? _GEN_2271 : _GEN_1855; // @[StoreSet.scala 542:70]
  wire [1:0] _GEN_2688 = io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore ? _GEN_2272 : _GEN_1856; // @[StoreSet.scala 542:70]
  wire [1:0] _GEN_2689 = io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore ? _GEN_2273 : _GEN_1857; // @[StoreSet.scala 542:70]
  wire [5:0] _flushItself_T_1 = {robIdxVec_0_0_flag,robIdxVec_0_0_value}; // @[CircularQueuePtr.scala 61:50]
  wire [5:0] _flushItself_T_2 = {io_redirect_bits_robIdx_flag,io_redirect_bits_robIdx_value}; // @[CircularQueuePtr.scala 61:70]
  wire  _flushItself_T_3 = _flushItself_T_1 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself = io_redirect_bits_level & _flushItself_T_3; // @[Rob.scala 122:51]
  wire  differentFlag = robIdxVec_0_0_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare = robIdxVec_0_0_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_26 = differentFlag ^ compare; // @[CircularQueuePtr.scala 88:19]
  wire  _T_28 = io_redirect_valid & (flushItself | _T_26); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_5 = {robIdxVec_0_1_flag,robIdxVec_0_1_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_7 = _flushItself_T_5 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_1 = io_redirect_bits_level & _flushItself_T_7; // @[Rob.scala 122:51]
  wire  differentFlag_1 = robIdxVec_0_1_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_1 = robIdxVec_0_1_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_30 = differentFlag_1 ^ compare_1; // @[CircularQueuePtr.scala 88:19]
  wire  _T_32 = io_redirect_valid & (flushItself_1 | _T_30); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_9 = {robIdxVec_0_2_flag,robIdxVec_0_2_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_11 = _flushItself_T_9 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_2 = io_redirect_bits_level & _flushItself_T_11; // @[Rob.scala 122:51]
  wire  differentFlag_2 = robIdxVec_0_2_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_2 = robIdxVec_0_2_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_34 = differentFlag_2 ^ compare_2; // @[CircularQueuePtr.scala 88:19]
  wire  _T_36 = io_redirect_valid & (flushItself_2 | _T_34); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_13 = {robIdxVec_0_3_flag,robIdxVec_0_3_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_15 = _flushItself_T_13 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_3 = io_redirect_bits_level & _flushItself_T_15; // @[Rob.scala 122:51]
  wire  differentFlag_3 = robIdxVec_0_3_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_3 = robIdxVec_0_3_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_38 = differentFlag_3 ^ compare_3; // @[CircularQueuePtr.scala 88:19]
  wire  _T_40 = io_redirect_valid & (flushItself_3 | _T_38); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_17 = {robIdxVec_1_0_flag,robIdxVec_1_0_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_19 = _flushItself_T_17 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_4 = io_redirect_bits_level & _flushItself_T_19; // @[Rob.scala 122:51]
  wire  differentFlag_4 = robIdxVec_1_0_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_4 = robIdxVec_1_0_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_42 = differentFlag_4 ^ compare_4; // @[CircularQueuePtr.scala 88:19]
  wire  _T_44 = io_redirect_valid & (flushItself_4 | _T_42); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_21 = {robIdxVec_1_1_flag,robIdxVec_1_1_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_23 = _flushItself_T_21 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_5 = io_redirect_bits_level & _flushItself_T_23; // @[Rob.scala 122:51]
  wire  differentFlag_5 = robIdxVec_1_1_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_5 = robIdxVec_1_1_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_46 = differentFlag_5 ^ compare_5; // @[CircularQueuePtr.scala 88:19]
  wire  _T_48 = io_redirect_valid & (flushItself_5 | _T_46); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_25 = {robIdxVec_1_2_flag,robIdxVec_1_2_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_27 = _flushItself_T_25 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_6 = io_redirect_bits_level & _flushItself_T_27; // @[Rob.scala 122:51]
  wire  differentFlag_6 = robIdxVec_1_2_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_6 = robIdxVec_1_2_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_50 = differentFlag_6 ^ compare_6; // @[CircularQueuePtr.scala 88:19]
  wire  _T_52 = io_redirect_valid & (flushItself_6 | _T_50); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_29 = {robIdxVec_1_3_flag,robIdxVec_1_3_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_31 = _flushItself_T_29 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_7 = io_redirect_bits_level & _flushItself_T_31; // @[Rob.scala 122:51]
  wire  differentFlag_7 = robIdxVec_1_3_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_7 = robIdxVec_1_3_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_54 = differentFlag_7 ^ compare_7; // @[CircularQueuePtr.scala 88:19]
  wire  _T_56 = io_redirect_valid & (flushItself_7 | _T_54); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_33 = {robIdxVec_2_0_flag,robIdxVec_2_0_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_35 = _flushItself_T_33 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_8 = io_redirect_bits_level & _flushItself_T_35; // @[Rob.scala 122:51]
  wire  differentFlag_8 = robIdxVec_2_0_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_8 = robIdxVec_2_0_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_58 = differentFlag_8 ^ compare_8; // @[CircularQueuePtr.scala 88:19]
  wire  _T_60 = io_redirect_valid & (flushItself_8 | _T_58); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_37 = {robIdxVec_2_1_flag,robIdxVec_2_1_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_39 = _flushItself_T_37 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_9 = io_redirect_bits_level & _flushItself_T_39; // @[Rob.scala 122:51]
  wire  differentFlag_9 = robIdxVec_2_1_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_9 = robIdxVec_2_1_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_62 = differentFlag_9 ^ compare_9; // @[CircularQueuePtr.scala 88:19]
  wire  _T_64 = io_redirect_valid & (flushItself_9 | _T_62); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_41 = {robIdxVec_2_2_flag,robIdxVec_2_2_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_43 = _flushItself_T_41 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_10 = io_redirect_bits_level & _flushItself_T_43; // @[Rob.scala 122:51]
  wire  differentFlag_10 = robIdxVec_2_2_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_10 = robIdxVec_2_2_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_66 = differentFlag_10 ^ compare_10; // @[CircularQueuePtr.scala 88:19]
  wire  _T_68 = io_redirect_valid & (flushItself_10 | _T_66); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_45 = {robIdxVec_2_3_flag,robIdxVec_2_3_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_47 = _flushItself_T_45 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_11 = io_redirect_bits_level & _flushItself_T_47; // @[Rob.scala 122:51]
  wire  differentFlag_11 = robIdxVec_2_3_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_11 = robIdxVec_2_3_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_70 = differentFlag_11 ^ compare_11; // @[CircularQueuePtr.scala 88:19]
  wire  _T_72 = io_redirect_valid & (flushItself_11 | _T_70); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_49 = {robIdxVec_3_0_flag,robIdxVec_3_0_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_51 = _flushItself_T_49 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_12 = io_redirect_bits_level & _flushItself_T_51; // @[Rob.scala 122:51]
  wire  differentFlag_12 = robIdxVec_3_0_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_12 = robIdxVec_3_0_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_74 = differentFlag_12 ^ compare_12; // @[CircularQueuePtr.scala 88:19]
  wire  _T_76 = io_redirect_valid & (flushItself_12 | _T_74); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_53 = {robIdxVec_3_1_flag,robIdxVec_3_1_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_55 = _flushItself_T_53 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_13 = io_redirect_bits_level & _flushItself_T_55; // @[Rob.scala 122:51]
  wire  differentFlag_13 = robIdxVec_3_1_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_13 = robIdxVec_3_1_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_78 = differentFlag_13 ^ compare_13; // @[CircularQueuePtr.scala 88:19]
  wire  _T_80 = io_redirect_valid & (flushItself_13 | _T_78); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_57 = {robIdxVec_3_2_flag,robIdxVec_3_2_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_59 = _flushItself_T_57 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_14 = io_redirect_bits_level & _flushItself_T_59; // @[Rob.scala 122:51]
  wire  differentFlag_14 = robIdxVec_3_2_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_14 = robIdxVec_3_2_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_82 = differentFlag_14 ^ compare_14; // @[CircularQueuePtr.scala 88:19]
  wire  _T_84 = io_redirect_valid & (flushItself_14 | _T_82); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_61 = {robIdxVec_3_3_flag,robIdxVec_3_3_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_63 = _flushItself_T_61 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_15 = io_redirect_bits_level & _flushItself_T_63; // @[Rob.scala 122:51]
  wire  differentFlag_15 = robIdxVec_3_3_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_15 = robIdxVec_3_3_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_86 = differentFlag_15 ^ compare_15; // @[CircularQueuePtr.scala 88:19]
  wire  _T_88 = io_redirect_valid & (flushItself_15 | _T_86); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_65 = {robIdxVec_4_0_flag,robIdxVec_4_0_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_67 = _flushItself_T_65 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_16 = io_redirect_bits_level & _flushItself_T_67; // @[Rob.scala 122:51]
  wire  differentFlag_16 = robIdxVec_4_0_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_16 = robIdxVec_4_0_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_90 = differentFlag_16 ^ compare_16; // @[CircularQueuePtr.scala 88:19]
  wire  _T_92 = io_redirect_valid & (flushItself_16 | _T_90); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_69 = {robIdxVec_4_1_flag,robIdxVec_4_1_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_71 = _flushItself_T_69 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_17 = io_redirect_bits_level & _flushItself_T_71; // @[Rob.scala 122:51]
  wire  differentFlag_17 = robIdxVec_4_1_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_17 = robIdxVec_4_1_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_94 = differentFlag_17 ^ compare_17; // @[CircularQueuePtr.scala 88:19]
  wire  _T_96 = io_redirect_valid & (flushItself_17 | _T_94); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_73 = {robIdxVec_4_2_flag,robIdxVec_4_2_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_75 = _flushItself_T_73 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_18 = io_redirect_bits_level & _flushItself_T_75; // @[Rob.scala 122:51]
  wire  differentFlag_18 = robIdxVec_4_2_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_18 = robIdxVec_4_2_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_98 = differentFlag_18 ^ compare_18; // @[CircularQueuePtr.scala 88:19]
  wire  _T_100 = io_redirect_valid & (flushItself_18 | _T_98); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_77 = {robIdxVec_4_3_flag,robIdxVec_4_3_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_79 = _flushItself_T_77 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_19 = io_redirect_bits_level & _flushItself_T_79; // @[Rob.scala 122:51]
  wire  differentFlag_19 = robIdxVec_4_3_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_19 = robIdxVec_4_3_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_102 = differentFlag_19 ^ compare_19; // @[CircularQueuePtr.scala 88:19]
  wire  _T_104 = io_redirect_valid & (flushItself_19 | _T_102); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_81 = {robIdxVec_5_0_flag,robIdxVec_5_0_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_83 = _flushItself_T_81 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_20 = io_redirect_bits_level & _flushItself_T_83; // @[Rob.scala 122:51]
  wire  differentFlag_20 = robIdxVec_5_0_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_20 = robIdxVec_5_0_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_106 = differentFlag_20 ^ compare_20; // @[CircularQueuePtr.scala 88:19]
  wire  _T_108 = io_redirect_valid & (flushItself_20 | _T_106); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_85 = {robIdxVec_5_1_flag,robIdxVec_5_1_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_87 = _flushItself_T_85 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_21 = io_redirect_bits_level & _flushItself_T_87; // @[Rob.scala 122:51]
  wire  differentFlag_21 = robIdxVec_5_1_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_21 = robIdxVec_5_1_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_110 = differentFlag_21 ^ compare_21; // @[CircularQueuePtr.scala 88:19]
  wire  _T_112 = io_redirect_valid & (flushItself_21 | _T_110); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_89 = {robIdxVec_5_2_flag,robIdxVec_5_2_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_91 = _flushItself_T_89 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_22 = io_redirect_bits_level & _flushItself_T_91; // @[Rob.scala 122:51]
  wire  differentFlag_22 = robIdxVec_5_2_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_22 = robIdxVec_5_2_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_114 = differentFlag_22 ^ compare_22; // @[CircularQueuePtr.scala 88:19]
  wire  _T_116 = io_redirect_valid & (flushItself_22 | _T_114); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_93 = {robIdxVec_5_3_flag,robIdxVec_5_3_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_95 = _flushItself_T_93 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_23 = io_redirect_bits_level & _flushItself_T_95; // @[Rob.scala 122:51]
  wire  differentFlag_23 = robIdxVec_5_3_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_23 = robIdxVec_5_3_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_118 = differentFlag_23 ^ compare_23; // @[CircularQueuePtr.scala 88:19]
  wire  _T_120 = io_redirect_valid & (flushItself_23 | _T_118); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_97 = {robIdxVec_6_0_flag,robIdxVec_6_0_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_99 = _flushItself_T_97 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_24 = io_redirect_bits_level & _flushItself_T_99; // @[Rob.scala 122:51]
  wire  differentFlag_24 = robIdxVec_6_0_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_24 = robIdxVec_6_0_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_122 = differentFlag_24 ^ compare_24; // @[CircularQueuePtr.scala 88:19]
  wire  _T_124 = io_redirect_valid & (flushItself_24 | _T_122); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_101 = {robIdxVec_6_1_flag,robIdxVec_6_1_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_103 = _flushItself_T_101 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_25 = io_redirect_bits_level & _flushItself_T_103; // @[Rob.scala 122:51]
  wire  differentFlag_25 = robIdxVec_6_1_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_25 = robIdxVec_6_1_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_126 = differentFlag_25 ^ compare_25; // @[CircularQueuePtr.scala 88:19]
  wire  _T_128 = io_redirect_valid & (flushItself_25 | _T_126); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_105 = {robIdxVec_6_2_flag,robIdxVec_6_2_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_107 = _flushItself_T_105 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_26 = io_redirect_bits_level & _flushItself_T_107; // @[Rob.scala 122:51]
  wire  differentFlag_26 = robIdxVec_6_2_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_26 = robIdxVec_6_2_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_130 = differentFlag_26 ^ compare_26; // @[CircularQueuePtr.scala 88:19]
  wire  _T_132 = io_redirect_valid & (flushItself_26 | _T_130); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_109 = {robIdxVec_6_3_flag,robIdxVec_6_3_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_111 = _flushItself_T_109 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_27 = io_redirect_bits_level & _flushItself_T_111; // @[Rob.scala 122:51]
  wire  differentFlag_27 = robIdxVec_6_3_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_27 = robIdxVec_6_3_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_134 = differentFlag_27 ^ compare_27; // @[CircularQueuePtr.scala 88:19]
  wire  _T_136 = io_redirect_valid & (flushItself_27 | _T_134); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_113 = {robIdxVec_7_0_flag,robIdxVec_7_0_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_115 = _flushItself_T_113 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_28 = io_redirect_bits_level & _flushItself_T_115; // @[Rob.scala 122:51]
  wire  differentFlag_28 = robIdxVec_7_0_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_28 = robIdxVec_7_0_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_138 = differentFlag_28 ^ compare_28; // @[CircularQueuePtr.scala 88:19]
  wire  _T_140 = io_redirect_valid & (flushItself_28 | _T_138); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_117 = {robIdxVec_7_1_flag,robIdxVec_7_1_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_119 = _flushItself_T_117 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_29 = io_redirect_bits_level & _flushItself_T_119; // @[Rob.scala 122:51]
  wire  differentFlag_29 = robIdxVec_7_1_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_29 = robIdxVec_7_1_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_142 = differentFlag_29 ^ compare_29; // @[CircularQueuePtr.scala 88:19]
  wire  _T_144 = io_redirect_valid & (flushItself_29 | _T_142); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_121 = {robIdxVec_7_2_flag,robIdxVec_7_2_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_123 = _flushItself_T_121 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_30 = io_redirect_bits_level & _flushItself_T_123; // @[Rob.scala 122:51]
  wire  differentFlag_30 = robIdxVec_7_2_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_30 = robIdxVec_7_2_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_146 = differentFlag_30 ^ compare_30; // @[CircularQueuePtr.scala 88:19]
  wire  _T_148 = io_redirect_valid & (flushItself_30 | _T_146); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_125 = {robIdxVec_7_3_flag,robIdxVec_7_3_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_127 = _flushItself_T_125 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_31 = io_redirect_bits_level & _flushItself_T_127; // @[Rob.scala 122:51]
  wire  differentFlag_31 = robIdxVec_7_3_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_31 = robIdxVec_7_3_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_150 = differentFlag_31 ^ compare_31; // @[CircularQueuePtr.scala 88:19]
  wire  _T_152 = io_redirect_valid & (flushItself_31 | _T_150); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_129 = {robIdxVec_8_0_flag,robIdxVec_8_0_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_131 = _flushItself_T_129 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_32 = io_redirect_bits_level & _flushItself_T_131; // @[Rob.scala 122:51]
  wire  differentFlag_32 = robIdxVec_8_0_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_32 = robIdxVec_8_0_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_154 = differentFlag_32 ^ compare_32; // @[CircularQueuePtr.scala 88:19]
  wire  _T_156 = io_redirect_valid & (flushItself_32 | _T_154); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_133 = {robIdxVec_8_1_flag,robIdxVec_8_1_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_135 = _flushItself_T_133 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_33 = io_redirect_bits_level & _flushItself_T_135; // @[Rob.scala 122:51]
  wire  differentFlag_33 = robIdxVec_8_1_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_33 = robIdxVec_8_1_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_158 = differentFlag_33 ^ compare_33; // @[CircularQueuePtr.scala 88:19]
  wire  _T_160 = io_redirect_valid & (flushItself_33 | _T_158); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_137 = {robIdxVec_8_2_flag,robIdxVec_8_2_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_139 = _flushItself_T_137 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_34 = io_redirect_bits_level & _flushItself_T_139; // @[Rob.scala 122:51]
  wire  differentFlag_34 = robIdxVec_8_2_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_34 = robIdxVec_8_2_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_162 = differentFlag_34 ^ compare_34; // @[CircularQueuePtr.scala 88:19]
  wire  _T_164 = io_redirect_valid & (flushItself_34 | _T_162); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_141 = {robIdxVec_8_3_flag,robIdxVec_8_3_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_143 = _flushItself_T_141 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_35 = io_redirect_bits_level & _flushItself_T_143; // @[Rob.scala 122:51]
  wire  differentFlag_35 = robIdxVec_8_3_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_35 = robIdxVec_8_3_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_166 = differentFlag_35 ^ compare_35; // @[CircularQueuePtr.scala 88:19]
  wire  _T_168 = io_redirect_valid & (flushItself_35 | _T_166); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_145 = {robIdxVec_9_0_flag,robIdxVec_9_0_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_147 = _flushItself_T_145 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_36 = io_redirect_bits_level & _flushItself_T_147; // @[Rob.scala 122:51]
  wire  differentFlag_36 = robIdxVec_9_0_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_36 = robIdxVec_9_0_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_170 = differentFlag_36 ^ compare_36; // @[CircularQueuePtr.scala 88:19]
  wire  _T_172 = io_redirect_valid & (flushItself_36 | _T_170); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_149 = {robIdxVec_9_1_flag,robIdxVec_9_1_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_151 = _flushItself_T_149 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_37 = io_redirect_bits_level & _flushItself_T_151; // @[Rob.scala 122:51]
  wire  differentFlag_37 = robIdxVec_9_1_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_37 = robIdxVec_9_1_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_174 = differentFlag_37 ^ compare_37; // @[CircularQueuePtr.scala 88:19]
  wire  _T_176 = io_redirect_valid & (flushItself_37 | _T_174); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_153 = {robIdxVec_9_2_flag,robIdxVec_9_2_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_155 = _flushItself_T_153 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_38 = io_redirect_bits_level & _flushItself_T_155; // @[Rob.scala 122:51]
  wire  differentFlag_38 = robIdxVec_9_2_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_38 = robIdxVec_9_2_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_178 = differentFlag_38 ^ compare_38; // @[CircularQueuePtr.scala 88:19]
  wire  _T_180 = io_redirect_valid & (flushItself_38 | _T_178); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_157 = {robIdxVec_9_3_flag,robIdxVec_9_3_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_159 = _flushItself_T_157 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_39 = io_redirect_bits_level & _flushItself_T_159; // @[Rob.scala 122:51]
  wire  differentFlag_39 = robIdxVec_9_3_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_39 = robIdxVec_9_3_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_182 = differentFlag_39 ^ compare_39; // @[CircularQueuePtr.scala 88:19]
  wire  _T_184 = io_redirect_valid & (flushItself_39 | _T_182); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_161 = {robIdxVec_10_0_flag,robIdxVec_10_0_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_163 = _flushItself_T_161 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_40 = io_redirect_bits_level & _flushItself_T_163; // @[Rob.scala 122:51]
  wire  differentFlag_40 = robIdxVec_10_0_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_40 = robIdxVec_10_0_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_186 = differentFlag_40 ^ compare_40; // @[CircularQueuePtr.scala 88:19]
  wire  _T_188 = io_redirect_valid & (flushItself_40 | _T_186); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_165 = {robIdxVec_10_1_flag,robIdxVec_10_1_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_167 = _flushItself_T_165 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_41 = io_redirect_bits_level & _flushItself_T_167; // @[Rob.scala 122:51]
  wire  differentFlag_41 = robIdxVec_10_1_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_41 = robIdxVec_10_1_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_190 = differentFlag_41 ^ compare_41; // @[CircularQueuePtr.scala 88:19]
  wire  _T_192 = io_redirect_valid & (flushItself_41 | _T_190); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_169 = {robIdxVec_10_2_flag,robIdxVec_10_2_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_171 = _flushItself_T_169 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_42 = io_redirect_bits_level & _flushItself_T_171; // @[Rob.scala 122:51]
  wire  differentFlag_42 = robIdxVec_10_2_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_42 = robIdxVec_10_2_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_194 = differentFlag_42 ^ compare_42; // @[CircularQueuePtr.scala 88:19]
  wire  _T_196 = io_redirect_valid & (flushItself_42 | _T_194); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_173 = {robIdxVec_10_3_flag,robIdxVec_10_3_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_175 = _flushItself_T_173 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_43 = io_redirect_bits_level & _flushItself_T_175; // @[Rob.scala 122:51]
  wire  differentFlag_43 = robIdxVec_10_3_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_43 = robIdxVec_10_3_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_198 = differentFlag_43 ^ compare_43; // @[CircularQueuePtr.scala 88:19]
  wire  _T_200 = io_redirect_valid & (flushItself_43 | _T_198); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_177 = {robIdxVec_11_0_flag,robIdxVec_11_0_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_179 = _flushItself_T_177 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_44 = io_redirect_bits_level & _flushItself_T_179; // @[Rob.scala 122:51]
  wire  differentFlag_44 = robIdxVec_11_0_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_44 = robIdxVec_11_0_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_202 = differentFlag_44 ^ compare_44; // @[CircularQueuePtr.scala 88:19]
  wire  _T_204 = io_redirect_valid & (flushItself_44 | _T_202); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_181 = {robIdxVec_11_1_flag,robIdxVec_11_1_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_183 = _flushItself_T_181 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_45 = io_redirect_bits_level & _flushItself_T_183; // @[Rob.scala 122:51]
  wire  differentFlag_45 = robIdxVec_11_1_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_45 = robIdxVec_11_1_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_206 = differentFlag_45 ^ compare_45; // @[CircularQueuePtr.scala 88:19]
  wire  _T_208 = io_redirect_valid & (flushItself_45 | _T_206); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_185 = {robIdxVec_11_2_flag,robIdxVec_11_2_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_187 = _flushItself_T_185 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_46 = io_redirect_bits_level & _flushItself_T_187; // @[Rob.scala 122:51]
  wire  differentFlag_46 = robIdxVec_11_2_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_46 = robIdxVec_11_2_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_210 = differentFlag_46 ^ compare_46; // @[CircularQueuePtr.scala 88:19]
  wire  _T_212 = io_redirect_valid & (flushItself_46 | _T_210); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_189 = {robIdxVec_11_3_flag,robIdxVec_11_3_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_191 = _flushItself_T_189 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_47 = io_redirect_bits_level & _flushItself_T_191; // @[Rob.scala 122:51]
  wire  differentFlag_47 = robIdxVec_11_3_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_47 = robIdxVec_11_3_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_214 = differentFlag_47 ^ compare_47; // @[CircularQueuePtr.scala 88:19]
  wire  _T_216 = io_redirect_valid & (flushItself_47 | _T_214); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_193 = {robIdxVec_12_0_flag,robIdxVec_12_0_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_195 = _flushItself_T_193 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_48 = io_redirect_bits_level & _flushItself_T_195; // @[Rob.scala 122:51]
  wire  differentFlag_48 = robIdxVec_12_0_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_48 = robIdxVec_12_0_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_218 = differentFlag_48 ^ compare_48; // @[CircularQueuePtr.scala 88:19]
  wire  _T_220 = io_redirect_valid & (flushItself_48 | _T_218); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_197 = {robIdxVec_12_1_flag,robIdxVec_12_1_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_199 = _flushItself_T_197 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_49 = io_redirect_bits_level & _flushItself_T_199; // @[Rob.scala 122:51]
  wire  differentFlag_49 = robIdxVec_12_1_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_49 = robIdxVec_12_1_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_222 = differentFlag_49 ^ compare_49; // @[CircularQueuePtr.scala 88:19]
  wire  _T_224 = io_redirect_valid & (flushItself_49 | _T_222); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_201 = {robIdxVec_12_2_flag,robIdxVec_12_2_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_203 = _flushItself_T_201 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_50 = io_redirect_bits_level & _flushItself_T_203; // @[Rob.scala 122:51]
  wire  differentFlag_50 = robIdxVec_12_2_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_50 = robIdxVec_12_2_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_226 = differentFlag_50 ^ compare_50; // @[CircularQueuePtr.scala 88:19]
  wire  _T_228 = io_redirect_valid & (flushItself_50 | _T_226); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_205 = {robIdxVec_12_3_flag,robIdxVec_12_3_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_207 = _flushItself_T_205 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_51 = io_redirect_bits_level & _flushItself_T_207; // @[Rob.scala 122:51]
  wire  differentFlag_51 = robIdxVec_12_3_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_51 = robIdxVec_12_3_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_230 = differentFlag_51 ^ compare_51; // @[CircularQueuePtr.scala 88:19]
  wire  _T_232 = io_redirect_valid & (flushItself_51 | _T_230); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_209 = {robIdxVec_13_0_flag,robIdxVec_13_0_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_211 = _flushItself_T_209 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_52 = io_redirect_bits_level & _flushItself_T_211; // @[Rob.scala 122:51]
  wire  differentFlag_52 = robIdxVec_13_0_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_52 = robIdxVec_13_0_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_234 = differentFlag_52 ^ compare_52; // @[CircularQueuePtr.scala 88:19]
  wire  _T_236 = io_redirect_valid & (flushItself_52 | _T_234); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_213 = {robIdxVec_13_1_flag,robIdxVec_13_1_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_215 = _flushItself_T_213 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_53 = io_redirect_bits_level & _flushItself_T_215; // @[Rob.scala 122:51]
  wire  differentFlag_53 = robIdxVec_13_1_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_53 = robIdxVec_13_1_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_238 = differentFlag_53 ^ compare_53; // @[CircularQueuePtr.scala 88:19]
  wire  _T_240 = io_redirect_valid & (flushItself_53 | _T_238); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_217 = {robIdxVec_13_2_flag,robIdxVec_13_2_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_219 = _flushItself_T_217 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_54 = io_redirect_bits_level & _flushItself_T_219; // @[Rob.scala 122:51]
  wire  differentFlag_54 = robIdxVec_13_2_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_54 = robIdxVec_13_2_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_242 = differentFlag_54 ^ compare_54; // @[CircularQueuePtr.scala 88:19]
  wire  _T_244 = io_redirect_valid & (flushItself_54 | _T_242); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_221 = {robIdxVec_13_3_flag,robIdxVec_13_3_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_223 = _flushItself_T_221 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_55 = io_redirect_bits_level & _flushItself_T_223; // @[Rob.scala 122:51]
  wire  differentFlag_55 = robIdxVec_13_3_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_55 = robIdxVec_13_3_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_246 = differentFlag_55 ^ compare_55; // @[CircularQueuePtr.scala 88:19]
  wire  _T_248 = io_redirect_valid & (flushItself_55 | _T_246); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_225 = {robIdxVec_14_0_flag,robIdxVec_14_0_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_227 = _flushItself_T_225 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_56 = io_redirect_bits_level & _flushItself_T_227; // @[Rob.scala 122:51]
  wire  differentFlag_56 = robIdxVec_14_0_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_56 = robIdxVec_14_0_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_250 = differentFlag_56 ^ compare_56; // @[CircularQueuePtr.scala 88:19]
  wire  _T_252 = io_redirect_valid & (flushItself_56 | _T_250); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_229 = {robIdxVec_14_1_flag,robIdxVec_14_1_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_231 = _flushItself_T_229 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_57 = io_redirect_bits_level & _flushItself_T_231; // @[Rob.scala 122:51]
  wire  differentFlag_57 = robIdxVec_14_1_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_57 = robIdxVec_14_1_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_254 = differentFlag_57 ^ compare_57; // @[CircularQueuePtr.scala 88:19]
  wire  _T_256 = io_redirect_valid & (flushItself_57 | _T_254); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_233 = {robIdxVec_14_2_flag,robIdxVec_14_2_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_235 = _flushItself_T_233 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_58 = io_redirect_bits_level & _flushItself_T_235; // @[Rob.scala 122:51]
  wire  differentFlag_58 = robIdxVec_14_2_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_58 = robIdxVec_14_2_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_258 = differentFlag_58 ^ compare_58; // @[CircularQueuePtr.scala 88:19]
  wire  _T_260 = io_redirect_valid & (flushItself_58 | _T_258); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_237 = {robIdxVec_14_3_flag,robIdxVec_14_3_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_239 = _flushItself_T_237 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_59 = io_redirect_bits_level & _flushItself_T_239; // @[Rob.scala 122:51]
  wire  differentFlag_59 = robIdxVec_14_3_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_59 = robIdxVec_14_3_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_262 = differentFlag_59 ^ compare_59; // @[CircularQueuePtr.scala 88:19]
  wire  _T_264 = io_redirect_valid & (flushItself_59 | _T_262); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_241 = {robIdxVec_15_0_flag,robIdxVec_15_0_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_243 = _flushItself_T_241 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_60 = io_redirect_bits_level & _flushItself_T_243; // @[Rob.scala 122:51]
  wire  differentFlag_60 = robIdxVec_15_0_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_60 = robIdxVec_15_0_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_266 = differentFlag_60 ^ compare_60; // @[CircularQueuePtr.scala 88:19]
  wire  _T_268 = io_redirect_valid & (flushItself_60 | _T_266); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_245 = {robIdxVec_15_1_flag,robIdxVec_15_1_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_247 = _flushItself_T_245 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_61 = io_redirect_bits_level & _flushItself_T_247; // @[Rob.scala 122:51]
  wire  differentFlag_61 = robIdxVec_15_1_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_61 = robIdxVec_15_1_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_270 = differentFlag_61 ^ compare_61; // @[CircularQueuePtr.scala 88:19]
  wire  _T_272 = io_redirect_valid & (flushItself_61 | _T_270); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_249 = {robIdxVec_15_2_flag,robIdxVec_15_2_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_251 = _flushItself_T_249 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_62 = io_redirect_bits_level & _flushItself_T_251; // @[Rob.scala 122:51]
  wire  differentFlag_62 = robIdxVec_15_2_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_62 = robIdxVec_15_2_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_274 = differentFlag_62 ^ compare_62; // @[CircularQueuePtr.scala 88:19]
  wire  _T_276 = io_redirect_valid & (flushItself_62 | _T_274); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_253 = {robIdxVec_15_3_flag,robIdxVec_15_3_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_255 = _flushItself_T_253 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_63 = io_redirect_bits_level & _flushItself_T_255; // @[Rob.scala 122:51]
  wire  differentFlag_63 = robIdxVec_15_3_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_63 = robIdxVec_15_3_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_278 = differentFlag_63 ^ compare_63; // @[CircularQueuePtr.scala 88:19]
  wire  _T_280 = io_redirect_valid & (flushItself_63 | _T_278); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_257 = {robIdxVec_16_0_flag,robIdxVec_16_0_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_259 = _flushItself_T_257 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_64 = io_redirect_bits_level & _flushItself_T_259; // @[Rob.scala 122:51]
  wire  differentFlag_64 = robIdxVec_16_0_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_64 = robIdxVec_16_0_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_282 = differentFlag_64 ^ compare_64; // @[CircularQueuePtr.scala 88:19]
  wire  _T_284 = io_redirect_valid & (flushItself_64 | _T_282); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_261 = {robIdxVec_16_1_flag,robIdxVec_16_1_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_263 = _flushItself_T_261 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_65 = io_redirect_bits_level & _flushItself_T_263; // @[Rob.scala 122:51]
  wire  differentFlag_65 = robIdxVec_16_1_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_65 = robIdxVec_16_1_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_286 = differentFlag_65 ^ compare_65; // @[CircularQueuePtr.scala 88:19]
  wire  _T_288 = io_redirect_valid & (flushItself_65 | _T_286); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_265 = {robIdxVec_16_2_flag,robIdxVec_16_2_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_267 = _flushItself_T_265 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_66 = io_redirect_bits_level & _flushItself_T_267; // @[Rob.scala 122:51]
  wire  differentFlag_66 = robIdxVec_16_2_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_66 = robIdxVec_16_2_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_290 = differentFlag_66 ^ compare_66; // @[CircularQueuePtr.scala 88:19]
  wire  _T_292 = io_redirect_valid & (flushItself_66 | _T_290); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_269 = {robIdxVec_16_3_flag,robIdxVec_16_3_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_271 = _flushItself_T_269 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_67 = io_redirect_bits_level & _flushItself_T_271; // @[Rob.scala 122:51]
  wire  differentFlag_67 = robIdxVec_16_3_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_67 = robIdxVec_16_3_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_294 = differentFlag_67 ^ compare_67; // @[CircularQueuePtr.scala 88:19]
  wire  _T_296 = io_redirect_valid & (flushItself_67 | _T_294); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_273 = {robIdxVec_17_0_flag,robIdxVec_17_0_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_275 = _flushItself_T_273 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_68 = io_redirect_bits_level & _flushItself_T_275; // @[Rob.scala 122:51]
  wire  differentFlag_68 = robIdxVec_17_0_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_68 = robIdxVec_17_0_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_298 = differentFlag_68 ^ compare_68; // @[CircularQueuePtr.scala 88:19]
  wire  _T_300 = io_redirect_valid & (flushItself_68 | _T_298); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_277 = {robIdxVec_17_1_flag,robIdxVec_17_1_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_279 = _flushItself_T_277 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_69 = io_redirect_bits_level & _flushItself_T_279; // @[Rob.scala 122:51]
  wire  differentFlag_69 = robIdxVec_17_1_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_69 = robIdxVec_17_1_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_302 = differentFlag_69 ^ compare_69; // @[CircularQueuePtr.scala 88:19]
  wire  _T_304 = io_redirect_valid & (flushItself_69 | _T_302); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_281 = {robIdxVec_17_2_flag,robIdxVec_17_2_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_283 = _flushItself_T_281 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_70 = io_redirect_bits_level & _flushItself_T_283; // @[Rob.scala 122:51]
  wire  differentFlag_70 = robIdxVec_17_2_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_70 = robIdxVec_17_2_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_306 = differentFlag_70 ^ compare_70; // @[CircularQueuePtr.scala 88:19]
  wire  _T_308 = io_redirect_valid & (flushItself_70 | _T_306); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_285 = {robIdxVec_17_3_flag,robIdxVec_17_3_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_287 = _flushItself_T_285 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_71 = io_redirect_bits_level & _flushItself_T_287; // @[Rob.scala 122:51]
  wire  differentFlag_71 = robIdxVec_17_3_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_71 = robIdxVec_17_3_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_310 = differentFlag_71 ^ compare_71; // @[CircularQueuePtr.scala 88:19]
  wire  _T_312 = io_redirect_valid & (flushItself_71 | _T_310); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_289 = {robIdxVec_18_0_flag,robIdxVec_18_0_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_291 = _flushItself_T_289 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_72 = io_redirect_bits_level & _flushItself_T_291; // @[Rob.scala 122:51]
  wire  differentFlag_72 = robIdxVec_18_0_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_72 = robIdxVec_18_0_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_314 = differentFlag_72 ^ compare_72; // @[CircularQueuePtr.scala 88:19]
  wire  _T_316 = io_redirect_valid & (flushItself_72 | _T_314); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_293 = {robIdxVec_18_1_flag,robIdxVec_18_1_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_295 = _flushItself_T_293 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_73 = io_redirect_bits_level & _flushItself_T_295; // @[Rob.scala 122:51]
  wire  differentFlag_73 = robIdxVec_18_1_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_73 = robIdxVec_18_1_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_318 = differentFlag_73 ^ compare_73; // @[CircularQueuePtr.scala 88:19]
  wire  _T_320 = io_redirect_valid & (flushItself_73 | _T_318); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_297 = {robIdxVec_18_2_flag,robIdxVec_18_2_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_299 = _flushItself_T_297 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_74 = io_redirect_bits_level & _flushItself_T_299; // @[Rob.scala 122:51]
  wire  differentFlag_74 = robIdxVec_18_2_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_74 = robIdxVec_18_2_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_322 = differentFlag_74 ^ compare_74; // @[CircularQueuePtr.scala 88:19]
  wire  _T_324 = io_redirect_valid & (flushItself_74 | _T_322); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_301 = {robIdxVec_18_3_flag,robIdxVec_18_3_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_303 = _flushItself_T_301 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_75 = io_redirect_bits_level & _flushItself_T_303; // @[Rob.scala 122:51]
  wire  differentFlag_75 = robIdxVec_18_3_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_75 = robIdxVec_18_3_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_326 = differentFlag_75 ^ compare_75; // @[CircularQueuePtr.scala 88:19]
  wire  _T_328 = io_redirect_valid & (flushItself_75 | _T_326); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_305 = {robIdxVec_19_0_flag,robIdxVec_19_0_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_307 = _flushItself_T_305 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_76 = io_redirect_bits_level & _flushItself_T_307; // @[Rob.scala 122:51]
  wire  differentFlag_76 = robIdxVec_19_0_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_76 = robIdxVec_19_0_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_330 = differentFlag_76 ^ compare_76; // @[CircularQueuePtr.scala 88:19]
  wire  _T_332 = io_redirect_valid & (flushItself_76 | _T_330); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_309 = {robIdxVec_19_1_flag,robIdxVec_19_1_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_311 = _flushItself_T_309 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_77 = io_redirect_bits_level & _flushItself_T_311; // @[Rob.scala 122:51]
  wire  differentFlag_77 = robIdxVec_19_1_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_77 = robIdxVec_19_1_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_334 = differentFlag_77 ^ compare_77; // @[CircularQueuePtr.scala 88:19]
  wire  _T_336 = io_redirect_valid & (flushItself_77 | _T_334); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_313 = {robIdxVec_19_2_flag,robIdxVec_19_2_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_315 = _flushItself_T_313 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_78 = io_redirect_bits_level & _flushItself_T_315; // @[Rob.scala 122:51]
  wire  differentFlag_78 = robIdxVec_19_2_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_78 = robIdxVec_19_2_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_338 = differentFlag_78 ^ compare_78; // @[CircularQueuePtr.scala 88:19]
  wire  _T_340 = io_redirect_valid & (flushItself_78 | _T_338); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_317 = {robIdxVec_19_3_flag,robIdxVec_19_3_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_319 = _flushItself_T_317 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_79 = io_redirect_bits_level & _flushItself_T_319; // @[Rob.scala 122:51]
  wire  differentFlag_79 = robIdxVec_19_3_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_79 = robIdxVec_19_3_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_342 = differentFlag_79 ^ compare_79; // @[CircularQueuePtr.scala 88:19]
  wire  _T_344 = io_redirect_valid & (flushItself_79 | _T_342); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_321 = {robIdxVec_20_0_flag,robIdxVec_20_0_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_323 = _flushItself_T_321 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_80 = io_redirect_bits_level & _flushItself_T_323; // @[Rob.scala 122:51]
  wire  differentFlag_80 = robIdxVec_20_0_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_80 = robIdxVec_20_0_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_346 = differentFlag_80 ^ compare_80; // @[CircularQueuePtr.scala 88:19]
  wire  _T_348 = io_redirect_valid & (flushItself_80 | _T_346); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_325 = {robIdxVec_20_1_flag,robIdxVec_20_1_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_327 = _flushItself_T_325 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_81 = io_redirect_bits_level & _flushItself_T_327; // @[Rob.scala 122:51]
  wire  differentFlag_81 = robIdxVec_20_1_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_81 = robIdxVec_20_1_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_350 = differentFlag_81 ^ compare_81; // @[CircularQueuePtr.scala 88:19]
  wire  _T_352 = io_redirect_valid & (flushItself_81 | _T_350); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_329 = {robIdxVec_20_2_flag,robIdxVec_20_2_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_331 = _flushItself_T_329 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_82 = io_redirect_bits_level & _flushItself_T_331; // @[Rob.scala 122:51]
  wire  differentFlag_82 = robIdxVec_20_2_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_82 = robIdxVec_20_2_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_354 = differentFlag_82 ^ compare_82; // @[CircularQueuePtr.scala 88:19]
  wire  _T_356 = io_redirect_valid & (flushItself_82 | _T_354); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_333 = {robIdxVec_20_3_flag,robIdxVec_20_3_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_335 = _flushItself_T_333 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_83 = io_redirect_bits_level & _flushItself_T_335; // @[Rob.scala 122:51]
  wire  differentFlag_83 = robIdxVec_20_3_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_83 = robIdxVec_20_3_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_358 = differentFlag_83 ^ compare_83; // @[CircularQueuePtr.scala 88:19]
  wire  _T_360 = io_redirect_valid & (flushItself_83 | _T_358); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_337 = {robIdxVec_21_0_flag,robIdxVec_21_0_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_339 = _flushItself_T_337 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_84 = io_redirect_bits_level & _flushItself_T_339; // @[Rob.scala 122:51]
  wire  differentFlag_84 = robIdxVec_21_0_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_84 = robIdxVec_21_0_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_362 = differentFlag_84 ^ compare_84; // @[CircularQueuePtr.scala 88:19]
  wire  _T_364 = io_redirect_valid & (flushItself_84 | _T_362); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_341 = {robIdxVec_21_1_flag,robIdxVec_21_1_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_343 = _flushItself_T_341 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_85 = io_redirect_bits_level & _flushItself_T_343; // @[Rob.scala 122:51]
  wire  differentFlag_85 = robIdxVec_21_1_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_85 = robIdxVec_21_1_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_366 = differentFlag_85 ^ compare_85; // @[CircularQueuePtr.scala 88:19]
  wire  _T_368 = io_redirect_valid & (flushItself_85 | _T_366); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_345 = {robIdxVec_21_2_flag,robIdxVec_21_2_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_347 = _flushItself_T_345 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_86 = io_redirect_bits_level & _flushItself_T_347; // @[Rob.scala 122:51]
  wire  differentFlag_86 = robIdxVec_21_2_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_86 = robIdxVec_21_2_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_370 = differentFlag_86 ^ compare_86; // @[CircularQueuePtr.scala 88:19]
  wire  _T_372 = io_redirect_valid & (flushItself_86 | _T_370); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_349 = {robIdxVec_21_3_flag,robIdxVec_21_3_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_351 = _flushItself_T_349 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_87 = io_redirect_bits_level & _flushItself_T_351; // @[Rob.scala 122:51]
  wire  differentFlag_87 = robIdxVec_21_3_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_87 = robIdxVec_21_3_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_374 = differentFlag_87 ^ compare_87; // @[CircularQueuePtr.scala 88:19]
  wire  _T_376 = io_redirect_valid & (flushItself_87 | _T_374); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_353 = {robIdxVec_22_0_flag,robIdxVec_22_0_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_355 = _flushItself_T_353 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_88 = io_redirect_bits_level & _flushItself_T_355; // @[Rob.scala 122:51]
  wire  differentFlag_88 = robIdxVec_22_0_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_88 = robIdxVec_22_0_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_378 = differentFlag_88 ^ compare_88; // @[CircularQueuePtr.scala 88:19]
  wire  _T_380 = io_redirect_valid & (flushItself_88 | _T_378); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_357 = {robIdxVec_22_1_flag,robIdxVec_22_1_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_359 = _flushItself_T_357 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_89 = io_redirect_bits_level & _flushItself_T_359; // @[Rob.scala 122:51]
  wire  differentFlag_89 = robIdxVec_22_1_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_89 = robIdxVec_22_1_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_382 = differentFlag_89 ^ compare_89; // @[CircularQueuePtr.scala 88:19]
  wire  _T_384 = io_redirect_valid & (flushItself_89 | _T_382); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_361 = {robIdxVec_22_2_flag,robIdxVec_22_2_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_363 = _flushItself_T_361 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_90 = io_redirect_bits_level & _flushItself_T_363; // @[Rob.scala 122:51]
  wire  differentFlag_90 = robIdxVec_22_2_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_90 = robIdxVec_22_2_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_386 = differentFlag_90 ^ compare_90; // @[CircularQueuePtr.scala 88:19]
  wire  _T_388 = io_redirect_valid & (flushItself_90 | _T_386); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_365 = {robIdxVec_22_3_flag,robIdxVec_22_3_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_367 = _flushItself_T_365 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_91 = io_redirect_bits_level & _flushItself_T_367; // @[Rob.scala 122:51]
  wire  differentFlag_91 = robIdxVec_22_3_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_91 = robIdxVec_22_3_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_390 = differentFlag_91 ^ compare_91; // @[CircularQueuePtr.scala 88:19]
  wire  _T_392 = io_redirect_valid & (flushItself_91 | _T_390); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_369 = {robIdxVec_23_0_flag,robIdxVec_23_0_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_371 = _flushItself_T_369 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_92 = io_redirect_bits_level & _flushItself_T_371; // @[Rob.scala 122:51]
  wire  differentFlag_92 = robIdxVec_23_0_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_92 = robIdxVec_23_0_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_394 = differentFlag_92 ^ compare_92; // @[CircularQueuePtr.scala 88:19]
  wire  _T_396 = io_redirect_valid & (flushItself_92 | _T_394); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_373 = {robIdxVec_23_1_flag,robIdxVec_23_1_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_375 = _flushItself_T_373 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_93 = io_redirect_bits_level & _flushItself_T_375; // @[Rob.scala 122:51]
  wire  differentFlag_93 = robIdxVec_23_1_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_93 = robIdxVec_23_1_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_398 = differentFlag_93 ^ compare_93; // @[CircularQueuePtr.scala 88:19]
  wire  _T_400 = io_redirect_valid & (flushItself_93 | _T_398); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_377 = {robIdxVec_23_2_flag,robIdxVec_23_2_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_379 = _flushItself_T_377 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_94 = io_redirect_bits_level & _flushItself_T_379; // @[Rob.scala 122:51]
  wire  differentFlag_94 = robIdxVec_23_2_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_94 = robIdxVec_23_2_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_402 = differentFlag_94 ^ compare_94; // @[CircularQueuePtr.scala 88:19]
  wire  _T_404 = io_redirect_valid & (flushItself_94 | _T_402); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_381 = {robIdxVec_23_3_flag,robIdxVec_23_3_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_383 = _flushItself_T_381 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_95 = io_redirect_bits_level & _flushItself_T_383; // @[Rob.scala 122:51]
  wire  differentFlag_95 = robIdxVec_23_3_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_95 = robIdxVec_23_3_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_406 = differentFlag_95 ^ compare_95; // @[CircularQueuePtr.scala 88:19]
  wire  _T_408 = io_redirect_valid & (flushItself_95 | _T_406); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_385 = {robIdxVec_24_0_flag,robIdxVec_24_0_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_387 = _flushItself_T_385 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_96 = io_redirect_bits_level & _flushItself_T_387; // @[Rob.scala 122:51]
  wire  differentFlag_96 = robIdxVec_24_0_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_96 = robIdxVec_24_0_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_410 = differentFlag_96 ^ compare_96; // @[CircularQueuePtr.scala 88:19]
  wire  _T_412 = io_redirect_valid & (flushItself_96 | _T_410); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_389 = {robIdxVec_24_1_flag,robIdxVec_24_1_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_391 = _flushItself_T_389 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_97 = io_redirect_bits_level & _flushItself_T_391; // @[Rob.scala 122:51]
  wire  differentFlag_97 = robIdxVec_24_1_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_97 = robIdxVec_24_1_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_414 = differentFlag_97 ^ compare_97; // @[CircularQueuePtr.scala 88:19]
  wire  _T_416 = io_redirect_valid & (flushItself_97 | _T_414); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_393 = {robIdxVec_24_2_flag,robIdxVec_24_2_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_395 = _flushItself_T_393 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_98 = io_redirect_bits_level & _flushItself_T_395; // @[Rob.scala 122:51]
  wire  differentFlag_98 = robIdxVec_24_2_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_98 = robIdxVec_24_2_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_418 = differentFlag_98 ^ compare_98; // @[CircularQueuePtr.scala 88:19]
  wire  _T_420 = io_redirect_valid & (flushItself_98 | _T_418); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_397 = {robIdxVec_24_3_flag,robIdxVec_24_3_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_399 = _flushItself_T_397 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_99 = io_redirect_bits_level & _flushItself_T_399; // @[Rob.scala 122:51]
  wire  differentFlag_99 = robIdxVec_24_3_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_99 = robIdxVec_24_3_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_422 = differentFlag_99 ^ compare_99; // @[CircularQueuePtr.scala 88:19]
  wire  _T_424 = io_redirect_valid & (flushItself_99 | _T_422); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_401 = {robIdxVec_25_0_flag,robIdxVec_25_0_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_403 = _flushItself_T_401 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_100 = io_redirect_bits_level & _flushItself_T_403; // @[Rob.scala 122:51]
  wire  differentFlag_100 = robIdxVec_25_0_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_100 = robIdxVec_25_0_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_426 = differentFlag_100 ^ compare_100; // @[CircularQueuePtr.scala 88:19]
  wire  _T_428 = io_redirect_valid & (flushItself_100 | _T_426); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_405 = {robIdxVec_25_1_flag,robIdxVec_25_1_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_407 = _flushItself_T_405 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_101 = io_redirect_bits_level & _flushItself_T_407; // @[Rob.scala 122:51]
  wire  differentFlag_101 = robIdxVec_25_1_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_101 = robIdxVec_25_1_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_430 = differentFlag_101 ^ compare_101; // @[CircularQueuePtr.scala 88:19]
  wire  _T_432 = io_redirect_valid & (flushItself_101 | _T_430); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_409 = {robIdxVec_25_2_flag,robIdxVec_25_2_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_411 = _flushItself_T_409 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_102 = io_redirect_bits_level & _flushItself_T_411; // @[Rob.scala 122:51]
  wire  differentFlag_102 = robIdxVec_25_2_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_102 = robIdxVec_25_2_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_434 = differentFlag_102 ^ compare_102; // @[CircularQueuePtr.scala 88:19]
  wire  _T_436 = io_redirect_valid & (flushItself_102 | _T_434); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_413 = {robIdxVec_25_3_flag,robIdxVec_25_3_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_415 = _flushItself_T_413 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_103 = io_redirect_bits_level & _flushItself_T_415; // @[Rob.scala 122:51]
  wire  differentFlag_103 = robIdxVec_25_3_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_103 = robIdxVec_25_3_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_438 = differentFlag_103 ^ compare_103; // @[CircularQueuePtr.scala 88:19]
  wire  _T_440 = io_redirect_valid & (flushItself_103 | _T_438); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_417 = {robIdxVec_26_0_flag,robIdxVec_26_0_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_419 = _flushItself_T_417 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_104 = io_redirect_bits_level & _flushItself_T_419; // @[Rob.scala 122:51]
  wire  differentFlag_104 = robIdxVec_26_0_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_104 = robIdxVec_26_0_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_442 = differentFlag_104 ^ compare_104; // @[CircularQueuePtr.scala 88:19]
  wire  _T_444 = io_redirect_valid & (flushItself_104 | _T_442); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_421 = {robIdxVec_26_1_flag,robIdxVec_26_1_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_423 = _flushItself_T_421 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_105 = io_redirect_bits_level & _flushItself_T_423; // @[Rob.scala 122:51]
  wire  differentFlag_105 = robIdxVec_26_1_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_105 = robIdxVec_26_1_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_446 = differentFlag_105 ^ compare_105; // @[CircularQueuePtr.scala 88:19]
  wire  _T_448 = io_redirect_valid & (flushItself_105 | _T_446); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_425 = {robIdxVec_26_2_flag,robIdxVec_26_2_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_427 = _flushItself_T_425 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_106 = io_redirect_bits_level & _flushItself_T_427; // @[Rob.scala 122:51]
  wire  differentFlag_106 = robIdxVec_26_2_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_106 = robIdxVec_26_2_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_450 = differentFlag_106 ^ compare_106; // @[CircularQueuePtr.scala 88:19]
  wire  _T_452 = io_redirect_valid & (flushItself_106 | _T_450); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_429 = {robIdxVec_26_3_flag,robIdxVec_26_3_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_431 = _flushItself_T_429 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_107 = io_redirect_bits_level & _flushItself_T_431; // @[Rob.scala 122:51]
  wire  differentFlag_107 = robIdxVec_26_3_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_107 = robIdxVec_26_3_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_454 = differentFlag_107 ^ compare_107; // @[CircularQueuePtr.scala 88:19]
  wire  _T_456 = io_redirect_valid & (flushItself_107 | _T_454); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_433 = {robIdxVec_27_0_flag,robIdxVec_27_0_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_435 = _flushItself_T_433 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_108 = io_redirect_bits_level & _flushItself_T_435; // @[Rob.scala 122:51]
  wire  differentFlag_108 = robIdxVec_27_0_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_108 = robIdxVec_27_0_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_458 = differentFlag_108 ^ compare_108; // @[CircularQueuePtr.scala 88:19]
  wire  _T_460 = io_redirect_valid & (flushItself_108 | _T_458); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_437 = {robIdxVec_27_1_flag,robIdxVec_27_1_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_439 = _flushItself_T_437 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_109 = io_redirect_bits_level & _flushItself_T_439; // @[Rob.scala 122:51]
  wire  differentFlag_109 = robIdxVec_27_1_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_109 = robIdxVec_27_1_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_462 = differentFlag_109 ^ compare_109; // @[CircularQueuePtr.scala 88:19]
  wire  _T_464 = io_redirect_valid & (flushItself_109 | _T_462); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_441 = {robIdxVec_27_2_flag,robIdxVec_27_2_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_443 = _flushItself_T_441 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_110 = io_redirect_bits_level & _flushItself_T_443; // @[Rob.scala 122:51]
  wire  differentFlag_110 = robIdxVec_27_2_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_110 = robIdxVec_27_2_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_466 = differentFlag_110 ^ compare_110; // @[CircularQueuePtr.scala 88:19]
  wire  _T_468 = io_redirect_valid & (flushItself_110 | _T_466); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_445 = {robIdxVec_27_3_flag,robIdxVec_27_3_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_447 = _flushItself_T_445 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_111 = io_redirect_bits_level & _flushItself_T_447; // @[Rob.scala 122:51]
  wire  differentFlag_111 = robIdxVec_27_3_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_111 = robIdxVec_27_3_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_470 = differentFlag_111 ^ compare_111; // @[CircularQueuePtr.scala 88:19]
  wire  _T_472 = io_redirect_valid & (flushItself_111 | _T_470); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_449 = {robIdxVec_28_0_flag,robIdxVec_28_0_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_451 = _flushItself_T_449 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_112 = io_redirect_bits_level & _flushItself_T_451; // @[Rob.scala 122:51]
  wire  differentFlag_112 = robIdxVec_28_0_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_112 = robIdxVec_28_0_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_474 = differentFlag_112 ^ compare_112; // @[CircularQueuePtr.scala 88:19]
  wire  _T_476 = io_redirect_valid & (flushItself_112 | _T_474); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_453 = {robIdxVec_28_1_flag,robIdxVec_28_1_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_455 = _flushItself_T_453 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_113 = io_redirect_bits_level & _flushItself_T_455; // @[Rob.scala 122:51]
  wire  differentFlag_113 = robIdxVec_28_1_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_113 = robIdxVec_28_1_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_478 = differentFlag_113 ^ compare_113; // @[CircularQueuePtr.scala 88:19]
  wire  _T_480 = io_redirect_valid & (flushItself_113 | _T_478); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_457 = {robIdxVec_28_2_flag,robIdxVec_28_2_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_459 = _flushItself_T_457 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_114 = io_redirect_bits_level & _flushItself_T_459; // @[Rob.scala 122:51]
  wire  differentFlag_114 = robIdxVec_28_2_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_114 = robIdxVec_28_2_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_482 = differentFlag_114 ^ compare_114; // @[CircularQueuePtr.scala 88:19]
  wire  _T_484 = io_redirect_valid & (flushItself_114 | _T_482); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_461 = {robIdxVec_28_3_flag,robIdxVec_28_3_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_463 = _flushItself_T_461 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_115 = io_redirect_bits_level & _flushItself_T_463; // @[Rob.scala 122:51]
  wire  differentFlag_115 = robIdxVec_28_3_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_115 = robIdxVec_28_3_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_486 = differentFlag_115 ^ compare_115; // @[CircularQueuePtr.scala 88:19]
  wire  _T_488 = io_redirect_valid & (flushItself_115 | _T_486); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_465 = {robIdxVec_29_0_flag,robIdxVec_29_0_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_467 = _flushItself_T_465 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_116 = io_redirect_bits_level & _flushItself_T_467; // @[Rob.scala 122:51]
  wire  differentFlag_116 = robIdxVec_29_0_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_116 = robIdxVec_29_0_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_490 = differentFlag_116 ^ compare_116; // @[CircularQueuePtr.scala 88:19]
  wire  _T_492 = io_redirect_valid & (flushItself_116 | _T_490); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_469 = {robIdxVec_29_1_flag,robIdxVec_29_1_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_471 = _flushItself_T_469 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_117 = io_redirect_bits_level & _flushItself_T_471; // @[Rob.scala 122:51]
  wire  differentFlag_117 = robIdxVec_29_1_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_117 = robIdxVec_29_1_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_494 = differentFlag_117 ^ compare_117; // @[CircularQueuePtr.scala 88:19]
  wire  _T_496 = io_redirect_valid & (flushItself_117 | _T_494); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_473 = {robIdxVec_29_2_flag,robIdxVec_29_2_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_475 = _flushItself_T_473 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_118 = io_redirect_bits_level & _flushItself_T_475; // @[Rob.scala 122:51]
  wire  differentFlag_118 = robIdxVec_29_2_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_118 = robIdxVec_29_2_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_498 = differentFlag_118 ^ compare_118; // @[CircularQueuePtr.scala 88:19]
  wire  _T_500 = io_redirect_valid & (flushItself_118 | _T_498); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_477 = {robIdxVec_29_3_flag,robIdxVec_29_3_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_479 = _flushItself_T_477 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_119 = io_redirect_bits_level & _flushItself_T_479; // @[Rob.scala 122:51]
  wire  differentFlag_119 = robIdxVec_29_3_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_119 = robIdxVec_29_3_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_502 = differentFlag_119 ^ compare_119; // @[CircularQueuePtr.scala 88:19]
  wire  _T_504 = io_redirect_valid & (flushItself_119 | _T_502); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_481 = {robIdxVec_30_0_flag,robIdxVec_30_0_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_483 = _flushItself_T_481 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_120 = io_redirect_bits_level & _flushItself_T_483; // @[Rob.scala 122:51]
  wire  differentFlag_120 = robIdxVec_30_0_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_120 = robIdxVec_30_0_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_506 = differentFlag_120 ^ compare_120; // @[CircularQueuePtr.scala 88:19]
  wire  _T_508 = io_redirect_valid & (flushItself_120 | _T_506); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_485 = {robIdxVec_30_1_flag,robIdxVec_30_1_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_487 = _flushItself_T_485 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_121 = io_redirect_bits_level & _flushItself_T_487; // @[Rob.scala 122:51]
  wire  differentFlag_121 = robIdxVec_30_1_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_121 = robIdxVec_30_1_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_510 = differentFlag_121 ^ compare_121; // @[CircularQueuePtr.scala 88:19]
  wire  _T_512 = io_redirect_valid & (flushItself_121 | _T_510); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_489 = {robIdxVec_30_2_flag,robIdxVec_30_2_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_491 = _flushItself_T_489 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_122 = io_redirect_bits_level & _flushItself_T_491; // @[Rob.scala 122:51]
  wire  differentFlag_122 = robIdxVec_30_2_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_122 = robIdxVec_30_2_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_514 = differentFlag_122 ^ compare_122; // @[CircularQueuePtr.scala 88:19]
  wire  _T_516 = io_redirect_valid & (flushItself_122 | _T_514); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_493 = {robIdxVec_30_3_flag,robIdxVec_30_3_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_495 = _flushItself_T_493 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_123 = io_redirect_bits_level & _flushItself_T_495; // @[Rob.scala 122:51]
  wire  differentFlag_123 = robIdxVec_30_3_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_123 = robIdxVec_30_3_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_518 = differentFlag_123 ^ compare_123; // @[CircularQueuePtr.scala 88:19]
  wire  _T_520 = io_redirect_valid & (flushItself_123 | _T_518); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_497 = {robIdxVec_31_0_flag,robIdxVec_31_0_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_499 = _flushItself_T_497 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_124 = io_redirect_bits_level & _flushItself_T_499; // @[Rob.scala 122:51]
  wire  differentFlag_124 = robIdxVec_31_0_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_124 = robIdxVec_31_0_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_522 = differentFlag_124 ^ compare_124; // @[CircularQueuePtr.scala 88:19]
  wire  _T_524 = io_redirect_valid & (flushItself_124 | _T_522); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_501 = {robIdxVec_31_1_flag,robIdxVec_31_1_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_503 = _flushItself_T_501 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_125 = io_redirect_bits_level & _flushItself_T_503; // @[Rob.scala 122:51]
  wire  differentFlag_125 = robIdxVec_31_1_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_125 = robIdxVec_31_1_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_526 = differentFlag_125 ^ compare_125; // @[CircularQueuePtr.scala 88:19]
  wire  _T_528 = io_redirect_valid & (flushItself_125 | _T_526); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_505 = {robIdxVec_31_2_flag,robIdxVec_31_2_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_507 = _flushItself_T_505 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_126 = io_redirect_bits_level & _flushItself_T_507; // @[Rob.scala 122:51]
  wire  differentFlag_126 = robIdxVec_31_2_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_126 = robIdxVec_31_2_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_530 = differentFlag_126 ^ compare_126; // @[CircularQueuePtr.scala 88:19]
  wire  _T_532 = io_redirect_valid & (flushItself_126 | _T_530); // @[Rob.scala 123:20]
  wire [5:0] _flushItself_T_509 = {robIdxVec_31_3_flag,robIdxVec_31_3_value}; // @[CircularQueuePtr.scala 61:50]
  wire  _flushItself_T_511 = _flushItself_T_509 == _flushItself_T_2; // @[CircularQueuePtr.scala 61:52]
  wire  flushItself_127 = io_redirect_bits_level & _flushItself_T_511; // @[Rob.scala 122:51]
  wire  differentFlag_127 = robIdxVec_31_3_flag ^ io_redirect_bits_robIdx_flag; // @[CircularQueuePtr.scala 86:35]
  wire  compare_127 = robIdxVec_31_3_value > io_redirect_bits_robIdx_value; // @[CircularQueuePtr.scala 87:30]
  wire  _T_534 = differentFlag_127 ^ compare_127; // @[CircularQueuePtr.scala 88:19]
  wire  _T_536 = io_redirect_valid & (flushItself_127 | _T_534); // @[Rob.scala 123:20]
  reg  REG; // @[StoreSet.scala 562:15]
  wire [1:0] check_position = allocPtr_0 + 2'h1; // @[StoreSet.scala 565:51]
  wire  _GEN_3203 = 2'h1 == check_position ? validVec_0_1 : validVec_0_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3204 = 2'h2 == check_position ? validVec_0_2 : _GEN_3203; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3205 = 2'h3 == check_position ? validVec_0_3 : _GEN_3204; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3206 = ~_GEN_3205 ? check_position : _GEN_2658; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_1 = allocPtr_0 + 2'h2; // @[StoreSet.scala 565:51]
  wire  _GEN_3208 = 2'h1 == check_position_1 ? validVec_0_1 : validVec_0_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3209 = 2'h2 == check_position_1 ? validVec_0_2 : _GEN_3208; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3210 = 2'h3 == check_position_1 ? validVec_0_3 : _GEN_3209; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3211 = ~_GEN_3210 ? check_position_1 : _GEN_3206; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_2 = allocPtr_0 + 2'h3; // @[StoreSet.scala 565:51]
  wire  _GEN_3213 = 2'h1 == check_position_2 ? validVec_0_1 : validVec_0_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3214 = 2'h2 == check_position_2 ? validVec_0_2 : _GEN_3213; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3215 = 2'h3 == check_position_2 ? validVec_0_3 : _GEN_3214; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3216 = ~_GEN_3215 ? check_position_2 : _GEN_3211; // @[StoreSet.scala 566:43 567:23]
  wire [2:0] _GEN_6682 = {{1'd0}, allocPtr_0}; // @[StoreSet.scala 565:51]
  wire [2:0] check_position_3 = _GEN_6682 + 3'h4; // @[StoreSet.scala 565:51]
  wire  _GEN_3218 = 2'h1 == check_position_3[1:0] ? validVec_0_1 : validVec_0_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3219 = 2'h2 == check_position_3[1:0] ? validVec_0_2 : _GEN_3218; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3220 = 2'h3 == check_position_3[1:0] ? validVec_0_3 : _GEN_3219; // @[StoreSet.scala 566:{14,14}]
  wire [2:0] _GEN_3221 = ~_GEN_3220 ? check_position_3 : {{1'd0}, _GEN_3216}; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_4 = allocPtr_1 + 2'h1; // @[StoreSet.scala 565:51]
  wire  _GEN_3223 = 2'h1 == check_position_4 ? validVec_1_1 : validVec_1_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3224 = 2'h2 == check_position_4 ? validVec_1_2 : _GEN_3223; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3225 = 2'h3 == check_position_4 ? validVec_1_3 : _GEN_3224; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3226 = ~_GEN_3225 ? check_position_4 : _GEN_2659; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_5 = allocPtr_1 + 2'h2; // @[StoreSet.scala 565:51]
  wire  _GEN_3228 = 2'h1 == check_position_5 ? validVec_1_1 : validVec_1_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3229 = 2'h2 == check_position_5 ? validVec_1_2 : _GEN_3228; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3230 = 2'h3 == check_position_5 ? validVec_1_3 : _GEN_3229; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3231 = ~_GEN_3230 ? check_position_5 : _GEN_3226; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_6 = allocPtr_1 + 2'h3; // @[StoreSet.scala 565:51]
  wire  _GEN_3233 = 2'h1 == check_position_6 ? validVec_1_1 : validVec_1_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3234 = 2'h2 == check_position_6 ? validVec_1_2 : _GEN_3233; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3235 = 2'h3 == check_position_6 ? validVec_1_3 : _GEN_3234; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3236 = ~_GEN_3235 ? check_position_6 : _GEN_3231; // @[StoreSet.scala 566:43 567:23]
  wire [2:0] _GEN_6683 = {{1'd0}, allocPtr_1}; // @[StoreSet.scala 565:51]
  wire [2:0] check_position_7 = _GEN_6683 + 3'h4; // @[StoreSet.scala 565:51]
  wire  _GEN_3238 = 2'h1 == check_position_7[1:0] ? validVec_1_1 : validVec_1_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3239 = 2'h2 == check_position_7[1:0] ? validVec_1_2 : _GEN_3238; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3240 = 2'h3 == check_position_7[1:0] ? validVec_1_3 : _GEN_3239; // @[StoreSet.scala 566:{14,14}]
  wire [2:0] _GEN_3241 = ~_GEN_3240 ? check_position_7 : {{1'd0}, _GEN_3236}; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_8 = allocPtr_2 + 2'h1; // @[StoreSet.scala 565:51]
  wire  _GEN_3243 = 2'h1 == check_position_8 ? validVec_2_1 : validVec_2_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3244 = 2'h2 == check_position_8 ? validVec_2_2 : _GEN_3243; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3245 = 2'h3 == check_position_8 ? validVec_2_3 : _GEN_3244; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3246 = ~_GEN_3245 ? check_position_8 : _GEN_2660; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_9 = allocPtr_2 + 2'h2; // @[StoreSet.scala 565:51]
  wire  _GEN_3248 = 2'h1 == check_position_9 ? validVec_2_1 : validVec_2_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3249 = 2'h2 == check_position_9 ? validVec_2_2 : _GEN_3248; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3250 = 2'h3 == check_position_9 ? validVec_2_3 : _GEN_3249; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3251 = ~_GEN_3250 ? check_position_9 : _GEN_3246; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_10 = allocPtr_2 + 2'h3; // @[StoreSet.scala 565:51]
  wire  _GEN_3253 = 2'h1 == check_position_10 ? validVec_2_1 : validVec_2_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3254 = 2'h2 == check_position_10 ? validVec_2_2 : _GEN_3253; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3255 = 2'h3 == check_position_10 ? validVec_2_3 : _GEN_3254; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3256 = ~_GEN_3255 ? check_position_10 : _GEN_3251; // @[StoreSet.scala 566:43 567:23]
  wire [2:0] _GEN_6684 = {{1'd0}, allocPtr_2}; // @[StoreSet.scala 565:51]
  wire [2:0] check_position_11 = _GEN_6684 + 3'h4; // @[StoreSet.scala 565:51]
  wire  _GEN_3258 = 2'h1 == check_position_11[1:0] ? validVec_2_1 : validVec_2_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3259 = 2'h2 == check_position_11[1:0] ? validVec_2_2 : _GEN_3258; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3260 = 2'h3 == check_position_11[1:0] ? validVec_2_3 : _GEN_3259; // @[StoreSet.scala 566:{14,14}]
  wire [2:0] _GEN_3261 = ~_GEN_3260 ? check_position_11 : {{1'd0}, _GEN_3256}; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_12 = allocPtr_3 + 2'h1; // @[StoreSet.scala 565:51]
  wire  _GEN_3263 = 2'h1 == check_position_12 ? validVec_3_1 : validVec_3_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3264 = 2'h2 == check_position_12 ? validVec_3_2 : _GEN_3263; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3265 = 2'h3 == check_position_12 ? validVec_3_3 : _GEN_3264; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3266 = ~_GEN_3265 ? check_position_12 : _GEN_2661; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_13 = allocPtr_3 + 2'h2; // @[StoreSet.scala 565:51]
  wire  _GEN_3268 = 2'h1 == check_position_13 ? validVec_3_1 : validVec_3_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3269 = 2'h2 == check_position_13 ? validVec_3_2 : _GEN_3268; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3270 = 2'h3 == check_position_13 ? validVec_3_3 : _GEN_3269; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3271 = ~_GEN_3270 ? check_position_13 : _GEN_3266; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_14 = allocPtr_3 + 2'h3; // @[StoreSet.scala 565:51]
  wire  _GEN_3273 = 2'h1 == check_position_14 ? validVec_3_1 : validVec_3_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3274 = 2'h2 == check_position_14 ? validVec_3_2 : _GEN_3273; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3275 = 2'h3 == check_position_14 ? validVec_3_3 : _GEN_3274; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3276 = ~_GEN_3275 ? check_position_14 : _GEN_3271; // @[StoreSet.scala 566:43 567:23]
  wire [2:0] _GEN_6685 = {{1'd0}, allocPtr_3}; // @[StoreSet.scala 565:51]
  wire [2:0] check_position_15 = _GEN_6685 + 3'h4; // @[StoreSet.scala 565:51]
  wire  _GEN_3278 = 2'h1 == check_position_15[1:0] ? validVec_3_1 : validVec_3_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3279 = 2'h2 == check_position_15[1:0] ? validVec_3_2 : _GEN_3278; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3280 = 2'h3 == check_position_15[1:0] ? validVec_3_3 : _GEN_3279; // @[StoreSet.scala 566:{14,14}]
  wire [2:0] _GEN_3281 = ~_GEN_3280 ? check_position_15 : {{1'd0}, _GEN_3276}; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_16 = allocPtr_4 + 2'h1; // @[StoreSet.scala 565:51]
  wire  _GEN_3283 = 2'h1 == check_position_16 ? validVec_4_1 : validVec_4_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3284 = 2'h2 == check_position_16 ? validVec_4_2 : _GEN_3283; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3285 = 2'h3 == check_position_16 ? validVec_4_3 : _GEN_3284; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3286 = ~_GEN_3285 ? check_position_16 : _GEN_2662; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_17 = allocPtr_4 + 2'h2; // @[StoreSet.scala 565:51]
  wire  _GEN_3288 = 2'h1 == check_position_17 ? validVec_4_1 : validVec_4_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3289 = 2'h2 == check_position_17 ? validVec_4_2 : _GEN_3288; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3290 = 2'h3 == check_position_17 ? validVec_4_3 : _GEN_3289; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3291 = ~_GEN_3290 ? check_position_17 : _GEN_3286; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_18 = allocPtr_4 + 2'h3; // @[StoreSet.scala 565:51]
  wire  _GEN_3293 = 2'h1 == check_position_18 ? validVec_4_1 : validVec_4_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3294 = 2'h2 == check_position_18 ? validVec_4_2 : _GEN_3293; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3295 = 2'h3 == check_position_18 ? validVec_4_3 : _GEN_3294; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3296 = ~_GEN_3295 ? check_position_18 : _GEN_3291; // @[StoreSet.scala 566:43 567:23]
  wire [2:0] _GEN_6686 = {{1'd0}, allocPtr_4}; // @[StoreSet.scala 565:51]
  wire [2:0] check_position_19 = _GEN_6686 + 3'h4; // @[StoreSet.scala 565:51]
  wire  _GEN_3298 = 2'h1 == check_position_19[1:0] ? validVec_4_1 : validVec_4_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3299 = 2'h2 == check_position_19[1:0] ? validVec_4_2 : _GEN_3298; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3300 = 2'h3 == check_position_19[1:0] ? validVec_4_3 : _GEN_3299; // @[StoreSet.scala 566:{14,14}]
  wire [2:0] _GEN_3301 = ~_GEN_3300 ? check_position_19 : {{1'd0}, _GEN_3296}; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_20 = allocPtr_5 + 2'h1; // @[StoreSet.scala 565:51]
  wire  _GEN_3303 = 2'h1 == check_position_20 ? validVec_5_1 : validVec_5_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3304 = 2'h2 == check_position_20 ? validVec_5_2 : _GEN_3303; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3305 = 2'h3 == check_position_20 ? validVec_5_3 : _GEN_3304; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3306 = ~_GEN_3305 ? check_position_20 : _GEN_2663; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_21 = allocPtr_5 + 2'h2; // @[StoreSet.scala 565:51]
  wire  _GEN_3308 = 2'h1 == check_position_21 ? validVec_5_1 : validVec_5_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3309 = 2'h2 == check_position_21 ? validVec_5_2 : _GEN_3308; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3310 = 2'h3 == check_position_21 ? validVec_5_3 : _GEN_3309; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3311 = ~_GEN_3310 ? check_position_21 : _GEN_3306; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_22 = allocPtr_5 + 2'h3; // @[StoreSet.scala 565:51]
  wire  _GEN_3313 = 2'h1 == check_position_22 ? validVec_5_1 : validVec_5_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3314 = 2'h2 == check_position_22 ? validVec_5_2 : _GEN_3313; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3315 = 2'h3 == check_position_22 ? validVec_5_3 : _GEN_3314; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3316 = ~_GEN_3315 ? check_position_22 : _GEN_3311; // @[StoreSet.scala 566:43 567:23]
  wire [2:0] _GEN_6687 = {{1'd0}, allocPtr_5}; // @[StoreSet.scala 565:51]
  wire [2:0] check_position_23 = _GEN_6687 + 3'h4; // @[StoreSet.scala 565:51]
  wire  _GEN_3318 = 2'h1 == check_position_23[1:0] ? validVec_5_1 : validVec_5_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3319 = 2'h2 == check_position_23[1:0] ? validVec_5_2 : _GEN_3318; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3320 = 2'h3 == check_position_23[1:0] ? validVec_5_3 : _GEN_3319; // @[StoreSet.scala 566:{14,14}]
  wire [2:0] _GEN_3321 = ~_GEN_3320 ? check_position_23 : {{1'd0}, _GEN_3316}; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_24 = allocPtr_6 + 2'h1; // @[StoreSet.scala 565:51]
  wire  _GEN_3323 = 2'h1 == check_position_24 ? validVec_6_1 : validVec_6_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3324 = 2'h2 == check_position_24 ? validVec_6_2 : _GEN_3323; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3325 = 2'h3 == check_position_24 ? validVec_6_3 : _GEN_3324; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3326 = ~_GEN_3325 ? check_position_24 : _GEN_2664; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_25 = allocPtr_6 + 2'h2; // @[StoreSet.scala 565:51]
  wire  _GEN_3328 = 2'h1 == check_position_25 ? validVec_6_1 : validVec_6_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3329 = 2'h2 == check_position_25 ? validVec_6_2 : _GEN_3328; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3330 = 2'h3 == check_position_25 ? validVec_6_3 : _GEN_3329; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3331 = ~_GEN_3330 ? check_position_25 : _GEN_3326; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_26 = allocPtr_6 + 2'h3; // @[StoreSet.scala 565:51]
  wire  _GEN_3333 = 2'h1 == check_position_26 ? validVec_6_1 : validVec_6_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3334 = 2'h2 == check_position_26 ? validVec_6_2 : _GEN_3333; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3335 = 2'h3 == check_position_26 ? validVec_6_3 : _GEN_3334; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3336 = ~_GEN_3335 ? check_position_26 : _GEN_3331; // @[StoreSet.scala 566:43 567:23]
  wire [2:0] _GEN_6688 = {{1'd0}, allocPtr_6}; // @[StoreSet.scala 565:51]
  wire [2:0] check_position_27 = _GEN_6688 + 3'h4; // @[StoreSet.scala 565:51]
  wire  _GEN_3338 = 2'h1 == check_position_27[1:0] ? validVec_6_1 : validVec_6_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3339 = 2'h2 == check_position_27[1:0] ? validVec_6_2 : _GEN_3338; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3340 = 2'h3 == check_position_27[1:0] ? validVec_6_3 : _GEN_3339; // @[StoreSet.scala 566:{14,14}]
  wire [2:0] _GEN_3341 = ~_GEN_3340 ? check_position_27 : {{1'd0}, _GEN_3336}; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_28 = allocPtr_7 + 2'h1; // @[StoreSet.scala 565:51]
  wire  _GEN_3343 = 2'h1 == check_position_28 ? validVec_7_1 : validVec_7_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3344 = 2'h2 == check_position_28 ? validVec_7_2 : _GEN_3343; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3345 = 2'h3 == check_position_28 ? validVec_7_3 : _GEN_3344; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3346 = ~_GEN_3345 ? check_position_28 : _GEN_2665; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_29 = allocPtr_7 + 2'h2; // @[StoreSet.scala 565:51]
  wire  _GEN_3348 = 2'h1 == check_position_29 ? validVec_7_1 : validVec_7_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3349 = 2'h2 == check_position_29 ? validVec_7_2 : _GEN_3348; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3350 = 2'h3 == check_position_29 ? validVec_7_3 : _GEN_3349; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3351 = ~_GEN_3350 ? check_position_29 : _GEN_3346; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_30 = allocPtr_7 + 2'h3; // @[StoreSet.scala 565:51]
  wire  _GEN_3353 = 2'h1 == check_position_30 ? validVec_7_1 : validVec_7_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3354 = 2'h2 == check_position_30 ? validVec_7_2 : _GEN_3353; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3355 = 2'h3 == check_position_30 ? validVec_7_3 : _GEN_3354; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3356 = ~_GEN_3355 ? check_position_30 : _GEN_3351; // @[StoreSet.scala 566:43 567:23]
  wire [2:0] _GEN_6689 = {{1'd0}, allocPtr_7}; // @[StoreSet.scala 565:51]
  wire [2:0] check_position_31 = _GEN_6689 + 3'h4; // @[StoreSet.scala 565:51]
  wire  _GEN_3358 = 2'h1 == check_position_31[1:0] ? validVec_7_1 : validVec_7_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3359 = 2'h2 == check_position_31[1:0] ? validVec_7_2 : _GEN_3358; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3360 = 2'h3 == check_position_31[1:0] ? validVec_7_3 : _GEN_3359; // @[StoreSet.scala 566:{14,14}]
  wire [2:0] _GEN_3361 = ~_GEN_3360 ? check_position_31 : {{1'd0}, _GEN_3356}; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_32 = allocPtr_8 + 2'h1; // @[StoreSet.scala 565:51]
  wire  _GEN_3363 = 2'h1 == check_position_32 ? validVec_8_1 : validVec_8_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3364 = 2'h2 == check_position_32 ? validVec_8_2 : _GEN_3363; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3365 = 2'h3 == check_position_32 ? validVec_8_3 : _GEN_3364; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3366 = ~_GEN_3365 ? check_position_32 : _GEN_2666; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_33 = allocPtr_8 + 2'h2; // @[StoreSet.scala 565:51]
  wire  _GEN_3368 = 2'h1 == check_position_33 ? validVec_8_1 : validVec_8_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3369 = 2'h2 == check_position_33 ? validVec_8_2 : _GEN_3368; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3370 = 2'h3 == check_position_33 ? validVec_8_3 : _GEN_3369; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3371 = ~_GEN_3370 ? check_position_33 : _GEN_3366; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_34 = allocPtr_8 + 2'h3; // @[StoreSet.scala 565:51]
  wire  _GEN_3373 = 2'h1 == check_position_34 ? validVec_8_1 : validVec_8_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3374 = 2'h2 == check_position_34 ? validVec_8_2 : _GEN_3373; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3375 = 2'h3 == check_position_34 ? validVec_8_3 : _GEN_3374; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3376 = ~_GEN_3375 ? check_position_34 : _GEN_3371; // @[StoreSet.scala 566:43 567:23]
  wire [2:0] _GEN_6690 = {{1'd0}, allocPtr_8}; // @[StoreSet.scala 565:51]
  wire [2:0] check_position_35 = _GEN_6690 + 3'h4; // @[StoreSet.scala 565:51]
  wire  _GEN_3378 = 2'h1 == check_position_35[1:0] ? validVec_8_1 : validVec_8_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3379 = 2'h2 == check_position_35[1:0] ? validVec_8_2 : _GEN_3378; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3380 = 2'h3 == check_position_35[1:0] ? validVec_8_3 : _GEN_3379; // @[StoreSet.scala 566:{14,14}]
  wire [2:0] _GEN_3381 = ~_GEN_3380 ? check_position_35 : {{1'd0}, _GEN_3376}; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_36 = allocPtr_9 + 2'h1; // @[StoreSet.scala 565:51]
  wire  _GEN_3383 = 2'h1 == check_position_36 ? validVec_9_1 : validVec_9_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3384 = 2'h2 == check_position_36 ? validVec_9_2 : _GEN_3383; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3385 = 2'h3 == check_position_36 ? validVec_9_3 : _GEN_3384; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3386 = ~_GEN_3385 ? check_position_36 : _GEN_2667; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_37 = allocPtr_9 + 2'h2; // @[StoreSet.scala 565:51]
  wire  _GEN_3388 = 2'h1 == check_position_37 ? validVec_9_1 : validVec_9_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3389 = 2'h2 == check_position_37 ? validVec_9_2 : _GEN_3388; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3390 = 2'h3 == check_position_37 ? validVec_9_3 : _GEN_3389; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3391 = ~_GEN_3390 ? check_position_37 : _GEN_3386; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_38 = allocPtr_9 + 2'h3; // @[StoreSet.scala 565:51]
  wire  _GEN_3393 = 2'h1 == check_position_38 ? validVec_9_1 : validVec_9_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3394 = 2'h2 == check_position_38 ? validVec_9_2 : _GEN_3393; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3395 = 2'h3 == check_position_38 ? validVec_9_3 : _GEN_3394; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3396 = ~_GEN_3395 ? check_position_38 : _GEN_3391; // @[StoreSet.scala 566:43 567:23]
  wire [2:0] _GEN_6691 = {{1'd0}, allocPtr_9}; // @[StoreSet.scala 565:51]
  wire [2:0] check_position_39 = _GEN_6691 + 3'h4; // @[StoreSet.scala 565:51]
  wire  _GEN_3398 = 2'h1 == check_position_39[1:0] ? validVec_9_1 : validVec_9_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3399 = 2'h2 == check_position_39[1:0] ? validVec_9_2 : _GEN_3398; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3400 = 2'h3 == check_position_39[1:0] ? validVec_9_3 : _GEN_3399; // @[StoreSet.scala 566:{14,14}]
  wire [2:0] _GEN_3401 = ~_GEN_3400 ? check_position_39 : {{1'd0}, _GEN_3396}; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_40 = allocPtr_10 + 2'h1; // @[StoreSet.scala 565:51]
  wire  _GEN_3403 = 2'h1 == check_position_40 ? validVec_10_1 : validVec_10_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3404 = 2'h2 == check_position_40 ? validVec_10_2 : _GEN_3403; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3405 = 2'h3 == check_position_40 ? validVec_10_3 : _GEN_3404; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3406 = ~_GEN_3405 ? check_position_40 : _GEN_2668; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_41 = allocPtr_10 + 2'h2; // @[StoreSet.scala 565:51]
  wire  _GEN_3408 = 2'h1 == check_position_41 ? validVec_10_1 : validVec_10_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3409 = 2'h2 == check_position_41 ? validVec_10_2 : _GEN_3408; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3410 = 2'h3 == check_position_41 ? validVec_10_3 : _GEN_3409; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3411 = ~_GEN_3410 ? check_position_41 : _GEN_3406; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_42 = allocPtr_10 + 2'h3; // @[StoreSet.scala 565:51]
  wire  _GEN_3413 = 2'h1 == check_position_42 ? validVec_10_1 : validVec_10_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3414 = 2'h2 == check_position_42 ? validVec_10_2 : _GEN_3413; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3415 = 2'h3 == check_position_42 ? validVec_10_3 : _GEN_3414; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3416 = ~_GEN_3415 ? check_position_42 : _GEN_3411; // @[StoreSet.scala 566:43 567:23]
  wire [2:0] _GEN_6692 = {{1'd0}, allocPtr_10}; // @[StoreSet.scala 565:51]
  wire [2:0] check_position_43 = _GEN_6692 + 3'h4; // @[StoreSet.scala 565:51]
  wire  _GEN_3418 = 2'h1 == check_position_43[1:0] ? validVec_10_1 : validVec_10_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3419 = 2'h2 == check_position_43[1:0] ? validVec_10_2 : _GEN_3418; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3420 = 2'h3 == check_position_43[1:0] ? validVec_10_3 : _GEN_3419; // @[StoreSet.scala 566:{14,14}]
  wire [2:0] _GEN_3421 = ~_GEN_3420 ? check_position_43 : {{1'd0}, _GEN_3416}; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_44 = allocPtr_11 + 2'h1; // @[StoreSet.scala 565:51]
  wire  _GEN_3423 = 2'h1 == check_position_44 ? validVec_11_1 : validVec_11_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3424 = 2'h2 == check_position_44 ? validVec_11_2 : _GEN_3423; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3425 = 2'h3 == check_position_44 ? validVec_11_3 : _GEN_3424; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3426 = ~_GEN_3425 ? check_position_44 : _GEN_2669; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_45 = allocPtr_11 + 2'h2; // @[StoreSet.scala 565:51]
  wire  _GEN_3428 = 2'h1 == check_position_45 ? validVec_11_1 : validVec_11_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3429 = 2'h2 == check_position_45 ? validVec_11_2 : _GEN_3428; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3430 = 2'h3 == check_position_45 ? validVec_11_3 : _GEN_3429; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3431 = ~_GEN_3430 ? check_position_45 : _GEN_3426; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_46 = allocPtr_11 + 2'h3; // @[StoreSet.scala 565:51]
  wire  _GEN_3433 = 2'h1 == check_position_46 ? validVec_11_1 : validVec_11_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3434 = 2'h2 == check_position_46 ? validVec_11_2 : _GEN_3433; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3435 = 2'h3 == check_position_46 ? validVec_11_3 : _GEN_3434; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3436 = ~_GEN_3435 ? check_position_46 : _GEN_3431; // @[StoreSet.scala 566:43 567:23]
  wire [2:0] _GEN_6693 = {{1'd0}, allocPtr_11}; // @[StoreSet.scala 565:51]
  wire [2:0] check_position_47 = _GEN_6693 + 3'h4; // @[StoreSet.scala 565:51]
  wire  _GEN_3438 = 2'h1 == check_position_47[1:0] ? validVec_11_1 : validVec_11_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3439 = 2'h2 == check_position_47[1:0] ? validVec_11_2 : _GEN_3438; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3440 = 2'h3 == check_position_47[1:0] ? validVec_11_3 : _GEN_3439; // @[StoreSet.scala 566:{14,14}]
  wire [2:0] _GEN_3441 = ~_GEN_3440 ? check_position_47 : {{1'd0}, _GEN_3436}; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_48 = allocPtr_12 + 2'h1; // @[StoreSet.scala 565:51]
  wire  _GEN_3443 = 2'h1 == check_position_48 ? validVec_12_1 : validVec_12_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3444 = 2'h2 == check_position_48 ? validVec_12_2 : _GEN_3443; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3445 = 2'h3 == check_position_48 ? validVec_12_3 : _GEN_3444; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3446 = ~_GEN_3445 ? check_position_48 : _GEN_2670; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_49 = allocPtr_12 + 2'h2; // @[StoreSet.scala 565:51]
  wire  _GEN_3448 = 2'h1 == check_position_49 ? validVec_12_1 : validVec_12_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3449 = 2'h2 == check_position_49 ? validVec_12_2 : _GEN_3448; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3450 = 2'h3 == check_position_49 ? validVec_12_3 : _GEN_3449; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3451 = ~_GEN_3450 ? check_position_49 : _GEN_3446; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_50 = allocPtr_12 + 2'h3; // @[StoreSet.scala 565:51]
  wire  _GEN_3453 = 2'h1 == check_position_50 ? validVec_12_1 : validVec_12_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3454 = 2'h2 == check_position_50 ? validVec_12_2 : _GEN_3453; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3455 = 2'h3 == check_position_50 ? validVec_12_3 : _GEN_3454; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3456 = ~_GEN_3455 ? check_position_50 : _GEN_3451; // @[StoreSet.scala 566:43 567:23]
  wire [2:0] _GEN_6694 = {{1'd0}, allocPtr_12}; // @[StoreSet.scala 565:51]
  wire [2:0] check_position_51 = _GEN_6694 + 3'h4; // @[StoreSet.scala 565:51]
  wire  _GEN_3458 = 2'h1 == check_position_51[1:0] ? validVec_12_1 : validVec_12_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3459 = 2'h2 == check_position_51[1:0] ? validVec_12_2 : _GEN_3458; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3460 = 2'h3 == check_position_51[1:0] ? validVec_12_3 : _GEN_3459; // @[StoreSet.scala 566:{14,14}]
  wire [2:0] _GEN_3461 = ~_GEN_3460 ? check_position_51 : {{1'd0}, _GEN_3456}; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_52 = allocPtr_13 + 2'h1; // @[StoreSet.scala 565:51]
  wire  _GEN_3463 = 2'h1 == check_position_52 ? validVec_13_1 : validVec_13_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3464 = 2'h2 == check_position_52 ? validVec_13_2 : _GEN_3463; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3465 = 2'h3 == check_position_52 ? validVec_13_3 : _GEN_3464; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3466 = ~_GEN_3465 ? check_position_52 : _GEN_2671; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_53 = allocPtr_13 + 2'h2; // @[StoreSet.scala 565:51]
  wire  _GEN_3468 = 2'h1 == check_position_53 ? validVec_13_1 : validVec_13_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3469 = 2'h2 == check_position_53 ? validVec_13_2 : _GEN_3468; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3470 = 2'h3 == check_position_53 ? validVec_13_3 : _GEN_3469; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3471 = ~_GEN_3470 ? check_position_53 : _GEN_3466; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_54 = allocPtr_13 + 2'h3; // @[StoreSet.scala 565:51]
  wire  _GEN_3473 = 2'h1 == check_position_54 ? validVec_13_1 : validVec_13_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3474 = 2'h2 == check_position_54 ? validVec_13_2 : _GEN_3473; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3475 = 2'h3 == check_position_54 ? validVec_13_3 : _GEN_3474; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3476 = ~_GEN_3475 ? check_position_54 : _GEN_3471; // @[StoreSet.scala 566:43 567:23]
  wire [2:0] _GEN_6695 = {{1'd0}, allocPtr_13}; // @[StoreSet.scala 565:51]
  wire [2:0] check_position_55 = _GEN_6695 + 3'h4; // @[StoreSet.scala 565:51]
  wire  _GEN_3478 = 2'h1 == check_position_55[1:0] ? validVec_13_1 : validVec_13_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3479 = 2'h2 == check_position_55[1:0] ? validVec_13_2 : _GEN_3478; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3480 = 2'h3 == check_position_55[1:0] ? validVec_13_3 : _GEN_3479; // @[StoreSet.scala 566:{14,14}]
  wire [2:0] _GEN_3481 = ~_GEN_3480 ? check_position_55 : {{1'd0}, _GEN_3476}; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_56 = allocPtr_14 + 2'h1; // @[StoreSet.scala 565:51]
  wire  _GEN_3483 = 2'h1 == check_position_56 ? validVec_14_1 : validVec_14_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3484 = 2'h2 == check_position_56 ? validVec_14_2 : _GEN_3483; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3485 = 2'h3 == check_position_56 ? validVec_14_3 : _GEN_3484; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3486 = ~_GEN_3485 ? check_position_56 : _GEN_2672; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_57 = allocPtr_14 + 2'h2; // @[StoreSet.scala 565:51]
  wire  _GEN_3488 = 2'h1 == check_position_57 ? validVec_14_1 : validVec_14_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3489 = 2'h2 == check_position_57 ? validVec_14_2 : _GEN_3488; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3490 = 2'h3 == check_position_57 ? validVec_14_3 : _GEN_3489; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3491 = ~_GEN_3490 ? check_position_57 : _GEN_3486; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_58 = allocPtr_14 + 2'h3; // @[StoreSet.scala 565:51]
  wire  _GEN_3493 = 2'h1 == check_position_58 ? validVec_14_1 : validVec_14_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3494 = 2'h2 == check_position_58 ? validVec_14_2 : _GEN_3493; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3495 = 2'h3 == check_position_58 ? validVec_14_3 : _GEN_3494; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3496 = ~_GEN_3495 ? check_position_58 : _GEN_3491; // @[StoreSet.scala 566:43 567:23]
  wire [2:0] _GEN_6696 = {{1'd0}, allocPtr_14}; // @[StoreSet.scala 565:51]
  wire [2:0] check_position_59 = _GEN_6696 + 3'h4; // @[StoreSet.scala 565:51]
  wire  _GEN_3498 = 2'h1 == check_position_59[1:0] ? validVec_14_1 : validVec_14_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3499 = 2'h2 == check_position_59[1:0] ? validVec_14_2 : _GEN_3498; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3500 = 2'h3 == check_position_59[1:0] ? validVec_14_3 : _GEN_3499; // @[StoreSet.scala 566:{14,14}]
  wire [2:0] _GEN_3501 = ~_GEN_3500 ? check_position_59 : {{1'd0}, _GEN_3496}; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_60 = allocPtr_15 + 2'h1; // @[StoreSet.scala 565:51]
  wire  _GEN_3503 = 2'h1 == check_position_60 ? validVec_15_1 : validVec_15_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3504 = 2'h2 == check_position_60 ? validVec_15_2 : _GEN_3503; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3505 = 2'h3 == check_position_60 ? validVec_15_3 : _GEN_3504; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3506 = ~_GEN_3505 ? check_position_60 : _GEN_2673; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_61 = allocPtr_15 + 2'h2; // @[StoreSet.scala 565:51]
  wire  _GEN_3508 = 2'h1 == check_position_61 ? validVec_15_1 : validVec_15_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3509 = 2'h2 == check_position_61 ? validVec_15_2 : _GEN_3508; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3510 = 2'h3 == check_position_61 ? validVec_15_3 : _GEN_3509; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3511 = ~_GEN_3510 ? check_position_61 : _GEN_3506; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_62 = allocPtr_15 + 2'h3; // @[StoreSet.scala 565:51]
  wire  _GEN_3513 = 2'h1 == check_position_62 ? validVec_15_1 : validVec_15_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3514 = 2'h2 == check_position_62 ? validVec_15_2 : _GEN_3513; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3515 = 2'h3 == check_position_62 ? validVec_15_3 : _GEN_3514; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3516 = ~_GEN_3515 ? check_position_62 : _GEN_3511; // @[StoreSet.scala 566:43 567:23]
  wire [2:0] _GEN_6697 = {{1'd0}, allocPtr_15}; // @[StoreSet.scala 565:51]
  wire [2:0] check_position_63 = _GEN_6697 + 3'h4; // @[StoreSet.scala 565:51]
  wire  _GEN_3518 = 2'h1 == check_position_63[1:0] ? validVec_15_1 : validVec_15_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3519 = 2'h2 == check_position_63[1:0] ? validVec_15_2 : _GEN_3518; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3520 = 2'h3 == check_position_63[1:0] ? validVec_15_3 : _GEN_3519; // @[StoreSet.scala 566:{14,14}]
  wire [2:0] _GEN_3521 = ~_GEN_3520 ? check_position_63 : {{1'd0}, _GEN_3516}; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_64 = allocPtr_16 + 2'h1; // @[StoreSet.scala 565:51]
  wire  _GEN_3523 = 2'h1 == check_position_64 ? validVec_16_1 : validVec_16_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3524 = 2'h2 == check_position_64 ? validVec_16_2 : _GEN_3523; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3525 = 2'h3 == check_position_64 ? validVec_16_3 : _GEN_3524; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3526 = ~_GEN_3525 ? check_position_64 : _GEN_2674; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_65 = allocPtr_16 + 2'h2; // @[StoreSet.scala 565:51]
  wire  _GEN_3528 = 2'h1 == check_position_65 ? validVec_16_1 : validVec_16_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3529 = 2'h2 == check_position_65 ? validVec_16_2 : _GEN_3528; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3530 = 2'h3 == check_position_65 ? validVec_16_3 : _GEN_3529; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3531 = ~_GEN_3530 ? check_position_65 : _GEN_3526; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_66 = allocPtr_16 + 2'h3; // @[StoreSet.scala 565:51]
  wire  _GEN_3533 = 2'h1 == check_position_66 ? validVec_16_1 : validVec_16_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3534 = 2'h2 == check_position_66 ? validVec_16_2 : _GEN_3533; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3535 = 2'h3 == check_position_66 ? validVec_16_3 : _GEN_3534; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3536 = ~_GEN_3535 ? check_position_66 : _GEN_3531; // @[StoreSet.scala 566:43 567:23]
  wire [2:0] _GEN_6698 = {{1'd0}, allocPtr_16}; // @[StoreSet.scala 565:51]
  wire [2:0] check_position_67 = _GEN_6698 + 3'h4; // @[StoreSet.scala 565:51]
  wire  _GEN_3538 = 2'h1 == check_position_67[1:0] ? validVec_16_1 : validVec_16_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3539 = 2'h2 == check_position_67[1:0] ? validVec_16_2 : _GEN_3538; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3540 = 2'h3 == check_position_67[1:0] ? validVec_16_3 : _GEN_3539; // @[StoreSet.scala 566:{14,14}]
  wire [2:0] _GEN_3541 = ~_GEN_3540 ? check_position_67 : {{1'd0}, _GEN_3536}; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_68 = allocPtr_17 + 2'h1; // @[StoreSet.scala 565:51]
  wire  _GEN_3543 = 2'h1 == check_position_68 ? validVec_17_1 : validVec_17_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3544 = 2'h2 == check_position_68 ? validVec_17_2 : _GEN_3543; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3545 = 2'h3 == check_position_68 ? validVec_17_3 : _GEN_3544; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3546 = ~_GEN_3545 ? check_position_68 : _GEN_2675; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_69 = allocPtr_17 + 2'h2; // @[StoreSet.scala 565:51]
  wire  _GEN_3548 = 2'h1 == check_position_69 ? validVec_17_1 : validVec_17_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3549 = 2'h2 == check_position_69 ? validVec_17_2 : _GEN_3548; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3550 = 2'h3 == check_position_69 ? validVec_17_3 : _GEN_3549; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3551 = ~_GEN_3550 ? check_position_69 : _GEN_3546; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_70 = allocPtr_17 + 2'h3; // @[StoreSet.scala 565:51]
  wire  _GEN_3553 = 2'h1 == check_position_70 ? validVec_17_1 : validVec_17_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3554 = 2'h2 == check_position_70 ? validVec_17_2 : _GEN_3553; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3555 = 2'h3 == check_position_70 ? validVec_17_3 : _GEN_3554; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3556 = ~_GEN_3555 ? check_position_70 : _GEN_3551; // @[StoreSet.scala 566:43 567:23]
  wire [2:0] _GEN_6699 = {{1'd0}, allocPtr_17}; // @[StoreSet.scala 565:51]
  wire [2:0] check_position_71 = _GEN_6699 + 3'h4; // @[StoreSet.scala 565:51]
  wire  _GEN_3558 = 2'h1 == check_position_71[1:0] ? validVec_17_1 : validVec_17_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3559 = 2'h2 == check_position_71[1:0] ? validVec_17_2 : _GEN_3558; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3560 = 2'h3 == check_position_71[1:0] ? validVec_17_3 : _GEN_3559; // @[StoreSet.scala 566:{14,14}]
  wire [2:0] _GEN_3561 = ~_GEN_3560 ? check_position_71 : {{1'd0}, _GEN_3556}; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_72 = allocPtr_18 + 2'h1; // @[StoreSet.scala 565:51]
  wire  _GEN_3563 = 2'h1 == check_position_72 ? validVec_18_1 : validVec_18_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3564 = 2'h2 == check_position_72 ? validVec_18_2 : _GEN_3563; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3565 = 2'h3 == check_position_72 ? validVec_18_3 : _GEN_3564; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3566 = ~_GEN_3565 ? check_position_72 : _GEN_2676; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_73 = allocPtr_18 + 2'h2; // @[StoreSet.scala 565:51]
  wire  _GEN_3568 = 2'h1 == check_position_73 ? validVec_18_1 : validVec_18_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3569 = 2'h2 == check_position_73 ? validVec_18_2 : _GEN_3568; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3570 = 2'h3 == check_position_73 ? validVec_18_3 : _GEN_3569; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3571 = ~_GEN_3570 ? check_position_73 : _GEN_3566; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_74 = allocPtr_18 + 2'h3; // @[StoreSet.scala 565:51]
  wire  _GEN_3573 = 2'h1 == check_position_74 ? validVec_18_1 : validVec_18_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3574 = 2'h2 == check_position_74 ? validVec_18_2 : _GEN_3573; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3575 = 2'h3 == check_position_74 ? validVec_18_3 : _GEN_3574; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3576 = ~_GEN_3575 ? check_position_74 : _GEN_3571; // @[StoreSet.scala 566:43 567:23]
  wire [2:0] _GEN_6700 = {{1'd0}, allocPtr_18}; // @[StoreSet.scala 565:51]
  wire [2:0] check_position_75 = _GEN_6700 + 3'h4; // @[StoreSet.scala 565:51]
  wire  _GEN_3578 = 2'h1 == check_position_75[1:0] ? validVec_18_1 : validVec_18_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3579 = 2'h2 == check_position_75[1:0] ? validVec_18_2 : _GEN_3578; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3580 = 2'h3 == check_position_75[1:0] ? validVec_18_3 : _GEN_3579; // @[StoreSet.scala 566:{14,14}]
  wire [2:0] _GEN_3581 = ~_GEN_3580 ? check_position_75 : {{1'd0}, _GEN_3576}; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_76 = allocPtr_19 + 2'h1; // @[StoreSet.scala 565:51]
  wire  _GEN_3583 = 2'h1 == check_position_76 ? validVec_19_1 : validVec_19_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3584 = 2'h2 == check_position_76 ? validVec_19_2 : _GEN_3583; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3585 = 2'h3 == check_position_76 ? validVec_19_3 : _GEN_3584; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3586 = ~_GEN_3585 ? check_position_76 : _GEN_2677; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_77 = allocPtr_19 + 2'h2; // @[StoreSet.scala 565:51]
  wire  _GEN_3588 = 2'h1 == check_position_77 ? validVec_19_1 : validVec_19_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3589 = 2'h2 == check_position_77 ? validVec_19_2 : _GEN_3588; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3590 = 2'h3 == check_position_77 ? validVec_19_3 : _GEN_3589; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3591 = ~_GEN_3590 ? check_position_77 : _GEN_3586; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_78 = allocPtr_19 + 2'h3; // @[StoreSet.scala 565:51]
  wire  _GEN_3593 = 2'h1 == check_position_78 ? validVec_19_1 : validVec_19_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3594 = 2'h2 == check_position_78 ? validVec_19_2 : _GEN_3593; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3595 = 2'h3 == check_position_78 ? validVec_19_3 : _GEN_3594; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3596 = ~_GEN_3595 ? check_position_78 : _GEN_3591; // @[StoreSet.scala 566:43 567:23]
  wire [2:0] _GEN_6701 = {{1'd0}, allocPtr_19}; // @[StoreSet.scala 565:51]
  wire [2:0] check_position_79 = _GEN_6701 + 3'h4; // @[StoreSet.scala 565:51]
  wire  _GEN_3598 = 2'h1 == check_position_79[1:0] ? validVec_19_1 : validVec_19_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3599 = 2'h2 == check_position_79[1:0] ? validVec_19_2 : _GEN_3598; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3600 = 2'h3 == check_position_79[1:0] ? validVec_19_3 : _GEN_3599; // @[StoreSet.scala 566:{14,14}]
  wire [2:0] _GEN_3601 = ~_GEN_3600 ? check_position_79 : {{1'd0}, _GEN_3596}; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_80 = allocPtr_20 + 2'h1; // @[StoreSet.scala 565:51]
  wire  _GEN_3603 = 2'h1 == check_position_80 ? validVec_20_1 : validVec_20_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3604 = 2'h2 == check_position_80 ? validVec_20_2 : _GEN_3603; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3605 = 2'h3 == check_position_80 ? validVec_20_3 : _GEN_3604; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3606 = ~_GEN_3605 ? check_position_80 : _GEN_2678; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_81 = allocPtr_20 + 2'h2; // @[StoreSet.scala 565:51]
  wire  _GEN_3608 = 2'h1 == check_position_81 ? validVec_20_1 : validVec_20_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3609 = 2'h2 == check_position_81 ? validVec_20_2 : _GEN_3608; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3610 = 2'h3 == check_position_81 ? validVec_20_3 : _GEN_3609; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3611 = ~_GEN_3610 ? check_position_81 : _GEN_3606; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_82 = allocPtr_20 + 2'h3; // @[StoreSet.scala 565:51]
  wire  _GEN_3613 = 2'h1 == check_position_82 ? validVec_20_1 : validVec_20_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3614 = 2'h2 == check_position_82 ? validVec_20_2 : _GEN_3613; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3615 = 2'h3 == check_position_82 ? validVec_20_3 : _GEN_3614; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3616 = ~_GEN_3615 ? check_position_82 : _GEN_3611; // @[StoreSet.scala 566:43 567:23]
  wire [2:0] _GEN_6702 = {{1'd0}, allocPtr_20}; // @[StoreSet.scala 565:51]
  wire [2:0] check_position_83 = _GEN_6702 + 3'h4; // @[StoreSet.scala 565:51]
  wire  _GEN_3618 = 2'h1 == check_position_83[1:0] ? validVec_20_1 : validVec_20_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3619 = 2'h2 == check_position_83[1:0] ? validVec_20_2 : _GEN_3618; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3620 = 2'h3 == check_position_83[1:0] ? validVec_20_3 : _GEN_3619; // @[StoreSet.scala 566:{14,14}]
  wire [2:0] _GEN_3621 = ~_GEN_3620 ? check_position_83 : {{1'd0}, _GEN_3616}; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_84 = allocPtr_21 + 2'h1; // @[StoreSet.scala 565:51]
  wire  _GEN_3623 = 2'h1 == check_position_84 ? validVec_21_1 : validVec_21_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3624 = 2'h2 == check_position_84 ? validVec_21_2 : _GEN_3623; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3625 = 2'h3 == check_position_84 ? validVec_21_3 : _GEN_3624; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3626 = ~_GEN_3625 ? check_position_84 : _GEN_2679; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_85 = allocPtr_21 + 2'h2; // @[StoreSet.scala 565:51]
  wire  _GEN_3628 = 2'h1 == check_position_85 ? validVec_21_1 : validVec_21_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3629 = 2'h2 == check_position_85 ? validVec_21_2 : _GEN_3628; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3630 = 2'h3 == check_position_85 ? validVec_21_3 : _GEN_3629; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3631 = ~_GEN_3630 ? check_position_85 : _GEN_3626; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_86 = allocPtr_21 + 2'h3; // @[StoreSet.scala 565:51]
  wire  _GEN_3633 = 2'h1 == check_position_86 ? validVec_21_1 : validVec_21_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3634 = 2'h2 == check_position_86 ? validVec_21_2 : _GEN_3633; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3635 = 2'h3 == check_position_86 ? validVec_21_3 : _GEN_3634; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3636 = ~_GEN_3635 ? check_position_86 : _GEN_3631; // @[StoreSet.scala 566:43 567:23]
  wire [2:0] _GEN_6703 = {{1'd0}, allocPtr_21}; // @[StoreSet.scala 565:51]
  wire [2:0] check_position_87 = _GEN_6703 + 3'h4; // @[StoreSet.scala 565:51]
  wire  _GEN_3638 = 2'h1 == check_position_87[1:0] ? validVec_21_1 : validVec_21_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3639 = 2'h2 == check_position_87[1:0] ? validVec_21_2 : _GEN_3638; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3640 = 2'h3 == check_position_87[1:0] ? validVec_21_3 : _GEN_3639; // @[StoreSet.scala 566:{14,14}]
  wire [2:0] _GEN_3641 = ~_GEN_3640 ? check_position_87 : {{1'd0}, _GEN_3636}; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_88 = allocPtr_22 + 2'h1; // @[StoreSet.scala 565:51]
  wire  _GEN_3643 = 2'h1 == check_position_88 ? validVec_22_1 : validVec_22_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3644 = 2'h2 == check_position_88 ? validVec_22_2 : _GEN_3643; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3645 = 2'h3 == check_position_88 ? validVec_22_3 : _GEN_3644; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3646 = ~_GEN_3645 ? check_position_88 : _GEN_2680; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_89 = allocPtr_22 + 2'h2; // @[StoreSet.scala 565:51]
  wire  _GEN_3648 = 2'h1 == check_position_89 ? validVec_22_1 : validVec_22_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3649 = 2'h2 == check_position_89 ? validVec_22_2 : _GEN_3648; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3650 = 2'h3 == check_position_89 ? validVec_22_3 : _GEN_3649; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3651 = ~_GEN_3650 ? check_position_89 : _GEN_3646; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_90 = allocPtr_22 + 2'h3; // @[StoreSet.scala 565:51]
  wire  _GEN_3653 = 2'h1 == check_position_90 ? validVec_22_1 : validVec_22_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3654 = 2'h2 == check_position_90 ? validVec_22_2 : _GEN_3653; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3655 = 2'h3 == check_position_90 ? validVec_22_3 : _GEN_3654; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3656 = ~_GEN_3655 ? check_position_90 : _GEN_3651; // @[StoreSet.scala 566:43 567:23]
  wire [2:0] _GEN_6704 = {{1'd0}, allocPtr_22}; // @[StoreSet.scala 565:51]
  wire [2:0] check_position_91 = _GEN_6704 + 3'h4; // @[StoreSet.scala 565:51]
  wire  _GEN_3658 = 2'h1 == check_position_91[1:0] ? validVec_22_1 : validVec_22_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3659 = 2'h2 == check_position_91[1:0] ? validVec_22_2 : _GEN_3658; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3660 = 2'h3 == check_position_91[1:0] ? validVec_22_3 : _GEN_3659; // @[StoreSet.scala 566:{14,14}]
  wire [2:0] _GEN_3661 = ~_GEN_3660 ? check_position_91 : {{1'd0}, _GEN_3656}; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_92 = allocPtr_23 + 2'h1; // @[StoreSet.scala 565:51]
  wire  _GEN_3663 = 2'h1 == check_position_92 ? validVec_23_1 : validVec_23_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3664 = 2'h2 == check_position_92 ? validVec_23_2 : _GEN_3663; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3665 = 2'h3 == check_position_92 ? validVec_23_3 : _GEN_3664; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3666 = ~_GEN_3665 ? check_position_92 : _GEN_2681; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_93 = allocPtr_23 + 2'h2; // @[StoreSet.scala 565:51]
  wire  _GEN_3668 = 2'h1 == check_position_93 ? validVec_23_1 : validVec_23_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3669 = 2'h2 == check_position_93 ? validVec_23_2 : _GEN_3668; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3670 = 2'h3 == check_position_93 ? validVec_23_3 : _GEN_3669; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3671 = ~_GEN_3670 ? check_position_93 : _GEN_3666; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_94 = allocPtr_23 + 2'h3; // @[StoreSet.scala 565:51]
  wire  _GEN_3673 = 2'h1 == check_position_94 ? validVec_23_1 : validVec_23_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3674 = 2'h2 == check_position_94 ? validVec_23_2 : _GEN_3673; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3675 = 2'h3 == check_position_94 ? validVec_23_3 : _GEN_3674; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3676 = ~_GEN_3675 ? check_position_94 : _GEN_3671; // @[StoreSet.scala 566:43 567:23]
  wire [2:0] _GEN_6705 = {{1'd0}, allocPtr_23}; // @[StoreSet.scala 565:51]
  wire [2:0] check_position_95 = _GEN_6705 + 3'h4; // @[StoreSet.scala 565:51]
  wire  _GEN_3678 = 2'h1 == check_position_95[1:0] ? validVec_23_1 : validVec_23_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3679 = 2'h2 == check_position_95[1:0] ? validVec_23_2 : _GEN_3678; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3680 = 2'h3 == check_position_95[1:0] ? validVec_23_3 : _GEN_3679; // @[StoreSet.scala 566:{14,14}]
  wire [2:0] _GEN_3681 = ~_GEN_3680 ? check_position_95 : {{1'd0}, _GEN_3676}; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_96 = allocPtr_24 + 2'h1; // @[StoreSet.scala 565:51]
  wire  _GEN_3683 = 2'h1 == check_position_96 ? validVec_24_1 : validVec_24_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3684 = 2'h2 == check_position_96 ? validVec_24_2 : _GEN_3683; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3685 = 2'h3 == check_position_96 ? validVec_24_3 : _GEN_3684; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3686 = ~_GEN_3685 ? check_position_96 : _GEN_2682; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_97 = allocPtr_24 + 2'h2; // @[StoreSet.scala 565:51]
  wire  _GEN_3688 = 2'h1 == check_position_97 ? validVec_24_1 : validVec_24_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3689 = 2'h2 == check_position_97 ? validVec_24_2 : _GEN_3688; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3690 = 2'h3 == check_position_97 ? validVec_24_3 : _GEN_3689; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3691 = ~_GEN_3690 ? check_position_97 : _GEN_3686; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_98 = allocPtr_24 + 2'h3; // @[StoreSet.scala 565:51]
  wire  _GEN_3693 = 2'h1 == check_position_98 ? validVec_24_1 : validVec_24_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3694 = 2'h2 == check_position_98 ? validVec_24_2 : _GEN_3693; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3695 = 2'h3 == check_position_98 ? validVec_24_3 : _GEN_3694; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3696 = ~_GEN_3695 ? check_position_98 : _GEN_3691; // @[StoreSet.scala 566:43 567:23]
  wire [2:0] _GEN_6706 = {{1'd0}, allocPtr_24}; // @[StoreSet.scala 565:51]
  wire [2:0] check_position_99 = _GEN_6706 + 3'h4; // @[StoreSet.scala 565:51]
  wire  _GEN_3698 = 2'h1 == check_position_99[1:0] ? validVec_24_1 : validVec_24_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3699 = 2'h2 == check_position_99[1:0] ? validVec_24_2 : _GEN_3698; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3700 = 2'h3 == check_position_99[1:0] ? validVec_24_3 : _GEN_3699; // @[StoreSet.scala 566:{14,14}]
  wire [2:0] _GEN_3701 = ~_GEN_3700 ? check_position_99 : {{1'd0}, _GEN_3696}; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_100 = allocPtr_25 + 2'h1; // @[StoreSet.scala 565:51]
  wire  _GEN_3703 = 2'h1 == check_position_100 ? validVec_25_1 : validVec_25_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3704 = 2'h2 == check_position_100 ? validVec_25_2 : _GEN_3703; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3705 = 2'h3 == check_position_100 ? validVec_25_3 : _GEN_3704; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3706 = ~_GEN_3705 ? check_position_100 : _GEN_2683; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_101 = allocPtr_25 + 2'h2; // @[StoreSet.scala 565:51]
  wire  _GEN_3708 = 2'h1 == check_position_101 ? validVec_25_1 : validVec_25_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3709 = 2'h2 == check_position_101 ? validVec_25_2 : _GEN_3708; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3710 = 2'h3 == check_position_101 ? validVec_25_3 : _GEN_3709; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3711 = ~_GEN_3710 ? check_position_101 : _GEN_3706; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_102 = allocPtr_25 + 2'h3; // @[StoreSet.scala 565:51]
  wire  _GEN_3713 = 2'h1 == check_position_102 ? validVec_25_1 : validVec_25_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3714 = 2'h2 == check_position_102 ? validVec_25_2 : _GEN_3713; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3715 = 2'h3 == check_position_102 ? validVec_25_3 : _GEN_3714; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3716 = ~_GEN_3715 ? check_position_102 : _GEN_3711; // @[StoreSet.scala 566:43 567:23]
  wire [2:0] _GEN_6707 = {{1'd0}, allocPtr_25}; // @[StoreSet.scala 565:51]
  wire [2:0] check_position_103 = _GEN_6707 + 3'h4; // @[StoreSet.scala 565:51]
  wire  _GEN_3718 = 2'h1 == check_position_103[1:0] ? validVec_25_1 : validVec_25_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3719 = 2'h2 == check_position_103[1:0] ? validVec_25_2 : _GEN_3718; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3720 = 2'h3 == check_position_103[1:0] ? validVec_25_3 : _GEN_3719; // @[StoreSet.scala 566:{14,14}]
  wire [2:0] _GEN_3721 = ~_GEN_3720 ? check_position_103 : {{1'd0}, _GEN_3716}; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_104 = allocPtr_26 + 2'h1; // @[StoreSet.scala 565:51]
  wire  _GEN_3723 = 2'h1 == check_position_104 ? validVec_26_1 : validVec_26_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3724 = 2'h2 == check_position_104 ? validVec_26_2 : _GEN_3723; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3725 = 2'h3 == check_position_104 ? validVec_26_3 : _GEN_3724; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3726 = ~_GEN_3725 ? check_position_104 : _GEN_2684; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_105 = allocPtr_26 + 2'h2; // @[StoreSet.scala 565:51]
  wire  _GEN_3728 = 2'h1 == check_position_105 ? validVec_26_1 : validVec_26_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3729 = 2'h2 == check_position_105 ? validVec_26_2 : _GEN_3728; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3730 = 2'h3 == check_position_105 ? validVec_26_3 : _GEN_3729; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3731 = ~_GEN_3730 ? check_position_105 : _GEN_3726; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_106 = allocPtr_26 + 2'h3; // @[StoreSet.scala 565:51]
  wire  _GEN_3733 = 2'h1 == check_position_106 ? validVec_26_1 : validVec_26_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3734 = 2'h2 == check_position_106 ? validVec_26_2 : _GEN_3733; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3735 = 2'h3 == check_position_106 ? validVec_26_3 : _GEN_3734; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3736 = ~_GEN_3735 ? check_position_106 : _GEN_3731; // @[StoreSet.scala 566:43 567:23]
  wire [2:0] _GEN_6708 = {{1'd0}, allocPtr_26}; // @[StoreSet.scala 565:51]
  wire [2:0] check_position_107 = _GEN_6708 + 3'h4; // @[StoreSet.scala 565:51]
  wire  _GEN_3738 = 2'h1 == check_position_107[1:0] ? validVec_26_1 : validVec_26_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3739 = 2'h2 == check_position_107[1:0] ? validVec_26_2 : _GEN_3738; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3740 = 2'h3 == check_position_107[1:0] ? validVec_26_3 : _GEN_3739; // @[StoreSet.scala 566:{14,14}]
  wire [2:0] _GEN_3741 = ~_GEN_3740 ? check_position_107 : {{1'd0}, _GEN_3736}; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_108 = allocPtr_27 + 2'h1; // @[StoreSet.scala 565:51]
  wire  _GEN_3743 = 2'h1 == check_position_108 ? validVec_27_1 : validVec_27_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3744 = 2'h2 == check_position_108 ? validVec_27_2 : _GEN_3743; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3745 = 2'h3 == check_position_108 ? validVec_27_3 : _GEN_3744; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3746 = ~_GEN_3745 ? check_position_108 : _GEN_2685; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_109 = allocPtr_27 + 2'h2; // @[StoreSet.scala 565:51]
  wire  _GEN_3748 = 2'h1 == check_position_109 ? validVec_27_1 : validVec_27_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3749 = 2'h2 == check_position_109 ? validVec_27_2 : _GEN_3748; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3750 = 2'h3 == check_position_109 ? validVec_27_3 : _GEN_3749; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3751 = ~_GEN_3750 ? check_position_109 : _GEN_3746; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_110 = allocPtr_27 + 2'h3; // @[StoreSet.scala 565:51]
  wire  _GEN_3753 = 2'h1 == check_position_110 ? validVec_27_1 : validVec_27_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3754 = 2'h2 == check_position_110 ? validVec_27_2 : _GEN_3753; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3755 = 2'h3 == check_position_110 ? validVec_27_3 : _GEN_3754; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3756 = ~_GEN_3755 ? check_position_110 : _GEN_3751; // @[StoreSet.scala 566:43 567:23]
  wire [2:0] _GEN_6709 = {{1'd0}, allocPtr_27}; // @[StoreSet.scala 565:51]
  wire [2:0] check_position_111 = _GEN_6709 + 3'h4; // @[StoreSet.scala 565:51]
  wire  _GEN_3758 = 2'h1 == check_position_111[1:0] ? validVec_27_1 : validVec_27_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3759 = 2'h2 == check_position_111[1:0] ? validVec_27_2 : _GEN_3758; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3760 = 2'h3 == check_position_111[1:0] ? validVec_27_3 : _GEN_3759; // @[StoreSet.scala 566:{14,14}]
  wire [2:0] _GEN_3761 = ~_GEN_3760 ? check_position_111 : {{1'd0}, _GEN_3756}; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_112 = allocPtr_28 + 2'h1; // @[StoreSet.scala 565:51]
  wire  _GEN_3763 = 2'h1 == check_position_112 ? validVec_28_1 : validVec_28_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3764 = 2'h2 == check_position_112 ? validVec_28_2 : _GEN_3763; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3765 = 2'h3 == check_position_112 ? validVec_28_3 : _GEN_3764; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3766 = ~_GEN_3765 ? check_position_112 : _GEN_2686; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_113 = allocPtr_28 + 2'h2; // @[StoreSet.scala 565:51]
  wire  _GEN_3768 = 2'h1 == check_position_113 ? validVec_28_1 : validVec_28_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3769 = 2'h2 == check_position_113 ? validVec_28_2 : _GEN_3768; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3770 = 2'h3 == check_position_113 ? validVec_28_3 : _GEN_3769; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3771 = ~_GEN_3770 ? check_position_113 : _GEN_3766; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_114 = allocPtr_28 + 2'h3; // @[StoreSet.scala 565:51]
  wire  _GEN_3773 = 2'h1 == check_position_114 ? validVec_28_1 : validVec_28_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3774 = 2'h2 == check_position_114 ? validVec_28_2 : _GEN_3773; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3775 = 2'h3 == check_position_114 ? validVec_28_3 : _GEN_3774; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3776 = ~_GEN_3775 ? check_position_114 : _GEN_3771; // @[StoreSet.scala 566:43 567:23]
  wire [2:0] _GEN_6710 = {{1'd0}, allocPtr_28}; // @[StoreSet.scala 565:51]
  wire [2:0] check_position_115 = _GEN_6710 + 3'h4; // @[StoreSet.scala 565:51]
  wire  _GEN_3778 = 2'h1 == check_position_115[1:0] ? validVec_28_1 : validVec_28_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3779 = 2'h2 == check_position_115[1:0] ? validVec_28_2 : _GEN_3778; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3780 = 2'h3 == check_position_115[1:0] ? validVec_28_3 : _GEN_3779; // @[StoreSet.scala 566:{14,14}]
  wire [2:0] _GEN_3781 = ~_GEN_3780 ? check_position_115 : {{1'd0}, _GEN_3776}; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_116 = allocPtr_29 + 2'h1; // @[StoreSet.scala 565:51]
  wire  _GEN_3783 = 2'h1 == check_position_116 ? validVec_29_1 : validVec_29_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3784 = 2'h2 == check_position_116 ? validVec_29_2 : _GEN_3783; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3785 = 2'h3 == check_position_116 ? validVec_29_3 : _GEN_3784; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3786 = ~_GEN_3785 ? check_position_116 : _GEN_2687; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_117 = allocPtr_29 + 2'h2; // @[StoreSet.scala 565:51]
  wire  _GEN_3788 = 2'h1 == check_position_117 ? validVec_29_1 : validVec_29_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3789 = 2'h2 == check_position_117 ? validVec_29_2 : _GEN_3788; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3790 = 2'h3 == check_position_117 ? validVec_29_3 : _GEN_3789; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3791 = ~_GEN_3790 ? check_position_117 : _GEN_3786; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_118 = allocPtr_29 + 2'h3; // @[StoreSet.scala 565:51]
  wire  _GEN_3793 = 2'h1 == check_position_118 ? validVec_29_1 : validVec_29_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3794 = 2'h2 == check_position_118 ? validVec_29_2 : _GEN_3793; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3795 = 2'h3 == check_position_118 ? validVec_29_3 : _GEN_3794; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3796 = ~_GEN_3795 ? check_position_118 : _GEN_3791; // @[StoreSet.scala 566:43 567:23]
  wire [2:0] _GEN_6711 = {{1'd0}, allocPtr_29}; // @[StoreSet.scala 565:51]
  wire [2:0] check_position_119 = _GEN_6711 + 3'h4; // @[StoreSet.scala 565:51]
  wire  _GEN_3798 = 2'h1 == check_position_119[1:0] ? validVec_29_1 : validVec_29_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3799 = 2'h2 == check_position_119[1:0] ? validVec_29_2 : _GEN_3798; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3800 = 2'h3 == check_position_119[1:0] ? validVec_29_3 : _GEN_3799; // @[StoreSet.scala 566:{14,14}]
  wire [2:0] _GEN_3801 = ~_GEN_3800 ? check_position_119 : {{1'd0}, _GEN_3796}; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_120 = allocPtr_30 + 2'h1; // @[StoreSet.scala 565:51]
  wire  _GEN_3803 = 2'h1 == check_position_120 ? validVec_30_1 : validVec_30_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3804 = 2'h2 == check_position_120 ? validVec_30_2 : _GEN_3803; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3805 = 2'h3 == check_position_120 ? validVec_30_3 : _GEN_3804; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3806 = ~_GEN_3805 ? check_position_120 : _GEN_2688; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_121 = allocPtr_30 + 2'h2; // @[StoreSet.scala 565:51]
  wire  _GEN_3808 = 2'h1 == check_position_121 ? validVec_30_1 : validVec_30_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3809 = 2'h2 == check_position_121 ? validVec_30_2 : _GEN_3808; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3810 = 2'h3 == check_position_121 ? validVec_30_3 : _GEN_3809; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3811 = ~_GEN_3810 ? check_position_121 : _GEN_3806; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_122 = allocPtr_30 + 2'h3; // @[StoreSet.scala 565:51]
  wire  _GEN_3813 = 2'h1 == check_position_122 ? validVec_30_1 : validVec_30_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3814 = 2'h2 == check_position_122 ? validVec_30_2 : _GEN_3813; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3815 = 2'h3 == check_position_122 ? validVec_30_3 : _GEN_3814; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3816 = ~_GEN_3815 ? check_position_122 : _GEN_3811; // @[StoreSet.scala 566:43 567:23]
  wire [2:0] _GEN_6712 = {{1'd0}, allocPtr_30}; // @[StoreSet.scala 565:51]
  wire [2:0] check_position_123 = _GEN_6712 + 3'h4; // @[StoreSet.scala 565:51]
  wire  _GEN_3818 = 2'h1 == check_position_123[1:0] ? validVec_30_1 : validVec_30_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3819 = 2'h2 == check_position_123[1:0] ? validVec_30_2 : _GEN_3818; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3820 = 2'h3 == check_position_123[1:0] ? validVec_30_3 : _GEN_3819; // @[StoreSet.scala 566:{14,14}]
  wire [2:0] _GEN_3821 = ~_GEN_3820 ? check_position_123 : {{1'd0}, _GEN_3816}; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_124 = allocPtr_31 + 2'h1; // @[StoreSet.scala 565:51]
  wire  _GEN_3823 = 2'h1 == check_position_124 ? validVec_31_1 : validVec_31_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3824 = 2'h2 == check_position_124 ? validVec_31_2 : _GEN_3823; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3825 = 2'h3 == check_position_124 ? validVec_31_3 : _GEN_3824; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3826 = ~_GEN_3825 ? check_position_124 : _GEN_2689; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_125 = allocPtr_31 + 2'h2; // @[StoreSet.scala 565:51]
  wire  _GEN_3828 = 2'h1 == check_position_125 ? validVec_31_1 : validVec_31_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3829 = 2'h2 == check_position_125 ? validVec_31_2 : _GEN_3828; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3830 = 2'h3 == check_position_125 ? validVec_31_3 : _GEN_3829; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3831 = ~_GEN_3830 ? check_position_125 : _GEN_3826; // @[StoreSet.scala 566:43 567:23]
  wire [1:0] check_position_126 = allocPtr_31 + 2'h3; // @[StoreSet.scala 565:51]
  wire  _GEN_3833 = 2'h1 == check_position_126 ? validVec_31_1 : validVec_31_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3834 = 2'h2 == check_position_126 ? validVec_31_2 : _GEN_3833; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3835 = 2'h3 == check_position_126 ? validVec_31_3 : _GEN_3834; // @[StoreSet.scala 566:{14,14}]
  wire [1:0] _GEN_3836 = ~_GEN_3835 ? check_position_126 : _GEN_3831; // @[StoreSet.scala 566:43 567:23]
  wire [2:0] _GEN_6713 = {{1'd0}, allocPtr_31}; // @[StoreSet.scala 565:51]
  wire [2:0] check_position_127 = _GEN_6713 + 3'h4; // @[StoreSet.scala 565:51]
  wire  _GEN_3838 = 2'h1 == check_position_127[1:0] ? validVec_31_1 : validVec_31_0; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3839 = 2'h2 == check_position_127[1:0] ? validVec_31_2 : _GEN_3838; // @[StoreSet.scala 566:{14,14}]
  wire  _GEN_3840 = 2'h3 == check_position_127[1:0] ? validVec_31_3 : _GEN_3839; // @[StoreSet.scala 566:{14,14}]
  wire [2:0] _GEN_3841 = ~_GEN_3840 ? check_position_127 : {{1'd0}, _GEN_3836}; // @[StoreSet.scala 566:43 567:23]
  wire [2:0] _GEN_3842 = REG ? _GEN_3221 : {{1'd0}, _GEN_2658}; // @[StoreSet.scala 562:37]
  wire [2:0] _GEN_3843 = REG ? _GEN_3241 : {{1'd0}, _GEN_2659}; // @[StoreSet.scala 562:37]
  wire [2:0] _GEN_3844 = REG ? _GEN_3261 : {{1'd0}, _GEN_2660}; // @[StoreSet.scala 562:37]
  wire [2:0] _GEN_3845 = REG ? _GEN_3281 : {{1'd0}, _GEN_2661}; // @[StoreSet.scala 562:37]
  wire [2:0] _GEN_3846 = REG ? _GEN_3301 : {{1'd0}, _GEN_2662}; // @[StoreSet.scala 562:37]
  wire [2:0] _GEN_3847 = REG ? _GEN_3321 : {{1'd0}, _GEN_2663}; // @[StoreSet.scala 562:37]
  wire [2:0] _GEN_3848 = REG ? _GEN_3341 : {{1'd0}, _GEN_2664}; // @[StoreSet.scala 562:37]
  wire [2:0] _GEN_3849 = REG ? _GEN_3361 : {{1'd0}, _GEN_2665}; // @[StoreSet.scala 562:37]
  wire [2:0] _GEN_3850 = REG ? _GEN_3381 : {{1'd0}, _GEN_2666}; // @[StoreSet.scala 562:37]
  wire [2:0] _GEN_3851 = REG ? _GEN_3401 : {{1'd0}, _GEN_2667}; // @[StoreSet.scala 562:37]
  wire [2:0] _GEN_3852 = REG ? _GEN_3421 : {{1'd0}, _GEN_2668}; // @[StoreSet.scala 562:37]
  wire [2:0] _GEN_3853 = REG ? _GEN_3441 : {{1'd0}, _GEN_2669}; // @[StoreSet.scala 562:37]
  wire [2:0] _GEN_3854 = REG ? _GEN_3461 : {{1'd0}, _GEN_2670}; // @[StoreSet.scala 562:37]
  wire [2:0] _GEN_3855 = REG ? _GEN_3481 : {{1'd0}, _GEN_2671}; // @[StoreSet.scala 562:37]
  wire [2:0] _GEN_3856 = REG ? _GEN_3501 : {{1'd0}, _GEN_2672}; // @[StoreSet.scala 562:37]
  wire [2:0] _GEN_3857 = REG ? _GEN_3521 : {{1'd0}, _GEN_2673}; // @[StoreSet.scala 562:37]
  wire [2:0] _GEN_3858 = REG ? _GEN_3541 : {{1'd0}, _GEN_2674}; // @[StoreSet.scala 562:37]
  wire [2:0] _GEN_3859 = REG ? _GEN_3561 : {{1'd0}, _GEN_2675}; // @[StoreSet.scala 562:37]
  wire [2:0] _GEN_3860 = REG ? _GEN_3581 : {{1'd0}, _GEN_2676}; // @[StoreSet.scala 562:37]
  wire [2:0] _GEN_3861 = REG ? _GEN_3601 : {{1'd0}, _GEN_2677}; // @[StoreSet.scala 562:37]
  wire [2:0] _GEN_3862 = REG ? _GEN_3621 : {{1'd0}, _GEN_2678}; // @[StoreSet.scala 562:37]
  wire [2:0] _GEN_3863 = REG ? _GEN_3641 : {{1'd0}, _GEN_2679}; // @[StoreSet.scala 562:37]
  wire [2:0] _GEN_3864 = REG ? _GEN_3661 : {{1'd0}, _GEN_2680}; // @[StoreSet.scala 562:37]
  wire [2:0] _GEN_3865 = REG ? _GEN_3681 : {{1'd0}, _GEN_2681}; // @[StoreSet.scala 562:37]
  wire [2:0] _GEN_3866 = REG ? _GEN_3701 : {{1'd0}, _GEN_2682}; // @[StoreSet.scala 562:37]
  wire [2:0] _GEN_3867 = REG ? _GEN_3721 : {{1'd0}, _GEN_2683}; // @[StoreSet.scala 562:37]
  wire [2:0] _GEN_3868 = REG ? _GEN_3741 : {{1'd0}, _GEN_2684}; // @[StoreSet.scala 562:37]
  wire [2:0] _GEN_3869 = REG ? _GEN_3761 : {{1'd0}, _GEN_2685}; // @[StoreSet.scala 562:37]
  wire [2:0] _GEN_3870 = REG ? _GEN_3781 : {{1'd0}, _GEN_2686}; // @[StoreSet.scala 562:37]
  wire [2:0] _GEN_3871 = REG ? _GEN_3801 : {{1'd0}, _GEN_2687}; // @[StoreSet.scala 562:37]
  wire [2:0] _GEN_3872 = REG ? _GEN_3821 : {{1'd0}, _GEN_2688}; // @[StoreSet.scala 562:37]
  wire [2:0] _GEN_3873 = REG ? _GEN_3841 : {{1'd0}, _GEN_2689}; // @[StoreSet.scala 562:37]
  assign io_dispatch_resp_0_bits_shouldWait = _io_dispatch_resp_0_bits_shouldWait_T_4 & ~io_csrCtrl_lvpred_disable |
    io_csrCtrl_no_spec_load; // @[StoreSet.scala 519:39]
  assign io_dispatch_resp_0_bits_robIdx_flag = 5'h1f == io_dispatch_req_0_bits_ssid & 2'h3 ==
    _io_dispatch_resp_0_bits_robIdx_T_1 ? robIdxVec_31_3_flag : _GEN_190; // @[StoreSet.scala 520:{37,37}]
  assign io_dispatch_resp_0_bits_robIdx_value = 5'h1f == io_dispatch_req_0_bits_ssid & 2'h3 ==
    _io_dispatch_resp_0_bits_robIdx_T_1 ? robIdxVec_31_3_value : _GEN_318; // @[StoreSet.scala 520:{37,37}]
  assign io_dispatch_resp_1_bits_shouldWait = _io_dispatch_resp_1_bits_shouldWait_T_4 & ~io_csrCtrl_lvpred_disable |
    io_csrCtrl_no_spec_load; // @[StoreSet.scala 519:39]
  assign io_dispatch_resp_1_bits_robIdx_flag = hitInDispatchBundleVec_1_0 ? io_dispatch_req_0_bits_robIdx_flag :
    _GEN_511; // @[StoreSet.scala 520:37 523:40 524:43]
  assign io_dispatch_resp_1_bits_robIdx_value = hitInDispatchBundleVec_1_0 ? io_dispatch_req_0_bits_robIdx_value :
    _GEN_639; // @[StoreSet.scala 520:37 523:40 524:43]
  always @(posedge clock) begin
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4382 & _GEN_5787) begin // @[StoreSet.scala 547:30]
        robIdxVec_0_0_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_0_0_flag <= _GEN_1986;
      end
    end else begin
      robIdxVec_0_0_flag <= _GEN_1986;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4382 & _GEN_5787) begin // @[StoreSet.scala 547:30]
        robIdxVec_0_0_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_0_0_value <= _GEN_2114;
      end
    end else begin
      robIdxVec_0_0_value <= _GEN_2114;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4382 & _GEN_5790) begin // @[StoreSet.scala 547:30]
        robIdxVec_0_1_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_0_1_flag <= _GEN_1987;
      end
    end else begin
      robIdxVec_0_1_flag <= _GEN_1987;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4382 & _GEN_5790) begin // @[StoreSet.scala 547:30]
        robIdxVec_0_1_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_0_1_value <= _GEN_2115;
      end
    end else begin
      robIdxVec_0_1_value <= _GEN_2115;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4382 & _GEN_5793) begin // @[StoreSet.scala 547:30]
        robIdxVec_0_2_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_0_2_flag <= _GEN_1988;
      end
    end else begin
      robIdxVec_0_2_flag <= _GEN_1988;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4382 & _GEN_5793) begin // @[StoreSet.scala 547:30]
        robIdxVec_0_2_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_0_2_value <= _GEN_2116;
      end
    end else begin
      robIdxVec_0_2_value <= _GEN_2116;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4382 & _GEN_5796) begin // @[StoreSet.scala 547:30]
        robIdxVec_0_3_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_0_3_flag <= _GEN_1989;
      end
    end else begin
      robIdxVec_0_3_flag <= _GEN_1989;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4382 & _GEN_5796) begin // @[StoreSet.scala 547:30]
        robIdxVec_0_3_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_0_3_value <= _GEN_2117;
      end
    end else begin
      robIdxVec_0_3_value <= _GEN_2117;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4388 & _GEN_5787) begin // @[StoreSet.scala 547:30]
        robIdxVec_1_0_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_1_0_flag <= _GEN_1990;
      end
    end else begin
      robIdxVec_1_0_flag <= _GEN_1990;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4388 & _GEN_5787) begin // @[StoreSet.scala 547:30]
        robIdxVec_1_0_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_1_0_value <= _GEN_2118;
      end
    end else begin
      robIdxVec_1_0_value <= _GEN_2118;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4388 & _GEN_5790) begin // @[StoreSet.scala 547:30]
        robIdxVec_1_1_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_1_1_flag <= _GEN_1991;
      end
    end else begin
      robIdxVec_1_1_flag <= _GEN_1991;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4388 & _GEN_5790) begin // @[StoreSet.scala 547:30]
        robIdxVec_1_1_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_1_1_value <= _GEN_2119;
      end
    end else begin
      robIdxVec_1_1_value <= _GEN_2119;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4388 & _GEN_5793) begin // @[StoreSet.scala 547:30]
        robIdxVec_1_2_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_1_2_flag <= _GEN_1992;
      end
    end else begin
      robIdxVec_1_2_flag <= _GEN_1992;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4388 & _GEN_5793) begin // @[StoreSet.scala 547:30]
        robIdxVec_1_2_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_1_2_value <= _GEN_2120;
      end
    end else begin
      robIdxVec_1_2_value <= _GEN_2120;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4388 & _GEN_5796) begin // @[StoreSet.scala 547:30]
        robIdxVec_1_3_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_1_3_flag <= _GEN_1993;
      end
    end else begin
      robIdxVec_1_3_flag <= _GEN_1993;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4388 & _GEN_5796) begin // @[StoreSet.scala 547:30]
        robIdxVec_1_3_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_1_3_value <= _GEN_2121;
      end
    end else begin
      robIdxVec_1_3_value <= _GEN_2121;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4396 & _GEN_5787) begin // @[StoreSet.scala 547:30]
        robIdxVec_2_0_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_2_0_flag <= _GEN_1994;
      end
    end else begin
      robIdxVec_2_0_flag <= _GEN_1994;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4396 & _GEN_5787) begin // @[StoreSet.scala 547:30]
        robIdxVec_2_0_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_2_0_value <= _GEN_2122;
      end
    end else begin
      robIdxVec_2_0_value <= _GEN_2122;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4396 & _GEN_5790) begin // @[StoreSet.scala 547:30]
        robIdxVec_2_1_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_2_1_flag <= _GEN_1995;
      end
    end else begin
      robIdxVec_2_1_flag <= _GEN_1995;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4396 & _GEN_5790) begin // @[StoreSet.scala 547:30]
        robIdxVec_2_1_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_2_1_value <= _GEN_2123;
      end
    end else begin
      robIdxVec_2_1_value <= _GEN_2123;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4396 & _GEN_5793) begin // @[StoreSet.scala 547:30]
        robIdxVec_2_2_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_2_2_flag <= _GEN_1996;
      end
    end else begin
      robIdxVec_2_2_flag <= _GEN_1996;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4396 & _GEN_5793) begin // @[StoreSet.scala 547:30]
        robIdxVec_2_2_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_2_2_value <= _GEN_2124;
      end
    end else begin
      robIdxVec_2_2_value <= _GEN_2124;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4396 & _GEN_5796) begin // @[StoreSet.scala 547:30]
        robIdxVec_2_3_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_2_3_flag <= _GEN_1997;
      end
    end else begin
      robIdxVec_2_3_flag <= _GEN_1997;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4396 & _GEN_5796) begin // @[StoreSet.scala 547:30]
        robIdxVec_2_3_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_2_3_value <= _GEN_2125;
      end
    end else begin
      robIdxVec_2_3_value <= _GEN_2125;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4404 & _GEN_5787) begin // @[StoreSet.scala 547:30]
        robIdxVec_3_0_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_3_0_flag <= _GEN_1998;
      end
    end else begin
      robIdxVec_3_0_flag <= _GEN_1998;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4404 & _GEN_5787) begin // @[StoreSet.scala 547:30]
        robIdxVec_3_0_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_3_0_value <= _GEN_2126;
      end
    end else begin
      robIdxVec_3_0_value <= _GEN_2126;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4404 & _GEN_5790) begin // @[StoreSet.scala 547:30]
        robIdxVec_3_1_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_3_1_flag <= _GEN_1999;
      end
    end else begin
      robIdxVec_3_1_flag <= _GEN_1999;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4404 & _GEN_5790) begin // @[StoreSet.scala 547:30]
        robIdxVec_3_1_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_3_1_value <= _GEN_2127;
      end
    end else begin
      robIdxVec_3_1_value <= _GEN_2127;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4404 & _GEN_5793) begin // @[StoreSet.scala 547:30]
        robIdxVec_3_2_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_3_2_flag <= _GEN_2000;
      end
    end else begin
      robIdxVec_3_2_flag <= _GEN_2000;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4404 & _GEN_5793) begin // @[StoreSet.scala 547:30]
        robIdxVec_3_2_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_3_2_value <= _GEN_2128;
      end
    end else begin
      robIdxVec_3_2_value <= _GEN_2128;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4404 & _GEN_5796) begin // @[StoreSet.scala 547:30]
        robIdxVec_3_3_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_3_3_flag <= _GEN_2001;
      end
    end else begin
      robIdxVec_3_3_flag <= _GEN_2001;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4404 & _GEN_5796) begin // @[StoreSet.scala 547:30]
        robIdxVec_3_3_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_3_3_value <= _GEN_2129;
      end
    end else begin
      robIdxVec_3_3_value <= _GEN_2129;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4412 & _GEN_5787) begin // @[StoreSet.scala 547:30]
        robIdxVec_4_0_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_4_0_flag <= _GEN_2002;
      end
    end else begin
      robIdxVec_4_0_flag <= _GEN_2002;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4412 & _GEN_5787) begin // @[StoreSet.scala 547:30]
        robIdxVec_4_0_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_4_0_value <= _GEN_2130;
      end
    end else begin
      robIdxVec_4_0_value <= _GEN_2130;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4412 & _GEN_5790) begin // @[StoreSet.scala 547:30]
        robIdxVec_4_1_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_4_1_flag <= _GEN_2003;
      end
    end else begin
      robIdxVec_4_1_flag <= _GEN_2003;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4412 & _GEN_5790) begin // @[StoreSet.scala 547:30]
        robIdxVec_4_1_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_4_1_value <= _GEN_2131;
      end
    end else begin
      robIdxVec_4_1_value <= _GEN_2131;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4412 & _GEN_5793) begin // @[StoreSet.scala 547:30]
        robIdxVec_4_2_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_4_2_flag <= _GEN_2004;
      end
    end else begin
      robIdxVec_4_2_flag <= _GEN_2004;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4412 & _GEN_5793) begin // @[StoreSet.scala 547:30]
        robIdxVec_4_2_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_4_2_value <= _GEN_2132;
      end
    end else begin
      robIdxVec_4_2_value <= _GEN_2132;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4412 & _GEN_5796) begin // @[StoreSet.scala 547:30]
        robIdxVec_4_3_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_4_3_flag <= _GEN_2005;
      end
    end else begin
      robIdxVec_4_3_flag <= _GEN_2005;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4412 & _GEN_5796) begin // @[StoreSet.scala 547:30]
        robIdxVec_4_3_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_4_3_value <= _GEN_2133;
      end
    end else begin
      robIdxVec_4_3_value <= _GEN_2133;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4420 & _GEN_5787) begin // @[StoreSet.scala 547:30]
        robIdxVec_5_0_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_5_0_flag <= _GEN_2006;
      end
    end else begin
      robIdxVec_5_0_flag <= _GEN_2006;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4420 & _GEN_5787) begin // @[StoreSet.scala 547:30]
        robIdxVec_5_0_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_5_0_value <= _GEN_2134;
      end
    end else begin
      robIdxVec_5_0_value <= _GEN_2134;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4420 & _GEN_5790) begin // @[StoreSet.scala 547:30]
        robIdxVec_5_1_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_5_1_flag <= _GEN_2007;
      end
    end else begin
      robIdxVec_5_1_flag <= _GEN_2007;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4420 & _GEN_5790) begin // @[StoreSet.scala 547:30]
        robIdxVec_5_1_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_5_1_value <= _GEN_2135;
      end
    end else begin
      robIdxVec_5_1_value <= _GEN_2135;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4420 & _GEN_5793) begin // @[StoreSet.scala 547:30]
        robIdxVec_5_2_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_5_2_flag <= _GEN_2008;
      end
    end else begin
      robIdxVec_5_2_flag <= _GEN_2008;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4420 & _GEN_5793) begin // @[StoreSet.scala 547:30]
        robIdxVec_5_2_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_5_2_value <= _GEN_2136;
      end
    end else begin
      robIdxVec_5_2_value <= _GEN_2136;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4420 & _GEN_5796) begin // @[StoreSet.scala 547:30]
        robIdxVec_5_3_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_5_3_flag <= _GEN_2009;
      end
    end else begin
      robIdxVec_5_3_flag <= _GEN_2009;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4420 & _GEN_5796) begin // @[StoreSet.scala 547:30]
        robIdxVec_5_3_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_5_3_value <= _GEN_2137;
      end
    end else begin
      robIdxVec_5_3_value <= _GEN_2137;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4428 & _GEN_5787) begin // @[StoreSet.scala 547:30]
        robIdxVec_6_0_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_6_0_flag <= _GEN_2010;
      end
    end else begin
      robIdxVec_6_0_flag <= _GEN_2010;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4428 & _GEN_5787) begin // @[StoreSet.scala 547:30]
        robIdxVec_6_0_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_6_0_value <= _GEN_2138;
      end
    end else begin
      robIdxVec_6_0_value <= _GEN_2138;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4428 & _GEN_5790) begin // @[StoreSet.scala 547:30]
        robIdxVec_6_1_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_6_1_flag <= _GEN_2011;
      end
    end else begin
      robIdxVec_6_1_flag <= _GEN_2011;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4428 & _GEN_5790) begin // @[StoreSet.scala 547:30]
        robIdxVec_6_1_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_6_1_value <= _GEN_2139;
      end
    end else begin
      robIdxVec_6_1_value <= _GEN_2139;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4428 & _GEN_5793) begin // @[StoreSet.scala 547:30]
        robIdxVec_6_2_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_6_2_flag <= _GEN_2012;
      end
    end else begin
      robIdxVec_6_2_flag <= _GEN_2012;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4428 & _GEN_5793) begin // @[StoreSet.scala 547:30]
        robIdxVec_6_2_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_6_2_value <= _GEN_2140;
      end
    end else begin
      robIdxVec_6_2_value <= _GEN_2140;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4428 & _GEN_5796) begin // @[StoreSet.scala 547:30]
        robIdxVec_6_3_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_6_3_flag <= _GEN_2013;
      end
    end else begin
      robIdxVec_6_3_flag <= _GEN_2013;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4428 & _GEN_5796) begin // @[StoreSet.scala 547:30]
        robIdxVec_6_3_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_6_3_value <= _GEN_2141;
      end
    end else begin
      robIdxVec_6_3_value <= _GEN_2141;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4436 & _GEN_5787) begin // @[StoreSet.scala 547:30]
        robIdxVec_7_0_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_7_0_flag <= _GEN_2014;
      end
    end else begin
      robIdxVec_7_0_flag <= _GEN_2014;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4436 & _GEN_5787) begin // @[StoreSet.scala 547:30]
        robIdxVec_7_0_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_7_0_value <= _GEN_2142;
      end
    end else begin
      robIdxVec_7_0_value <= _GEN_2142;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4436 & _GEN_5790) begin // @[StoreSet.scala 547:30]
        robIdxVec_7_1_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_7_1_flag <= _GEN_2015;
      end
    end else begin
      robIdxVec_7_1_flag <= _GEN_2015;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4436 & _GEN_5790) begin // @[StoreSet.scala 547:30]
        robIdxVec_7_1_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_7_1_value <= _GEN_2143;
      end
    end else begin
      robIdxVec_7_1_value <= _GEN_2143;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4436 & _GEN_5793) begin // @[StoreSet.scala 547:30]
        robIdxVec_7_2_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_7_2_flag <= _GEN_2016;
      end
    end else begin
      robIdxVec_7_2_flag <= _GEN_2016;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4436 & _GEN_5793) begin // @[StoreSet.scala 547:30]
        robIdxVec_7_2_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_7_2_value <= _GEN_2144;
      end
    end else begin
      robIdxVec_7_2_value <= _GEN_2144;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4436 & _GEN_5796) begin // @[StoreSet.scala 547:30]
        robIdxVec_7_3_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_7_3_flag <= _GEN_2017;
      end
    end else begin
      robIdxVec_7_3_flag <= _GEN_2017;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4436 & _GEN_5796) begin // @[StoreSet.scala 547:30]
        robIdxVec_7_3_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_7_3_value <= _GEN_2145;
      end
    end else begin
      robIdxVec_7_3_value <= _GEN_2145;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4444 & _GEN_5787) begin // @[StoreSet.scala 547:30]
        robIdxVec_8_0_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_8_0_flag <= _GEN_2018;
      end
    end else begin
      robIdxVec_8_0_flag <= _GEN_2018;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4444 & _GEN_5787) begin // @[StoreSet.scala 547:30]
        robIdxVec_8_0_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_8_0_value <= _GEN_2146;
      end
    end else begin
      robIdxVec_8_0_value <= _GEN_2146;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4444 & _GEN_5790) begin // @[StoreSet.scala 547:30]
        robIdxVec_8_1_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_8_1_flag <= _GEN_2019;
      end
    end else begin
      robIdxVec_8_1_flag <= _GEN_2019;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4444 & _GEN_5790) begin // @[StoreSet.scala 547:30]
        robIdxVec_8_1_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_8_1_value <= _GEN_2147;
      end
    end else begin
      robIdxVec_8_1_value <= _GEN_2147;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4444 & _GEN_5793) begin // @[StoreSet.scala 547:30]
        robIdxVec_8_2_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_8_2_flag <= _GEN_2020;
      end
    end else begin
      robIdxVec_8_2_flag <= _GEN_2020;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4444 & _GEN_5793) begin // @[StoreSet.scala 547:30]
        robIdxVec_8_2_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_8_2_value <= _GEN_2148;
      end
    end else begin
      robIdxVec_8_2_value <= _GEN_2148;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4444 & _GEN_5796) begin // @[StoreSet.scala 547:30]
        robIdxVec_8_3_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_8_3_flag <= _GEN_2021;
      end
    end else begin
      robIdxVec_8_3_flag <= _GEN_2021;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4444 & _GEN_5796) begin // @[StoreSet.scala 547:30]
        robIdxVec_8_3_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_8_3_value <= _GEN_2149;
      end
    end else begin
      robIdxVec_8_3_value <= _GEN_2149;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4452 & _GEN_5787) begin // @[StoreSet.scala 547:30]
        robIdxVec_9_0_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_9_0_flag <= _GEN_2022;
      end
    end else begin
      robIdxVec_9_0_flag <= _GEN_2022;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4452 & _GEN_5787) begin // @[StoreSet.scala 547:30]
        robIdxVec_9_0_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_9_0_value <= _GEN_2150;
      end
    end else begin
      robIdxVec_9_0_value <= _GEN_2150;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4452 & _GEN_5790) begin // @[StoreSet.scala 547:30]
        robIdxVec_9_1_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_9_1_flag <= _GEN_2023;
      end
    end else begin
      robIdxVec_9_1_flag <= _GEN_2023;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4452 & _GEN_5790) begin // @[StoreSet.scala 547:30]
        robIdxVec_9_1_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_9_1_value <= _GEN_2151;
      end
    end else begin
      robIdxVec_9_1_value <= _GEN_2151;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4452 & _GEN_5793) begin // @[StoreSet.scala 547:30]
        robIdxVec_9_2_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_9_2_flag <= _GEN_2024;
      end
    end else begin
      robIdxVec_9_2_flag <= _GEN_2024;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4452 & _GEN_5793) begin // @[StoreSet.scala 547:30]
        robIdxVec_9_2_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_9_2_value <= _GEN_2152;
      end
    end else begin
      robIdxVec_9_2_value <= _GEN_2152;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4452 & _GEN_5796) begin // @[StoreSet.scala 547:30]
        robIdxVec_9_3_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_9_3_flag <= _GEN_2025;
      end
    end else begin
      robIdxVec_9_3_flag <= _GEN_2025;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4452 & _GEN_5796) begin // @[StoreSet.scala 547:30]
        robIdxVec_9_3_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_9_3_value <= _GEN_2153;
      end
    end else begin
      robIdxVec_9_3_value <= _GEN_2153;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4460 & _GEN_5787) begin // @[StoreSet.scala 547:30]
        robIdxVec_10_0_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_10_0_flag <= _GEN_2026;
      end
    end else begin
      robIdxVec_10_0_flag <= _GEN_2026;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4460 & _GEN_5787) begin // @[StoreSet.scala 547:30]
        robIdxVec_10_0_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_10_0_value <= _GEN_2154;
      end
    end else begin
      robIdxVec_10_0_value <= _GEN_2154;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4460 & _GEN_5790) begin // @[StoreSet.scala 547:30]
        robIdxVec_10_1_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_10_1_flag <= _GEN_2027;
      end
    end else begin
      robIdxVec_10_1_flag <= _GEN_2027;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4460 & _GEN_5790) begin // @[StoreSet.scala 547:30]
        robIdxVec_10_1_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_10_1_value <= _GEN_2155;
      end
    end else begin
      robIdxVec_10_1_value <= _GEN_2155;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4460 & _GEN_5793) begin // @[StoreSet.scala 547:30]
        robIdxVec_10_2_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_10_2_flag <= _GEN_2028;
      end
    end else begin
      robIdxVec_10_2_flag <= _GEN_2028;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4460 & _GEN_5793) begin // @[StoreSet.scala 547:30]
        robIdxVec_10_2_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_10_2_value <= _GEN_2156;
      end
    end else begin
      robIdxVec_10_2_value <= _GEN_2156;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4460 & _GEN_5796) begin // @[StoreSet.scala 547:30]
        robIdxVec_10_3_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_10_3_flag <= _GEN_2029;
      end
    end else begin
      robIdxVec_10_3_flag <= _GEN_2029;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4460 & _GEN_5796) begin // @[StoreSet.scala 547:30]
        robIdxVec_10_3_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_10_3_value <= _GEN_2157;
      end
    end else begin
      robIdxVec_10_3_value <= _GEN_2157;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4468 & _GEN_5787) begin // @[StoreSet.scala 547:30]
        robIdxVec_11_0_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_11_0_flag <= _GEN_2030;
      end
    end else begin
      robIdxVec_11_0_flag <= _GEN_2030;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4468 & _GEN_5787) begin // @[StoreSet.scala 547:30]
        robIdxVec_11_0_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_11_0_value <= _GEN_2158;
      end
    end else begin
      robIdxVec_11_0_value <= _GEN_2158;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4468 & _GEN_5790) begin // @[StoreSet.scala 547:30]
        robIdxVec_11_1_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_11_1_flag <= _GEN_2031;
      end
    end else begin
      robIdxVec_11_1_flag <= _GEN_2031;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4468 & _GEN_5790) begin // @[StoreSet.scala 547:30]
        robIdxVec_11_1_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_11_1_value <= _GEN_2159;
      end
    end else begin
      robIdxVec_11_1_value <= _GEN_2159;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4468 & _GEN_5793) begin // @[StoreSet.scala 547:30]
        robIdxVec_11_2_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_11_2_flag <= _GEN_2032;
      end
    end else begin
      robIdxVec_11_2_flag <= _GEN_2032;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4468 & _GEN_5793) begin // @[StoreSet.scala 547:30]
        robIdxVec_11_2_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_11_2_value <= _GEN_2160;
      end
    end else begin
      robIdxVec_11_2_value <= _GEN_2160;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4468 & _GEN_5796) begin // @[StoreSet.scala 547:30]
        robIdxVec_11_3_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_11_3_flag <= _GEN_2033;
      end
    end else begin
      robIdxVec_11_3_flag <= _GEN_2033;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4468 & _GEN_5796) begin // @[StoreSet.scala 547:30]
        robIdxVec_11_3_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_11_3_value <= _GEN_2161;
      end
    end else begin
      robIdxVec_11_3_value <= _GEN_2161;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4476 & _GEN_5787) begin // @[StoreSet.scala 547:30]
        robIdxVec_12_0_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_12_0_flag <= _GEN_2034;
      end
    end else begin
      robIdxVec_12_0_flag <= _GEN_2034;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4476 & _GEN_5787) begin // @[StoreSet.scala 547:30]
        robIdxVec_12_0_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_12_0_value <= _GEN_2162;
      end
    end else begin
      robIdxVec_12_0_value <= _GEN_2162;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4476 & _GEN_5790) begin // @[StoreSet.scala 547:30]
        robIdxVec_12_1_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_12_1_flag <= _GEN_2035;
      end
    end else begin
      robIdxVec_12_1_flag <= _GEN_2035;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4476 & _GEN_5790) begin // @[StoreSet.scala 547:30]
        robIdxVec_12_1_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_12_1_value <= _GEN_2163;
      end
    end else begin
      robIdxVec_12_1_value <= _GEN_2163;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4476 & _GEN_5793) begin // @[StoreSet.scala 547:30]
        robIdxVec_12_2_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_12_2_flag <= _GEN_2036;
      end
    end else begin
      robIdxVec_12_2_flag <= _GEN_2036;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4476 & _GEN_5793) begin // @[StoreSet.scala 547:30]
        robIdxVec_12_2_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_12_2_value <= _GEN_2164;
      end
    end else begin
      robIdxVec_12_2_value <= _GEN_2164;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4476 & _GEN_5796) begin // @[StoreSet.scala 547:30]
        robIdxVec_12_3_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_12_3_flag <= _GEN_2037;
      end
    end else begin
      robIdxVec_12_3_flag <= _GEN_2037;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4476 & _GEN_5796) begin // @[StoreSet.scala 547:30]
        robIdxVec_12_3_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_12_3_value <= _GEN_2165;
      end
    end else begin
      robIdxVec_12_3_value <= _GEN_2165;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4484 & _GEN_5787) begin // @[StoreSet.scala 547:30]
        robIdxVec_13_0_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_13_0_flag <= _GEN_2038;
      end
    end else begin
      robIdxVec_13_0_flag <= _GEN_2038;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4484 & _GEN_5787) begin // @[StoreSet.scala 547:30]
        robIdxVec_13_0_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_13_0_value <= _GEN_2166;
      end
    end else begin
      robIdxVec_13_0_value <= _GEN_2166;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4484 & _GEN_5790) begin // @[StoreSet.scala 547:30]
        robIdxVec_13_1_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_13_1_flag <= _GEN_2039;
      end
    end else begin
      robIdxVec_13_1_flag <= _GEN_2039;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4484 & _GEN_5790) begin // @[StoreSet.scala 547:30]
        robIdxVec_13_1_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_13_1_value <= _GEN_2167;
      end
    end else begin
      robIdxVec_13_1_value <= _GEN_2167;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4484 & _GEN_5793) begin // @[StoreSet.scala 547:30]
        robIdxVec_13_2_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_13_2_flag <= _GEN_2040;
      end
    end else begin
      robIdxVec_13_2_flag <= _GEN_2040;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4484 & _GEN_5793) begin // @[StoreSet.scala 547:30]
        robIdxVec_13_2_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_13_2_value <= _GEN_2168;
      end
    end else begin
      robIdxVec_13_2_value <= _GEN_2168;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4484 & _GEN_5796) begin // @[StoreSet.scala 547:30]
        robIdxVec_13_3_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_13_3_flag <= _GEN_2041;
      end
    end else begin
      robIdxVec_13_3_flag <= _GEN_2041;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4484 & _GEN_5796) begin // @[StoreSet.scala 547:30]
        robIdxVec_13_3_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_13_3_value <= _GEN_2169;
      end
    end else begin
      robIdxVec_13_3_value <= _GEN_2169;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4492 & _GEN_5787) begin // @[StoreSet.scala 547:30]
        robIdxVec_14_0_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_14_0_flag <= _GEN_2042;
      end
    end else begin
      robIdxVec_14_0_flag <= _GEN_2042;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4492 & _GEN_5787) begin // @[StoreSet.scala 547:30]
        robIdxVec_14_0_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_14_0_value <= _GEN_2170;
      end
    end else begin
      robIdxVec_14_0_value <= _GEN_2170;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4492 & _GEN_5790) begin // @[StoreSet.scala 547:30]
        robIdxVec_14_1_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_14_1_flag <= _GEN_2043;
      end
    end else begin
      robIdxVec_14_1_flag <= _GEN_2043;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4492 & _GEN_5790) begin // @[StoreSet.scala 547:30]
        robIdxVec_14_1_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_14_1_value <= _GEN_2171;
      end
    end else begin
      robIdxVec_14_1_value <= _GEN_2171;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4492 & _GEN_5793) begin // @[StoreSet.scala 547:30]
        robIdxVec_14_2_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_14_2_flag <= _GEN_2044;
      end
    end else begin
      robIdxVec_14_2_flag <= _GEN_2044;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4492 & _GEN_5793) begin // @[StoreSet.scala 547:30]
        robIdxVec_14_2_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_14_2_value <= _GEN_2172;
      end
    end else begin
      robIdxVec_14_2_value <= _GEN_2172;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4492 & _GEN_5796) begin // @[StoreSet.scala 547:30]
        robIdxVec_14_3_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_14_3_flag <= _GEN_2045;
      end
    end else begin
      robIdxVec_14_3_flag <= _GEN_2045;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4492 & _GEN_5796) begin // @[StoreSet.scala 547:30]
        robIdxVec_14_3_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_14_3_value <= _GEN_2173;
      end
    end else begin
      robIdxVec_14_3_value <= _GEN_2173;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4500 & _GEN_5787) begin // @[StoreSet.scala 547:30]
        robIdxVec_15_0_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_15_0_flag <= _GEN_2046;
      end
    end else begin
      robIdxVec_15_0_flag <= _GEN_2046;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4500 & _GEN_5787) begin // @[StoreSet.scala 547:30]
        robIdxVec_15_0_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_15_0_value <= _GEN_2174;
      end
    end else begin
      robIdxVec_15_0_value <= _GEN_2174;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4500 & _GEN_5790) begin // @[StoreSet.scala 547:30]
        robIdxVec_15_1_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_15_1_flag <= _GEN_2047;
      end
    end else begin
      robIdxVec_15_1_flag <= _GEN_2047;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4500 & _GEN_5790) begin // @[StoreSet.scala 547:30]
        robIdxVec_15_1_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_15_1_value <= _GEN_2175;
      end
    end else begin
      robIdxVec_15_1_value <= _GEN_2175;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4500 & _GEN_5793) begin // @[StoreSet.scala 547:30]
        robIdxVec_15_2_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_15_2_flag <= _GEN_2048;
      end
    end else begin
      robIdxVec_15_2_flag <= _GEN_2048;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4500 & _GEN_5793) begin // @[StoreSet.scala 547:30]
        robIdxVec_15_2_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_15_2_value <= _GEN_2176;
      end
    end else begin
      robIdxVec_15_2_value <= _GEN_2176;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4500 & _GEN_5796) begin // @[StoreSet.scala 547:30]
        robIdxVec_15_3_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_15_3_flag <= _GEN_2049;
      end
    end else begin
      robIdxVec_15_3_flag <= _GEN_2049;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4500 & _GEN_5796) begin // @[StoreSet.scala 547:30]
        robIdxVec_15_3_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_15_3_value <= _GEN_2177;
      end
    end else begin
      robIdxVec_15_3_value <= _GEN_2177;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4508 & _GEN_5787) begin // @[StoreSet.scala 547:30]
        robIdxVec_16_0_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_16_0_flag <= _GEN_2050;
      end
    end else begin
      robIdxVec_16_0_flag <= _GEN_2050;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4508 & _GEN_5787) begin // @[StoreSet.scala 547:30]
        robIdxVec_16_0_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_16_0_value <= _GEN_2178;
      end
    end else begin
      robIdxVec_16_0_value <= _GEN_2178;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4508 & _GEN_5790) begin // @[StoreSet.scala 547:30]
        robIdxVec_16_1_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_16_1_flag <= _GEN_2051;
      end
    end else begin
      robIdxVec_16_1_flag <= _GEN_2051;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4508 & _GEN_5790) begin // @[StoreSet.scala 547:30]
        robIdxVec_16_1_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_16_1_value <= _GEN_2179;
      end
    end else begin
      robIdxVec_16_1_value <= _GEN_2179;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4508 & _GEN_5793) begin // @[StoreSet.scala 547:30]
        robIdxVec_16_2_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_16_2_flag <= _GEN_2052;
      end
    end else begin
      robIdxVec_16_2_flag <= _GEN_2052;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4508 & _GEN_5793) begin // @[StoreSet.scala 547:30]
        robIdxVec_16_2_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_16_2_value <= _GEN_2180;
      end
    end else begin
      robIdxVec_16_2_value <= _GEN_2180;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4508 & _GEN_5796) begin // @[StoreSet.scala 547:30]
        robIdxVec_16_3_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_16_3_flag <= _GEN_2053;
      end
    end else begin
      robIdxVec_16_3_flag <= _GEN_2053;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4508 & _GEN_5796) begin // @[StoreSet.scala 547:30]
        robIdxVec_16_3_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_16_3_value <= _GEN_2181;
      end
    end else begin
      robIdxVec_16_3_value <= _GEN_2181;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4516 & _GEN_5787) begin // @[StoreSet.scala 547:30]
        robIdxVec_17_0_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_17_0_flag <= _GEN_2054;
      end
    end else begin
      robIdxVec_17_0_flag <= _GEN_2054;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4516 & _GEN_5787) begin // @[StoreSet.scala 547:30]
        robIdxVec_17_0_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_17_0_value <= _GEN_2182;
      end
    end else begin
      robIdxVec_17_0_value <= _GEN_2182;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4516 & _GEN_5790) begin // @[StoreSet.scala 547:30]
        robIdxVec_17_1_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_17_1_flag <= _GEN_2055;
      end
    end else begin
      robIdxVec_17_1_flag <= _GEN_2055;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4516 & _GEN_5790) begin // @[StoreSet.scala 547:30]
        robIdxVec_17_1_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_17_1_value <= _GEN_2183;
      end
    end else begin
      robIdxVec_17_1_value <= _GEN_2183;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4516 & _GEN_5793) begin // @[StoreSet.scala 547:30]
        robIdxVec_17_2_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_17_2_flag <= _GEN_2056;
      end
    end else begin
      robIdxVec_17_2_flag <= _GEN_2056;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4516 & _GEN_5793) begin // @[StoreSet.scala 547:30]
        robIdxVec_17_2_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_17_2_value <= _GEN_2184;
      end
    end else begin
      robIdxVec_17_2_value <= _GEN_2184;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4516 & _GEN_5796) begin // @[StoreSet.scala 547:30]
        robIdxVec_17_3_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_17_3_flag <= _GEN_2057;
      end
    end else begin
      robIdxVec_17_3_flag <= _GEN_2057;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4516 & _GEN_5796) begin // @[StoreSet.scala 547:30]
        robIdxVec_17_3_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_17_3_value <= _GEN_2185;
      end
    end else begin
      robIdxVec_17_3_value <= _GEN_2185;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4524 & _GEN_5787) begin // @[StoreSet.scala 547:30]
        robIdxVec_18_0_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_18_0_flag <= _GEN_2058;
      end
    end else begin
      robIdxVec_18_0_flag <= _GEN_2058;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4524 & _GEN_5787) begin // @[StoreSet.scala 547:30]
        robIdxVec_18_0_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_18_0_value <= _GEN_2186;
      end
    end else begin
      robIdxVec_18_0_value <= _GEN_2186;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4524 & _GEN_5790) begin // @[StoreSet.scala 547:30]
        robIdxVec_18_1_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_18_1_flag <= _GEN_2059;
      end
    end else begin
      robIdxVec_18_1_flag <= _GEN_2059;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4524 & _GEN_5790) begin // @[StoreSet.scala 547:30]
        robIdxVec_18_1_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_18_1_value <= _GEN_2187;
      end
    end else begin
      robIdxVec_18_1_value <= _GEN_2187;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4524 & _GEN_5793) begin // @[StoreSet.scala 547:30]
        robIdxVec_18_2_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_18_2_flag <= _GEN_2060;
      end
    end else begin
      robIdxVec_18_2_flag <= _GEN_2060;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4524 & _GEN_5793) begin // @[StoreSet.scala 547:30]
        robIdxVec_18_2_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_18_2_value <= _GEN_2188;
      end
    end else begin
      robIdxVec_18_2_value <= _GEN_2188;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4524 & _GEN_5796) begin // @[StoreSet.scala 547:30]
        robIdxVec_18_3_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_18_3_flag <= _GEN_2061;
      end
    end else begin
      robIdxVec_18_3_flag <= _GEN_2061;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4524 & _GEN_5796) begin // @[StoreSet.scala 547:30]
        robIdxVec_18_3_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_18_3_value <= _GEN_2189;
      end
    end else begin
      robIdxVec_18_3_value <= _GEN_2189;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4532 & _GEN_5787) begin // @[StoreSet.scala 547:30]
        robIdxVec_19_0_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_19_0_flag <= _GEN_2062;
      end
    end else begin
      robIdxVec_19_0_flag <= _GEN_2062;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4532 & _GEN_5787) begin // @[StoreSet.scala 547:30]
        robIdxVec_19_0_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_19_0_value <= _GEN_2190;
      end
    end else begin
      robIdxVec_19_0_value <= _GEN_2190;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4532 & _GEN_5790) begin // @[StoreSet.scala 547:30]
        robIdxVec_19_1_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_19_1_flag <= _GEN_2063;
      end
    end else begin
      robIdxVec_19_1_flag <= _GEN_2063;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4532 & _GEN_5790) begin // @[StoreSet.scala 547:30]
        robIdxVec_19_1_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_19_1_value <= _GEN_2191;
      end
    end else begin
      robIdxVec_19_1_value <= _GEN_2191;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4532 & _GEN_5793) begin // @[StoreSet.scala 547:30]
        robIdxVec_19_2_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_19_2_flag <= _GEN_2064;
      end
    end else begin
      robIdxVec_19_2_flag <= _GEN_2064;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4532 & _GEN_5793) begin // @[StoreSet.scala 547:30]
        robIdxVec_19_2_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_19_2_value <= _GEN_2192;
      end
    end else begin
      robIdxVec_19_2_value <= _GEN_2192;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4532 & _GEN_5796) begin // @[StoreSet.scala 547:30]
        robIdxVec_19_3_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_19_3_flag <= _GEN_2065;
      end
    end else begin
      robIdxVec_19_3_flag <= _GEN_2065;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4532 & _GEN_5796) begin // @[StoreSet.scala 547:30]
        robIdxVec_19_3_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_19_3_value <= _GEN_2193;
      end
    end else begin
      robIdxVec_19_3_value <= _GEN_2193;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4540 & _GEN_5787) begin // @[StoreSet.scala 547:30]
        robIdxVec_20_0_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_20_0_flag <= _GEN_2066;
      end
    end else begin
      robIdxVec_20_0_flag <= _GEN_2066;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4540 & _GEN_5787) begin // @[StoreSet.scala 547:30]
        robIdxVec_20_0_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_20_0_value <= _GEN_2194;
      end
    end else begin
      robIdxVec_20_0_value <= _GEN_2194;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4540 & _GEN_5790) begin // @[StoreSet.scala 547:30]
        robIdxVec_20_1_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_20_1_flag <= _GEN_2067;
      end
    end else begin
      robIdxVec_20_1_flag <= _GEN_2067;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4540 & _GEN_5790) begin // @[StoreSet.scala 547:30]
        robIdxVec_20_1_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_20_1_value <= _GEN_2195;
      end
    end else begin
      robIdxVec_20_1_value <= _GEN_2195;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4540 & _GEN_5793) begin // @[StoreSet.scala 547:30]
        robIdxVec_20_2_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_20_2_flag <= _GEN_2068;
      end
    end else begin
      robIdxVec_20_2_flag <= _GEN_2068;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4540 & _GEN_5793) begin // @[StoreSet.scala 547:30]
        robIdxVec_20_2_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_20_2_value <= _GEN_2196;
      end
    end else begin
      robIdxVec_20_2_value <= _GEN_2196;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4540 & _GEN_5796) begin // @[StoreSet.scala 547:30]
        robIdxVec_20_3_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_20_3_flag <= _GEN_2069;
      end
    end else begin
      robIdxVec_20_3_flag <= _GEN_2069;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4540 & _GEN_5796) begin // @[StoreSet.scala 547:30]
        robIdxVec_20_3_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_20_3_value <= _GEN_2197;
      end
    end else begin
      robIdxVec_20_3_value <= _GEN_2197;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4548 & _GEN_5787) begin // @[StoreSet.scala 547:30]
        robIdxVec_21_0_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_21_0_flag <= _GEN_2070;
      end
    end else begin
      robIdxVec_21_0_flag <= _GEN_2070;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4548 & _GEN_5787) begin // @[StoreSet.scala 547:30]
        robIdxVec_21_0_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_21_0_value <= _GEN_2198;
      end
    end else begin
      robIdxVec_21_0_value <= _GEN_2198;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4548 & _GEN_5790) begin // @[StoreSet.scala 547:30]
        robIdxVec_21_1_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_21_1_flag <= _GEN_2071;
      end
    end else begin
      robIdxVec_21_1_flag <= _GEN_2071;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4548 & _GEN_5790) begin // @[StoreSet.scala 547:30]
        robIdxVec_21_1_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_21_1_value <= _GEN_2199;
      end
    end else begin
      robIdxVec_21_1_value <= _GEN_2199;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4548 & _GEN_5793) begin // @[StoreSet.scala 547:30]
        robIdxVec_21_2_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_21_2_flag <= _GEN_2072;
      end
    end else begin
      robIdxVec_21_2_flag <= _GEN_2072;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4548 & _GEN_5793) begin // @[StoreSet.scala 547:30]
        robIdxVec_21_2_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_21_2_value <= _GEN_2200;
      end
    end else begin
      robIdxVec_21_2_value <= _GEN_2200;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4548 & _GEN_5796) begin // @[StoreSet.scala 547:30]
        robIdxVec_21_3_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_21_3_flag <= _GEN_2073;
      end
    end else begin
      robIdxVec_21_3_flag <= _GEN_2073;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4548 & _GEN_5796) begin // @[StoreSet.scala 547:30]
        robIdxVec_21_3_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_21_3_value <= _GEN_2201;
      end
    end else begin
      robIdxVec_21_3_value <= _GEN_2201;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4556 & _GEN_5787) begin // @[StoreSet.scala 547:30]
        robIdxVec_22_0_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_22_0_flag <= _GEN_2074;
      end
    end else begin
      robIdxVec_22_0_flag <= _GEN_2074;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4556 & _GEN_5787) begin // @[StoreSet.scala 547:30]
        robIdxVec_22_0_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_22_0_value <= _GEN_2202;
      end
    end else begin
      robIdxVec_22_0_value <= _GEN_2202;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4556 & _GEN_5790) begin // @[StoreSet.scala 547:30]
        robIdxVec_22_1_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_22_1_flag <= _GEN_2075;
      end
    end else begin
      robIdxVec_22_1_flag <= _GEN_2075;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4556 & _GEN_5790) begin // @[StoreSet.scala 547:30]
        robIdxVec_22_1_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_22_1_value <= _GEN_2203;
      end
    end else begin
      robIdxVec_22_1_value <= _GEN_2203;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4556 & _GEN_5793) begin // @[StoreSet.scala 547:30]
        robIdxVec_22_2_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_22_2_flag <= _GEN_2076;
      end
    end else begin
      robIdxVec_22_2_flag <= _GEN_2076;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4556 & _GEN_5793) begin // @[StoreSet.scala 547:30]
        robIdxVec_22_2_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_22_2_value <= _GEN_2204;
      end
    end else begin
      robIdxVec_22_2_value <= _GEN_2204;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4556 & _GEN_5796) begin // @[StoreSet.scala 547:30]
        robIdxVec_22_3_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_22_3_flag <= _GEN_2077;
      end
    end else begin
      robIdxVec_22_3_flag <= _GEN_2077;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4556 & _GEN_5796) begin // @[StoreSet.scala 547:30]
        robIdxVec_22_3_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_22_3_value <= _GEN_2205;
      end
    end else begin
      robIdxVec_22_3_value <= _GEN_2205;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4564 & _GEN_5787) begin // @[StoreSet.scala 547:30]
        robIdxVec_23_0_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_23_0_flag <= _GEN_2078;
      end
    end else begin
      robIdxVec_23_0_flag <= _GEN_2078;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4564 & _GEN_5787) begin // @[StoreSet.scala 547:30]
        robIdxVec_23_0_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_23_0_value <= _GEN_2206;
      end
    end else begin
      robIdxVec_23_0_value <= _GEN_2206;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4564 & _GEN_5790) begin // @[StoreSet.scala 547:30]
        robIdxVec_23_1_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_23_1_flag <= _GEN_2079;
      end
    end else begin
      robIdxVec_23_1_flag <= _GEN_2079;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4564 & _GEN_5790) begin // @[StoreSet.scala 547:30]
        robIdxVec_23_1_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_23_1_value <= _GEN_2207;
      end
    end else begin
      robIdxVec_23_1_value <= _GEN_2207;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4564 & _GEN_5793) begin // @[StoreSet.scala 547:30]
        robIdxVec_23_2_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_23_2_flag <= _GEN_2080;
      end
    end else begin
      robIdxVec_23_2_flag <= _GEN_2080;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4564 & _GEN_5793) begin // @[StoreSet.scala 547:30]
        robIdxVec_23_2_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_23_2_value <= _GEN_2208;
      end
    end else begin
      robIdxVec_23_2_value <= _GEN_2208;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4564 & _GEN_5796) begin // @[StoreSet.scala 547:30]
        robIdxVec_23_3_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_23_3_flag <= _GEN_2081;
      end
    end else begin
      robIdxVec_23_3_flag <= _GEN_2081;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4564 & _GEN_5796) begin // @[StoreSet.scala 547:30]
        robIdxVec_23_3_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_23_3_value <= _GEN_2209;
      end
    end else begin
      robIdxVec_23_3_value <= _GEN_2209;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4572 & _GEN_5787) begin // @[StoreSet.scala 547:30]
        robIdxVec_24_0_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_24_0_flag <= _GEN_2082;
      end
    end else begin
      robIdxVec_24_0_flag <= _GEN_2082;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4572 & _GEN_5787) begin // @[StoreSet.scala 547:30]
        robIdxVec_24_0_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_24_0_value <= _GEN_2210;
      end
    end else begin
      robIdxVec_24_0_value <= _GEN_2210;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4572 & _GEN_5790) begin // @[StoreSet.scala 547:30]
        robIdxVec_24_1_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_24_1_flag <= _GEN_2083;
      end
    end else begin
      robIdxVec_24_1_flag <= _GEN_2083;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4572 & _GEN_5790) begin // @[StoreSet.scala 547:30]
        robIdxVec_24_1_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_24_1_value <= _GEN_2211;
      end
    end else begin
      robIdxVec_24_1_value <= _GEN_2211;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4572 & _GEN_5793) begin // @[StoreSet.scala 547:30]
        robIdxVec_24_2_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_24_2_flag <= _GEN_2084;
      end
    end else begin
      robIdxVec_24_2_flag <= _GEN_2084;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4572 & _GEN_5793) begin // @[StoreSet.scala 547:30]
        robIdxVec_24_2_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_24_2_value <= _GEN_2212;
      end
    end else begin
      robIdxVec_24_2_value <= _GEN_2212;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4572 & _GEN_5796) begin // @[StoreSet.scala 547:30]
        robIdxVec_24_3_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_24_3_flag <= _GEN_2085;
      end
    end else begin
      robIdxVec_24_3_flag <= _GEN_2085;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4572 & _GEN_5796) begin // @[StoreSet.scala 547:30]
        robIdxVec_24_3_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_24_3_value <= _GEN_2213;
      end
    end else begin
      robIdxVec_24_3_value <= _GEN_2213;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4580 & _GEN_5787) begin // @[StoreSet.scala 547:30]
        robIdxVec_25_0_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_25_0_flag <= _GEN_2086;
      end
    end else begin
      robIdxVec_25_0_flag <= _GEN_2086;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4580 & _GEN_5787) begin // @[StoreSet.scala 547:30]
        robIdxVec_25_0_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_25_0_value <= _GEN_2214;
      end
    end else begin
      robIdxVec_25_0_value <= _GEN_2214;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4580 & _GEN_5790) begin // @[StoreSet.scala 547:30]
        robIdxVec_25_1_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_25_1_flag <= _GEN_2087;
      end
    end else begin
      robIdxVec_25_1_flag <= _GEN_2087;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4580 & _GEN_5790) begin // @[StoreSet.scala 547:30]
        robIdxVec_25_1_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_25_1_value <= _GEN_2215;
      end
    end else begin
      robIdxVec_25_1_value <= _GEN_2215;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4580 & _GEN_5793) begin // @[StoreSet.scala 547:30]
        robIdxVec_25_2_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_25_2_flag <= _GEN_2088;
      end
    end else begin
      robIdxVec_25_2_flag <= _GEN_2088;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4580 & _GEN_5793) begin // @[StoreSet.scala 547:30]
        robIdxVec_25_2_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_25_2_value <= _GEN_2216;
      end
    end else begin
      robIdxVec_25_2_value <= _GEN_2216;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4580 & _GEN_5796) begin // @[StoreSet.scala 547:30]
        robIdxVec_25_3_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_25_3_flag <= _GEN_2089;
      end
    end else begin
      robIdxVec_25_3_flag <= _GEN_2089;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4580 & _GEN_5796) begin // @[StoreSet.scala 547:30]
        robIdxVec_25_3_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_25_3_value <= _GEN_2217;
      end
    end else begin
      robIdxVec_25_3_value <= _GEN_2217;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4588 & _GEN_5787) begin // @[StoreSet.scala 547:30]
        robIdxVec_26_0_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_26_0_flag <= _GEN_2090;
      end
    end else begin
      robIdxVec_26_0_flag <= _GEN_2090;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4588 & _GEN_5787) begin // @[StoreSet.scala 547:30]
        robIdxVec_26_0_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_26_0_value <= _GEN_2218;
      end
    end else begin
      robIdxVec_26_0_value <= _GEN_2218;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4588 & _GEN_5790) begin // @[StoreSet.scala 547:30]
        robIdxVec_26_1_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_26_1_flag <= _GEN_2091;
      end
    end else begin
      robIdxVec_26_1_flag <= _GEN_2091;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4588 & _GEN_5790) begin // @[StoreSet.scala 547:30]
        robIdxVec_26_1_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_26_1_value <= _GEN_2219;
      end
    end else begin
      robIdxVec_26_1_value <= _GEN_2219;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4588 & _GEN_5793) begin // @[StoreSet.scala 547:30]
        robIdxVec_26_2_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_26_2_flag <= _GEN_2092;
      end
    end else begin
      robIdxVec_26_2_flag <= _GEN_2092;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4588 & _GEN_5793) begin // @[StoreSet.scala 547:30]
        robIdxVec_26_2_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_26_2_value <= _GEN_2220;
      end
    end else begin
      robIdxVec_26_2_value <= _GEN_2220;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4588 & _GEN_5796) begin // @[StoreSet.scala 547:30]
        robIdxVec_26_3_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_26_3_flag <= _GEN_2093;
      end
    end else begin
      robIdxVec_26_3_flag <= _GEN_2093;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4588 & _GEN_5796) begin // @[StoreSet.scala 547:30]
        robIdxVec_26_3_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_26_3_value <= _GEN_2221;
      end
    end else begin
      robIdxVec_26_3_value <= _GEN_2221;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4596 & _GEN_5787) begin // @[StoreSet.scala 547:30]
        robIdxVec_27_0_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_27_0_flag <= _GEN_2094;
      end
    end else begin
      robIdxVec_27_0_flag <= _GEN_2094;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4596 & _GEN_5787) begin // @[StoreSet.scala 547:30]
        robIdxVec_27_0_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_27_0_value <= _GEN_2222;
      end
    end else begin
      robIdxVec_27_0_value <= _GEN_2222;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4596 & _GEN_5790) begin // @[StoreSet.scala 547:30]
        robIdxVec_27_1_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_27_1_flag <= _GEN_2095;
      end
    end else begin
      robIdxVec_27_1_flag <= _GEN_2095;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4596 & _GEN_5790) begin // @[StoreSet.scala 547:30]
        robIdxVec_27_1_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_27_1_value <= _GEN_2223;
      end
    end else begin
      robIdxVec_27_1_value <= _GEN_2223;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4596 & _GEN_5793) begin // @[StoreSet.scala 547:30]
        robIdxVec_27_2_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_27_2_flag <= _GEN_2096;
      end
    end else begin
      robIdxVec_27_2_flag <= _GEN_2096;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4596 & _GEN_5793) begin // @[StoreSet.scala 547:30]
        robIdxVec_27_2_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_27_2_value <= _GEN_2224;
      end
    end else begin
      robIdxVec_27_2_value <= _GEN_2224;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4596 & _GEN_5796) begin // @[StoreSet.scala 547:30]
        robIdxVec_27_3_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_27_3_flag <= _GEN_2097;
      end
    end else begin
      robIdxVec_27_3_flag <= _GEN_2097;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4596 & _GEN_5796) begin // @[StoreSet.scala 547:30]
        robIdxVec_27_3_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_27_3_value <= _GEN_2225;
      end
    end else begin
      robIdxVec_27_3_value <= _GEN_2225;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4604 & _GEN_5787) begin // @[StoreSet.scala 547:30]
        robIdxVec_28_0_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_28_0_flag <= _GEN_2098;
      end
    end else begin
      robIdxVec_28_0_flag <= _GEN_2098;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4604 & _GEN_5787) begin // @[StoreSet.scala 547:30]
        robIdxVec_28_0_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_28_0_value <= _GEN_2226;
      end
    end else begin
      robIdxVec_28_0_value <= _GEN_2226;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4604 & _GEN_5790) begin // @[StoreSet.scala 547:30]
        robIdxVec_28_1_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_28_1_flag <= _GEN_2099;
      end
    end else begin
      robIdxVec_28_1_flag <= _GEN_2099;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4604 & _GEN_5790) begin // @[StoreSet.scala 547:30]
        robIdxVec_28_1_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_28_1_value <= _GEN_2227;
      end
    end else begin
      robIdxVec_28_1_value <= _GEN_2227;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4604 & _GEN_5793) begin // @[StoreSet.scala 547:30]
        robIdxVec_28_2_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_28_2_flag <= _GEN_2100;
      end
    end else begin
      robIdxVec_28_2_flag <= _GEN_2100;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4604 & _GEN_5793) begin // @[StoreSet.scala 547:30]
        robIdxVec_28_2_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_28_2_value <= _GEN_2228;
      end
    end else begin
      robIdxVec_28_2_value <= _GEN_2228;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4604 & _GEN_5796) begin // @[StoreSet.scala 547:30]
        robIdxVec_28_3_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_28_3_flag <= _GEN_2101;
      end
    end else begin
      robIdxVec_28_3_flag <= _GEN_2101;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4604 & _GEN_5796) begin // @[StoreSet.scala 547:30]
        robIdxVec_28_3_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_28_3_value <= _GEN_2229;
      end
    end else begin
      robIdxVec_28_3_value <= _GEN_2229;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4612 & _GEN_5787) begin // @[StoreSet.scala 547:30]
        robIdxVec_29_0_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_29_0_flag <= _GEN_2102;
      end
    end else begin
      robIdxVec_29_0_flag <= _GEN_2102;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4612 & _GEN_5787) begin // @[StoreSet.scala 547:30]
        robIdxVec_29_0_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_29_0_value <= _GEN_2230;
      end
    end else begin
      robIdxVec_29_0_value <= _GEN_2230;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4612 & _GEN_5790) begin // @[StoreSet.scala 547:30]
        robIdxVec_29_1_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_29_1_flag <= _GEN_2103;
      end
    end else begin
      robIdxVec_29_1_flag <= _GEN_2103;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4612 & _GEN_5790) begin // @[StoreSet.scala 547:30]
        robIdxVec_29_1_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_29_1_value <= _GEN_2231;
      end
    end else begin
      robIdxVec_29_1_value <= _GEN_2231;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4612 & _GEN_5793) begin // @[StoreSet.scala 547:30]
        robIdxVec_29_2_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_29_2_flag <= _GEN_2104;
      end
    end else begin
      robIdxVec_29_2_flag <= _GEN_2104;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4612 & _GEN_5793) begin // @[StoreSet.scala 547:30]
        robIdxVec_29_2_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_29_2_value <= _GEN_2232;
      end
    end else begin
      robIdxVec_29_2_value <= _GEN_2232;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4612 & _GEN_5796) begin // @[StoreSet.scala 547:30]
        robIdxVec_29_3_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_29_3_flag <= _GEN_2105;
      end
    end else begin
      robIdxVec_29_3_flag <= _GEN_2105;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4612 & _GEN_5796) begin // @[StoreSet.scala 547:30]
        robIdxVec_29_3_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_29_3_value <= _GEN_2233;
      end
    end else begin
      robIdxVec_29_3_value <= _GEN_2233;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4620 & _GEN_5787) begin // @[StoreSet.scala 547:30]
        robIdxVec_30_0_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_30_0_flag <= _GEN_2106;
      end
    end else begin
      robIdxVec_30_0_flag <= _GEN_2106;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4620 & _GEN_5787) begin // @[StoreSet.scala 547:30]
        robIdxVec_30_0_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_30_0_value <= _GEN_2234;
      end
    end else begin
      robIdxVec_30_0_value <= _GEN_2234;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4620 & _GEN_5790) begin // @[StoreSet.scala 547:30]
        robIdxVec_30_1_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_30_1_flag <= _GEN_2107;
      end
    end else begin
      robIdxVec_30_1_flag <= _GEN_2107;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4620 & _GEN_5790) begin // @[StoreSet.scala 547:30]
        robIdxVec_30_1_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_30_1_value <= _GEN_2235;
      end
    end else begin
      robIdxVec_30_1_value <= _GEN_2235;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4620 & _GEN_5793) begin // @[StoreSet.scala 547:30]
        robIdxVec_30_2_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_30_2_flag <= _GEN_2108;
      end
    end else begin
      robIdxVec_30_2_flag <= _GEN_2108;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4620 & _GEN_5793) begin // @[StoreSet.scala 547:30]
        robIdxVec_30_2_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_30_2_value <= _GEN_2236;
      end
    end else begin
      robIdxVec_30_2_value <= _GEN_2236;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4620 & _GEN_5796) begin // @[StoreSet.scala 547:30]
        robIdxVec_30_3_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_30_3_flag <= _GEN_2109;
      end
    end else begin
      robIdxVec_30_3_flag <= _GEN_2109;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4620 & _GEN_5796) begin // @[StoreSet.scala 547:30]
        robIdxVec_30_3_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_30_3_value <= _GEN_2237;
      end
    end else begin
      robIdxVec_30_3_value <= _GEN_2237;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4628 & _GEN_5787) begin // @[StoreSet.scala 547:30]
        robIdxVec_31_0_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_31_0_flag <= _GEN_2110;
      end
    end else begin
      robIdxVec_31_0_flag <= _GEN_2110;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4628 & _GEN_5787) begin // @[StoreSet.scala 547:30]
        robIdxVec_31_0_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_31_0_value <= _GEN_2238;
      end
    end else begin
      robIdxVec_31_0_value <= _GEN_2238;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4628 & _GEN_5790) begin // @[StoreSet.scala 547:30]
        robIdxVec_31_1_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_31_1_flag <= _GEN_2111;
      end
    end else begin
      robIdxVec_31_1_flag <= _GEN_2111;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4628 & _GEN_5790) begin // @[StoreSet.scala 547:30]
        robIdxVec_31_1_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_31_1_value <= _GEN_2239;
      end
    end else begin
      robIdxVec_31_1_value <= _GEN_2239;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4628 & _GEN_5793) begin // @[StoreSet.scala 547:30]
        robIdxVec_31_2_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_31_2_flag <= _GEN_2112;
      end
    end else begin
      robIdxVec_31_2_flag <= _GEN_2112;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4628 & _GEN_5793) begin // @[StoreSet.scala 547:30]
        robIdxVec_31_2_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_31_2_value <= _GEN_2240;
      end
    end else begin
      robIdxVec_31_2_value <= _GEN_2240;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4628 & _GEN_5796) begin // @[StoreSet.scala 547:30]
        robIdxVec_31_3_flag <= io_dispatch_req_1_bits_robIdx_flag; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_31_3_flag <= _GEN_2113;
      end
    end else begin
      robIdxVec_31_3_flag <= _GEN_2113;
    end
    if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      if (_GEN_4628 & _GEN_5796) begin // @[StoreSet.scala 547:30]
        robIdxVec_31_3_value <= io_dispatch_req_1_bits_robIdx_value; // @[StoreSet.scala 547:30]
      end else begin
        robIdxVec_31_3_value <= _GEN_2241;
      end
    end else begin
      robIdxVec_31_3_value <= _GEN_2241;
    end
    REG <= io_redirect_valid; // @[StoreSet.scala 562:15]
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_0_0 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_0_0 & _T_28) begin // @[StoreSet.scala 542:70]
      validVec_0_0 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_0_0 <= _GEN_2274;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_0_0 <= _GEN_1442;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1057) begin
      validVec_0_0 <= _GEN_1058;
    end else begin
      validVec_0_0 <= _GEN_706;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_0_1 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_0_1 & _T_32) begin // @[StoreSet.scala 542:70]
      validVec_0_1 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_0_1 <= _GEN_2275;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_0_1 <= _GEN_1443;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1153) begin
      validVec_0_1 <= _GEN_1154;
    end else begin
      validVec_0_1 <= _GEN_802;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_0_2 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_0_2 & _T_36) begin // @[StoreSet.scala 542:70]
      validVec_0_2 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_0_2 <= _GEN_2276;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_0_2 <= _GEN_1444;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1249) begin
      validVec_0_2 <= _GEN_1250;
    end else begin
      validVec_0_2 <= _GEN_898;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_0_3 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_0_3 & _T_40) begin // @[StoreSet.scala 542:70]
      validVec_0_3 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_0_3 <= _GEN_2277;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_0_3 <= _GEN_1445;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1345) begin
      validVec_0_3 <= _GEN_1346;
    end else begin
      validVec_0_3 <= _GEN_994;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_1_0 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_1_0 & _T_44) begin // @[StoreSet.scala 542:70]
      validVec_1_0 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_1_0 <= _GEN_2278;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_1_0 <= _GEN_1446;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1057) begin
      validVec_1_0 <= _GEN_1059;
    end else begin
      validVec_1_0 <= _GEN_707;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_1_1 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_1_1 & _T_48) begin // @[StoreSet.scala 542:70]
      validVec_1_1 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_1_1 <= _GEN_2279;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_1_1 <= _GEN_1447;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1153) begin
      validVec_1_1 <= _GEN_1155;
    end else begin
      validVec_1_1 <= _GEN_803;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_1_2 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_1_2 & _T_52) begin // @[StoreSet.scala 542:70]
      validVec_1_2 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_1_2 <= _GEN_2280;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_1_2 <= _GEN_1448;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1249) begin
      validVec_1_2 <= _GEN_1251;
    end else begin
      validVec_1_2 <= _GEN_899;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_1_3 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_1_3 & _T_56) begin // @[StoreSet.scala 542:70]
      validVec_1_3 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_1_3 <= _GEN_2281;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_1_3 <= _GEN_1449;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1345) begin
      validVec_1_3 <= _GEN_1347;
    end else begin
      validVec_1_3 <= _GEN_995;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_2_0 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_2_0 & _T_60) begin // @[StoreSet.scala 542:70]
      validVec_2_0 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_2_0 <= _GEN_2282;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_2_0 <= _GEN_1450;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1057) begin
      validVec_2_0 <= _GEN_1060;
    end else begin
      validVec_2_0 <= _GEN_708;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_2_1 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_2_1 & _T_64) begin // @[StoreSet.scala 542:70]
      validVec_2_1 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_2_1 <= _GEN_2283;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_2_1 <= _GEN_1451;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1153) begin
      validVec_2_1 <= _GEN_1156;
    end else begin
      validVec_2_1 <= _GEN_804;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_2_2 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_2_2 & _T_68) begin // @[StoreSet.scala 542:70]
      validVec_2_2 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_2_2 <= _GEN_2284;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_2_2 <= _GEN_1452;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1249) begin
      validVec_2_2 <= _GEN_1252;
    end else begin
      validVec_2_2 <= _GEN_900;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_2_3 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_2_3 & _T_72) begin // @[StoreSet.scala 542:70]
      validVec_2_3 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_2_3 <= _GEN_2285;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_2_3 <= _GEN_1453;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1345) begin
      validVec_2_3 <= _GEN_1348;
    end else begin
      validVec_2_3 <= _GEN_996;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_3_0 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_3_0 & _T_76) begin // @[StoreSet.scala 542:70]
      validVec_3_0 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_3_0 <= _GEN_2286;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_3_0 <= _GEN_1454;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1057) begin
      validVec_3_0 <= _GEN_1061;
    end else begin
      validVec_3_0 <= _GEN_709;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_3_1 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_3_1 & _T_80) begin // @[StoreSet.scala 542:70]
      validVec_3_1 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_3_1 <= _GEN_2287;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_3_1 <= _GEN_1455;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1153) begin
      validVec_3_1 <= _GEN_1157;
    end else begin
      validVec_3_1 <= _GEN_805;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_3_2 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_3_2 & _T_84) begin // @[StoreSet.scala 542:70]
      validVec_3_2 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_3_2 <= _GEN_2288;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_3_2 <= _GEN_1456;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1249) begin
      validVec_3_2 <= _GEN_1253;
    end else begin
      validVec_3_2 <= _GEN_901;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_3_3 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_3_3 & _T_88) begin // @[StoreSet.scala 542:70]
      validVec_3_3 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_3_3 <= _GEN_2289;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_3_3 <= _GEN_1457;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1345) begin
      validVec_3_3 <= _GEN_1349;
    end else begin
      validVec_3_3 <= _GEN_997;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_4_0 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_4_0 & _T_92) begin // @[StoreSet.scala 542:70]
      validVec_4_0 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_4_0 <= _GEN_2290;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_4_0 <= _GEN_1458;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1057) begin
      validVec_4_0 <= _GEN_1062;
    end else begin
      validVec_4_0 <= _GEN_710;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_4_1 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_4_1 & _T_96) begin // @[StoreSet.scala 542:70]
      validVec_4_1 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_4_1 <= _GEN_2291;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_4_1 <= _GEN_1459;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1153) begin
      validVec_4_1 <= _GEN_1158;
    end else begin
      validVec_4_1 <= _GEN_806;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_4_2 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_4_2 & _T_100) begin // @[StoreSet.scala 542:70]
      validVec_4_2 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_4_2 <= _GEN_2292;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_4_2 <= _GEN_1460;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1249) begin
      validVec_4_2 <= _GEN_1254;
    end else begin
      validVec_4_2 <= _GEN_902;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_4_3 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_4_3 & _T_104) begin // @[StoreSet.scala 542:70]
      validVec_4_3 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_4_3 <= _GEN_2293;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_4_3 <= _GEN_1461;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1345) begin
      validVec_4_3 <= _GEN_1350;
    end else begin
      validVec_4_3 <= _GEN_998;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_5_0 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_5_0 & _T_108) begin // @[StoreSet.scala 542:70]
      validVec_5_0 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_5_0 <= _GEN_2294;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_5_0 <= _GEN_1462;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1057) begin
      validVec_5_0 <= _GEN_1063;
    end else begin
      validVec_5_0 <= _GEN_711;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_5_1 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_5_1 & _T_112) begin // @[StoreSet.scala 542:70]
      validVec_5_1 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_5_1 <= _GEN_2295;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_5_1 <= _GEN_1463;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1153) begin
      validVec_5_1 <= _GEN_1159;
    end else begin
      validVec_5_1 <= _GEN_807;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_5_2 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_5_2 & _T_116) begin // @[StoreSet.scala 542:70]
      validVec_5_2 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_5_2 <= _GEN_2296;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_5_2 <= _GEN_1464;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1249) begin
      validVec_5_2 <= _GEN_1255;
    end else begin
      validVec_5_2 <= _GEN_903;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_5_3 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_5_3 & _T_120) begin // @[StoreSet.scala 542:70]
      validVec_5_3 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_5_3 <= _GEN_2297;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_5_3 <= _GEN_1465;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1345) begin
      validVec_5_3 <= _GEN_1351;
    end else begin
      validVec_5_3 <= _GEN_999;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_6_0 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_6_0 & _T_124) begin // @[StoreSet.scala 542:70]
      validVec_6_0 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_6_0 <= _GEN_2298;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_6_0 <= _GEN_1466;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1057) begin
      validVec_6_0 <= _GEN_1064;
    end else begin
      validVec_6_0 <= _GEN_712;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_6_1 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_6_1 & _T_128) begin // @[StoreSet.scala 542:70]
      validVec_6_1 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_6_1 <= _GEN_2299;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_6_1 <= _GEN_1467;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1153) begin
      validVec_6_1 <= _GEN_1160;
    end else begin
      validVec_6_1 <= _GEN_808;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_6_2 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_6_2 & _T_132) begin // @[StoreSet.scala 542:70]
      validVec_6_2 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_6_2 <= _GEN_2300;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_6_2 <= _GEN_1468;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1249) begin
      validVec_6_2 <= _GEN_1256;
    end else begin
      validVec_6_2 <= _GEN_904;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_6_3 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_6_3 & _T_136) begin // @[StoreSet.scala 542:70]
      validVec_6_3 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_6_3 <= _GEN_2301;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_6_3 <= _GEN_1469;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1345) begin
      validVec_6_3 <= _GEN_1352;
    end else begin
      validVec_6_3 <= _GEN_1000;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_7_0 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_7_0 & _T_140) begin // @[StoreSet.scala 542:70]
      validVec_7_0 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_7_0 <= _GEN_2302;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_7_0 <= _GEN_1470;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1057) begin
      validVec_7_0 <= _GEN_1065;
    end else begin
      validVec_7_0 <= _GEN_713;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_7_1 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_7_1 & _T_144) begin // @[StoreSet.scala 542:70]
      validVec_7_1 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_7_1 <= _GEN_2303;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_7_1 <= _GEN_1471;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1153) begin
      validVec_7_1 <= _GEN_1161;
    end else begin
      validVec_7_1 <= _GEN_809;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_7_2 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_7_2 & _T_148) begin // @[StoreSet.scala 542:70]
      validVec_7_2 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_7_2 <= _GEN_2304;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_7_2 <= _GEN_1472;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1249) begin
      validVec_7_2 <= _GEN_1257;
    end else begin
      validVec_7_2 <= _GEN_905;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_7_3 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_7_3 & _T_152) begin // @[StoreSet.scala 542:70]
      validVec_7_3 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_7_3 <= _GEN_2305;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_7_3 <= _GEN_1473;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1345) begin
      validVec_7_3 <= _GEN_1353;
    end else begin
      validVec_7_3 <= _GEN_1001;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_8_0 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_8_0 & _T_156) begin // @[StoreSet.scala 542:70]
      validVec_8_0 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_8_0 <= _GEN_2306;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_8_0 <= _GEN_1474;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1057) begin
      validVec_8_0 <= _GEN_1066;
    end else begin
      validVec_8_0 <= _GEN_714;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_8_1 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_8_1 & _T_160) begin // @[StoreSet.scala 542:70]
      validVec_8_1 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_8_1 <= _GEN_2307;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_8_1 <= _GEN_1475;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1153) begin
      validVec_8_1 <= _GEN_1162;
    end else begin
      validVec_8_1 <= _GEN_810;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_8_2 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_8_2 & _T_164) begin // @[StoreSet.scala 542:70]
      validVec_8_2 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_8_2 <= _GEN_2308;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_8_2 <= _GEN_1476;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1249) begin
      validVec_8_2 <= _GEN_1258;
    end else begin
      validVec_8_2 <= _GEN_906;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_8_3 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_8_3 & _T_168) begin // @[StoreSet.scala 542:70]
      validVec_8_3 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_8_3 <= _GEN_2309;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_8_3 <= _GEN_1477;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1345) begin
      validVec_8_3 <= _GEN_1354;
    end else begin
      validVec_8_3 <= _GEN_1002;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_9_0 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_9_0 & _T_172) begin // @[StoreSet.scala 542:70]
      validVec_9_0 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_9_0 <= _GEN_2310;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_9_0 <= _GEN_1478;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1057) begin
      validVec_9_0 <= _GEN_1067;
    end else begin
      validVec_9_0 <= _GEN_715;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_9_1 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_9_1 & _T_176) begin // @[StoreSet.scala 542:70]
      validVec_9_1 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_9_1 <= _GEN_2311;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_9_1 <= _GEN_1479;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1153) begin
      validVec_9_1 <= _GEN_1163;
    end else begin
      validVec_9_1 <= _GEN_811;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_9_2 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_9_2 & _T_180) begin // @[StoreSet.scala 542:70]
      validVec_9_2 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_9_2 <= _GEN_2312;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_9_2 <= _GEN_1480;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1249) begin
      validVec_9_2 <= _GEN_1259;
    end else begin
      validVec_9_2 <= _GEN_907;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_9_3 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_9_3 & _T_184) begin // @[StoreSet.scala 542:70]
      validVec_9_3 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_9_3 <= _GEN_2313;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_9_3 <= _GEN_1481;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1345) begin
      validVec_9_3 <= _GEN_1355;
    end else begin
      validVec_9_3 <= _GEN_1003;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_10_0 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_10_0 & _T_188) begin // @[StoreSet.scala 542:70]
      validVec_10_0 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_10_0 <= _GEN_2314;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_10_0 <= _GEN_1482;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1057) begin
      validVec_10_0 <= _GEN_1068;
    end else begin
      validVec_10_0 <= _GEN_716;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_10_1 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_10_1 & _T_192) begin // @[StoreSet.scala 542:70]
      validVec_10_1 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_10_1 <= _GEN_2315;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_10_1 <= _GEN_1483;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1153) begin
      validVec_10_1 <= _GEN_1164;
    end else begin
      validVec_10_1 <= _GEN_812;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_10_2 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_10_2 & _T_196) begin // @[StoreSet.scala 542:70]
      validVec_10_2 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_10_2 <= _GEN_2316;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_10_2 <= _GEN_1484;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1249) begin
      validVec_10_2 <= _GEN_1260;
    end else begin
      validVec_10_2 <= _GEN_908;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_10_3 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_10_3 & _T_200) begin // @[StoreSet.scala 542:70]
      validVec_10_3 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_10_3 <= _GEN_2317;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_10_3 <= _GEN_1485;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1345) begin
      validVec_10_3 <= _GEN_1356;
    end else begin
      validVec_10_3 <= _GEN_1004;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_11_0 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_11_0 & _T_204) begin // @[StoreSet.scala 542:70]
      validVec_11_0 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_11_0 <= _GEN_2318;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_11_0 <= _GEN_1486;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1057) begin
      validVec_11_0 <= _GEN_1069;
    end else begin
      validVec_11_0 <= _GEN_717;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_11_1 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_11_1 & _T_208) begin // @[StoreSet.scala 542:70]
      validVec_11_1 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_11_1 <= _GEN_2319;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_11_1 <= _GEN_1487;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1153) begin
      validVec_11_1 <= _GEN_1165;
    end else begin
      validVec_11_1 <= _GEN_813;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_11_2 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_11_2 & _T_212) begin // @[StoreSet.scala 542:70]
      validVec_11_2 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_11_2 <= _GEN_2320;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_11_2 <= _GEN_1488;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1249) begin
      validVec_11_2 <= _GEN_1261;
    end else begin
      validVec_11_2 <= _GEN_909;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_11_3 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_11_3 & _T_216) begin // @[StoreSet.scala 542:70]
      validVec_11_3 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_11_3 <= _GEN_2321;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_11_3 <= _GEN_1489;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1345) begin
      validVec_11_3 <= _GEN_1357;
    end else begin
      validVec_11_3 <= _GEN_1005;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_12_0 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_12_0 & _T_220) begin // @[StoreSet.scala 542:70]
      validVec_12_0 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_12_0 <= _GEN_2322;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_12_0 <= _GEN_1490;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1057) begin
      validVec_12_0 <= _GEN_1070;
    end else begin
      validVec_12_0 <= _GEN_718;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_12_1 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_12_1 & _T_224) begin // @[StoreSet.scala 542:70]
      validVec_12_1 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_12_1 <= _GEN_2323;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_12_1 <= _GEN_1491;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1153) begin
      validVec_12_1 <= _GEN_1166;
    end else begin
      validVec_12_1 <= _GEN_814;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_12_2 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_12_2 & _T_228) begin // @[StoreSet.scala 542:70]
      validVec_12_2 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_12_2 <= _GEN_2324;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_12_2 <= _GEN_1492;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1249) begin
      validVec_12_2 <= _GEN_1262;
    end else begin
      validVec_12_2 <= _GEN_910;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_12_3 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_12_3 & _T_232) begin // @[StoreSet.scala 542:70]
      validVec_12_3 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_12_3 <= _GEN_2325;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_12_3 <= _GEN_1493;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1345) begin
      validVec_12_3 <= _GEN_1358;
    end else begin
      validVec_12_3 <= _GEN_1006;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_13_0 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_13_0 & _T_236) begin // @[StoreSet.scala 542:70]
      validVec_13_0 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_13_0 <= _GEN_2326;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_13_0 <= _GEN_1494;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1057) begin
      validVec_13_0 <= _GEN_1071;
    end else begin
      validVec_13_0 <= _GEN_719;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_13_1 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_13_1 & _T_240) begin // @[StoreSet.scala 542:70]
      validVec_13_1 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_13_1 <= _GEN_2327;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_13_1 <= _GEN_1495;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1153) begin
      validVec_13_1 <= _GEN_1167;
    end else begin
      validVec_13_1 <= _GEN_815;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_13_2 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_13_2 & _T_244) begin // @[StoreSet.scala 542:70]
      validVec_13_2 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_13_2 <= _GEN_2328;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_13_2 <= _GEN_1496;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1249) begin
      validVec_13_2 <= _GEN_1263;
    end else begin
      validVec_13_2 <= _GEN_911;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_13_3 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_13_3 & _T_248) begin // @[StoreSet.scala 542:70]
      validVec_13_3 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_13_3 <= _GEN_2329;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_13_3 <= _GEN_1497;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1345) begin
      validVec_13_3 <= _GEN_1359;
    end else begin
      validVec_13_3 <= _GEN_1007;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_14_0 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_14_0 & _T_252) begin // @[StoreSet.scala 542:70]
      validVec_14_0 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_14_0 <= _GEN_2330;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_14_0 <= _GEN_1498;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1057) begin
      validVec_14_0 <= _GEN_1072;
    end else begin
      validVec_14_0 <= _GEN_720;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_14_1 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_14_1 & _T_256) begin // @[StoreSet.scala 542:70]
      validVec_14_1 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_14_1 <= _GEN_2331;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_14_1 <= _GEN_1499;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1153) begin
      validVec_14_1 <= _GEN_1168;
    end else begin
      validVec_14_1 <= _GEN_816;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_14_2 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_14_2 & _T_260) begin // @[StoreSet.scala 542:70]
      validVec_14_2 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_14_2 <= _GEN_2332;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_14_2 <= _GEN_1500;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1249) begin
      validVec_14_2 <= _GEN_1264;
    end else begin
      validVec_14_2 <= _GEN_912;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_14_3 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_14_3 & _T_264) begin // @[StoreSet.scala 542:70]
      validVec_14_3 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_14_3 <= _GEN_2333;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_14_3 <= _GEN_1501;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1345) begin
      validVec_14_3 <= _GEN_1360;
    end else begin
      validVec_14_3 <= _GEN_1008;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_15_0 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_15_0 & _T_268) begin // @[StoreSet.scala 542:70]
      validVec_15_0 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_15_0 <= _GEN_2334;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_15_0 <= _GEN_1502;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1057) begin
      validVec_15_0 <= _GEN_1073;
    end else begin
      validVec_15_0 <= _GEN_721;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_15_1 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_15_1 & _T_272) begin // @[StoreSet.scala 542:70]
      validVec_15_1 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_15_1 <= _GEN_2335;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_15_1 <= _GEN_1503;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1153) begin
      validVec_15_1 <= _GEN_1169;
    end else begin
      validVec_15_1 <= _GEN_817;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_15_2 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_15_2 & _T_276) begin // @[StoreSet.scala 542:70]
      validVec_15_2 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_15_2 <= _GEN_2336;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_15_2 <= _GEN_1504;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1249) begin
      validVec_15_2 <= _GEN_1265;
    end else begin
      validVec_15_2 <= _GEN_913;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_15_3 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_15_3 & _T_280) begin // @[StoreSet.scala 542:70]
      validVec_15_3 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_15_3 <= _GEN_2337;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_15_3 <= _GEN_1505;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1345) begin
      validVec_15_3 <= _GEN_1361;
    end else begin
      validVec_15_3 <= _GEN_1009;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_16_0 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_16_0 & _T_284) begin // @[StoreSet.scala 542:70]
      validVec_16_0 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_16_0 <= _GEN_2338;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_16_0 <= _GEN_1506;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1057) begin
      validVec_16_0 <= _GEN_1074;
    end else begin
      validVec_16_0 <= _GEN_722;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_16_1 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_16_1 & _T_288) begin // @[StoreSet.scala 542:70]
      validVec_16_1 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_16_1 <= _GEN_2339;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_16_1 <= _GEN_1507;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1153) begin
      validVec_16_1 <= _GEN_1170;
    end else begin
      validVec_16_1 <= _GEN_818;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_16_2 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_16_2 & _T_292) begin // @[StoreSet.scala 542:70]
      validVec_16_2 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_16_2 <= _GEN_2340;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_16_2 <= _GEN_1508;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1249) begin
      validVec_16_2 <= _GEN_1266;
    end else begin
      validVec_16_2 <= _GEN_914;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_16_3 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_16_3 & _T_296) begin // @[StoreSet.scala 542:70]
      validVec_16_3 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_16_3 <= _GEN_2341;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_16_3 <= _GEN_1509;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1345) begin
      validVec_16_3 <= _GEN_1362;
    end else begin
      validVec_16_3 <= _GEN_1010;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_17_0 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_17_0 & _T_300) begin // @[StoreSet.scala 542:70]
      validVec_17_0 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_17_0 <= _GEN_2342;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_17_0 <= _GEN_1510;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1057) begin
      validVec_17_0 <= _GEN_1075;
    end else begin
      validVec_17_0 <= _GEN_723;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_17_1 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_17_1 & _T_304) begin // @[StoreSet.scala 542:70]
      validVec_17_1 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_17_1 <= _GEN_2343;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_17_1 <= _GEN_1511;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1153) begin
      validVec_17_1 <= _GEN_1171;
    end else begin
      validVec_17_1 <= _GEN_819;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_17_2 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_17_2 & _T_308) begin // @[StoreSet.scala 542:70]
      validVec_17_2 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_17_2 <= _GEN_2344;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_17_2 <= _GEN_1512;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1249) begin
      validVec_17_2 <= _GEN_1267;
    end else begin
      validVec_17_2 <= _GEN_915;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_17_3 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_17_3 & _T_312) begin // @[StoreSet.scala 542:70]
      validVec_17_3 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_17_3 <= _GEN_2345;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_17_3 <= _GEN_1513;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1345) begin
      validVec_17_3 <= _GEN_1363;
    end else begin
      validVec_17_3 <= _GEN_1011;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_18_0 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_18_0 & _T_316) begin // @[StoreSet.scala 542:70]
      validVec_18_0 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_18_0 <= _GEN_2346;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_18_0 <= _GEN_1514;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1057) begin
      validVec_18_0 <= _GEN_1076;
    end else begin
      validVec_18_0 <= _GEN_724;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_18_1 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_18_1 & _T_320) begin // @[StoreSet.scala 542:70]
      validVec_18_1 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_18_1 <= _GEN_2347;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_18_1 <= _GEN_1515;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1153) begin
      validVec_18_1 <= _GEN_1172;
    end else begin
      validVec_18_1 <= _GEN_820;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_18_2 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_18_2 & _T_324) begin // @[StoreSet.scala 542:70]
      validVec_18_2 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_18_2 <= _GEN_2348;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_18_2 <= _GEN_1516;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1249) begin
      validVec_18_2 <= _GEN_1268;
    end else begin
      validVec_18_2 <= _GEN_916;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_18_3 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_18_3 & _T_328) begin // @[StoreSet.scala 542:70]
      validVec_18_3 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_18_3 <= _GEN_2349;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_18_3 <= _GEN_1517;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1345) begin
      validVec_18_3 <= _GEN_1364;
    end else begin
      validVec_18_3 <= _GEN_1012;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_19_0 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_19_0 & _T_332) begin // @[StoreSet.scala 542:70]
      validVec_19_0 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_19_0 <= _GEN_2350;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_19_0 <= _GEN_1518;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1057) begin
      validVec_19_0 <= _GEN_1077;
    end else begin
      validVec_19_0 <= _GEN_725;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_19_1 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_19_1 & _T_336) begin // @[StoreSet.scala 542:70]
      validVec_19_1 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_19_1 <= _GEN_2351;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_19_1 <= _GEN_1519;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1153) begin
      validVec_19_1 <= _GEN_1173;
    end else begin
      validVec_19_1 <= _GEN_821;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_19_2 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_19_2 & _T_340) begin // @[StoreSet.scala 542:70]
      validVec_19_2 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_19_2 <= _GEN_2352;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_19_2 <= _GEN_1520;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1249) begin
      validVec_19_2 <= _GEN_1269;
    end else begin
      validVec_19_2 <= _GEN_917;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_19_3 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_19_3 & _T_344) begin // @[StoreSet.scala 542:70]
      validVec_19_3 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_19_3 <= _GEN_2353;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_19_3 <= _GEN_1521;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1345) begin
      validVec_19_3 <= _GEN_1365;
    end else begin
      validVec_19_3 <= _GEN_1013;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_20_0 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_20_0 & _T_348) begin // @[StoreSet.scala 542:70]
      validVec_20_0 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_20_0 <= _GEN_2354;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_20_0 <= _GEN_1522;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1057) begin
      validVec_20_0 <= _GEN_1078;
    end else begin
      validVec_20_0 <= _GEN_726;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_20_1 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_20_1 & _T_352) begin // @[StoreSet.scala 542:70]
      validVec_20_1 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_20_1 <= _GEN_2355;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_20_1 <= _GEN_1523;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1153) begin
      validVec_20_1 <= _GEN_1174;
    end else begin
      validVec_20_1 <= _GEN_822;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_20_2 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_20_2 & _T_356) begin // @[StoreSet.scala 542:70]
      validVec_20_2 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_20_2 <= _GEN_2356;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_20_2 <= _GEN_1524;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1249) begin
      validVec_20_2 <= _GEN_1270;
    end else begin
      validVec_20_2 <= _GEN_918;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_20_3 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_20_3 & _T_360) begin // @[StoreSet.scala 542:70]
      validVec_20_3 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_20_3 <= _GEN_2357;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_20_3 <= _GEN_1525;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1345) begin
      validVec_20_3 <= _GEN_1366;
    end else begin
      validVec_20_3 <= _GEN_1014;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_21_0 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_21_0 & _T_364) begin // @[StoreSet.scala 542:70]
      validVec_21_0 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_21_0 <= _GEN_2358;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_21_0 <= _GEN_1526;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1057) begin
      validVec_21_0 <= _GEN_1079;
    end else begin
      validVec_21_0 <= _GEN_727;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_21_1 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_21_1 & _T_368) begin // @[StoreSet.scala 542:70]
      validVec_21_1 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_21_1 <= _GEN_2359;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_21_1 <= _GEN_1527;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1153) begin
      validVec_21_1 <= _GEN_1175;
    end else begin
      validVec_21_1 <= _GEN_823;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_21_2 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_21_2 & _T_372) begin // @[StoreSet.scala 542:70]
      validVec_21_2 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_21_2 <= _GEN_2360;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_21_2 <= _GEN_1528;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1249) begin
      validVec_21_2 <= _GEN_1271;
    end else begin
      validVec_21_2 <= _GEN_919;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_21_3 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_21_3 & _T_376) begin // @[StoreSet.scala 542:70]
      validVec_21_3 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_21_3 <= _GEN_2361;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_21_3 <= _GEN_1529;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1345) begin
      validVec_21_3 <= _GEN_1367;
    end else begin
      validVec_21_3 <= _GEN_1015;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_22_0 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_22_0 & _T_380) begin // @[StoreSet.scala 542:70]
      validVec_22_0 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_22_0 <= _GEN_2362;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_22_0 <= _GEN_1530;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1057) begin
      validVec_22_0 <= _GEN_1080;
    end else begin
      validVec_22_0 <= _GEN_728;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_22_1 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_22_1 & _T_384) begin // @[StoreSet.scala 542:70]
      validVec_22_1 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_22_1 <= _GEN_2363;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_22_1 <= _GEN_1531;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1153) begin
      validVec_22_1 <= _GEN_1176;
    end else begin
      validVec_22_1 <= _GEN_824;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_22_2 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_22_2 & _T_388) begin // @[StoreSet.scala 542:70]
      validVec_22_2 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_22_2 <= _GEN_2364;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_22_2 <= _GEN_1532;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1249) begin
      validVec_22_2 <= _GEN_1272;
    end else begin
      validVec_22_2 <= _GEN_920;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_22_3 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_22_3 & _T_392) begin // @[StoreSet.scala 542:70]
      validVec_22_3 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_22_3 <= _GEN_2365;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_22_3 <= _GEN_1533;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1345) begin
      validVec_22_3 <= _GEN_1368;
    end else begin
      validVec_22_3 <= _GEN_1016;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_23_0 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_23_0 & _T_396) begin // @[StoreSet.scala 542:70]
      validVec_23_0 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_23_0 <= _GEN_2366;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_23_0 <= _GEN_1534;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1057) begin
      validVec_23_0 <= _GEN_1081;
    end else begin
      validVec_23_0 <= _GEN_729;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_23_1 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_23_1 & _T_400) begin // @[StoreSet.scala 542:70]
      validVec_23_1 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_23_1 <= _GEN_2367;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_23_1 <= _GEN_1535;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1153) begin
      validVec_23_1 <= _GEN_1177;
    end else begin
      validVec_23_1 <= _GEN_825;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_23_2 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_23_2 & _T_404) begin // @[StoreSet.scala 542:70]
      validVec_23_2 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_23_2 <= _GEN_2368;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_23_2 <= _GEN_1536;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1249) begin
      validVec_23_2 <= _GEN_1273;
    end else begin
      validVec_23_2 <= _GEN_921;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_23_3 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_23_3 & _T_408) begin // @[StoreSet.scala 542:70]
      validVec_23_3 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_23_3 <= _GEN_2369;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_23_3 <= _GEN_1537;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1345) begin
      validVec_23_3 <= _GEN_1369;
    end else begin
      validVec_23_3 <= _GEN_1017;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_24_0 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_24_0 & _T_412) begin // @[StoreSet.scala 542:70]
      validVec_24_0 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_24_0 <= _GEN_2370;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_24_0 <= _GEN_1538;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1057) begin
      validVec_24_0 <= _GEN_1082;
    end else begin
      validVec_24_0 <= _GEN_730;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_24_1 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_24_1 & _T_416) begin // @[StoreSet.scala 542:70]
      validVec_24_1 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_24_1 <= _GEN_2371;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_24_1 <= _GEN_1539;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1153) begin
      validVec_24_1 <= _GEN_1178;
    end else begin
      validVec_24_1 <= _GEN_826;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_24_2 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_24_2 & _T_420) begin // @[StoreSet.scala 542:70]
      validVec_24_2 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_24_2 <= _GEN_2372;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_24_2 <= _GEN_1540;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1249) begin
      validVec_24_2 <= _GEN_1274;
    end else begin
      validVec_24_2 <= _GEN_922;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_24_3 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_24_3 & _T_424) begin // @[StoreSet.scala 542:70]
      validVec_24_3 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_24_3 <= _GEN_2373;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_24_3 <= _GEN_1541;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1345) begin
      validVec_24_3 <= _GEN_1370;
    end else begin
      validVec_24_3 <= _GEN_1018;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_25_0 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_25_0 & _T_428) begin // @[StoreSet.scala 542:70]
      validVec_25_0 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_25_0 <= _GEN_2374;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_25_0 <= _GEN_1542;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1057) begin
      validVec_25_0 <= _GEN_1083;
    end else begin
      validVec_25_0 <= _GEN_731;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_25_1 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_25_1 & _T_432) begin // @[StoreSet.scala 542:70]
      validVec_25_1 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_25_1 <= _GEN_2375;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_25_1 <= _GEN_1543;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1153) begin
      validVec_25_1 <= _GEN_1179;
    end else begin
      validVec_25_1 <= _GEN_827;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_25_2 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_25_2 & _T_436) begin // @[StoreSet.scala 542:70]
      validVec_25_2 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_25_2 <= _GEN_2376;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_25_2 <= _GEN_1544;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1249) begin
      validVec_25_2 <= _GEN_1275;
    end else begin
      validVec_25_2 <= _GEN_923;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_25_3 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_25_3 & _T_440) begin // @[StoreSet.scala 542:70]
      validVec_25_3 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_25_3 <= _GEN_2377;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_25_3 <= _GEN_1545;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1345) begin
      validVec_25_3 <= _GEN_1371;
    end else begin
      validVec_25_3 <= _GEN_1019;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_26_0 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_26_0 & _T_444) begin // @[StoreSet.scala 542:70]
      validVec_26_0 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_26_0 <= _GEN_2378;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_26_0 <= _GEN_1546;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1057) begin
      validVec_26_0 <= _GEN_1084;
    end else begin
      validVec_26_0 <= _GEN_732;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_26_1 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_26_1 & _T_448) begin // @[StoreSet.scala 542:70]
      validVec_26_1 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_26_1 <= _GEN_2379;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_26_1 <= _GEN_1547;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1153) begin
      validVec_26_1 <= _GEN_1180;
    end else begin
      validVec_26_1 <= _GEN_828;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_26_2 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_26_2 & _T_452) begin // @[StoreSet.scala 542:70]
      validVec_26_2 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_26_2 <= _GEN_2380;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_26_2 <= _GEN_1548;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1249) begin
      validVec_26_2 <= _GEN_1276;
    end else begin
      validVec_26_2 <= _GEN_924;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_26_3 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_26_3 & _T_456) begin // @[StoreSet.scala 542:70]
      validVec_26_3 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_26_3 <= _GEN_2381;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_26_3 <= _GEN_1549;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1345) begin
      validVec_26_3 <= _GEN_1372;
    end else begin
      validVec_26_3 <= _GEN_1020;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_27_0 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_27_0 & _T_460) begin // @[StoreSet.scala 542:70]
      validVec_27_0 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_27_0 <= _GEN_2382;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_27_0 <= _GEN_1550;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1057) begin
      validVec_27_0 <= _GEN_1085;
    end else begin
      validVec_27_0 <= _GEN_733;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_27_1 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_27_1 & _T_464) begin // @[StoreSet.scala 542:70]
      validVec_27_1 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_27_1 <= _GEN_2383;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_27_1 <= _GEN_1551;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1153) begin
      validVec_27_1 <= _GEN_1181;
    end else begin
      validVec_27_1 <= _GEN_829;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_27_2 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_27_2 & _T_468) begin // @[StoreSet.scala 542:70]
      validVec_27_2 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_27_2 <= _GEN_2384;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_27_2 <= _GEN_1552;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1249) begin
      validVec_27_2 <= _GEN_1277;
    end else begin
      validVec_27_2 <= _GEN_925;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_27_3 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_27_3 & _T_472) begin // @[StoreSet.scala 542:70]
      validVec_27_3 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_27_3 <= _GEN_2385;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_27_3 <= _GEN_1553;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1345) begin
      validVec_27_3 <= _GEN_1373;
    end else begin
      validVec_27_3 <= _GEN_1021;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_28_0 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_28_0 & _T_476) begin // @[StoreSet.scala 542:70]
      validVec_28_0 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_28_0 <= _GEN_2386;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_28_0 <= _GEN_1554;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1057) begin
      validVec_28_0 <= _GEN_1086;
    end else begin
      validVec_28_0 <= _GEN_734;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_28_1 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_28_1 & _T_480) begin // @[StoreSet.scala 542:70]
      validVec_28_1 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_28_1 <= _GEN_2387;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_28_1 <= _GEN_1555;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1153) begin
      validVec_28_1 <= _GEN_1182;
    end else begin
      validVec_28_1 <= _GEN_830;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_28_2 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_28_2 & _T_484) begin // @[StoreSet.scala 542:70]
      validVec_28_2 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_28_2 <= _GEN_2388;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_28_2 <= _GEN_1556;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1249) begin
      validVec_28_2 <= _GEN_1278;
    end else begin
      validVec_28_2 <= _GEN_926;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_28_3 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_28_3 & _T_488) begin // @[StoreSet.scala 542:70]
      validVec_28_3 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_28_3 <= _GEN_2389;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_28_3 <= _GEN_1557;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1345) begin
      validVec_28_3 <= _GEN_1374;
    end else begin
      validVec_28_3 <= _GEN_1022;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_29_0 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_29_0 & _T_492) begin // @[StoreSet.scala 542:70]
      validVec_29_0 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_29_0 <= _GEN_2390;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_29_0 <= _GEN_1558;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1057) begin
      validVec_29_0 <= _GEN_1087;
    end else begin
      validVec_29_0 <= _GEN_735;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_29_1 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_29_1 & _T_496) begin // @[StoreSet.scala 542:70]
      validVec_29_1 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_29_1 <= _GEN_2391;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_29_1 <= _GEN_1559;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1153) begin
      validVec_29_1 <= _GEN_1183;
    end else begin
      validVec_29_1 <= _GEN_831;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_29_2 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_29_2 & _T_500) begin // @[StoreSet.scala 542:70]
      validVec_29_2 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_29_2 <= _GEN_2392;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_29_2 <= _GEN_1560;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1249) begin
      validVec_29_2 <= _GEN_1279;
    end else begin
      validVec_29_2 <= _GEN_927;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_29_3 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_29_3 & _T_504) begin // @[StoreSet.scala 542:70]
      validVec_29_3 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_29_3 <= _GEN_2393;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_29_3 <= _GEN_1561;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1345) begin
      validVec_29_3 <= _GEN_1375;
    end else begin
      validVec_29_3 <= _GEN_1023;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_30_0 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_30_0 & _T_508) begin // @[StoreSet.scala 542:70]
      validVec_30_0 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_30_0 <= _GEN_2394;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_30_0 <= _GEN_1562;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1057) begin
      validVec_30_0 <= _GEN_1088;
    end else begin
      validVec_30_0 <= _GEN_736;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_30_1 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_30_1 & _T_512) begin // @[StoreSet.scala 542:70]
      validVec_30_1 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_30_1 <= _GEN_2395;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_30_1 <= _GEN_1563;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1153) begin
      validVec_30_1 <= _GEN_1184;
    end else begin
      validVec_30_1 <= _GEN_832;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_30_2 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_30_2 & _T_516) begin // @[StoreSet.scala 542:70]
      validVec_30_2 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_30_2 <= _GEN_2396;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_30_2 <= _GEN_1564;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1249) begin
      validVec_30_2 <= _GEN_1280;
    end else begin
      validVec_30_2 <= _GEN_928;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_30_3 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_30_3 & _T_520) begin // @[StoreSet.scala 542:70]
      validVec_30_3 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_30_3 <= _GEN_2397;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_30_3 <= _GEN_1565;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1345) begin
      validVec_30_3 <= _GEN_1376;
    end else begin
      validVec_30_3 <= _GEN_1024;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_31_0 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_31_0 & _T_524) begin // @[StoreSet.scala 542:70]
      validVec_31_0 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_31_0 <= _GEN_2398;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_31_0 <= _GEN_1566;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1057) begin
      validVec_31_0 <= _GEN_1089;
    end else begin
      validVec_31_0 <= _GEN_737;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_31_1 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_31_1 & _T_528) begin // @[StoreSet.scala 542:70]
      validVec_31_1 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_31_1 <= _GEN_2399;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_31_1 <= _GEN_1567;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1153) begin
      validVec_31_1 <= _GEN_1185;
    end else begin
      validVec_31_1 <= _GEN_833;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_31_2 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_31_2 & _T_532) begin // @[StoreSet.scala 542:70]
      validVec_31_2 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_31_2 <= _GEN_2400;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_31_2 <= _GEN_1568;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1249) begin
      validVec_31_2 <= _GEN_1281;
    end else begin
      validVec_31_2 <= _GEN_929;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 554:69]
      validVec_31_3 <= 1'h0; // @[StoreSet.scala 555:24]
    end else if (validVec_31_3 & _T_536) begin // @[StoreSet.scala 542:70]
      validVec_31_3 <= 1'h0;
    end else if (io_dispatch_req_1_valid & io_dispatch_req_1_bits_isstore) begin // @[StoreSet.scala 542:70]
      validVec_31_3 <= _GEN_2401;
    end else if (_hitInDispatchBundleVec_T) begin // @[StoreSet.scala 534:179]
      validVec_31_3 <= _GEN_1569;
    end else if (io_storeIssue_1_valid & io_storeIssue_1_bits_uop_cf_storeSetHit & io_storeIssue_1_bits_uop_robIdx_value
       == _GEN_1345) begin
      validVec_31_3 <= _GEN_1377;
    end else begin
      validVec_31_3 <= _GEN_1025;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 493:25]
      allocPtr_0 <= 2'h0; // @[StoreSet.scala 493:25]
    end else begin
      allocPtr_0 <= _GEN_3842[1:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 493:25]
      allocPtr_1 <= 2'h0; // @[StoreSet.scala 493:25]
    end else begin
      allocPtr_1 <= _GEN_3843[1:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 493:25]
      allocPtr_2 <= 2'h0; // @[StoreSet.scala 493:25]
    end else begin
      allocPtr_2 <= _GEN_3844[1:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 493:25]
      allocPtr_3 <= 2'h0; // @[StoreSet.scala 493:25]
    end else begin
      allocPtr_3 <= _GEN_3845[1:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 493:25]
      allocPtr_4 <= 2'h0; // @[StoreSet.scala 493:25]
    end else begin
      allocPtr_4 <= _GEN_3846[1:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 493:25]
      allocPtr_5 <= 2'h0; // @[StoreSet.scala 493:25]
    end else begin
      allocPtr_5 <= _GEN_3847[1:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 493:25]
      allocPtr_6 <= 2'h0; // @[StoreSet.scala 493:25]
    end else begin
      allocPtr_6 <= _GEN_3848[1:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 493:25]
      allocPtr_7 <= 2'h0; // @[StoreSet.scala 493:25]
    end else begin
      allocPtr_7 <= _GEN_3849[1:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 493:25]
      allocPtr_8 <= 2'h0; // @[StoreSet.scala 493:25]
    end else begin
      allocPtr_8 <= _GEN_3850[1:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 493:25]
      allocPtr_9 <= 2'h0; // @[StoreSet.scala 493:25]
    end else begin
      allocPtr_9 <= _GEN_3851[1:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 493:25]
      allocPtr_10 <= 2'h0; // @[StoreSet.scala 493:25]
    end else begin
      allocPtr_10 <= _GEN_3852[1:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 493:25]
      allocPtr_11 <= 2'h0; // @[StoreSet.scala 493:25]
    end else begin
      allocPtr_11 <= _GEN_3853[1:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 493:25]
      allocPtr_12 <= 2'h0; // @[StoreSet.scala 493:25]
    end else begin
      allocPtr_12 <= _GEN_3854[1:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 493:25]
      allocPtr_13 <= 2'h0; // @[StoreSet.scala 493:25]
    end else begin
      allocPtr_13 <= _GEN_3855[1:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 493:25]
      allocPtr_14 <= 2'h0; // @[StoreSet.scala 493:25]
    end else begin
      allocPtr_14 <= _GEN_3856[1:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 493:25]
      allocPtr_15 <= 2'h0; // @[StoreSet.scala 493:25]
    end else begin
      allocPtr_15 <= _GEN_3857[1:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 493:25]
      allocPtr_16 <= 2'h0; // @[StoreSet.scala 493:25]
    end else begin
      allocPtr_16 <= _GEN_3858[1:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 493:25]
      allocPtr_17 <= 2'h0; // @[StoreSet.scala 493:25]
    end else begin
      allocPtr_17 <= _GEN_3859[1:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 493:25]
      allocPtr_18 <= 2'h0; // @[StoreSet.scala 493:25]
    end else begin
      allocPtr_18 <= _GEN_3860[1:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 493:25]
      allocPtr_19 <= 2'h0; // @[StoreSet.scala 493:25]
    end else begin
      allocPtr_19 <= _GEN_3861[1:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 493:25]
      allocPtr_20 <= 2'h0; // @[StoreSet.scala 493:25]
    end else begin
      allocPtr_20 <= _GEN_3862[1:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 493:25]
      allocPtr_21 <= 2'h0; // @[StoreSet.scala 493:25]
    end else begin
      allocPtr_21 <= _GEN_3863[1:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 493:25]
      allocPtr_22 <= 2'h0; // @[StoreSet.scala 493:25]
    end else begin
      allocPtr_22 <= _GEN_3864[1:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 493:25]
      allocPtr_23 <= 2'h0; // @[StoreSet.scala 493:25]
    end else begin
      allocPtr_23 <= _GEN_3865[1:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 493:25]
      allocPtr_24 <= 2'h0; // @[StoreSet.scala 493:25]
    end else begin
      allocPtr_24 <= _GEN_3866[1:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 493:25]
      allocPtr_25 <= 2'h0; // @[StoreSet.scala 493:25]
    end else begin
      allocPtr_25 <= _GEN_3867[1:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 493:25]
      allocPtr_26 <= 2'h0; // @[StoreSet.scala 493:25]
    end else begin
      allocPtr_26 <= _GEN_3868[1:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 493:25]
      allocPtr_27 <= 2'h0; // @[StoreSet.scala 493:25]
    end else begin
      allocPtr_27 <= _GEN_3869[1:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 493:25]
      allocPtr_28 <= 2'h0; // @[StoreSet.scala 493:25]
    end else begin
      allocPtr_28 <= _GEN_3870[1:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 493:25]
      allocPtr_29 <= 2'h0; // @[StoreSet.scala 493:25]
    end else begin
      allocPtr_29 <= _GEN_3871[1:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 493:25]
      allocPtr_30 <= 2'h0; // @[StoreSet.scala 493:25]
    end else begin
      allocPtr_30 <= _GEN_3872[1:0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[StoreSet.scala 493:25]
      allocPtr_31 <= 2'h0; // @[StoreSet.scala 493:25]
    end else begin
      allocPtr_31 <= _GEN_3873[1:0];
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  validVec_0_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  validVec_0_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  validVec_0_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  validVec_0_3 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  validVec_1_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  validVec_1_1 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  validVec_1_2 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  validVec_1_3 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  validVec_2_0 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  validVec_2_1 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  validVec_2_2 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  validVec_2_3 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  validVec_3_0 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  validVec_3_1 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  validVec_3_2 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  validVec_3_3 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  validVec_4_0 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  validVec_4_1 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  validVec_4_2 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  validVec_4_3 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  validVec_5_0 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  validVec_5_1 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  validVec_5_2 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  validVec_5_3 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  validVec_6_0 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  validVec_6_1 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  validVec_6_2 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  validVec_6_3 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  validVec_7_0 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  validVec_7_1 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  validVec_7_2 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  validVec_7_3 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  validVec_8_0 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  validVec_8_1 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  validVec_8_2 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  validVec_8_3 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  validVec_9_0 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  validVec_9_1 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  validVec_9_2 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  validVec_9_3 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  validVec_10_0 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  validVec_10_1 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  validVec_10_2 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  validVec_10_3 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  validVec_11_0 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  validVec_11_1 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  validVec_11_2 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  validVec_11_3 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  validVec_12_0 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  validVec_12_1 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  validVec_12_2 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  validVec_12_3 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  validVec_13_0 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  validVec_13_1 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  validVec_13_2 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  validVec_13_3 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  validVec_14_0 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  validVec_14_1 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  validVec_14_2 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  validVec_14_3 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  validVec_15_0 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  validVec_15_1 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  validVec_15_2 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  validVec_15_3 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  validVec_16_0 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  validVec_16_1 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  validVec_16_2 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  validVec_16_3 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  validVec_17_0 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  validVec_17_1 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  validVec_17_2 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  validVec_17_3 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  validVec_18_0 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  validVec_18_1 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  validVec_18_2 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  validVec_18_3 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  validVec_19_0 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  validVec_19_1 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  validVec_19_2 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  validVec_19_3 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  validVec_20_0 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  validVec_20_1 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  validVec_20_2 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  validVec_20_3 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  validVec_21_0 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  validVec_21_1 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  validVec_21_2 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  validVec_21_3 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  validVec_22_0 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  validVec_22_1 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  validVec_22_2 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  validVec_22_3 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  validVec_23_0 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  validVec_23_1 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  validVec_23_2 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  validVec_23_3 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  validVec_24_0 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  validVec_24_1 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  validVec_24_2 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  validVec_24_3 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  validVec_25_0 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  validVec_25_1 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  validVec_25_2 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  validVec_25_3 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  validVec_26_0 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  validVec_26_1 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  validVec_26_2 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  validVec_26_3 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  validVec_27_0 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  validVec_27_1 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  validVec_27_2 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  validVec_27_3 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  validVec_28_0 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  validVec_28_1 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  validVec_28_2 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  validVec_28_3 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  validVec_29_0 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  validVec_29_1 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  validVec_29_2 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  validVec_29_3 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  validVec_30_0 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  validVec_30_1 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  validVec_30_2 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  validVec_30_3 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  validVec_31_0 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  validVec_31_1 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  validVec_31_2 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  validVec_31_3 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  robIdxVec_0_0_flag = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  robIdxVec_0_0_value = _RAND_129[4:0];
  _RAND_130 = {1{`RANDOM}};
  robIdxVec_0_1_flag = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  robIdxVec_0_1_value = _RAND_131[4:0];
  _RAND_132 = {1{`RANDOM}};
  robIdxVec_0_2_flag = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  robIdxVec_0_2_value = _RAND_133[4:0];
  _RAND_134 = {1{`RANDOM}};
  robIdxVec_0_3_flag = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  robIdxVec_0_3_value = _RAND_135[4:0];
  _RAND_136 = {1{`RANDOM}};
  robIdxVec_1_0_flag = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  robIdxVec_1_0_value = _RAND_137[4:0];
  _RAND_138 = {1{`RANDOM}};
  robIdxVec_1_1_flag = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  robIdxVec_1_1_value = _RAND_139[4:0];
  _RAND_140 = {1{`RANDOM}};
  robIdxVec_1_2_flag = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  robIdxVec_1_2_value = _RAND_141[4:0];
  _RAND_142 = {1{`RANDOM}};
  robIdxVec_1_3_flag = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  robIdxVec_1_3_value = _RAND_143[4:0];
  _RAND_144 = {1{`RANDOM}};
  robIdxVec_2_0_flag = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  robIdxVec_2_0_value = _RAND_145[4:0];
  _RAND_146 = {1{`RANDOM}};
  robIdxVec_2_1_flag = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  robIdxVec_2_1_value = _RAND_147[4:0];
  _RAND_148 = {1{`RANDOM}};
  robIdxVec_2_2_flag = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  robIdxVec_2_2_value = _RAND_149[4:0];
  _RAND_150 = {1{`RANDOM}};
  robIdxVec_2_3_flag = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  robIdxVec_2_3_value = _RAND_151[4:0];
  _RAND_152 = {1{`RANDOM}};
  robIdxVec_3_0_flag = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  robIdxVec_3_0_value = _RAND_153[4:0];
  _RAND_154 = {1{`RANDOM}};
  robIdxVec_3_1_flag = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  robIdxVec_3_1_value = _RAND_155[4:0];
  _RAND_156 = {1{`RANDOM}};
  robIdxVec_3_2_flag = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  robIdxVec_3_2_value = _RAND_157[4:0];
  _RAND_158 = {1{`RANDOM}};
  robIdxVec_3_3_flag = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  robIdxVec_3_3_value = _RAND_159[4:0];
  _RAND_160 = {1{`RANDOM}};
  robIdxVec_4_0_flag = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  robIdxVec_4_0_value = _RAND_161[4:0];
  _RAND_162 = {1{`RANDOM}};
  robIdxVec_4_1_flag = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  robIdxVec_4_1_value = _RAND_163[4:0];
  _RAND_164 = {1{`RANDOM}};
  robIdxVec_4_2_flag = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  robIdxVec_4_2_value = _RAND_165[4:0];
  _RAND_166 = {1{`RANDOM}};
  robIdxVec_4_3_flag = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  robIdxVec_4_3_value = _RAND_167[4:0];
  _RAND_168 = {1{`RANDOM}};
  robIdxVec_5_0_flag = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  robIdxVec_5_0_value = _RAND_169[4:0];
  _RAND_170 = {1{`RANDOM}};
  robIdxVec_5_1_flag = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  robIdxVec_5_1_value = _RAND_171[4:0];
  _RAND_172 = {1{`RANDOM}};
  robIdxVec_5_2_flag = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  robIdxVec_5_2_value = _RAND_173[4:0];
  _RAND_174 = {1{`RANDOM}};
  robIdxVec_5_3_flag = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  robIdxVec_5_3_value = _RAND_175[4:0];
  _RAND_176 = {1{`RANDOM}};
  robIdxVec_6_0_flag = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  robIdxVec_6_0_value = _RAND_177[4:0];
  _RAND_178 = {1{`RANDOM}};
  robIdxVec_6_1_flag = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  robIdxVec_6_1_value = _RAND_179[4:0];
  _RAND_180 = {1{`RANDOM}};
  robIdxVec_6_2_flag = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  robIdxVec_6_2_value = _RAND_181[4:0];
  _RAND_182 = {1{`RANDOM}};
  robIdxVec_6_3_flag = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  robIdxVec_6_3_value = _RAND_183[4:0];
  _RAND_184 = {1{`RANDOM}};
  robIdxVec_7_0_flag = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  robIdxVec_7_0_value = _RAND_185[4:0];
  _RAND_186 = {1{`RANDOM}};
  robIdxVec_7_1_flag = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  robIdxVec_7_1_value = _RAND_187[4:0];
  _RAND_188 = {1{`RANDOM}};
  robIdxVec_7_2_flag = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  robIdxVec_7_2_value = _RAND_189[4:0];
  _RAND_190 = {1{`RANDOM}};
  robIdxVec_7_3_flag = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  robIdxVec_7_3_value = _RAND_191[4:0];
  _RAND_192 = {1{`RANDOM}};
  robIdxVec_8_0_flag = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  robIdxVec_8_0_value = _RAND_193[4:0];
  _RAND_194 = {1{`RANDOM}};
  robIdxVec_8_1_flag = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  robIdxVec_8_1_value = _RAND_195[4:0];
  _RAND_196 = {1{`RANDOM}};
  robIdxVec_8_2_flag = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  robIdxVec_8_2_value = _RAND_197[4:0];
  _RAND_198 = {1{`RANDOM}};
  robIdxVec_8_3_flag = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  robIdxVec_8_3_value = _RAND_199[4:0];
  _RAND_200 = {1{`RANDOM}};
  robIdxVec_9_0_flag = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  robIdxVec_9_0_value = _RAND_201[4:0];
  _RAND_202 = {1{`RANDOM}};
  robIdxVec_9_1_flag = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  robIdxVec_9_1_value = _RAND_203[4:0];
  _RAND_204 = {1{`RANDOM}};
  robIdxVec_9_2_flag = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  robIdxVec_9_2_value = _RAND_205[4:0];
  _RAND_206 = {1{`RANDOM}};
  robIdxVec_9_3_flag = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  robIdxVec_9_3_value = _RAND_207[4:0];
  _RAND_208 = {1{`RANDOM}};
  robIdxVec_10_0_flag = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  robIdxVec_10_0_value = _RAND_209[4:0];
  _RAND_210 = {1{`RANDOM}};
  robIdxVec_10_1_flag = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  robIdxVec_10_1_value = _RAND_211[4:0];
  _RAND_212 = {1{`RANDOM}};
  robIdxVec_10_2_flag = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  robIdxVec_10_2_value = _RAND_213[4:0];
  _RAND_214 = {1{`RANDOM}};
  robIdxVec_10_3_flag = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  robIdxVec_10_3_value = _RAND_215[4:0];
  _RAND_216 = {1{`RANDOM}};
  robIdxVec_11_0_flag = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  robIdxVec_11_0_value = _RAND_217[4:0];
  _RAND_218 = {1{`RANDOM}};
  robIdxVec_11_1_flag = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  robIdxVec_11_1_value = _RAND_219[4:0];
  _RAND_220 = {1{`RANDOM}};
  robIdxVec_11_2_flag = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  robIdxVec_11_2_value = _RAND_221[4:0];
  _RAND_222 = {1{`RANDOM}};
  robIdxVec_11_3_flag = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  robIdxVec_11_3_value = _RAND_223[4:0];
  _RAND_224 = {1{`RANDOM}};
  robIdxVec_12_0_flag = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  robIdxVec_12_0_value = _RAND_225[4:0];
  _RAND_226 = {1{`RANDOM}};
  robIdxVec_12_1_flag = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  robIdxVec_12_1_value = _RAND_227[4:0];
  _RAND_228 = {1{`RANDOM}};
  robIdxVec_12_2_flag = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  robIdxVec_12_2_value = _RAND_229[4:0];
  _RAND_230 = {1{`RANDOM}};
  robIdxVec_12_3_flag = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  robIdxVec_12_3_value = _RAND_231[4:0];
  _RAND_232 = {1{`RANDOM}};
  robIdxVec_13_0_flag = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  robIdxVec_13_0_value = _RAND_233[4:0];
  _RAND_234 = {1{`RANDOM}};
  robIdxVec_13_1_flag = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  robIdxVec_13_1_value = _RAND_235[4:0];
  _RAND_236 = {1{`RANDOM}};
  robIdxVec_13_2_flag = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  robIdxVec_13_2_value = _RAND_237[4:0];
  _RAND_238 = {1{`RANDOM}};
  robIdxVec_13_3_flag = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  robIdxVec_13_3_value = _RAND_239[4:0];
  _RAND_240 = {1{`RANDOM}};
  robIdxVec_14_0_flag = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  robIdxVec_14_0_value = _RAND_241[4:0];
  _RAND_242 = {1{`RANDOM}};
  robIdxVec_14_1_flag = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  robIdxVec_14_1_value = _RAND_243[4:0];
  _RAND_244 = {1{`RANDOM}};
  robIdxVec_14_2_flag = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  robIdxVec_14_2_value = _RAND_245[4:0];
  _RAND_246 = {1{`RANDOM}};
  robIdxVec_14_3_flag = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  robIdxVec_14_3_value = _RAND_247[4:0];
  _RAND_248 = {1{`RANDOM}};
  robIdxVec_15_0_flag = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  robIdxVec_15_0_value = _RAND_249[4:0];
  _RAND_250 = {1{`RANDOM}};
  robIdxVec_15_1_flag = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  robIdxVec_15_1_value = _RAND_251[4:0];
  _RAND_252 = {1{`RANDOM}};
  robIdxVec_15_2_flag = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  robIdxVec_15_2_value = _RAND_253[4:0];
  _RAND_254 = {1{`RANDOM}};
  robIdxVec_15_3_flag = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  robIdxVec_15_3_value = _RAND_255[4:0];
  _RAND_256 = {1{`RANDOM}};
  robIdxVec_16_0_flag = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  robIdxVec_16_0_value = _RAND_257[4:0];
  _RAND_258 = {1{`RANDOM}};
  robIdxVec_16_1_flag = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  robIdxVec_16_1_value = _RAND_259[4:0];
  _RAND_260 = {1{`RANDOM}};
  robIdxVec_16_2_flag = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  robIdxVec_16_2_value = _RAND_261[4:0];
  _RAND_262 = {1{`RANDOM}};
  robIdxVec_16_3_flag = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  robIdxVec_16_3_value = _RAND_263[4:0];
  _RAND_264 = {1{`RANDOM}};
  robIdxVec_17_0_flag = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  robIdxVec_17_0_value = _RAND_265[4:0];
  _RAND_266 = {1{`RANDOM}};
  robIdxVec_17_1_flag = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  robIdxVec_17_1_value = _RAND_267[4:0];
  _RAND_268 = {1{`RANDOM}};
  robIdxVec_17_2_flag = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  robIdxVec_17_2_value = _RAND_269[4:0];
  _RAND_270 = {1{`RANDOM}};
  robIdxVec_17_3_flag = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  robIdxVec_17_3_value = _RAND_271[4:0];
  _RAND_272 = {1{`RANDOM}};
  robIdxVec_18_0_flag = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  robIdxVec_18_0_value = _RAND_273[4:0];
  _RAND_274 = {1{`RANDOM}};
  robIdxVec_18_1_flag = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  robIdxVec_18_1_value = _RAND_275[4:0];
  _RAND_276 = {1{`RANDOM}};
  robIdxVec_18_2_flag = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  robIdxVec_18_2_value = _RAND_277[4:0];
  _RAND_278 = {1{`RANDOM}};
  robIdxVec_18_3_flag = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  robIdxVec_18_3_value = _RAND_279[4:0];
  _RAND_280 = {1{`RANDOM}};
  robIdxVec_19_0_flag = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  robIdxVec_19_0_value = _RAND_281[4:0];
  _RAND_282 = {1{`RANDOM}};
  robIdxVec_19_1_flag = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  robIdxVec_19_1_value = _RAND_283[4:0];
  _RAND_284 = {1{`RANDOM}};
  robIdxVec_19_2_flag = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  robIdxVec_19_2_value = _RAND_285[4:0];
  _RAND_286 = {1{`RANDOM}};
  robIdxVec_19_3_flag = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  robIdxVec_19_3_value = _RAND_287[4:0];
  _RAND_288 = {1{`RANDOM}};
  robIdxVec_20_0_flag = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  robIdxVec_20_0_value = _RAND_289[4:0];
  _RAND_290 = {1{`RANDOM}};
  robIdxVec_20_1_flag = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  robIdxVec_20_1_value = _RAND_291[4:0];
  _RAND_292 = {1{`RANDOM}};
  robIdxVec_20_2_flag = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  robIdxVec_20_2_value = _RAND_293[4:0];
  _RAND_294 = {1{`RANDOM}};
  robIdxVec_20_3_flag = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  robIdxVec_20_3_value = _RAND_295[4:0];
  _RAND_296 = {1{`RANDOM}};
  robIdxVec_21_0_flag = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  robIdxVec_21_0_value = _RAND_297[4:0];
  _RAND_298 = {1{`RANDOM}};
  robIdxVec_21_1_flag = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  robIdxVec_21_1_value = _RAND_299[4:0];
  _RAND_300 = {1{`RANDOM}};
  robIdxVec_21_2_flag = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  robIdxVec_21_2_value = _RAND_301[4:0];
  _RAND_302 = {1{`RANDOM}};
  robIdxVec_21_3_flag = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  robIdxVec_21_3_value = _RAND_303[4:0];
  _RAND_304 = {1{`RANDOM}};
  robIdxVec_22_0_flag = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  robIdxVec_22_0_value = _RAND_305[4:0];
  _RAND_306 = {1{`RANDOM}};
  robIdxVec_22_1_flag = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  robIdxVec_22_1_value = _RAND_307[4:0];
  _RAND_308 = {1{`RANDOM}};
  robIdxVec_22_2_flag = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  robIdxVec_22_2_value = _RAND_309[4:0];
  _RAND_310 = {1{`RANDOM}};
  robIdxVec_22_3_flag = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  robIdxVec_22_3_value = _RAND_311[4:0];
  _RAND_312 = {1{`RANDOM}};
  robIdxVec_23_0_flag = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  robIdxVec_23_0_value = _RAND_313[4:0];
  _RAND_314 = {1{`RANDOM}};
  robIdxVec_23_1_flag = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  robIdxVec_23_1_value = _RAND_315[4:0];
  _RAND_316 = {1{`RANDOM}};
  robIdxVec_23_2_flag = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  robIdxVec_23_2_value = _RAND_317[4:0];
  _RAND_318 = {1{`RANDOM}};
  robIdxVec_23_3_flag = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  robIdxVec_23_3_value = _RAND_319[4:0];
  _RAND_320 = {1{`RANDOM}};
  robIdxVec_24_0_flag = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  robIdxVec_24_0_value = _RAND_321[4:0];
  _RAND_322 = {1{`RANDOM}};
  robIdxVec_24_1_flag = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  robIdxVec_24_1_value = _RAND_323[4:0];
  _RAND_324 = {1{`RANDOM}};
  robIdxVec_24_2_flag = _RAND_324[0:0];
  _RAND_325 = {1{`RANDOM}};
  robIdxVec_24_2_value = _RAND_325[4:0];
  _RAND_326 = {1{`RANDOM}};
  robIdxVec_24_3_flag = _RAND_326[0:0];
  _RAND_327 = {1{`RANDOM}};
  robIdxVec_24_3_value = _RAND_327[4:0];
  _RAND_328 = {1{`RANDOM}};
  robIdxVec_25_0_flag = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  robIdxVec_25_0_value = _RAND_329[4:0];
  _RAND_330 = {1{`RANDOM}};
  robIdxVec_25_1_flag = _RAND_330[0:0];
  _RAND_331 = {1{`RANDOM}};
  robIdxVec_25_1_value = _RAND_331[4:0];
  _RAND_332 = {1{`RANDOM}};
  robIdxVec_25_2_flag = _RAND_332[0:0];
  _RAND_333 = {1{`RANDOM}};
  robIdxVec_25_2_value = _RAND_333[4:0];
  _RAND_334 = {1{`RANDOM}};
  robIdxVec_25_3_flag = _RAND_334[0:0];
  _RAND_335 = {1{`RANDOM}};
  robIdxVec_25_3_value = _RAND_335[4:0];
  _RAND_336 = {1{`RANDOM}};
  robIdxVec_26_0_flag = _RAND_336[0:0];
  _RAND_337 = {1{`RANDOM}};
  robIdxVec_26_0_value = _RAND_337[4:0];
  _RAND_338 = {1{`RANDOM}};
  robIdxVec_26_1_flag = _RAND_338[0:0];
  _RAND_339 = {1{`RANDOM}};
  robIdxVec_26_1_value = _RAND_339[4:0];
  _RAND_340 = {1{`RANDOM}};
  robIdxVec_26_2_flag = _RAND_340[0:0];
  _RAND_341 = {1{`RANDOM}};
  robIdxVec_26_2_value = _RAND_341[4:0];
  _RAND_342 = {1{`RANDOM}};
  robIdxVec_26_3_flag = _RAND_342[0:0];
  _RAND_343 = {1{`RANDOM}};
  robIdxVec_26_3_value = _RAND_343[4:0];
  _RAND_344 = {1{`RANDOM}};
  robIdxVec_27_0_flag = _RAND_344[0:0];
  _RAND_345 = {1{`RANDOM}};
  robIdxVec_27_0_value = _RAND_345[4:0];
  _RAND_346 = {1{`RANDOM}};
  robIdxVec_27_1_flag = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  robIdxVec_27_1_value = _RAND_347[4:0];
  _RAND_348 = {1{`RANDOM}};
  robIdxVec_27_2_flag = _RAND_348[0:0];
  _RAND_349 = {1{`RANDOM}};
  robIdxVec_27_2_value = _RAND_349[4:0];
  _RAND_350 = {1{`RANDOM}};
  robIdxVec_27_3_flag = _RAND_350[0:0];
  _RAND_351 = {1{`RANDOM}};
  robIdxVec_27_3_value = _RAND_351[4:0];
  _RAND_352 = {1{`RANDOM}};
  robIdxVec_28_0_flag = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  robIdxVec_28_0_value = _RAND_353[4:0];
  _RAND_354 = {1{`RANDOM}};
  robIdxVec_28_1_flag = _RAND_354[0:0];
  _RAND_355 = {1{`RANDOM}};
  robIdxVec_28_1_value = _RAND_355[4:0];
  _RAND_356 = {1{`RANDOM}};
  robIdxVec_28_2_flag = _RAND_356[0:0];
  _RAND_357 = {1{`RANDOM}};
  robIdxVec_28_2_value = _RAND_357[4:0];
  _RAND_358 = {1{`RANDOM}};
  robIdxVec_28_3_flag = _RAND_358[0:0];
  _RAND_359 = {1{`RANDOM}};
  robIdxVec_28_3_value = _RAND_359[4:0];
  _RAND_360 = {1{`RANDOM}};
  robIdxVec_29_0_flag = _RAND_360[0:0];
  _RAND_361 = {1{`RANDOM}};
  robIdxVec_29_0_value = _RAND_361[4:0];
  _RAND_362 = {1{`RANDOM}};
  robIdxVec_29_1_flag = _RAND_362[0:0];
  _RAND_363 = {1{`RANDOM}};
  robIdxVec_29_1_value = _RAND_363[4:0];
  _RAND_364 = {1{`RANDOM}};
  robIdxVec_29_2_flag = _RAND_364[0:0];
  _RAND_365 = {1{`RANDOM}};
  robIdxVec_29_2_value = _RAND_365[4:0];
  _RAND_366 = {1{`RANDOM}};
  robIdxVec_29_3_flag = _RAND_366[0:0];
  _RAND_367 = {1{`RANDOM}};
  robIdxVec_29_3_value = _RAND_367[4:0];
  _RAND_368 = {1{`RANDOM}};
  robIdxVec_30_0_flag = _RAND_368[0:0];
  _RAND_369 = {1{`RANDOM}};
  robIdxVec_30_0_value = _RAND_369[4:0];
  _RAND_370 = {1{`RANDOM}};
  robIdxVec_30_1_flag = _RAND_370[0:0];
  _RAND_371 = {1{`RANDOM}};
  robIdxVec_30_1_value = _RAND_371[4:0];
  _RAND_372 = {1{`RANDOM}};
  robIdxVec_30_2_flag = _RAND_372[0:0];
  _RAND_373 = {1{`RANDOM}};
  robIdxVec_30_2_value = _RAND_373[4:0];
  _RAND_374 = {1{`RANDOM}};
  robIdxVec_30_3_flag = _RAND_374[0:0];
  _RAND_375 = {1{`RANDOM}};
  robIdxVec_30_3_value = _RAND_375[4:0];
  _RAND_376 = {1{`RANDOM}};
  robIdxVec_31_0_flag = _RAND_376[0:0];
  _RAND_377 = {1{`RANDOM}};
  robIdxVec_31_0_value = _RAND_377[4:0];
  _RAND_378 = {1{`RANDOM}};
  robIdxVec_31_1_flag = _RAND_378[0:0];
  _RAND_379 = {1{`RANDOM}};
  robIdxVec_31_1_value = _RAND_379[4:0];
  _RAND_380 = {1{`RANDOM}};
  robIdxVec_31_2_flag = _RAND_380[0:0];
  _RAND_381 = {1{`RANDOM}};
  robIdxVec_31_2_value = _RAND_381[4:0];
  _RAND_382 = {1{`RANDOM}};
  robIdxVec_31_3_flag = _RAND_382[0:0];
  _RAND_383 = {1{`RANDOM}};
  robIdxVec_31_3_value = _RAND_383[4:0];
  _RAND_384 = {1{`RANDOM}};
  allocPtr_0 = _RAND_384[1:0];
  _RAND_385 = {1{`RANDOM}};
  allocPtr_1 = _RAND_385[1:0];
  _RAND_386 = {1{`RANDOM}};
  allocPtr_2 = _RAND_386[1:0];
  _RAND_387 = {1{`RANDOM}};
  allocPtr_3 = _RAND_387[1:0];
  _RAND_388 = {1{`RANDOM}};
  allocPtr_4 = _RAND_388[1:0];
  _RAND_389 = {1{`RANDOM}};
  allocPtr_5 = _RAND_389[1:0];
  _RAND_390 = {1{`RANDOM}};
  allocPtr_6 = _RAND_390[1:0];
  _RAND_391 = {1{`RANDOM}};
  allocPtr_7 = _RAND_391[1:0];
  _RAND_392 = {1{`RANDOM}};
  allocPtr_8 = _RAND_392[1:0];
  _RAND_393 = {1{`RANDOM}};
  allocPtr_9 = _RAND_393[1:0];
  _RAND_394 = {1{`RANDOM}};
  allocPtr_10 = _RAND_394[1:0];
  _RAND_395 = {1{`RANDOM}};
  allocPtr_11 = _RAND_395[1:0];
  _RAND_396 = {1{`RANDOM}};
  allocPtr_12 = _RAND_396[1:0];
  _RAND_397 = {1{`RANDOM}};
  allocPtr_13 = _RAND_397[1:0];
  _RAND_398 = {1{`RANDOM}};
  allocPtr_14 = _RAND_398[1:0];
  _RAND_399 = {1{`RANDOM}};
  allocPtr_15 = _RAND_399[1:0];
  _RAND_400 = {1{`RANDOM}};
  allocPtr_16 = _RAND_400[1:0];
  _RAND_401 = {1{`RANDOM}};
  allocPtr_17 = _RAND_401[1:0];
  _RAND_402 = {1{`RANDOM}};
  allocPtr_18 = _RAND_402[1:0];
  _RAND_403 = {1{`RANDOM}};
  allocPtr_19 = _RAND_403[1:0];
  _RAND_404 = {1{`RANDOM}};
  allocPtr_20 = _RAND_404[1:0];
  _RAND_405 = {1{`RANDOM}};
  allocPtr_21 = _RAND_405[1:0];
  _RAND_406 = {1{`RANDOM}};
  allocPtr_22 = _RAND_406[1:0];
  _RAND_407 = {1{`RANDOM}};
  allocPtr_23 = _RAND_407[1:0];
  _RAND_408 = {1{`RANDOM}};
  allocPtr_24 = _RAND_408[1:0];
  _RAND_409 = {1{`RANDOM}};
  allocPtr_25 = _RAND_409[1:0];
  _RAND_410 = {1{`RANDOM}};
  allocPtr_26 = _RAND_410[1:0];
  _RAND_411 = {1{`RANDOM}};
  allocPtr_27 = _RAND_411[1:0];
  _RAND_412 = {1{`RANDOM}};
  allocPtr_28 = _RAND_412[1:0];
  _RAND_413 = {1{`RANDOM}};
  allocPtr_29 = _RAND_413[1:0];
  _RAND_414 = {1{`RANDOM}};
  allocPtr_30 = _RAND_414[1:0];
  _RAND_415 = {1{`RANDOM}};
  allocPtr_31 = _RAND_415[1:0];
  _RAND_416 = {1{`RANDOM}};
  REG = _RAND_416[0:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    validVec_0_0 = 1'h0;
  end
  if (reset) begin
    validVec_0_1 = 1'h0;
  end
  if (reset) begin
    validVec_0_2 = 1'h0;
  end
  if (reset) begin
    validVec_0_3 = 1'h0;
  end
  if (reset) begin
    validVec_1_0 = 1'h0;
  end
  if (reset) begin
    validVec_1_1 = 1'h0;
  end
  if (reset) begin
    validVec_1_2 = 1'h0;
  end
  if (reset) begin
    validVec_1_3 = 1'h0;
  end
  if (reset) begin
    validVec_2_0 = 1'h0;
  end
  if (reset) begin
    validVec_2_1 = 1'h0;
  end
  if (reset) begin
    validVec_2_2 = 1'h0;
  end
  if (reset) begin
    validVec_2_3 = 1'h0;
  end
  if (reset) begin
    validVec_3_0 = 1'h0;
  end
  if (reset) begin
    validVec_3_1 = 1'h0;
  end
  if (reset) begin
    validVec_3_2 = 1'h0;
  end
  if (reset) begin
    validVec_3_3 = 1'h0;
  end
  if (reset) begin
    validVec_4_0 = 1'h0;
  end
  if (reset) begin
    validVec_4_1 = 1'h0;
  end
  if (reset) begin
    validVec_4_2 = 1'h0;
  end
  if (reset) begin
    validVec_4_3 = 1'h0;
  end
  if (reset) begin
    validVec_5_0 = 1'h0;
  end
  if (reset) begin
    validVec_5_1 = 1'h0;
  end
  if (reset) begin
    validVec_5_2 = 1'h0;
  end
  if (reset) begin
    validVec_5_3 = 1'h0;
  end
  if (reset) begin
    validVec_6_0 = 1'h0;
  end
  if (reset) begin
    validVec_6_1 = 1'h0;
  end
  if (reset) begin
    validVec_6_2 = 1'h0;
  end
  if (reset) begin
    validVec_6_3 = 1'h0;
  end
  if (reset) begin
    validVec_7_0 = 1'h0;
  end
  if (reset) begin
    validVec_7_1 = 1'h0;
  end
  if (reset) begin
    validVec_7_2 = 1'h0;
  end
  if (reset) begin
    validVec_7_3 = 1'h0;
  end
  if (reset) begin
    validVec_8_0 = 1'h0;
  end
  if (reset) begin
    validVec_8_1 = 1'h0;
  end
  if (reset) begin
    validVec_8_2 = 1'h0;
  end
  if (reset) begin
    validVec_8_3 = 1'h0;
  end
  if (reset) begin
    validVec_9_0 = 1'h0;
  end
  if (reset) begin
    validVec_9_1 = 1'h0;
  end
  if (reset) begin
    validVec_9_2 = 1'h0;
  end
  if (reset) begin
    validVec_9_3 = 1'h0;
  end
  if (reset) begin
    validVec_10_0 = 1'h0;
  end
  if (reset) begin
    validVec_10_1 = 1'h0;
  end
  if (reset) begin
    validVec_10_2 = 1'h0;
  end
  if (reset) begin
    validVec_10_3 = 1'h0;
  end
  if (reset) begin
    validVec_11_0 = 1'h0;
  end
  if (reset) begin
    validVec_11_1 = 1'h0;
  end
  if (reset) begin
    validVec_11_2 = 1'h0;
  end
  if (reset) begin
    validVec_11_3 = 1'h0;
  end
  if (reset) begin
    validVec_12_0 = 1'h0;
  end
  if (reset) begin
    validVec_12_1 = 1'h0;
  end
  if (reset) begin
    validVec_12_2 = 1'h0;
  end
  if (reset) begin
    validVec_12_3 = 1'h0;
  end
  if (reset) begin
    validVec_13_0 = 1'h0;
  end
  if (reset) begin
    validVec_13_1 = 1'h0;
  end
  if (reset) begin
    validVec_13_2 = 1'h0;
  end
  if (reset) begin
    validVec_13_3 = 1'h0;
  end
  if (reset) begin
    validVec_14_0 = 1'h0;
  end
  if (reset) begin
    validVec_14_1 = 1'h0;
  end
  if (reset) begin
    validVec_14_2 = 1'h0;
  end
  if (reset) begin
    validVec_14_3 = 1'h0;
  end
  if (reset) begin
    validVec_15_0 = 1'h0;
  end
  if (reset) begin
    validVec_15_1 = 1'h0;
  end
  if (reset) begin
    validVec_15_2 = 1'h0;
  end
  if (reset) begin
    validVec_15_3 = 1'h0;
  end
  if (reset) begin
    validVec_16_0 = 1'h0;
  end
  if (reset) begin
    validVec_16_1 = 1'h0;
  end
  if (reset) begin
    validVec_16_2 = 1'h0;
  end
  if (reset) begin
    validVec_16_3 = 1'h0;
  end
  if (reset) begin
    validVec_17_0 = 1'h0;
  end
  if (reset) begin
    validVec_17_1 = 1'h0;
  end
  if (reset) begin
    validVec_17_2 = 1'h0;
  end
  if (reset) begin
    validVec_17_3 = 1'h0;
  end
  if (reset) begin
    validVec_18_0 = 1'h0;
  end
  if (reset) begin
    validVec_18_1 = 1'h0;
  end
  if (reset) begin
    validVec_18_2 = 1'h0;
  end
  if (reset) begin
    validVec_18_3 = 1'h0;
  end
  if (reset) begin
    validVec_19_0 = 1'h0;
  end
  if (reset) begin
    validVec_19_1 = 1'h0;
  end
  if (reset) begin
    validVec_19_2 = 1'h0;
  end
  if (reset) begin
    validVec_19_3 = 1'h0;
  end
  if (reset) begin
    validVec_20_0 = 1'h0;
  end
  if (reset) begin
    validVec_20_1 = 1'h0;
  end
  if (reset) begin
    validVec_20_2 = 1'h0;
  end
  if (reset) begin
    validVec_20_3 = 1'h0;
  end
  if (reset) begin
    validVec_21_0 = 1'h0;
  end
  if (reset) begin
    validVec_21_1 = 1'h0;
  end
  if (reset) begin
    validVec_21_2 = 1'h0;
  end
  if (reset) begin
    validVec_21_3 = 1'h0;
  end
  if (reset) begin
    validVec_22_0 = 1'h0;
  end
  if (reset) begin
    validVec_22_1 = 1'h0;
  end
  if (reset) begin
    validVec_22_2 = 1'h0;
  end
  if (reset) begin
    validVec_22_3 = 1'h0;
  end
  if (reset) begin
    validVec_23_0 = 1'h0;
  end
  if (reset) begin
    validVec_23_1 = 1'h0;
  end
  if (reset) begin
    validVec_23_2 = 1'h0;
  end
  if (reset) begin
    validVec_23_3 = 1'h0;
  end
  if (reset) begin
    validVec_24_0 = 1'h0;
  end
  if (reset) begin
    validVec_24_1 = 1'h0;
  end
  if (reset) begin
    validVec_24_2 = 1'h0;
  end
  if (reset) begin
    validVec_24_3 = 1'h0;
  end
  if (reset) begin
    validVec_25_0 = 1'h0;
  end
  if (reset) begin
    validVec_25_1 = 1'h0;
  end
  if (reset) begin
    validVec_25_2 = 1'h0;
  end
  if (reset) begin
    validVec_25_3 = 1'h0;
  end
  if (reset) begin
    validVec_26_0 = 1'h0;
  end
  if (reset) begin
    validVec_26_1 = 1'h0;
  end
  if (reset) begin
    validVec_26_2 = 1'h0;
  end
  if (reset) begin
    validVec_26_3 = 1'h0;
  end
  if (reset) begin
    validVec_27_0 = 1'h0;
  end
  if (reset) begin
    validVec_27_1 = 1'h0;
  end
  if (reset) begin
    validVec_27_2 = 1'h0;
  end
  if (reset) begin
    validVec_27_3 = 1'h0;
  end
  if (reset) begin
    validVec_28_0 = 1'h0;
  end
  if (reset) begin
    validVec_28_1 = 1'h0;
  end
  if (reset) begin
    validVec_28_2 = 1'h0;
  end
  if (reset) begin
    validVec_28_3 = 1'h0;
  end
  if (reset) begin
    validVec_29_0 = 1'h0;
  end
  if (reset) begin
    validVec_29_1 = 1'h0;
  end
  if (reset) begin
    validVec_29_2 = 1'h0;
  end
  if (reset) begin
    validVec_29_3 = 1'h0;
  end
  if (reset) begin
    validVec_30_0 = 1'h0;
  end
  if (reset) begin
    validVec_30_1 = 1'h0;
  end
  if (reset) begin
    validVec_30_2 = 1'h0;
  end
  if (reset) begin
    validVec_30_3 = 1'h0;
  end
  if (reset) begin
    validVec_31_0 = 1'h0;
  end
  if (reset) begin
    validVec_31_1 = 1'h0;
  end
  if (reset) begin
    validVec_31_2 = 1'h0;
  end
  if (reset) begin
    validVec_31_3 = 1'h0;
  end
  if (reset) begin
    allocPtr_0 = 2'h0;
  end
  if (reset) begin
    allocPtr_1 = 2'h0;
  end
  if (reset) begin
    allocPtr_2 = 2'h0;
  end
  if (reset) begin
    allocPtr_3 = 2'h0;
  end
  if (reset) begin
    allocPtr_4 = 2'h0;
  end
  if (reset) begin
    allocPtr_5 = 2'h0;
  end
  if (reset) begin
    allocPtr_6 = 2'h0;
  end
  if (reset) begin
    allocPtr_7 = 2'h0;
  end
  if (reset) begin
    allocPtr_8 = 2'h0;
  end
  if (reset) begin
    allocPtr_9 = 2'h0;
  end
  if (reset) begin
    allocPtr_10 = 2'h0;
  end
  if (reset) begin
    allocPtr_11 = 2'h0;
  end
  if (reset) begin
    allocPtr_12 = 2'h0;
  end
  if (reset) begin
    allocPtr_13 = 2'h0;
  end
  if (reset) begin
    allocPtr_14 = 2'h0;
  end
  if (reset) begin
    allocPtr_15 = 2'h0;
  end
  if (reset) begin
    allocPtr_16 = 2'h0;
  end
  if (reset) begin
    allocPtr_17 = 2'h0;
  end
  if (reset) begin
    allocPtr_18 = 2'h0;
  end
  if (reset) begin
    allocPtr_19 = 2'h0;
  end
  if (reset) begin
    allocPtr_20 = 2'h0;
  end
  if (reset) begin
    allocPtr_21 = 2'h0;
  end
  if (reset) begin
    allocPtr_22 = 2'h0;
  end
  if (reset) begin
    allocPtr_23 = 2'h0;
  end
  if (reset) begin
    allocPtr_24 = 2'h0;
  end
  if (reset) begin
    allocPtr_25 = 2'h0;
  end
  if (reset) begin
    allocPtr_26 = 2'h0;
  end
  if (reset) begin
    allocPtr_27 = 2'h0;
  end
  if (reset) begin
    allocPtr_28 = 2'h0;
  end
  if (reset) begin
    allocPtr_29 = 2'h0;
  end
  if (reset) begin
    allocPtr_30 = 2'h0;
  end
  if (reset) begin
    allocPtr_31 = 2'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule

