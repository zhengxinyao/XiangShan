module PMPCheckerv2(
  input         clock,
  input         reset,
  input  [1:0]  io_check_env_mode,
  input         io_check_env_pmp_0_cfg_l,
  input  [1:0]  io_check_env_pmp_0_cfg_a,
  input         io_check_env_pmp_0_cfg_x,
  input         io_check_env_pmp_0_cfg_w,
  input         io_check_env_pmp_0_cfg_r,
  input  [33:0] io_check_env_pmp_0_addr,
  input  [35:0] io_check_env_pmp_0_mask,
  input         io_check_env_pmp_1_cfg_l,
  input  [1:0]  io_check_env_pmp_1_cfg_a,
  input         io_check_env_pmp_1_cfg_x,
  input         io_check_env_pmp_1_cfg_w,
  input         io_check_env_pmp_1_cfg_r,
  input  [33:0] io_check_env_pmp_1_addr,
  input  [35:0] io_check_env_pmp_1_mask,
  input         io_check_env_pmp_2_cfg_l,
  input  [1:0]  io_check_env_pmp_2_cfg_a,
  input         io_check_env_pmp_2_cfg_x,
  input         io_check_env_pmp_2_cfg_w,
  input         io_check_env_pmp_2_cfg_r,
  input  [33:0] io_check_env_pmp_2_addr,
  input  [35:0] io_check_env_pmp_2_mask,
  input         io_check_env_pmp_3_cfg_l,
  input  [1:0]  io_check_env_pmp_3_cfg_a,
  input         io_check_env_pmp_3_cfg_x,
  input         io_check_env_pmp_3_cfg_w,
  input         io_check_env_pmp_3_cfg_r,
  input  [33:0] io_check_env_pmp_3_addr,
  input  [35:0] io_check_env_pmp_3_mask,
  input         io_check_env_pmp_4_cfg_l,
  input  [1:0]  io_check_env_pmp_4_cfg_a,
  input         io_check_env_pmp_4_cfg_x,
  input         io_check_env_pmp_4_cfg_w,
  input         io_check_env_pmp_4_cfg_r,
  input  [33:0] io_check_env_pmp_4_addr,
  input  [35:0] io_check_env_pmp_4_mask,
  input         io_check_env_pmp_5_cfg_l,
  input  [1:0]  io_check_env_pmp_5_cfg_a,
  input         io_check_env_pmp_5_cfg_x,
  input         io_check_env_pmp_5_cfg_w,
  input         io_check_env_pmp_5_cfg_r,
  input  [33:0] io_check_env_pmp_5_addr,
  input  [35:0] io_check_env_pmp_5_mask,
  input         io_check_env_pmp_6_cfg_l,
  input  [1:0]  io_check_env_pmp_6_cfg_a,
  input         io_check_env_pmp_6_cfg_x,
  input         io_check_env_pmp_6_cfg_w,
  input         io_check_env_pmp_6_cfg_r,
  input  [33:0] io_check_env_pmp_6_addr,
  input  [35:0] io_check_env_pmp_6_mask,
  input         io_check_env_pmp_7_cfg_l,
  input  [1:0]  io_check_env_pmp_7_cfg_a,
  input         io_check_env_pmp_7_cfg_x,
  input         io_check_env_pmp_7_cfg_w,
  input         io_check_env_pmp_7_cfg_r,
  input  [33:0] io_check_env_pmp_7_addr,
  input  [35:0] io_check_env_pmp_7_mask,
  input         io_check_env_pmp_8_cfg_l,
  input  [1:0]  io_check_env_pmp_8_cfg_a,
  input         io_check_env_pmp_8_cfg_x,
  input         io_check_env_pmp_8_cfg_w,
  input         io_check_env_pmp_8_cfg_r,
  input  [33:0] io_check_env_pmp_8_addr,
  input  [35:0] io_check_env_pmp_8_mask,
  input         io_check_env_pmp_9_cfg_l,
  input  [1:0]  io_check_env_pmp_9_cfg_a,
  input         io_check_env_pmp_9_cfg_x,
  input         io_check_env_pmp_9_cfg_w,
  input         io_check_env_pmp_9_cfg_r,
  input  [33:0] io_check_env_pmp_9_addr,
  input  [35:0] io_check_env_pmp_9_mask,
  input         io_check_env_pmp_10_cfg_l,
  input  [1:0]  io_check_env_pmp_10_cfg_a,
  input         io_check_env_pmp_10_cfg_x,
  input         io_check_env_pmp_10_cfg_w,
  input         io_check_env_pmp_10_cfg_r,
  input  [33:0] io_check_env_pmp_10_addr,
  input  [35:0] io_check_env_pmp_10_mask,
  input         io_check_env_pmp_11_cfg_l,
  input  [1:0]  io_check_env_pmp_11_cfg_a,
  input         io_check_env_pmp_11_cfg_x,
  input         io_check_env_pmp_11_cfg_w,
  input         io_check_env_pmp_11_cfg_r,
  input  [33:0] io_check_env_pmp_11_addr,
  input  [35:0] io_check_env_pmp_11_mask,
  input         io_check_env_pmp_12_cfg_l,
  input  [1:0]  io_check_env_pmp_12_cfg_a,
  input         io_check_env_pmp_12_cfg_x,
  input         io_check_env_pmp_12_cfg_w,
  input         io_check_env_pmp_12_cfg_r,
  input  [33:0] io_check_env_pmp_12_addr,
  input  [35:0] io_check_env_pmp_12_mask,
  input         io_check_env_pmp_13_cfg_l,
  input  [1:0]  io_check_env_pmp_13_cfg_a,
  input         io_check_env_pmp_13_cfg_x,
  input         io_check_env_pmp_13_cfg_w,
  input         io_check_env_pmp_13_cfg_r,
  input  [33:0] io_check_env_pmp_13_addr,
  input  [35:0] io_check_env_pmp_13_mask,
  input         io_check_env_pmp_14_cfg_l,
  input  [1:0]  io_check_env_pmp_14_cfg_a,
  input         io_check_env_pmp_14_cfg_x,
  input         io_check_env_pmp_14_cfg_w,
  input         io_check_env_pmp_14_cfg_r,
  input  [33:0] io_check_env_pmp_14_addr,
  input  [35:0] io_check_env_pmp_14_mask,
  input         io_check_env_pmp_15_cfg_l,
  input  [1:0]  io_check_env_pmp_15_cfg_a,
  input         io_check_env_pmp_15_cfg_x,
  input         io_check_env_pmp_15_cfg_w,
  input         io_check_env_pmp_15_cfg_r,
  input  [33:0] io_check_env_pmp_15_addr,
  input  [35:0] io_check_env_pmp_15_mask,
  input         io_check_env_pma_0_cfg_c,
  input         io_check_env_pma_0_cfg_atomic,
  input  [1:0]  io_check_env_pma_0_cfg_a,
  input         io_check_env_pma_0_cfg_x,
  input         io_check_env_pma_0_cfg_w,
  input         io_check_env_pma_0_cfg_r,
  input  [33:0] io_check_env_pma_0_addr,
  input  [35:0] io_check_env_pma_0_mask,
  input         io_check_env_pma_1_cfg_c,
  input         io_check_env_pma_1_cfg_atomic,
  input  [1:0]  io_check_env_pma_1_cfg_a,
  input         io_check_env_pma_1_cfg_x,
  input         io_check_env_pma_1_cfg_w,
  input         io_check_env_pma_1_cfg_r,
  input  [33:0] io_check_env_pma_1_addr,
  input  [35:0] io_check_env_pma_1_mask,
  input         io_check_env_pma_2_cfg_c,
  input         io_check_env_pma_2_cfg_atomic,
  input  [1:0]  io_check_env_pma_2_cfg_a,
  input         io_check_env_pma_2_cfg_x,
  input         io_check_env_pma_2_cfg_w,
  input         io_check_env_pma_2_cfg_r,
  input  [33:0] io_check_env_pma_2_addr,
  input  [35:0] io_check_env_pma_2_mask,
  input         io_check_env_pma_3_cfg_c,
  input         io_check_env_pma_3_cfg_atomic,
  input  [1:0]  io_check_env_pma_3_cfg_a,
  input         io_check_env_pma_3_cfg_x,
  input         io_check_env_pma_3_cfg_w,
  input         io_check_env_pma_3_cfg_r,
  input  [33:0] io_check_env_pma_3_addr,
  input  [35:0] io_check_env_pma_3_mask,
  input         io_check_env_pma_4_cfg_c,
  input         io_check_env_pma_4_cfg_atomic,
  input  [1:0]  io_check_env_pma_4_cfg_a,
  input         io_check_env_pma_4_cfg_x,
  input         io_check_env_pma_4_cfg_w,
  input         io_check_env_pma_4_cfg_r,
  input  [33:0] io_check_env_pma_4_addr,
  input  [35:0] io_check_env_pma_4_mask,
  input         io_check_env_pma_5_cfg_c,
  input         io_check_env_pma_5_cfg_atomic,
  input  [1:0]  io_check_env_pma_5_cfg_a,
  input         io_check_env_pma_5_cfg_x,
  input         io_check_env_pma_5_cfg_w,
  input         io_check_env_pma_5_cfg_r,
  input  [33:0] io_check_env_pma_5_addr,
  input  [35:0] io_check_env_pma_5_mask,
  input         io_check_env_pma_6_cfg_c,
  input         io_check_env_pma_6_cfg_atomic,
  input  [1:0]  io_check_env_pma_6_cfg_a,
  input         io_check_env_pma_6_cfg_x,
  input         io_check_env_pma_6_cfg_w,
  input         io_check_env_pma_6_cfg_r,
  input  [33:0] io_check_env_pma_6_addr,
  input  [35:0] io_check_env_pma_6_mask,
  input         io_check_env_pma_7_cfg_c,
  input         io_check_env_pma_7_cfg_atomic,
  input  [1:0]  io_check_env_pma_7_cfg_a,
  input         io_check_env_pma_7_cfg_x,
  input         io_check_env_pma_7_cfg_w,
  input         io_check_env_pma_7_cfg_r,
  input  [33:0] io_check_env_pma_7_addr,
  input  [35:0] io_check_env_pma_7_mask,
  input         io_check_env_pma_8_cfg_c,
  input         io_check_env_pma_8_cfg_atomic,
  input  [1:0]  io_check_env_pma_8_cfg_a,
  input         io_check_env_pma_8_cfg_x,
  input         io_check_env_pma_8_cfg_w,
  input         io_check_env_pma_8_cfg_r,
  input  [33:0] io_check_env_pma_8_addr,
  input  [35:0] io_check_env_pma_8_mask,
  input         io_check_env_pma_9_cfg_c,
  input         io_check_env_pma_9_cfg_atomic,
  input  [1:0]  io_check_env_pma_9_cfg_a,
  input         io_check_env_pma_9_cfg_x,
  input         io_check_env_pma_9_cfg_w,
  input         io_check_env_pma_9_cfg_r,
  input  [33:0] io_check_env_pma_9_addr,
  input  [35:0] io_check_env_pma_9_mask,
  input         io_check_env_pma_10_cfg_c,
  input         io_check_env_pma_10_cfg_atomic,
  input  [1:0]  io_check_env_pma_10_cfg_a,
  input         io_check_env_pma_10_cfg_x,
  input         io_check_env_pma_10_cfg_w,
  input         io_check_env_pma_10_cfg_r,
  input  [33:0] io_check_env_pma_10_addr,
  input  [35:0] io_check_env_pma_10_mask,
  input         io_check_env_pma_11_cfg_c,
  input         io_check_env_pma_11_cfg_atomic,
  input  [1:0]  io_check_env_pma_11_cfg_a,
  input         io_check_env_pma_11_cfg_x,
  input         io_check_env_pma_11_cfg_w,
  input         io_check_env_pma_11_cfg_r,
  input  [33:0] io_check_env_pma_11_addr,
  input  [35:0] io_check_env_pma_11_mask,
  input         io_check_env_pma_12_cfg_c,
  input         io_check_env_pma_12_cfg_atomic,
  input  [1:0]  io_check_env_pma_12_cfg_a,
  input         io_check_env_pma_12_cfg_x,
  input         io_check_env_pma_12_cfg_w,
  input         io_check_env_pma_12_cfg_r,
  input  [33:0] io_check_env_pma_12_addr,
  input  [35:0] io_check_env_pma_12_mask,
  input         io_check_env_pma_13_cfg_c,
  input         io_check_env_pma_13_cfg_atomic,
  input  [1:0]  io_check_env_pma_13_cfg_a,
  input         io_check_env_pma_13_cfg_x,
  input         io_check_env_pma_13_cfg_w,
  input         io_check_env_pma_13_cfg_r,
  input  [33:0] io_check_env_pma_13_addr,
  input  [35:0] io_check_env_pma_13_mask,
  input         io_check_env_pma_14_cfg_c,
  input         io_check_env_pma_14_cfg_atomic,
  input  [1:0]  io_check_env_pma_14_cfg_a,
  input         io_check_env_pma_14_cfg_x,
  input         io_check_env_pma_14_cfg_w,
  input         io_check_env_pma_14_cfg_r,
  input  [33:0] io_check_env_pma_14_addr,
  input  [35:0] io_check_env_pma_14_mask,
  input         io_check_env_pma_15_cfg_c,
  input         io_check_env_pma_15_cfg_atomic,
  input  [1:0]  io_check_env_pma_15_cfg_a,
  input         io_check_env_pma_15_cfg_x,
  input         io_check_env_pma_15_cfg_w,
  input         io_check_env_pma_15_cfg_r,
  input  [33:0] io_check_env_pma_15_addr,
  input  [35:0] io_check_env_pma_15_mask,
  input         io_req_valid,
  input  [35:0] io_req_bits_addr,
  output        io_resp_c,
  output        io_resp_atomic,
  output        io_resp_x,
  output        io_resp_w,
  output        io_resp_r
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
`endif // RANDOMIZE_REG_INIT
  wire  res_pmp_passThrough = io_check_env_mode > 2'h1; // @[PMP.scala 423:65]
  wire [35:0] _res_pmp_is_match_T_1 = {io_check_env_pmp_0_addr, 2'h0}; // @[PMP.scala 190:35]
  wire [35:0] _res_pmp_is_match_T_3 = _res_pmp_is_match_T_1 & 36'hffffff000; // @[PMP.scala 190:50]
  wire [35:0] _res_pmp_is_match_T_4 = ~io_check_env_pmp_0_mask; // @[PMP.scala 232:10]
  wire [35:0] _res_pmp_is_match_T_5 = io_req_bits_addr & _res_pmp_is_match_T_4; // @[PMP.scala 232:8]
  wire [35:0] _res_pmp_is_match_T_7 = _res_pmp_is_match_T_3 & _res_pmp_is_match_T_4; // @[PMP.scala 232:21]
  wire  _res_pmp_is_match_T_8 = _res_pmp_is_match_T_5 == _res_pmp_is_match_T_7; // @[PMP.scala 232:14]
  wire  _res_pmp_is_match_T_9 = io_check_env_pmp_0_cfg_a == 2'h1; // @[PMP.scala 53:15]
  wire  _res_pmp_is_match_T_18 = io_req_bits_addr < _res_pmp_is_match_T_3; // @[PMP.scala 210:14]
  wire  _res_pmp_is_match_T_20 = _res_pmp_is_match_T_9 & _res_pmp_is_match_T_18; // @[PMP.scala 200:10]
  wire  res_pmp_ignore = res_pmp_passThrough & ~io_check_env_pmp_0_cfg_l; // @[PMP.scala 434:32]
  wire  res_pmp_cur_cfg_r = io_check_env_pmp_0_cfg_r | res_pmp_ignore; // @[PMP.scala 438:42]
  wire  res_pmp_cur_cfg_w = io_check_env_pmp_0_cfg_w | res_pmp_ignore; // @[PMP.scala 439:42]
  wire  res_pmp_cur_cfg_x = io_check_env_pmp_0_cfg_x | res_pmp_ignore; // @[PMP.scala 440:42]
  wire [35:0] _res_pmp_is_match_T_22 = {io_check_env_pmp_1_addr, 2'h0}; // @[PMP.scala 190:35]
  wire [35:0] _res_pmp_is_match_T_24 = _res_pmp_is_match_T_22 & 36'hffffff000; // @[PMP.scala 190:50]
  wire [35:0] _res_pmp_is_match_T_25 = ~io_check_env_pmp_1_mask; // @[PMP.scala 232:10]
  wire [35:0] _res_pmp_is_match_T_26 = io_req_bits_addr & _res_pmp_is_match_T_25; // @[PMP.scala 232:8]
  wire [35:0] _res_pmp_is_match_T_28 = _res_pmp_is_match_T_24 & _res_pmp_is_match_T_25; // @[PMP.scala 232:21]
  wire  _res_pmp_is_match_T_29 = _res_pmp_is_match_T_26 == _res_pmp_is_match_T_28; // @[PMP.scala 232:14]
  wire  _res_pmp_is_match_T_30 = io_check_env_pmp_1_cfg_a == 2'h1; // @[PMP.scala 53:15]
  wire  _res_pmp_is_match_T_35 = ~_res_pmp_is_match_T_18; // @[PMP.scala 220:5]
  wire  _res_pmp_is_match_T_39 = io_req_bits_addr < _res_pmp_is_match_T_24; // @[PMP.scala 210:14]
  wire  _res_pmp_is_match_T_40 = _res_pmp_is_match_T_35 & _res_pmp_is_match_T_39; // @[PMP.scala 228:56]
  wire  _res_pmp_is_match_T_41 = _res_pmp_is_match_T_30 & _res_pmp_is_match_T_40; // @[PMP.scala 200:10]
  wire  res_pmp_ignore_1 = res_pmp_passThrough & ~io_check_env_pmp_1_cfg_l; // @[PMP.scala 434:32]
  wire  res_pmp_cur_1_cfg_r = io_check_env_pmp_1_cfg_r | res_pmp_ignore_1; // @[PMP.scala 438:42]
  wire  res_pmp_cur_1_cfg_w = io_check_env_pmp_1_cfg_w | res_pmp_ignore_1; // @[PMP.scala 439:42]
  wire  res_pmp_cur_1_cfg_x = io_check_env_pmp_1_cfg_x | res_pmp_ignore_1; // @[PMP.scala 440:42]
  wire [35:0] _res_pmp_is_match_T_43 = {io_check_env_pmp_2_addr, 2'h0}; // @[PMP.scala 190:35]
  wire [35:0] _res_pmp_is_match_T_45 = _res_pmp_is_match_T_43 & 36'hffffff000; // @[PMP.scala 190:50]
  wire [35:0] _res_pmp_is_match_T_46 = ~io_check_env_pmp_2_mask; // @[PMP.scala 232:10]
  wire [35:0] _res_pmp_is_match_T_47 = io_req_bits_addr & _res_pmp_is_match_T_46; // @[PMP.scala 232:8]
  wire [35:0] _res_pmp_is_match_T_49 = _res_pmp_is_match_T_45 & _res_pmp_is_match_T_46; // @[PMP.scala 232:21]
  wire  _res_pmp_is_match_T_50 = _res_pmp_is_match_T_47 == _res_pmp_is_match_T_49; // @[PMP.scala 232:14]
  wire  _res_pmp_is_match_T_51 = io_check_env_pmp_2_cfg_a == 2'h1; // @[PMP.scala 53:15]
  wire  _res_pmp_is_match_T_56 = ~_res_pmp_is_match_T_39; // @[PMP.scala 220:5]
  wire  _res_pmp_is_match_T_60 = io_req_bits_addr < _res_pmp_is_match_T_45; // @[PMP.scala 210:14]
  wire  _res_pmp_is_match_T_61 = _res_pmp_is_match_T_56 & _res_pmp_is_match_T_60; // @[PMP.scala 228:56]
  wire  _res_pmp_is_match_T_62 = _res_pmp_is_match_T_51 & _res_pmp_is_match_T_61; // @[PMP.scala 200:10]
  wire  res_pmp_ignore_2 = res_pmp_passThrough & ~io_check_env_pmp_2_cfg_l; // @[PMP.scala 434:32]
  wire  res_pmp_cur_2_cfg_r = io_check_env_pmp_2_cfg_r | res_pmp_ignore_2; // @[PMP.scala 438:42]
  wire  res_pmp_cur_2_cfg_w = io_check_env_pmp_2_cfg_w | res_pmp_ignore_2; // @[PMP.scala 439:42]
  wire  res_pmp_cur_2_cfg_x = io_check_env_pmp_2_cfg_x | res_pmp_ignore_2; // @[PMP.scala 440:42]
  wire [35:0] _res_pmp_is_match_T_64 = {io_check_env_pmp_3_addr, 2'h0}; // @[PMP.scala 190:35]
  wire [35:0] _res_pmp_is_match_T_66 = _res_pmp_is_match_T_64 & 36'hffffff000; // @[PMP.scala 190:50]
  wire [35:0] _res_pmp_is_match_T_67 = ~io_check_env_pmp_3_mask; // @[PMP.scala 232:10]
  wire [35:0] _res_pmp_is_match_T_68 = io_req_bits_addr & _res_pmp_is_match_T_67; // @[PMP.scala 232:8]
  wire [35:0] _res_pmp_is_match_T_70 = _res_pmp_is_match_T_66 & _res_pmp_is_match_T_67; // @[PMP.scala 232:21]
  wire  _res_pmp_is_match_T_71 = _res_pmp_is_match_T_68 == _res_pmp_is_match_T_70; // @[PMP.scala 232:14]
  wire  _res_pmp_is_match_T_72 = io_check_env_pmp_3_cfg_a == 2'h1; // @[PMP.scala 53:15]
  wire  _res_pmp_is_match_T_77 = ~_res_pmp_is_match_T_60; // @[PMP.scala 220:5]
  wire  _res_pmp_is_match_T_81 = io_req_bits_addr < _res_pmp_is_match_T_66; // @[PMP.scala 210:14]
  wire  _res_pmp_is_match_T_82 = _res_pmp_is_match_T_77 & _res_pmp_is_match_T_81; // @[PMP.scala 228:56]
  wire  _res_pmp_is_match_T_83 = _res_pmp_is_match_T_72 & _res_pmp_is_match_T_82; // @[PMP.scala 200:10]
  wire  res_pmp_ignore_3 = res_pmp_passThrough & ~io_check_env_pmp_3_cfg_l; // @[PMP.scala 434:32]
  wire  res_pmp_cur_3_cfg_r = io_check_env_pmp_3_cfg_r | res_pmp_ignore_3; // @[PMP.scala 438:42]
  wire  res_pmp_cur_3_cfg_w = io_check_env_pmp_3_cfg_w | res_pmp_ignore_3; // @[PMP.scala 439:42]
  wire  res_pmp_cur_3_cfg_x = io_check_env_pmp_3_cfg_x | res_pmp_ignore_3; // @[PMP.scala 440:42]
  wire [35:0] _res_pmp_is_match_T_85 = {io_check_env_pmp_4_addr, 2'h0}; // @[PMP.scala 190:35]
  wire [35:0] _res_pmp_is_match_T_87 = _res_pmp_is_match_T_85 & 36'hffffff000; // @[PMP.scala 190:50]
  wire [35:0] _res_pmp_is_match_T_88 = ~io_check_env_pmp_4_mask; // @[PMP.scala 232:10]
  wire [35:0] _res_pmp_is_match_T_89 = io_req_bits_addr & _res_pmp_is_match_T_88; // @[PMP.scala 232:8]
  wire [35:0] _res_pmp_is_match_T_91 = _res_pmp_is_match_T_87 & _res_pmp_is_match_T_88; // @[PMP.scala 232:21]
  wire  _res_pmp_is_match_T_92 = _res_pmp_is_match_T_89 == _res_pmp_is_match_T_91; // @[PMP.scala 232:14]
  wire  _res_pmp_is_match_T_93 = io_check_env_pmp_4_cfg_a == 2'h1; // @[PMP.scala 53:15]
  wire  _res_pmp_is_match_T_98 = ~_res_pmp_is_match_T_81; // @[PMP.scala 220:5]
  wire  _res_pmp_is_match_T_102 = io_req_bits_addr < _res_pmp_is_match_T_87; // @[PMP.scala 210:14]
  wire  _res_pmp_is_match_T_103 = _res_pmp_is_match_T_98 & _res_pmp_is_match_T_102; // @[PMP.scala 228:56]
  wire  _res_pmp_is_match_T_104 = _res_pmp_is_match_T_93 & _res_pmp_is_match_T_103; // @[PMP.scala 200:10]
  wire  res_pmp_ignore_4 = res_pmp_passThrough & ~io_check_env_pmp_4_cfg_l; // @[PMP.scala 434:32]
  wire  res_pmp_cur_4_cfg_r = io_check_env_pmp_4_cfg_r | res_pmp_ignore_4; // @[PMP.scala 438:42]
  wire  res_pmp_cur_4_cfg_w = io_check_env_pmp_4_cfg_w | res_pmp_ignore_4; // @[PMP.scala 439:42]
  wire  res_pmp_cur_4_cfg_x = io_check_env_pmp_4_cfg_x | res_pmp_ignore_4; // @[PMP.scala 440:42]
  wire [35:0] _res_pmp_is_match_T_106 = {io_check_env_pmp_5_addr, 2'h0}; // @[PMP.scala 190:35]
  wire [35:0] _res_pmp_is_match_T_108 = _res_pmp_is_match_T_106 & 36'hffffff000; // @[PMP.scala 190:50]
  wire [35:0] _res_pmp_is_match_T_109 = ~io_check_env_pmp_5_mask; // @[PMP.scala 232:10]
  wire [35:0] _res_pmp_is_match_T_110 = io_req_bits_addr & _res_pmp_is_match_T_109; // @[PMP.scala 232:8]
  wire [35:0] _res_pmp_is_match_T_112 = _res_pmp_is_match_T_108 & _res_pmp_is_match_T_109; // @[PMP.scala 232:21]
  wire  _res_pmp_is_match_T_113 = _res_pmp_is_match_T_110 == _res_pmp_is_match_T_112; // @[PMP.scala 232:14]
  wire  _res_pmp_is_match_T_114 = io_check_env_pmp_5_cfg_a == 2'h1; // @[PMP.scala 53:15]
  wire  _res_pmp_is_match_T_119 = ~_res_pmp_is_match_T_102; // @[PMP.scala 220:5]
  wire  _res_pmp_is_match_T_123 = io_req_bits_addr < _res_pmp_is_match_T_108; // @[PMP.scala 210:14]
  wire  _res_pmp_is_match_T_124 = _res_pmp_is_match_T_119 & _res_pmp_is_match_T_123; // @[PMP.scala 228:56]
  wire  _res_pmp_is_match_T_125 = _res_pmp_is_match_T_114 & _res_pmp_is_match_T_124; // @[PMP.scala 200:10]
  wire  res_pmp_ignore_5 = res_pmp_passThrough & ~io_check_env_pmp_5_cfg_l; // @[PMP.scala 434:32]
  wire  res_pmp_cur_5_cfg_r = io_check_env_pmp_5_cfg_r | res_pmp_ignore_5; // @[PMP.scala 438:42]
  wire  res_pmp_cur_5_cfg_w = io_check_env_pmp_5_cfg_w | res_pmp_ignore_5; // @[PMP.scala 439:42]
  wire  res_pmp_cur_5_cfg_x = io_check_env_pmp_5_cfg_x | res_pmp_ignore_5; // @[PMP.scala 440:42]
  wire [35:0] _res_pmp_is_match_T_127 = {io_check_env_pmp_6_addr, 2'h0}; // @[PMP.scala 190:35]
  wire [35:0] _res_pmp_is_match_T_129 = _res_pmp_is_match_T_127 & 36'hffffff000; // @[PMP.scala 190:50]
  wire [35:0] _res_pmp_is_match_T_130 = ~io_check_env_pmp_6_mask; // @[PMP.scala 232:10]
  wire [35:0] _res_pmp_is_match_T_131 = io_req_bits_addr & _res_pmp_is_match_T_130; // @[PMP.scala 232:8]
  wire [35:0] _res_pmp_is_match_T_133 = _res_pmp_is_match_T_129 & _res_pmp_is_match_T_130; // @[PMP.scala 232:21]
  wire  _res_pmp_is_match_T_134 = _res_pmp_is_match_T_131 == _res_pmp_is_match_T_133; // @[PMP.scala 232:14]
  wire  _res_pmp_is_match_T_135 = io_check_env_pmp_6_cfg_a == 2'h1; // @[PMP.scala 53:15]
  wire  _res_pmp_is_match_T_140 = ~_res_pmp_is_match_T_123; // @[PMP.scala 220:5]
  wire  _res_pmp_is_match_T_144 = io_req_bits_addr < _res_pmp_is_match_T_129; // @[PMP.scala 210:14]
  wire  _res_pmp_is_match_T_145 = _res_pmp_is_match_T_140 & _res_pmp_is_match_T_144; // @[PMP.scala 228:56]
  wire  _res_pmp_is_match_T_146 = _res_pmp_is_match_T_135 & _res_pmp_is_match_T_145; // @[PMP.scala 200:10]
  wire  res_pmp_ignore_6 = res_pmp_passThrough & ~io_check_env_pmp_6_cfg_l; // @[PMP.scala 434:32]
  wire  res_pmp_cur_6_cfg_r = io_check_env_pmp_6_cfg_r | res_pmp_ignore_6; // @[PMP.scala 438:42]
  wire  res_pmp_cur_6_cfg_w = io_check_env_pmp_6_cfg_w | res_pmp_ignore_6; // @[PMP.scala 439:42]
  wire  res_pmp_cur_6_cfg_x = io_check_env_pmp_6_cfg_x | res_pmp_ignore_6; // @[PMP.scala 440:42]
  wire [35:0] _res_pmp_is_match_T_148 = {io_check_env_pmp_7_addr, 2'h0}; // @[PMP.scala 190:35]
  wire [35:0] _res_pmp_is_match_T_150 = _res_pmp_is_match_T_148 & 36'hffffff000; // @[PMP.scala 190:50]
  wire [35:0] _res_pmp_is_match_T_151 = ~io_check_env_pmp_7_mask; // @[PMP.scala 232:10]
  wire [35:0] _res_pmp_is_match_T_152 = io_req_bits_addr & _res_pmp_is_match_T_151; // @[PMP.scala 232:8]
  wire [35:0] _res_pmp_is_match_T_154 = _res_pmp_is_match_T_150 & _res_pmp_is_match_T_151; // @[PMP.scala 232:21]
  wire  _res_pmp_is_match_T_155 = _res_pmp_is_match_T_152 == _res_pmp_is_match_T_154; // @[PMP.scala 232:14]
  wire  _res_pmp_is_match_T_156 = io_check_env_pmp_7_cfg_a == 2'h1; // @[PMP.scala 53:15]
  wire  _res_pmp_is_match_T_161 = ~_res_pmp_is_match_T_144; // @[PMP.scala 220:5]
  wire  _res_pmp_is_match_T_165 = io_req_bits_addr < _res_pmp_is_match_T_150; // @[PMP.scala 210:14]
  wire  _res_pmp_is_match_T_166 = _res_pmp_is_match_T_161 & _res_pmp_is_match_T_165; // @[PMP.scala 228:56]
  wire  _res_pmp_is_match_T_167 = _res_pmp_is_match_T_156 & _res_pmp_is_match_T_166; // @[PMP.scala 200:10]
  wire  res_pmp_ignore_7 = res_pmp_passThrough & ~io_check_env_pmp_7_cfg_l; // @[PMP.scala 434:32]
  wire  res_pmp_cur_7_cfg_r = io_check_env_pmp_7_cfg_r | res_pmp_ignore_7; // @[PMP.scala 438:42]
  wire  res_pmp_cur_7_cfg_w = io_check_env_pmp_7_cfg_w | res_pmp_ignore_7; // @[PMP.scala 439:42]
  wire  res_pmp_cur_7_cfg_x = io_check_env_pmp_7_cfg_x | res_pmp_ignore_7; // @[PMP.scala 440:42]
  wire [35:0] _res_pmp_is_match_T_169 = {io_check_env_pmp_8_addr, 2'h0}; // @[PMP.scala 190:35]
  wire [35:0] _res_pmp_is_match_T_171 = _res_pmp_is_match_T_169 & 36'hffffff000; // @[PMP.scala 190:50]
  wire [35:0] _res_pmp_is_match_T_172 = ~io_check_env_pmp_8_mask; // @[PMP.scala 232:10]
  wire [35:0] _res_pmp_is_match_T_173 = io_req_bits_addr & _res_pmp_is_match_T_172; // @[PMP.scala 232:8]
  wire [35:0] _res_pmp_is_match_T_175 = _res_pmp_is_match_T_171 & _res_pmp_is_match_T_172; // @[PMP.scala 232:21]
  wire  _res_pmp_is_match_T_176 = _res_pmp_is_match_T_173 == _res_pmp_is_match_T_175; // @[PMP.scala 232:14]
  wire  _res_pmp_is_match_T_177 = io_check_env_pmp_8_cfg_a == 2'h1; // @[PMP.scala 53:15]
  wire  _res_pmp_is_match_T_182 = ~_res_pmp_is_match_T_165; // @[PMP.scala 220:5]
  wire  _res_pmp_is_match_T_186 = io_req_bits_addr < _res_pmp_is_match_T_171; // @[PMP.scala 210:14]
  wire  _res_pmp_is_match_T_187 = _res_pmp_is_match_T_182 & _res_pmp_is_match_T_186; // @[PMP.scala 228:56]
  wire  _res_pmp_is_match_T_188 = _res_pmp_is_match_T_177 & _res_pmp_is_match_T_187; // @[PMP.scala 200:10]
  wire  res_pmp_ignore_8 = res_pmp_passThrough & ~io_check_env_pmp_8_cfg_l; // @[PMP.scala 434:32]
  wire  res_pmp_cur_8_cfg_r = io_check_env_pmp_8_cfg_r | res_pmp_ignore_8; // @[PMP.scala 438:42]
  wire  res_pmp_cur_8_cfg_w = io_check_env_pmp_8_cfg_w | res_pmp_ignore_8; // @[PMP.scala 439:42]
  wire  res_pmp_cur_8_cfg_x = io_check_env_pmp_8_cfg_x | res_pmp_ignore_8; // @[PMP.scala 440:42]
  wire [35:0] _res_pmp_is_match_T_190 = {io_check_env_pmp_9_addr, 2'h0}; // @[PMP.scala 190:35]
  wire [35:0] _res_pmp_is_match_T_192 = _res_pmp_is_match_T_190 & 36'hffffff000; // @[PMP.scala 190:50]
  wire [35:0] _res_pmp_is_match_T_193 = ~io_check_env_pmp_9_mask; // @[PMP.scala 232:10]
  wire [35:0] _res_pmp_is_match_T_194 = io_req_bits_addr & _res_pmp_is_match_T_193; // @[PMP.scala 232:8]
  wire [35:0] _res_pmp_is_match_T_196 = _res_pmp_is_match_T_192 & _res_pmp_is_match_T_193; // @[PMP.scala 232:21]
  wire  _res_pmp_is_match_T_197 = _res_pmp_is_match_T_194 == _res_pmp_is_match_T_196; // @[PMP.scala 232:14]
  wire  _res_pmp_is_match_T_198 = io_check_env_pmp_9_cfg_a == 2'h1; // @[PMP.scala 53:15]
  wire  _res_pmp_is_match_T_203 = ~_res_pmp_is_match_T_186; // @[PMP.scala 220:5]
  wire  _res_pmp_is_match_T_207 = io_req_bits_addr < _res_pmp_is_match_T_192; // @[PMP.scala 210:14]
  wire  _res_pmp_is_match_T_208 = _res_pmp_is_match_T_203 & _res_pmp_is_match_T_207; // @[PMP.scala 228:56]
  wire  _res_pmp_is_match_T_209 = _res_pmp_is_match_T_198 & _res_pmp_is_match_T_208; // @[PMP.scala 200:10]
  wire  res_pmp_ignore_9 = res_pmp_passThrough & ~io_check_env_pmp_9_cfg_l; // @[PMP.scala 434:32]
  wire  res_pmp_cur_9_cfg_r = io_check_env_pmp_9_cfg_r | res_pmp_ignore_9; // @[PMP.scala 438:42]
  wire  res_pmp_cur_9_cfg_w = io_check_env_pmp_9_cfg_w | res_pmp_ignore_9; // @[PMP.scala 439:42]
  wire  res_pmp_cur_9_cfg_x = io_check_env_pmp_9_cfg_x | res_pmp_ignore_9; // @[PMP.scala 440:42]
  wire [35:0] _res_pmp_is_match_T_211 = {io_check_env_pmp_10_addr, 2'h0}; // @[PMP.scala 190:35]
  wire [35:0] _res_pmp_is_match_T_213 = _res_pmp_is_match_T_211 & 36'hffffff000; // @[PMP.scala 190:50]
  wire [35:0] _res_pmp_is_match_T_214 = ~io_check_env_pmp_10_mask; // @[PMP.scala 232:10]
  wire [35:0] _res_pmp_is_match_T_215 = io_req_bits_addr & _res_pmp_is_match_T_214; // @[PMP.scala 232:8]
  wire [35:0] _res_pmp_is_match_T_217 = _res_pmp_is_match_T_213 & _res_pmp_is_match_T_214; // @[PMP.scala 232:21]
  wire  _res_pmp_is_match_T_218 = _res_pmp_is_match_T_215 == _res_pmp_is_match_T_217; // @[PMP.scala 232:14]
  wire  _res_pmp_is_match_T_219 = io_check_env_pmp_10_cfg_a == 2'h1; // @[PMP.scala 53:15]
  wire  _res_pmp_is_match_T_224 = ~_res_pmp_is_match_T_207; // @[PMP.scala 220:5]
  wire  _res_pmp_is_match_T_228 = io_req_bits_addr < _res_pmp_is_match_T_213; // @[PMP.scala 210:14]
  wire  _res_pmp_is_match_T_229 = _res_pmp_is_match_T_224 & _res_pmp_is_match_T_228; // @[PMP.scala 228:56]
  wire  _res_pmp_is_match_T_230 = _res_pmp_is_match_T_219 & _res_pmp_is_match_T_229; // @[PMP.scala 200:10]
  wire  res_pmp_ignore_10 = res_pmp_passThrough & ~io_check_env_pmp_10_cfg_l; // @[PMP.scala 434:32]
  wire  res_pmp_cur_10_cfg_r = io_check_env_pmp_10_cfg_r | res_pmp_ignore_10; // @[PMP.scala 438:42]
  wire  res_pmp_cur_10_cfg_w = io_check_env_pmp_10_cfg_w | res_pmp_ignore_10; // @[PMP.scala 439:42]
  wire  res_pmp_cur_10_cfg_x = io_check_env_pmp_10_cfg_x | res_pmp_ignore_10; // @[PMP.scala 440:42]
  wire [35:0] _res_pmp_is_match_T_232 = {io_check_env_pmp_11_addr, 2'h0}; // @[PMP.scala 190:35]
  wire [35:0] _res_pmp_is_match_T_234 = _res_pmp_is_match_T_232 & 36'hffffff000; // @[PMP.scala 190:50]
  wire [35:0] _res_pmp_is_match_T_235 = ~io_check_env_pmp_11_mask; // @[PMP.scala 232:10]
  wire [35:0] _res_pmp_is_match_T_236 = io_req_bits_addr & _res_pmp_is_match_T_235; // @[PMP.scala 232:8]
  wire [35:0] _res_pmp_is_match_T_238 = _res_pmp_is_match_T_234 & _res_pmp_is_match_T_235; // @[PMP.scala 232:21]
  wire  _res_pmp_is_match_T_239 = _res_pmp_is_match_T_236 == _res_pmp_is_match_T_238; // @[PMP.scala 232:14]
  wire  _res_pmp_is_match_T_240 = io_check_env_pmp_11_cfg_a == 2'h1; // @[PMP.scala 53:15]
  wire  _res_pmp_is_match_T_245 = ~_res_pmp_is_match_T_228; // @[PMP.scala 220:5]
  wire  _res_pmp_is_match_T_249 = io_req_bits_addr < _res_pmp_is_match_T_234; // @[PMP.scala 210:14]
  wire  _res_pmp_is_match_T_250 = _res_pmp_is_match_T_245 & _res_pmp_is_match_T_249; // @[PMP.scala 228:56]
  wire  _res_pmp_is_match_T_251 = _res_pmp_is_match_T_240 & _res_pmp_is_match_T_250; // @[PMP.scala 200:10]
  wire  res_pmp_ignore_11 = res_pmp_passThrough & ~io_check_env_pmp_11_cfg_l; // @[PMP.scala 434:32]
  wire  res_pmp_cur_11_cfg_r = io_check_env_pmp_11_cfg_r | res_pmp_ignore_11; // @[PMP.scala 438:42]
  wire  res_pmp_cur_11_cfg_w = io_check_env_pmp_11_cfg_w | res_pmp_ignore_11; // @[PMP.scala 439:42]
  wire  res_pmp_cur_11_cfg_x = io_check_env_pmp_11_cfg_x | res_pmp_ignore_11; // @[PMP.scala 440:42]
  wire [35:0] _res_pmp_is_match_T_253 = {io_check_env_pmp_12_addr, 2'h0}; // @[PMP.scala 190:35]
  wire [35:0] _res_pmp_is_match_T_255 = _res_pmp_is_match_T_253 & 36'hffffff000; // @[PMP.scala 190:50]
  wire [35:0] _res_pmp_is_match_T_256 = ~io_check_env_pmp_12_mask; // @[PMP.scala 232:10]
  wire [35:0] _res_pmp_is_match_T_257 = io_req_bits_addr & _res_pmp_is_match_T_256; // @[PMP.scala 232:8]
  wire [35:0] _res_pmp_is_match_T_259 = _res_pmp_is_match_T_255 & _res_pmp_is_match_T_256; // @[PMP.scala 232:21]
  wire  _res_pmp_is_match_T_260 = _res_pmp_is_match_T_257 == _res_pmp_is_match_T_259; // @[PMP.scala 232:14]
  wire  _res_pmp_is_match_T_261 = io_check_env_pmp_12_cfg_a == 2'h1; // @[PMP.scala 53:15]
  wire  _res_pmp_is_match_T_266 = ~_res_pmp_is_match_T_249; // @[PMP.scala 220:5]
  wire  _res_pmp_is_match_T_270 = io_req_bits_addr < _res_pmp_is_match_T_255; // @[PMP.scala 210:14]
  wire  _res_pmp_is_match_T_271 = _res_pmp_is_match_T_266 & _res_pmp_is_match_T_270; // @[PMP.scala 228:56]
  wire  _res_pmp_is_match_T_272 = _res_pmp_is_match_T_261 & _res_pmp_is_match_T_271; // @[PMP.scala 200:10]
  wire  res_pmp_ignore_12 = res_pmp_passThrough & ~io_check_env_pmp_12_cfg_l; // @[PMP.scala 434:32]
  wire  res_pmp_cur_12_cfg_r = io_check_env_pmp_12_cfg_r | res_pmp_ignore_12; // @[PMP.scala 438:42]
  wire  res_pmp_cur_12_cfg_w = io_check_env_pmp_12_cfg_w | res_pmp_ignore_12; // @[PMP.scala 439:42]
  wire  res_pmp_cur_12_cfg_x = io_check_env_pmp_12_cfg_x | res_pmp_ignore_12; // @[PMP.scala 440:42]
  wire [35:0] _res_pmp_is_match_T_274 = {io_check_env_pmp_13_addr, 2'h0}; // @[PMP.scala 190:35]
  wire [35:0] _res_pmp_is_match_T_276 = _res_pmp_is_match_T_274 & 36'hffffff000; // @[PMP.scala 190:50]
  wire [35:0] _res_pmp_is_match_T_277 = ~io_check_env_pmp_13_mask; // @[PMP.scala 232:10]
  wire [35:0] _res_pmp_is_match_T_278 = io_req_bits_addr & _res_pmp_is_match_T_277; // @[PMP.scala 232:8]
  wire [35:0] _res_pmp_is_match_T_280 = _res_pmp_is_match_T_276 & _res_pmp_is_match_T_277; // @[PMP.scala 232:21]
  wire  _res_pmp_is_match_T_281 = _res_pmp_is_match_T_278 == _res_pmp_is_match_T_280; // @[PMP.scala 232:14]
  wire  _res_pmp_is_match_T_282 = io_check_env_pmp_13_cfg_a == 2'h1; // @[PMP.scala 53:15]
  wire  _res_pmp_is_match_T_287 = ~_res_pmp_is_match_T_270; // @[PMP.scala 220:5]
  wire  _res_pmp_is_match_T_291 = io_req_bits_addr < _res_pmp_is_match_T_276; // @[PMP.scala 210:14]
  wire  _res_pmp_is_match_T_292 = _res_pmp_is_match_T_287 & _res_pmp_is_match_T_291; // @[PMP.scala 228:56]
  wire  _res_pmp_is_match_T_293 = _res_pmp_is_match_T_282 & _res_pmp_is_match_T_292; // @[PMP.scala 200:10]
  wire  res_pmp_ignore_13 = res_pmp_passThrough & ~io_check_env_pmp_13_cfg_l; // @[PMP.scala 434:32]
  wire  res_pmp_cur_13_cfg_r = io_check_env_pmp_13_cfg_r | res_pmp_ignore_13; // @[PMP.scala 438:42]
  wire  res_pmp_cur_13_cfg_w = io_check_env_pmp_13_cfg_w | res_pmp_ignore_13; // @[PMP.scala 439:42]
  wire  res_pmp_cur_13_cfg_x = io_check_env_pmp_13_cfg_x | res_pmp_ignore_13; // @[PMP.scala 440:42]
  wire [35:0] _res_pmp_is_match_T_295 = {io_check_env_pmp_14_addr, 2'h0}; // @[PMP.scala 190:35]
  wire [35:0] _res_pmp_is_match_T_297 = _res_pmp_is_match_T_295 & 36'hffffff000; // @[PMP.scala 190:50]
  wire [35:0] _res_pmp_is_match_T_298 = ~io_check_env_pmp_14_mask; // @[PMP.scala 232:10]
  wire [35:0] _res_pmp_is_match_T_299 = io_req_bits_addr & _res_pmp_is_match_T_298; // @[PMP.scala 232:8]
  wire [35:0] _res_pmp_is_match_T_301 = _res_pmp_is_match_T_297 & _res_pmp_is_match_T_298; // @[PMP.scala 232:21]
  wire  _res_pmp_is_match_T_302 = _res_pmp_is_match_T_299 == _res_pmp_is_match_T_301; // @[PMP.scala 232:14]
  wire  _res_pmp_is_match_T_303 = io_check_env_pmp_14_cfg_a == 2'h1; // @[PMP.scala 53:15]
  wire  _res_pmp_is_match_T_308 = ~_res_pmp_is_match_T_291; // @[PMP.scala 220:5]
  wire  _res_pmp_is_match_T_312 = io_req_bits_addr < _res_pmp_is_match_T_297; // @[PMP.scala 210:14]
  wire  _res_pmp_is_match_T_313 = _res_pmp_is_match_T_308 & _res_pmp_is_match_T_312; // @[PMP.scala 228:56]
  wire  _res_pmp_is_match_T_314 = _res_pmp_is_match_T_303 & _res_pmp_is_match_T_313; // @[PMP.scala 200:10]
  wire  res_pmp_ignore_14 = res_pmp_passThrough & ~io_check_env_pmp_14_cfg_l; // @[PMP.scala 434:32]
  wire  res_pmp_cur_14_cfg_r = io_check_env_pmp_14_cfg_r | res_pmp_ignore_14; // @[PMP.scala 438:42]
  wire  res_pmp_cur_14_cfg_w = io_check_env_pmp_14_cfg_w | res_pmp_ignore_14; // @[PMP.scala 439:42]
  wire  res_pmp_cur_14_cfg_x = io_check_env_pmp_14_cfg_x | res_pmp_ignore_14; // @[PMP.scala 440:42]
  wire [35:0] _res_pmp_is_match_T_316 = {io_check_env_pmp_15_addr, 2'h0}; // @[PMP.scala 190:35]
  wire [35:0] _res_pmp_is_match_T_318 = _res_pmp_is_match_T_316 & 36'hffffff000; // @[PMP.scala 190:50]
  wire [35:0] _res_pmp_is_match_T_319 = ~io_check_env_pmp_15_mask; // @[PMP.scala 232:10]
  wire [35:0] _res_pmp_is_match_T_320 = io_req_bits_addr & _res_pmp_is_match_T_319; // @[PMP.scala 232:8]
  wire [35:0] _res_pmp_is_match_T_322 = _res_pmp_is_match_T_318 & _res_pmp_is_match_T_319; // @[PMP.scala 232:21]
  wire  _res_pmp_is_match_T_323 = _res_pmp_is_match_T_320 == _res_pmp_is_match_T_322; // @[PMP.scala 232:14]
  wire  _res_pmp_is_match_T_324 = io_check_env_pmp_15_cfg_a == 2'h1; // @[PMP.scala 53:15]
  wire  _res_pmp_is_match_T_329 = ~_res_pmp_is_match_T_312; // @[PMP.scala 220:5]
  wire  _res_pmp_is_match_T_333 = io_req_bits_addr < _res_pmp_is_match_T_318; // @[PMP.scala 210:14]
  wire  _res_pmp_is_match_T_334 = _res_pmp_is_match_T_329 & _res_pmp_is_match_T_333; // @[PMP.scala 228:56]
  wire  _res_pmp_is_match_T_335 = _res_pmp_is_match_T_324 & _res_pmp_is_match_T_334; // @[PMP.scala 200:10]
  wire  res_pmp_ignore_15 = res_pmp_passThrough & ~io_check_env_pmp_15_cfg_l; // @[PMP.scala 434:32]
  wire  res_pmp_cur_15_cfg_r = io_check_env_pmp_15_cfg_r | res_pmp_ignore_15; // @[PMP.scala 438:42]
  wire  res_pmp_cur_15_cfg_w = io_check_env_pmp_15_cfg_w | res_pmp_ignore_15; // @[PMP.scala 439:42]
  wire  res_pmp_cur_15_cfg_x = io_check_env_pmp_15_cfg_x | res_pmp_ignore_15; // @[PMP.scala 440:42]
  reg  res_pmp_r; // @[Reg.scala 28:20]
  reg  res_pmp_r1; // @[Reg.scala 28:20]
  reg  res_pmp_r2; // @[Reg.scala 28:20]
  reg  res_pmp_r3; // @[Reg.scala 28:20]
  reg  res_pmp_r4; // @[Reg.scala 28:20]
  reg  res_pmp_r5; // @[Reg.scala 28:20]
  reg  res_pmp_r6; // @[Reg.scala 28:20]
  reg  res_pmp_r7; // @[Reg.scala 28:20]
  reg  res_pmp_r8; // @[Reg.scala 28:20]
  reg  res_pmp_r9; // @[Reg.scala 28:20]
  reg  res_pmp_r10; // @[Reg.scala 28:20]
  reg  res_pmp_r11; // @[Reg.scala 28:20]
  reg  res_pmp_r12; // @[Reg.scala 28:20]
  reg  res_pmp_r13; // @[Reg.scala 28:20]
  reg  res_pmp_r14; // @[Reg.scala 28:20]
  reg  res_pmp_r15; // @[Reg.scala 28:20]
  reg  res_pmp_r17_0_cfg_x; // @[Reg.scala 16:16]
  reg  res_pmp_r17_0_cfg_w; // @[Reg.scala 16:16]
  reg  res_pmp_r17_0_cfg_r; // @[Reg.scala 16:16]
  reg  res_pmp_r17_1_cfg_x; // @[Reg.scala 16:16]
  reg  res_pmp_r17_1_cfg_w; // @[Reg.scala 16:16]
  reg  res_pmp_r17_1_cfg_r; // @[Reg.scala 16:16]
  reg  res_pmp_r17_2_cfg_x; // @[Reg.scala 16:16]
  reg  res_pmp_r17_2_cfg_w; // @[Reg.scala 16:16]
  reg  res_pmp_r17_2_cfg_r; // @[Reg.scala 16:16]
  reg  res_pmp_r17_3_cfg_x; // @[Reg.scala 16:16]
  reg  res_pmp_r17_3_cfg_w; // @[Reg.scala 16:16]
  reg  res_pmp_r17_3_cfg_r; // @[Reg.scala 16:16]
  reg  res_pmp_r17_4_cfg_x; // @[Reg.scala 16:16]
  reg  res_pmp_r17_4_cfg_w; // @[Reg.scala 16:16]
  reg  res_pmp_r17_4_cfg_r; // @[Reg.scala 16:16]
  reg  res_pmp_r17_5_cfg_x; // @[Reg.scala 16:16]
  reg  res_pmp_r17_5_cfg_w; // @[Reg.scala 16:16]
  reg  res_pmp_r17_5_cfg_r; // @[Reg.scala 16:16]
  reg  res_pmp_r17_6_cfg_x; // @[Reg.scala 16:16]
  reg  res_pmp_r17_6_cfg_w; // @[Reg.scala 16:16]
  reg  res_pmp_r17_6_cfg_r; // @[Reg.scala 16:16]
  reg  res_pmp_r17_7_cfg_x; // @[Reg.scala 16:16]
  reg  res_pmp_r17_7_cfg_w; // @[Reg.scala 16:16]
  reg  res_pmp_r17_7_cfg_r; // @[Reg.scala 16:16]
  reg  res_pmp_r17_8_cfg_x; // @[Reg.scala 16:16]
  reg  res_pmp_r17_8_cfg_w; // @[Reg.scala 16:16]
  reg  res_pmp_r17_8_cfg_r; // @[Reg.scala 16:16]
  reg  res_pmp_r17_9_cfg_x; // @[Reg.scala 16:16]
  reg  res_pmp_r17_9_cfg_w; // @[Reg.scala 16:16]
  reg  res_pmp_r17_9_cfg_r; // @[Reg.scala 16:16]
  reg  res_pmp_r17_10_cfg_x; // @[Reg.scala 16:16]
  reg  res_pmp_r17_10_cfg_w; // @[Reg.scala 16:16]
  reg  res_pmp_r17_10_cfg_r; // @[Reg.scala 16:16]
  reg  res_pmp_r17_11_cfg_x; // @[Reg.scala 16:16]
  reg  res_pmp_r17_11_cfg_w; // @[Reg.scala 16:16]
  reg  res_pmp_r17_11_cfg_r; // @[Reg.scala 16:16]
  reg  res_pmp_r17_12_cfg_x; // @[Reg.scala 16:16]
  reg  res_pmp_r17_12_cfg_w; // @[Reg.scala 16:16]
  reg  res_pmp_r17_12_cfg_r; // @[Reg.scala 16:16]
  reg  res_pmp_r17_13_cfg_x; // @[Reg.scala 16:16]
  reg  res_pmp_r17_13_cfg_w; // @[Reg.scala 16:16]
  reg  res_pmp_r17_13_cfg_r; // @[Reg.scala 16:16]
  reg  res_pmp_r17_14_cfg_x; // @[Reg.scala 16:16]
  reg  res_pmp_r17_14_cfg_w; // @[Reg.scala 16:16]
  reg  res_pmp_r17_14_cfg_r; // @[Reg.scala 16:16]
  reg  res_pmp_r17_15_cfg_x; // @[Reg.scala 16:16]
  reg  res_pmp_r17_15_cfg_w; // @[Reg.scala 16:16]
  reg  res_pmp_r17_15_cfg_r; // @[Reg.scala 16:16]
  reg  res_pmp_r17_16_cfg_x; // @[Reg.scala 16:16]
  reg  res_pmp_r17_16_cfg_w; // @[Reg.scala 16:16]
  reg  res_pmp_r17_16_cfg_r; // @[Reg.scala 16:16]
  wire  _res_pmp_T_1_cfg_x = res_pmp_r ? res_pmp_r17_0_cfg_x : res_pmp_r17_1_cfg_x; // @[ParallelMux.scala 90:77]
  wire  _res_pmp_T_1_cfg_w = res_pmp_r ? res_pmp_r17_0_cfg_w : res_pmp_r17_1_cfg_w; // @[ParallelMux.scala 90:77]
  wire  _res_pmp_T_1_cfg_r = res_pmp_r ? res_pmp_r17_0_cfg_r : res_pmp_r17_1_cfg_r; // @[ParallelMux.scala 90:77]
  wire  _res_pmp_T_3_cfg_x = res_pmp_r2 ? res_pmp_r17_2_cfg_x : res_pmp_r17_3_cfg_x; // @[ParallelMux.scala 90:77]
  wire  _res_pmp_T_3_cfg_w = res_pmp_r2 ? res_pmp_r17_2_cfg_w : res_pmp_r17_3_cfg_w; // @[ParallelMux.scala 90:77]
  wire  _res_pmp_T_3_cfg_r = res_pmp_r2 ? res_pmp_r17_2_cfg_r : res_pmp_r17_3_cfg_r; // @[ParallelMux.scala 90:77]
  wire  _res_pmp_T_5_cfg_x = res_pmp_r | res_pmp_r1 ? _res_pmp_T_1_cfg_x : _res_pmp_T_3_cfg_x; // @[ParallelMux.scala 90:77]
  wire  _res_pmp_T_5_cfg_w = res_pmp_r | res_pmp_r1 ? _res_pmp_T_1_cfg_w : _res_pmp_T_3_cfg_w; // @[ParallelMux.scala 90:77]
  wire  _res_pmp_T_5_cfg_r = res_pmp_r | res_pmp_r1 ? _res_pmp_T_1_cfg_r : _res_pmp_T_3_cfg_r; // @[ParallelMux.scala 90:77]
  wire  _res_pmp_T_7_cfg_x = res_pmp_r4 ? res_pmp_r17_4_cfg_x : res_pmp_r17_5_cfg_x; // @[ParallelMux.scala 90:77]
  wire  _res_pmp_T_7_cfg_w = res_pmp_r4 ? res_pmp_r17_4_cfg_w : res_pmp_r17_5_cfg_w; // @[ParallelMux.scala 90:77]
  wire  _res_pmp_T_7_cfg_r = res_pmp_r4 ? res_pmp_r17_4_cfg_r : res_pmp_r17_5_cfg_r; // @[ParallelMux.scala 90:77]
  wire  _res_pmp_T_9_cfg_x = res_pmp_r6 ? res_pmp_r17_6_cfg_x : res_pmp_r17_7_cfg_x; // @[ParallelMux.scala 90:77]
  wire  _res_pmp_T_9_cfg_w = res_pmp_r6 ? res_pmp_r17_6_cfg_w : res_pmp_r17_7_cfg_w; // @[ParallelMux.scala 90:77]
  wire  _res_pmp_T_9_cfg_r = res_pmp_r6 ? res_pmp_r17_6_cfg_r : res_pmp_r17_7_cfg_r; // @[ParallelMux.scala 90:77]
  wire  _res_pmp_T_11_cfg_x = res_pmp_r4 | res_pmp_r5 ? _res_pmp_T_7_cfg_x : _res_pmp_T_9_cfg_x; // @[ParallelMux.scala 90:77]
  wire  _res_pmp_T_11_cfg_w = res_pmp_r4 | res_pmp_r5 ? _res_pmp_T_7_cfg_w : _res_pmp_T_9_cfg_w; // @[ParallelMux.scala 90:77]
  wire  _res_pmp_T_11_cfg_r = res_pmp_r4 | res_pmp_r5 ? _res_pmp_T_7_cfg_r : _res_pmp_T_9_cfg_r; // @[ParallelMux.scala 90:77]
  wire  _res_pmp_T_13_cfg_x = res_pmp_r | res_pmp_r1 | (res_pmp_r2 | res_pmp_r3) ? _res_pmp_T_5_cfg_x :
    _res_pmp_T_11_cfg_x; // @[ParallelMux.scala 90:77]
  wire  _res_pmp_T_13_cfg_w = res_pmp_r | res_pmp_r1 | (res_pmp_r2 | res_pmp_r3) ? _res_pmp_T_5_cfg_w :
    _res_pmp_T_11_cfg_w; // @[ParallelMux.scala 90:77]
  wire  _res_pmp_T_13_cfg_r = res_pmp_r | res_pmp_r1 | (res_pmp_r2 | res_pmp_r3) ? _res_pmp_T_5_cfg_r :
    _res_pmp_T_11_cfg_r; // @[ParallelMux.scala 90:77]
  wire  _res_pmp_T_15_cfg_x = res_pmp_r8 ? res_pmp_r17_8_cfg_x : res_pmp_r17_9_cfg_x; // @[ParallelMux.scala 90:77]
  wire  _res_pmp_T_15_cfg_w = res_pmp_r8 ? res_pmp_r17_8_cfg_w : res_pmp_r17_9_cfg_w; // @[ParallelMux.scala 90:77]
  wire  _res_pmp_T_15_cfg_r = res_pmp_r8 ? res_pmp_r17_8_cfg_r : res_pmp_r17_9_cfg_r; // @[ParallelMux.scala 90:77]
  wire  _res_pmp_T_17_cfg_x = res_pmp_r10 ? res_pmp_r17_10_cfg_x : res_pmp_r17_11_cfg_x; // @[ParallelMux.scala 90:77]
  wire  _res_pmp_T_17_cfg_w = res_pmp_r10 ? res_pmp_r17_10_cfg_w : res_pmp_r17_11_cfg_w; // @[ParallelMux.scala 90:77]
  wire  _res_pmp_T_17_cfg_r = res_pmp_r10 ? res_pmp_r17_10_cfg_r : res_pmp_r17_11_cfg_r; // @[ParallelMux.scala 90:77]
  wire  _res_pmp_T_19_cfg_x = res_pmp_r8 | res_pmp_r9 ? _res_pmp_T_15_cfg_x : _res_pmp_T_17_cfg_x; // @[ParallelMux.scala 90:77]
  wire  _res_pmp_T_19_cfg_w = res_pmp_r8 | res_pmp_r9 ? _res_pmp_T_15_cfg_w : _res_pmp_T_17_cfg_w; // @[ParallelMux.scala 90:77]
  wire  _res_pmp_T_19_cfg_r = res_pmp_r8 | res_pmp_r9 ? _res_pmp_T_15_cfg_r : _res_pmp_T_17_cfg_r; // @[ParallelMux.scala 90:77]
  wire  _res_pmp_T_21_cfg_x = res_pmp_r12 ? res_pmp_r17_12_cfg_x : res_pmp_r17_13_cfg_x; // @[ParallelMux.scala 90:77]
  wire  _res_pmp_T_21_cfg_w = res_pmp_r12 ? res_pmp_r17_12_cfg_w : res_pmp_r17_13_cfg_w; // @[ParallelMux.scala 90:77]
  wire  _res_pmp_T_21_cfg_r = res_pmp_r12 ? res_pmp_r17_12_cfg_r : res_pmp_r17_13_cfg_r; // @[ParallelMux.scala 90:77]
  wire  _res_pmp_T_23_cfg_x = res_pmp_r15 ? res_pmp_r17_15_cfg_x : res_pmp_r17_16_cfg_x; // @[ParallelMux.scala 90:77]
  wire  _res_pmp_T_23_cfg_w = res_pmp_r15 ? res_pmp_r17_15_cfg_w : res_pmp_r17_16_cfg_w; // @[ParallelMux.scala 90:77]
  wire  _res_pmp_T_23_cfg_r = res_pmp_r15 ? res_pmp_r17_15_cfg_r : res_pmp_r17_16_cfg_r; // @[ParallelMux.scala 90:77]
  wire  _res_pmp_T_25_cfg_x = res_pmp_r14 ? res_pmp_r17_14_cfg_x : _res_pmp_T_23_cfg_x; // @[ParallelMux.scala 90:77]
  wire  _res_pmp_T_25_cfg_w = res_pmp_r14 ? res_pmp_r17_14_cfg_w : _res_pmp_T_23_cfg_w; // @[ParallelMux.scala 90:77]
  wire  _res_pmp_T_25_cfg_r = res_pmp_r14 ? res_pmp_r17_14_cfg_r : _res_pmp_T_23_cfg_r; // @[ParallelMux.scala 90:77]
  wire  _res_pmp_T_27_cfg_x = res_pmp_r12 | res_pmp_r13 ? _res_pmp_T_21_cfg_x : _res_pmp_T_25_cfg_x; // @[ParallelMux.scala 90:77]
  wire  _res_pmp_T_27_cfg_w = res_pmp_r12 | res_pmp_r13 ? _res_pmp_T_21_cfg_w : _res_pmp_T_25_cfg_w; // @[ParallelMux.scala 90:77]
  wire  _res_pmp_T_27_cfg_r = res_pmp_r12 | res_pmp_r13 ? _res_pmp_T_21_cfg_r : _res_pmp_T_25_cfg_r; // @[ParallelMux.scala 90:77]
  wire  _res_pmp_T_29_cfg_x = res_pmp_r8 | res_pmp_r9 | (res_pmp_r10 | res_pmp_r11) ? _res_pmp_T_19_cfg_x :
    _res_pmp_T_27_cfg_x; // @[ParallelMux.scala 90:77]
  wire  _res_pmp_T_29_cfg_w = res_pmp_r8 | res_pmp_r9 | (res_pmp_r10 | res_pmp_r11) ? _res_pmp_T_19_cfg_w :
    _res_pmp_T_27_cfg_w; // @[ParallelMux.scala 90:77]
  wire  _res_pmp_T_29_cfg_r = res_pmp_r8 | res_pmp_r9 | (res_pmp_r10 | res_pmp_r11) ? _res_pmp_T_19_cfg_r :
    _res_pmp_T_27_cfg_r; // @[ParallelMux.scala 90:77]
  wire  res_pmp_cfg_x = res_pmp_r | res_pmp_r1 | (res_pmp_r2 | res_pmp_r3) | (res_pmp_r4 | res_pmp_r5 | (
    res_pmp_r6 | res_pmp_r7)) ? _res_pmp_T_13_cfg_x : _res_pmp_T_29_cfg_x; // @[ParallelMux.scala 90:77]
  wire  res_pmp_cfg_w = res_pmp_r | res_pmp_r1 | (res_pmp_r2 | res_pmp_r3) | (res_pmp_r4 | res_pmp_r5 | (
    res_pmp_r6 | res_pmp_r7)) ? _res_pmp_T_13_cfg_w : _res_pmp_T_29_cfg_w; // @[ParallelMux.scala 90:77]
  wire  res_pmp_cfg_r = res_pmp_r | res_pmp_r1 | (res_pmp_r2 | res_pmp_r3) | (res_pmp_r4 | res_pmp_r5 | (
    res_pmp_r6 | res_pmp_r7)) ? _res_pmp_T_13_cfg_r : _res_pmp_T_29_cfg_r; // @[ParallelMux.scala 90:77]
  wire [35:0] _res_pma_is_match_T_1 = {io_check_env_pma_0_addr, 2'h0}; // @[PMP.scala 190:35]
  wire [35:0] _res_pma_is_match_T_3 = _res_pma_is_match_T_1 & 36'hffffff000; // @[PMP.scala 190:50]
  wire [35:0] _res_pma_is_match_T_4 = ~io_check_env_pma_0_mask; // @[PMP.scala 232:10]
  wire [35:0] _res_pma_is_match_T_5 = io_req_bits_addr & _res_pma_is_match_T_4; // @[PMP.scala 232:8]
  wire [35:0] _res_pma_is_match_T_7 = _res_pma_is_match_T_3 & _res_pma_is_match_T_4; // @[PMP.scala 232:21]
  wire  _res_pma_is_match_T_8 = _res_pma_is_match_T_5 == _res_pma_is_match_T_7; // @[PMP.scala 232:14]
  wire  _res_pma_is_match_T_9 = io_check_env_pma_0_cfg_a == 2'h1; // @[PMP.scala 53:15]
  wire  _res_pma_is_match_T_18 = io_req_bits_addr < _res_pma_is_match_T_3; // @[PMP.scala 210:14]
  wire  _res_pma_is_match_T_20 = _res_pma_is_match_T_9 & _res_pma_is_match_T_18; // @[PMP.scala 200:10]
  wire [35:0] _res_pma_is_match_T_22 = {io_check_env_pma_1_addr, 2'h0}; // @[PMP.scala 190:35]
  wire [35:0] _res_pma_is_match_T_24 = _res_pma_is_match_T_22 & 36'hffffff000; // @[PMP.scala 190:50]
  wire [35:0] _res_pma_is_match_T_25 = ~io_check_env_pma_1_mask; // @[PMP.scala 232:10]
  wire [35:0] _res_pma_is_match_T_26 = io_req_bits_addr & _res_pma_is_match_T_25; // @[PMP.scala 232:8]
  wire [35:0] _res_pma_is_match_T_28 = _res_pma_is_match_T_24 & _res_pma_is_match_T_25; // @[PMP.scala 232:21]
  wire  _res_pma_is_match_T_29 = _res_pma_is_match_T_26 == _res_pma_is_match_T_28; // @[PMP.scala 232:14]
  wire  _res_pma_is_match_T_30 = io_check_env_pma_1_cfg_a == 2'h1; // @[PMP.scala 53:15]
  wire  _res_pma_is_match_T_35 = ~_res_pma_is_match_T_18; // @[PMP.scala 220:5]
  wire  _res_pma_is_match_T_39 = io_req_bits_addr < _res_pma_is_match_T_24; // @[PMP.scala 210:14]
  wire  _res_pma_is_match_T_40 = _res_pma_is_match_T_35 & _res_pma_is_match_T_39; // @[PMP.scala 228:56]
  wire  _res_pma_is_match_T_41 = _res_pma_is_match_T_30 & _res_pma_is_match_T_40; // @[PMP.scala 200:10]
  wire [35:0] _res_pma_is_match_T_43 = {io_check_env_pma_2_addr, 2'h0}; // @[PMP.scala 190:35]
  wire [35:0] _res_pma_is_match_T_45 = _res_pma_is_match_T_43 & 36'hffffff000; // @[PMP.scala 190:50]
  wire [35:0] _res_pma_is_match_T_46 = ~io_check_env_pma_2_mask; // @[PMP.scala 232:10]
  wire [35:0] _res_pma_is_match_T_47 = io_req_bits_addr & _res_pma_is_match_T_46; // @[PMP.scala 232:8]
  wire [35:0] _res_pma_is_match_T_49 = _res_pma_is_match_T_45 & _res_pma_is_match_T_46; // @[PMP.scala 232:21]
  wire  _res_pma_is_match_T_50 = _res_pma_is_match_T_47 == _res_pma_is_match_T_49; // @[PMP.scala 232:14]
  wire  _res_pma_is_match_T_51 = io_check_env_pma_2_cfg_a == 2'h1; // @[PMP.scala 53:15]
  wire  _res_pma_is_match_T_56 = ~_res_pma_is_match_T_39; // @[PMP.scala 220:5]
  wire  _res_pma_is_match_T_60 = io_req_bits_addr < _res_pma_is_match_T_45; // @[PMP.scala 210:14]
  wire  _res_pma_is_match_T_61 = _res_pma_is_match_T_56 & _res_pma_is_match_T_60; // @[PMP.scala 228:56]
  wire  _res_pma_is_match_T_62 = _res_pma_is_match_T_51 & _res_pma_is_match_T_61; // @[PMP.scala 200:10]
  wire [35:0] _res_pma_is_match_T_64 = {io_check_env_pma_3_addr, 2'h0}; // @[PMP.scala 190:35]
  wire [35:0] _res_pma_is_match_T_66 = _res_pma_is_match_T_64 & 36'hffffff000; // @[PMP.scala 190:50]
  wire [35:0] _res_pma_is_match_T_67 = ~io_check_env_pma_3_mask; // @[PMP.scala 232:10]
  wire [35:0] _res_pma_is_match_T_68 = io_req_bits_addr & _res_pma_is_match_T_67; // @[PMP.scala 232:8]
  wire [35:0] _res_pma_is_match_T_70 = _res_pma_is_match_T_66 & _res_pma_is_match_T_67; // @[PMP.scala 232:21]
  wire  _res_pma_is_match_T_71 = _res_pma_is_match_T_68 == _res_pma_is_match_T_70; // @[PMP.scala 232:14]
  wire  _res_pma_is_match_T_72 = io_check_env_pma_3_cfg_a == 2'h1; // @[PMP.scala 53:15]
  wire  _res_pma_is_match_T_77 = ~_res_pma_is_match_T_60; // @[PMP.scala 220:5]
  wire  _res_pma_is_match_T_81 = io_req_bits_addr < _res_pma_is_match_T_66; // @[PMP.scala 210:14]
  wire  _res_pma_is_match_T_82 = _res_pma_is_match_T_77 & _res_pma_is_match_T_81; // @[PMP.scala 228:56]
  wire  _res_pma_is_match_T_83 = _res_pma_is_match_T_72 & _res_pma_is_match_T_82; // @[PMP.scala 200:10]
  wire [35:0] _res_pma_is_match_T_85 = {io_check_env_pma_4_addr, 2'h0}; // @[PMP.scala 190:35]
  wire [35:0] _res_pma_is_match_T_87 = _res_pma_is_match_T_85 & 36'hffffff000; // @[PMP.scala 190:50]
  wire [35:0] _res_pma_is_match_T_88 = ~io_check_env_pma_4_mask; // @[PMP.scala 232:10]
  wire [35:0] _res_pma_is_match_T_89 = io_req_bits_addr & _res_pma_is_match_T_88; // @[PMP.scala 232:8]
  wire [35:0] _res_pma_is_match_T_91 = _res_pma_is_match_T_87 & _res_pma_is_match_T_88; // @[PMP.scala 232:21]
  wire  _res_pma_is_match_T_92 = _res_pma_is_match_T_89 == _res_pma_is_match_T_91; // @[PMP.scala 232:14]
  wire  _res_pma_is_match_T_93 = io_check_env_pma_4_cfg_a == 2'h1; // @[PMP.scala 53:15]
  wire  _res_pma_is_match_T_98 = ~_res_pma_is_match_T_81; // @[PMP.scala 220:5]
  wire  _res_pma_is_match_T_102 = io_req_bits_addr < _res_pma_is_match_T_87; // @[PMP.scala 210:14]
  wire  _res_pma_is_match_T_103 = _res_pma_is_match_T_98 & _res_pma_is_match_T_102; // @[PMP.scala 228:56]
  wire  _res_pma_is_match_T_104 = _res_pma_is_match_T_93 & _res_pma_is_match_T_103; // @[PMP.scala 200:10]
  wire [35:0] _res_pma_is_match_T_106 = {io_check_env_pma_5_addr, 2'h0}; // @[PMP.scala 190:35]
  wire [35:0] _res_pma_is_match_T_108 = _res_pma_is_match_T_106 & 36'hffffff000; // @[PMP.scala 190:50]
  wire [35:0] _res_pma_is_match_T_109 = ~io_check_env_pma_5_mask; // @[PMP.scala 232:10]
  wire [35:0] _res_pma_is_match_T_110 = io_req_bits_addr & _res_pma_is_match_T_109; // @[PMP.scala 232:8]
  wire [35:0] _res_pma_is_match_T_112 = _res_pma_is_match_T_108 & _res_pma_is_match_T_109; // @[PMP.scala 232:21]
  wire  _res_pma_is_match_T_113 = _res_pma_is_match_T_110 == _res_pma_is_match_T_112; // @[PMP.scala 232:14]
  wire  _res_pma_is_match_T_114 = io_check_env_pma_5_cfg_a == 2'h1; // @[PMP.scala 53:15]
  wire  _res_pma_is_match_T_119 = ~_res_pma_is_match_T_102; // @[PMP.scala 220:5]
  wire  _res_pma_is_match_T_123 = io_req_bits_addr < _res_pma_is_match_T_108; // @[PMP.scala 210:14]
  wire  _res_pma_is_match_T_124 = _res_pma_is_match_T_119 & _res_pma_is_match_T_123; // @[PMP.scala 228:56]
  wire  _res_pma_is_match_T_125 = _res_pma_is_match_T_114 & _res_pma_is_match_T_124; // @[PMP.scala 200:10]
  wire [35:0] _res_pma_is_match_T_127 = {io_check_env_pma_6_addr, 2'h0}; // @[PMP.scala 190:35]
  wire [35:0] _res_pma_is_match_T_129 = _res_pma_is_match_T_127 & 36'hffffff000; // @[PMP.scala 190:50]
  wire [35:0] _res_pma_is_match_T_130 = ~io_check_env_pma_6_mask; // @[PMP.scala 232:10]
  wire [35:0] _res_pma_is_match_T_131 = io_req_bits_addr & _res_pma_is_match_T_130; // @[PMP.scala 232:8]
  wire [35:0] _res_pma_is_match_T_133 = _res_pma_is_match_T_129 & _res_pma_is_match_T_130; // @[PMP.scala 232:21]
  wire  _res_pma_is_match_T_134 = _res_pma_is_match_T_131 == _res_pma_is_match_T_133; // @[PMP.scala 232:14]
  wire  _res_pma_is_match_T_135 = io_check_env_pma_6_cfg_a == 2'h1; // @[PMP.scala 53:15]
  wire  _res_pma_is_match_T_140 = ~_res_pma_is_match_T_123; // @[PMP.scala 220:5]
  wire  _res_pma_is_match_T_144 = io_req_bits_addr < _res_pma_is_match_T_129; // @[PMP.scala 210:14]
  wire  _res_pma_is_match_T_145 = _res_pma_is_match_T_140 & _res_pma_is_match_T_144; // @[PMP.scala 228:56]
  wire  _res_pma_is_match_T_146 = _res_pma_is_match_T_135 & _res_pma_is_match_T_145; // @[PMP.scala 200:10]
  wire [35:0] _res_pma_is_match_T_148 = {io_check_env_pma_7_addr, 2'h0}; // @[PMP.scala 190:35]
  wire [35:0] _res_pma_is_match_T_150 = _res_pma_is_match_T_148 & 36'hffffff000; // @[PMP.scala 190:50]
  wire [35:0] _res_pma_is_match_T_151 = ~io_check_env_pma_7_mask; // @[PMP.scala 232:10]
  wire [35:0] _res_pma_is_match_T_152 = io_req_bits_addr & _res_pma_is_match_T_151; // @[PMP.scala 232:8]
  wire [35:0] _res_pma_is_match_T_154 = _res_pma_is_match_T_150 & _res_pma_is_match_T_151; // @[PMP.scala 232:21]
  wire  _res_pma_is_match_T_155 = _res_pma_is_match_T_152 == _res_pma_is_match_T_154; // @[PMP.scala 232:14]
  wire  _res_pma_is_match_T_156 = io_check_env_pma_7_cfg_a == 2'h1; // @[PMP.scala 53:15]
  wire  _res_pma_is_match_T_161 = ~_res_pma_is_match_T_144; // @[PMP.scala 220:5]
  wire  _res_pma_is_match_T_165 = io_req_bits_addr < _res_pma_is_match_T_150; // @[PMP.scala 210:14]
  wire  _res_pma_is_match_T_166 = _res_pma_is_match_T_161 & _res_pma_is_match_T_165; // @[PMP.scala 228:56]
  wire  _res_pma_is_match_T_167 = _res_pma_is_match_T_156 & _res_pma_is_match_T_166; // @[PMP.scala 200:10]
  wire [35:0] _res_pma_is_match_T_169 = {io_check_env_pma_8_addr, 2'h0}; // @[PMP.scala 190:35]
  wire [35:0] _res_pma_is_match_T_171 = _res_pma_is_match_T_169 & 36'hffffff000; // @[PMP.scala 190:50]
  wire [35:0] _res_pma_is_match_T_172 = ~io_check_env_pma_8_mask; // @[PMP.scala 232:10]
  wire [35:0] _res_pma_is_match_T_173 = io_req_bits_addr & _res_pma_is_match_T_172; // @[PMP.scala 232:8]
  wire [35:0] _res_pma_is_match_T_175 = _res_pma_is_match_T_171 & _res_pma_is_match_T_172; // @[PMP.scala 232:21]
  wire  _res_pma_is_match_T_176 = _res_pma_is_match_T_173 == _res_pma_is_match_T_175; // @[PMP.scala 232:14]
  wire  _res_pma_is_match_T_177 = io_check_env_pma_8_cfg_a == 2'h1; // @[PMP.scala 53:15]
  wire  _res_pma_is_match_T_182 = ~_res_pma_is_match_T_165; // @[PMP.scala 220:5]
  wire  _res_pma_is_match_T_186 = io_req_bits_addr < _res_pma_is_match_T_171; // @[PMP.scala 210:14]
  wire  _res_pma_is_match_T_187 = _res_pma_is_match_T_182 & _res_pma_is_match_T_186; // @[PMP.scala 228:56]
  wire  _res_pma_is_match_T_188 = _res_pma_is_match_T_177 & _res_pma_is_match_T_187; // @[PMP.scala 200:10]
  wire [35:0] _res_pma_is_match_T_190 = {io_check_env_pma_9_addr, 2'h0}; // @[PMP.scala 190:35]
  wire [35:0] _res_pma_is_match_T_192 = _res_pma_is_match_T_190 & 36'hffffff000; // @[PMP.scala 190:50]
  wire [35:0] _res_pma_is_match_T_193 = ~io_check_env_pma_9_mask; // @[PMP.scala 232:10]
  wire [35:0] _res_pma_is_match_T_194 = io_req_bits_addr & _res_pma_is_match_T_193; // @[PMP.scala 232:8]
  wire [35:0] _res_pma_is_match_T_196 = _res_pma_is_match_T_192 & _res_pma_is_match_T_193; // @[PMP.scala 232:21]
  wire  _res_pma_is_match_T_197 = _res_pma_is_match_T_194 == _res_pma_is_match_T_196; // @[PMP.scala 232:14]
  wire  _res_pma_is_match_T_198 = io_check_env_pma_9_cfg_a == 2'h1; // @[PMP.scala 53:15]
  wire  _res_pma_is_match_T_203 = ~_res_pma_is_match_T_186; // @[PMP.scala 220:5]
  wire  _res_pma_is_match_T_207 = io_req_bits_addr < _res_pma_is_match_T_192; // @[PMP.scala 210:14]
  wire  _res_pma_is_match_T_208 = _res_pma_is_match_T_203 & _res_pma_is_match_T_207; // @[PMP.scala 228:56]
  wire  _res_pma_is_match_T_209 = _res_pma_is_match_T_198 & _res_pma_is_match_T_208; // @[PMP.scala 200:10]
  wire [35:0] _res_pma_is_match_T_211 = {io_check_env_pma_10_addr, 2'h0}; // @[PMP.scala 190:35]
  wire [35:0] _res_pma_is_match_T_213 = _res_pma_is_match_T_211 & 36'hffffff000; // @[PMP.scala 190:50]
  wire [35:0] _res_pma_is_match_T_214 = ~io_check_env_pma_10_mask; // @[PMP.scala 232:10]
  wire [35:0] _res_pma_is_match_T_215 = io_req_bits_addr & _res_pma_is_match_T_214; // @[PMP.scala 232:8]
  wire [35:0] _res_pma_is_match_T_217 = _res_pma_is_match_T_213 & _res_pma_is_match_T_214; // @[PMP.scala 232:21]
  wire  _res_pma_is_match_T_218 = _res_pma_is_match_T_215 == _res_pma_is_match_T_217; // @[PMP.scala 232:14]
  wire  _res_pma_is_match_T_219 = io_check_env_pma_10_cfg_a == 2'h1; // @[PMP.scala 53:15]
  wire  _res_pma_is_match_T_224 = ~_res_pma_is_match_T_207; // @[PMP.scala 220:5]
  wire  _res_pma_is_match_T_228 = io_req_bits_addr < _res_pma_is_match_T_213; // @[PMP.scala 210:14]
  wire  _res_pma_is_match_T_229 = _res_pma_is_match_T_224 & _res_pma_is_match_T_228; // @[PMP.scala 228:56]
  wire  _res_pma_is_match_T_230 = _res_pma_is_match_T_219 & _res_pma_is_match_T_229; // @[PMP.scala 200:10]
  wire [35:0] _res_pma_is_match_T_232 = {io_check_env_pma_11_addr, 2'h0}; // @[PMP.scala 190:35]
  wire [35:0] _res_pma_is_match_T_234 = _res_pma_is_match_T_232 & 36'hffffff000; // @[PMP.scala 190:50]
  wire [35:0] _res_pma_is_match_T_235 = ~io_check_env_pma_11_mask; // @[PMP.scala 232:10]
  wire [35:0] _res_pma_is_match_T_236 = io_req_bits_addr & _res_pma_is_match_T_235; // @[PMP.scala 232:8]
  wire [35:0] _res_pma_is_match_T_238 = _res_pma_is_match_T_234 & _res_pma_is_match_T_235; // @[PMP.scala 232:21]
  wire  _res_pma_is_match_T_239 = _res_pma_is_match_T_236 == _res_pma_is_match_T_238; // @[PMP.scala 232:14]
  wire  _res_pma_is_match_T_240 = io_check_env_pma_11_cfg_a == 2'h1; // @[PMP.scala 53:15]
  wire  _res_pma_is_match_T_245 = ~_res_pma_is_match_T_228; // @[PMP.scala 220:5]
  wire  _res_pma_is_match_T_249 = io_req_bits_addr < _res_pma_is_match_T_234; // @[PMP.scala 210:14]
  wire  _res_pma_is_match_T_250 = _res_pma_is_match_T_245 & _res_pma_is_match_T_249; // @[PMP.scala 228:56]
  wire  _res_pma_is_match_T_251 = _res_pma_is_match_T_240 & _res_pma_is_match_T_250; // @[PMP.scala 200:10]
  wire [35:0] _res_pma_is_match_T_253 = {io_check_env_pma_12_addr, 2'h0}; // @[PMP.scala 190:35]
  wire [35:0] _res_pma_is_match_T_255 = _res_pma_is_match_T_253 & 36'hffffff000; // @[PMP.scala 190:50]
  wire [35:0] _res_pma_is_match_T_256 = ~io_check_env_pma_12_mask; // @[PMP.scala 232:10]
  wire [35:0] _res_pma_is_match_T_257 = io_req_bits_addr & _res_pma_is_match_T_256; // @[PMP.scala 232:8]
  wire [35:0] _res_pma_is_match_T_259 = _res_pma_is_match_T_255 & _res_pma_is_match_T_256; // @[PMP.scala 232:21]
  wire  _res_pma_is_match_T_260 = _res_pma_is_match_T_257 == _res_pma_is_match_T_259; // @[PMP.scala 232:14]
  wire  _res_pma_is_match_T_261 = io_check_env_pma_12_cfg_a == 2'h1; // @[PMP.scala 53:15]
  wire  _res_pma_is_match_T_266 = ~_res_pma_is_match_T_249; // @[PMP.scala 220:5]
  wire  _res_pma_is_match_T_270 = io_req_bits_addr < _res_pma_is_match_T_255; // @[PMP.scala 210:14]
  wire  _res_pma_is_match_T_271 = _res_pma_is_match_T_266 & _res_pma_is_match_T_270; // @[PMP.scala 228:56]
  wire  _res_pma_is_match_T_272 = _res_pma_is_match_T_261 & _res_pma_is_match_T_271; // @[PMP.scala 200:10]
  wire [35:0] _res_pma_is_match_T_274 = {io_check_env_pma_13_addr, 2'h0}; // @[PMP.scala 190:35]
  wire [35:0] _res_pma_is_match_T_276 = _res_pma_is_match_T_274 & 36'hffffff000; // @[PMP.scala 190:50]
  wire [35:0] _res_pma_is_match_T_277 = ~io_check_env_pma_13_mask; // @[PMP.scala 232:10]
  wire [35:0] _res_pma_is_match_T_278 = io_req_bits_addr & _res_pma_is_match_T_277; // @[PMP.scala 232:8]
  wire [35:0] _res_pma_is_match_T_280 = _res_pma_is_match_T_276 & _res_pma_is_match_T_277; // @[PMP.scala 232:21]
  wire  _res_pma_is_match_T_281 = _res_pma_is_match_T_278 == _res_pma_is_match_T_280; // @[PMP.scala 232:14]
  wire  _res_pma_is_match_T_282 = io_check_env_pma_13_cfg_a == 2'h1; // @[PMP.scala 53:15]
  wire  _res_pma_is_match_T_287 = ~_res_pma_is_match_T_270; // @[PMP.scala 220:5]
  wire  _res_pma_is_match_T_291 = io_req_bits_addr < _res_pma_is_match_T_276; // @[PMP.scala 210:14]
  wire  _res_pma_is_match_T_292 = _res_pma_is_match_T_287 & _res_pma_is_match_T_291; // @[PMP.scala 228:56]
  wire  _res_pma_is_match_T_293 = _res_pma_is_match_T_282 & _res_pma_is_match_T_292; // @[PMP.scala 200:10]
  wire [35:0] _res_pma_is_match_T_295 = {io_check_env_pma_14_addr, 2'h0}; // @[PMP.scala 190:35]
  wire [35:0] _res_pma_is_match_T_297 = _res_pma_is_match_T_295 & 36'hffffff000; // @[PMP.scala 190:50]
  wire [35:0] _res_pma_is_match_T_298 = ~io_check_env_pma_14_mask; // @[PMP.scala 232:10]
  wire [35:0] _res_pma_is_match_T_299 = io_req_bits_addr & _res_pma_is_match_T_298; // @[PMP.scala 232:8]
  wire [35:0] _res_pma_is_match_T_301 = _res_pma_is_match_T_297 & _res_pma_is_match_T_298; // @[PMP.scala 232:21]
  wire  _res_pma_is_match_T_302 = _res_pma_is_match_T_299 == _res_pma_is_match_T_301; // @[PMP.scala 232:14]
  wire  _res_pma_is_match_T_303 = io_check_env_pma_14_cfg_a == 2'h1; // @[PMP.scala 53:15]
  wire  _res_pma_is_match_T_308 = ~_res_pma_is_match_T_291; // @[PMP.scala 220:5]
  wire  _res_pma_is_match_T_312 = io_req_bits_addr < _res_pma_is_match_T_297; // @[PMP.scala 210:14]
  wire  _res_pma_is_match_T_313 = _res_pma_is_match_T_308 & _res_pma_is_match_T_312; // @[PMP.scala 228:56]
  wire  _res_pma_is_match_T_314 = _res_pma_is_match_T_303 & _res_pma_is_match_T_313; // @[PMP.scala 200:10]
  wire [35:0] _res_pma_is_match_T_316 = {io_check_env_pma_15_addr, 2'h0}; // @[PMP.scala 190:35]
  wire [35:0] _res_pma_is_match_T_318 = _res_pma_is_match_T_316 & 36'hffffff000; // @[PMP.scala 190:50]
  wire [35:0] _res_pma_is_match_T_319 = ~io_check_env_pma_15_mask; // @[PMP.scala 232:10]
  wire [35:0] _res_pma_is_match_T_320 = io_req_bits_addr & _res_pma_is_match_T_319; // @[PMP.scala 232:8]
  wire [35:0] _res_pma_is_match_T_322 = _res_pma_is_match_T_318 & _res_pma_is_match_T_319; // @[PMP.scala 232:21]
  wire  _res_pma_is_match_T_323 = _res_pma_is_match_T_320 == _res_pma_is_match_T_322; // @[PMP.scala 232:14]
  wire  _res_pma_is_match_T_324 = io_check_env_pma_15_cfg_a == 2'h1; // @[PMP.scala 53:15]
  wire  _res_pma_is_match_T_329 = ~_res_pma_is_match_T_312; // @[PMP.scala 220:5]
  wire  _res_pma_is_match_T_333 = io_req_bits_addr < _res_pma_is_match_T_318; // @[PMP.scala 210:14]
  wire  _res_pma_is_match_T_334 = _res_pma_is_match_T_329 & _res_pma_is_match_T_333; // @[PMP.scala 228:56]
  wire  _res_pma_is_match_T_335 = _res_pma_is_match_T_324 & _res_pma_is_match_T_334; // @[PMP.scala 200:10]
  reg  res_pma_r; // @[Reg.scala 28:20]
  reg  res_pma_r1; // @[Reg.scala 28:20]
  reg  res_pma_r2; // @[Reg.scala 28:20]
  reg  res_pma_r3; // @[Reg.scala 28:20]
  reg  res_pma_r4; // @[Reg.scala 28:20]
  reg  res_pma_r5; // @[Reg.scala 28:20]
  reg  res_pma_r6; // @[Reg.scala 28:20]
  reg  res_pma_r7; // @[Reg.scala 28:20]
  reg  res_pma_r8; // @[Reg.scala 28:20]
  reg  res_pma_r9; // @[Reg.scala 28:20]
  reg  res_pma_r10; // @[Reg.scala 28:20]
  reg  res_pma_r11; // @[Reg.scala 28:20]
  reg  res_pma_r12; // @[Reg.scala 28:20]
  reg  res_pma_r13; // @[Reg.scala 28:20]
  reg  res_pma_r14; // @[Reg.scala 28:20]
  reg  res_pma_r15; // @[Reg.scala 28:20]
  reg  res_pma_r17_0_cfg_c; // @[Reg.scala 16:16]
  reg  res_pma_r17_0_cfg_atomic; // @[Reg.scala 16:16]
  reg  res_pma_r17_0_cfg_x; // @[Reg.scala 16:16]
  reg  res_pma_r17_0_cfg_w; // @[Reg.scala 16:16]
  reg  res_pma_r17_0_cfg_r; // @[Reg.scala 16:16]
  reg  res_pma_r17_1_cfg_c; // @[Reg.scala 16:16]
  reg  res_pma_r17_1_cfg_atomic; // @[Reg.scala 16:16]
  reg  res_pma_r17_1_cfg_x; // @[Reg.scala 16:16]
  reg  res_pma_r17_1_cfg_w; // @[Reg.scala 16:16]
  reg  res_pma_r17_1_cfg_r; // @[Reg.scala 16:16]
  reg  res_pma_r17_2_cfg_c; // @[Reg.scala 16:16]
  reg  res_pma_r17_2_cfg_atomic; // @[Reg.scala 16:16]
  reg  res_pma_r17_2_cfg_x; // @[Reg.scala 16:16]
  reg  res_pma_r17_2_cfg_w; // @[Reg.scala 16:16]
  reg  res_pma_r17_2_cfg_r; // @[Reg.scala 16:16]
  reg  res_pma_r17_3_cfg_c; // @[Reg.scala 16:16]
  reg  res_pma_r17_3_cfg_atomic; // @[Reg.scala 16:16]
  reg  res_pma_r17_3_cfg_x; // @[Reg.scala 16:16]
  reg  res_pma_r17_3_cfg_w; // @[Reg.scala 16:16]
  reg  res_pma_r17_3_cfg_r; // @[Reg.scala 16:16]
  reg  res_pma_r17_4_cfg_c; // @[Reg.scala 16:16]
  reg  res_pma_r17_4_cfg_atomic; // @[Reg.scala 16:16]
  reg  res_pma_r17_4_cfg_x; // @[Reg.scala 16:16]
  reg  res_pma_r17_4_cfg_w; // @[Reg.scala 16:16]
  reg  res_pma_r17_4_cfg_r; // @[Reg.scala 16:16]
  reg  res_pma_r17_5_cfg_c; // @[Reg.scala 16:16]
  reg  res_pma_r17_5_cfg_atomic; // @[Reg.scala 16:16]
  reg  res_pma_r17_5_cfg_x; // @[Reg.scala 16:16]
  reg  res_pma_r17_5_cfg_w; // @[Reg.scala 16:16]
  reg  res_pma_r17_5_cfg_r; // @[Reg.scala 16:16]
  reg  res_pma_r17_6_cfg_c; // @[Reg.scala 16:16]
  reg  res_pma_r17_6_cfg_atomic; // @[Reg.scala 16:16]
  reg  res_pma_r17_6_cfg_x; // @[Reg.scala 16:16]
  reg  res_pma_r17_6_cfg_w; // @[Reg.scala 16:16]
  reg  res_pma_r17_6_cfg_r; // @[Reg.scala 16:16]
  reg  res_pma_r17_7_cfg_c; // @[Reg.scala 16:16]
  reg  res_pma_r17_7_cfg_atomic; // @[Reg.scala 16:16]
  reg  res_pma_r17_7_cfg_x; // @[Reg.scala 16:16]
  reg  res_pma_r17_7_cfg_w; // @[Reg.scala 16:16]
  reg  res_pma_r17_7_cfg_r; // @[Reg.scala 16:16]
  reg  res_pma_r17_8_cfg_c; // @[Reg.scala 16:16]
  reg  res_pma_r17_8_cfg_atomic; // @[Reg.scala 16:16]
  reg  res_pma_r17_8_cfg_x; // @[Reg.scala 16:16]
  reg  res_pma_r17_8_cfg_w; // @[Reg.scala 16:16]
  reg  res_pma_r17_8_cfg_r; // @[Reg.scala 16:16]
  reg  res_pma_r17_9_cfg_c; // @[Reg.scala 16:16]
  reg  res_pma_r17_9_cfg_atomic; // @[Reg.scala 16:16]
  reg  res_pma_r17_9_cfg_x; // @[Reg.scala 16:16]
  reg  res_pma_r17_9_cfg_w; // @[Reg.scala 16:16]
  reg  res_pma_r17_9_cfg_r; // @[Reg.scala 16:16]
  reg  res_pma_r17_10_cfg_c; // @[Reg.scala 16:16]
  reg  res_pma_r17_10_cfg_atomic; // @[Reg.scala 16:16]
  reg  res_pma_r17_10_cfg_x; // @[Reg.scala 16:16]
  reg  res_pma_r17_10_cfg_w; // @[Reg.scala 16:16]
  reg  res_pma_r17_10_cfg_r; // @[Reg.scala 16:16]
  reg  res_pma_r17_11_cfg_c; // @[Reg.scala 16:16]
  reg  res_pma_r17_11_cfg_atomic; // @[Reg.scala 16:16]
  reg  res_pma_r17_11_cfg_x; // @[Reg.scala 16:16]
  reg  res_pma_r17_11_cfg_w; // @[Reg.scala 16:16]
  reg  res_pma_r17_11_cfg_r; // @[Reg.scala 16:16]
  reg  res_pma_r17_12_cfg_c; // @[Reg.scala 16:16]
  reg  res_pma_r17_12_cfg_atomic; // @[Reg.scala 16:16]
  reg  res_pma_r17_12_cfg_x; // @[Reg.scala 16:16]
  reg  res_pma_r17_12_cfg_w; // @[Reg.scala 16:16]
  reg  res_pma_r17_12_cfg_r; // @[Reg.scala 16:16]
  reg  res_pma_r17_13_cfg_c; // @[Reg.scala 16:16]
  reg  res_pma_r17_13_cfg_atomic; // @[Reg.scala 16:16]
  reg  res_pma_r17_13_cfg_x; // @[Reg.scala 16:16]
  reg  res_pma_r17_13_cfg_w; // @[Reg.scala 16:16]
  reg  res_pma_r17_13_cfg_r; // @[Reg.scala 16:16]
  reg  res_pma_r17_14_cfg_c; // @[Reg.scala 16:16]
  reg  res_pma_r17_14_cfg_atomic; // @[Reg.scala 16:16]
  reg  res_pma_r17_14_cfg_x; // @[Reg.scala 16:16]
  reg  res_pma_r17_14_cfg_w; // @[Reg.scala 16:16]
  reg  res_pma_r17_14_cfg_r; // @[Reg.scala 16:16]
  reg  res_pma_r17_15_cfg_c; // @[Reg.scala 16:16]
  reg  res_pma_r17_15_cfg_atomic; // @[Reg.scala 16:16]
  reg  res_pma_r17_15_cfg_x; // @[Reg.scala 16:16]
  reg  res_pma_r17_15_cfg_w; // @[Reg.scala 16:16]
  reg  res_pma_r17_15_cfg_r; // @[Reg.scala 16:16]
  wire  _res_pma_T_1_cfg_c = res_pma_r ? res_pma_r17_0_cfg_c : res_pma_r17_1_cfg_c; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_1_cfg_atomic = res_pma_r ? res_pma_r17_0_cfg_atomic : res_pma_r17_1_cfg_atomic; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_1_cfg_x = res_pma_r ? res_pma_r17_0_cfg_x : res_pma_r17_1_cfg_x; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_1_cfg_w = res_pma_r ? res_pma_r17_0_cfg_w : res_pma_r17_1_cfg_w; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_1_cfg_r = res_pma_r ? res_pma_r17_0_cfg_r : res_pma_r17_1_cfg_r; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_3_cfg_c = res_pma_r2 ? res_pma_r17_2_cfg_c : res_pma_r17_3_cfg_c; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_3_cfg_atomic = res_pma_r2 ? res_pma_r17_2_cfg_atomic : res_pma_r17_3_cfg_atomic; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_3_cfg_x = res_pma_r2 ? res_pma_r17_2_cfg_x : res_pma_r17_3_cfg_x; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_3_cfg_w = res_pma_r2 ? res_pma_r17_2_cfg_w : res_pma_r17_3_cfg_w; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_3_cfg_r = res_pma_r2 ? res_pma_r17_2_cfg_r : res_pma_r17_3_cfg_r; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_5_cfg_c = res_pma_r | res_pma_r1 ? _res_pma_T_1_cfg_c : _res_pma_T_3_cfg_c; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_5_cfg_atomic = res_pma_r | res_pma_r1 ? _res_pma_T_1_cfg_atomic : _res_pma_T_3_cfg_atomic; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_5_cfg_x = res_pma_r | res_pma_r1 ? _res_pma_T_1_cfg_x : _res_pma_T_3_cfg_x; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_5_cfg_w = res_pma_r | res_pma_r1 ? _res_pma_T_1_cfg_w : _res_pma_T_3_cfg_w; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_5_cfg_r = res_pma_r | res_pma_r1 ? _res_pma_T_1_cfg_r : _res_pma_T_3_cfg_r; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_7_cfg_c = res_pma_r4 ? res_pma_r17_4_cfg_c : res_pma_r17_5_cfg_c; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_7_cfg_atomic = res_pma_r4 ? res_pma_r17_4_cfg_atomic : res_pma_r17_5_cfg_atomic; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_7_cfg_x = res_pma_r4 ? res_pma_r17_4_cfg_x : res_pma_r17_5_cfg_x; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_7_cfg_w = res_pma_r4 ? res_pma_r17_4_cfg_w : res_pma_r17_5_cfg_w; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_7_cfg_r = res_pma_r4 ? res_pma_r17_4_cfg_r : res_pma_r17_5_cfg_r; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_9_cfg_c = res_pma_r6 ? res_pma_r17_6_cfg_c : res_pma_r17_7_cfg_c; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_9_cfg_atomic = res_pma_r6 ? res_pma_r17_6_cfg_atomic : res_pma_r17_7_cfg_atomic; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_9_cfg_x = res_pma_r6 ? res_pma_r17_6_cfg_x : res_pma_r17_7_cfg_x; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_9_cfg_w = res_pma_r6 ? res_pma_r17_6_cfg_w : res_pma_r17_7_cfg_w; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_9_cfg_r = res_pma_r6 ? res_pma_r17_6_cfg_r : res_pma_r17_7_cfg_r; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_11_cfg_c = res_pma_r4 | res_pma_r5 ? _res_pma_T_7_cfg_c : _res_pma_T_9_cfg_c; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_11_cfg_atomic = res_pma_r4 | res_pma_r5 ? _res_pma_T_7_cfg_atomic : _res_pma_T_9_cfg_atomic; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_11_cfg_x = res_pma_r4 | res_pma_r5 ? _res_pma_T_7_cfg_x : _res_pma_T_9_cfg_x; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_11_cfg_w = res_pma_r4 | res_pma_r5 ? _res_pma_T_7_cfg_w : _res_pma_T_9_cfg_w; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_11_cfg_r = res_pma_r4 | res_pma_r5 ? _res_pma_T_7_cfg_r : _res_pma_T_9_cfg_r; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_13_cfg_c = res_pma_r | res_pma_r1 | (res_pma_r2 | res_pma_r3) ? _res_pma_T_5_cfg_c :
    _res_pma_T_11_cfg_c; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_13_cfg_atomic = res_pma_r | res_pma_r1 | (res_pma_r2 | res_pma_r3) ? _res_pma_T_5_cfg_atomic :
    _res_pma_T_11_cfg_atomic; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_13_cfg_x = res_pma_r | res_pma_r1 | (res_pma_r2 | res_pma_r3) ? _res_pma_T_5_cfg_x :
    _res_pma_T_11_cfg_x; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_13_cfg_w = res_pma_r | res_pma_r1 | (res_pma_r2 | res_pma_r3) ? _res_pma_T_5_cfg_w :
    _res_pma_T_11_cfg_w; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_13_cfg_r = res_pma_r | res_pma_r1 | (res_pma_r2 | res_pma_r3) ? _res_pma_T_5_cfg_r :
    _res_pma_T_11_cfg_r; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_15_cfg_c = res_pma_r8 ? res_pma_r17_8_cfg_c : res_pma_r17_9_cfg_c; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_15_cfg_atomic = res_pma_r8 ? res_pma_r17_8_cfg_atomic : res_pma_r17_9_cfg_atomic; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_15_cfg_x = res_pma_r8 ? res_pma_r17_8_cfg_x : res_pma_r17_9_cfg_x; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_15_cfg_w = res_pma_r8 ? res_pma_r17_8_cfg_w : res_pma_r17_9_cfg_w; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_15_cfg_r = res_pma_r8 ? res_pma_r17_8_cfg_r : res_pma_r17_9_cfg_r; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_17_cfg_c = res_pma_r10 ? res_pma_r17_10_cfg_c : res_pma_r17_11_cfg_c; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_17_cfg_atomic = res_pma_r10 ? res_pma_r17_10_cfg_atomic : res_pma_r17_11_cfg_atomic; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_17_cfg_x = res_pma_r10 ? res_pma_r17_10_cfg_x : res_pma_r17_11_cfg_x; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_17_cfg_w = res_pma_r10 ? res_pma_r17_10_cfg_w : res_pma_r17_11_cfg_w; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_17_cfg_r = res_pma_r10 ? res_pma_r17_10_cfg_r : res_pma_r17_11_cfg_r; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_19_cfg_c = res_pma_r8 | res_pma_r9 ? _res_pma_T_15_cfg_c : _res_pma_T_17_cfg_c; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_19_cfg_atomic = res_pma_r8 | res_pma_r9 ? _res_pma_T_15_cfg_atomic : _res_pma_T_17_cfg_atomic; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_19_cfg_x = res_pma_r8 | res_pma_r9 ? _res_pma_T_15_cfg_x : _res_pma_T_17_cfg_x; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_19_cfg_w = res_pma_r8 | res_pma_r9 ? _res_pma_T_15_cfg_w : _res_pma_T_17_cfg_w; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_19_cfg_r = res_pma_r8 | res_pma_r9 ? _res_pma_T_15_cfg_r : _res_pma_T_17_cfg_r; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_21_cfg_c = res_pma_r12 ? res_pma_r17_12_cfg_c : res_pma_r17_13_cfg_c; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_21_cfg_atomic = res_pma_r12 ? res_pma_r17_12_cfg_atomic : res_pma_r17_13_cfg_atomic; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_21_cfg_x = res_pma_r12 ? res_pma_r17_12_cfg_x : res_pma_r17_13_cfg_x; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_21_cfg_w = res_pma_r12 ? res_pma_r17_12_cfg_w : res_pma_r17_13_cfg_w; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_21_cfg_r = res_pma_r12 ? res_pma_r17_12_cfg_r : res_pma_r17_13_cfg_r; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_25_cfg_c = res_pma_r14 ? res_pma_r17_14_cfg_c : res_pma_r15 & res_pma_r17_15_cfg_c; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_25_cfg_atomic = res_pma_r14 ? res_pma_r17_14_cfg_atomic : res_pma_r15 & res_pma_r17_15_cfg_atomic
    ; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_25_cfg_x = res_pma_r14 ? res_pma_r17_14_cfg_x : res_pma_r15 & res_pma_r17_15_cfg_x; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_25_cfg_w = res_pma_r14 ? res_pma_r17_14_cfg_w : res_pma_r15 & res_pma_r17_15_cfg_w; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_25_cfg_r = res_pma_r14 ? res_pma_r17_14_cfg_r : res_pma_r15 & res_pma_r17_15_cfg_r; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_27_cfg_c = res_pma_r12 | res_pma_r13 ? _res_pma_T_21_cfg_c : _res_pma_T_25_cfg_c; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_27_cfg_atomic = res_pma_r12 | res_pma_r13 ? _res_pma_T_21_cfg_atomic : _res_pma_T_25_cfg_atomic; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_27_cfg_x = res_pma_r12 | res_pma_r13 ? _res_pma_T_21_cfg_x : _res_pma_T_25_cfg_x; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_27_cfg_w = res_pma_r12 | res_pma_r13 ? _res_pma_T_21_cfg_w : _res_pma_T_25_cfg_w; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_27_cfg_r = res_pma_r12 | res_pma_r13 ? _res_pma_T_21_cfg_r : _res_pma_T_25_cfg_r; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_29_cfg_c = res_pma_r8 | res_pma_r9 | (res_pma_r10 | res_pma_r11) ? _res_pma_T_19_cfg_c :
    _res_pma_T_27_cfg_c; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_29_cfg_atomic = res_pma_r8 | res_pma_r9 | (res_pma_r10 | res_pma_r11) ? _res_pma_T_19_cfg_atomic
     : _res_pma_T_27_cfg_atomic; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_29_cfg_x = res_pma_r8 | res_pma_r9 | (res_pma_r10 | res_pma_r11) ? _res_pma_T_19_cfg_x :
    _res_pma_T_27_cfg_x; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_29_cfg_w = res_pma_r8 | res_pma_r9 | (res_pma_r10 | res_pma_r11) ? _res_pma_T_19_cfg_w :
    _res_pma_T_27_cfg_w; // @[ParallelMux.scala 90:77]
  wire  _res_pma_T_29_cfg_r = res_pma_r8 | res_pma_r9 | (res_pma_r10 | res_pma_r11) ? _res_pma_T_19_cfg_r :
    _res_pma_T_27_cfg_r; // @[ParallelMux.scala 90:77]
  wire  res_pma_cfg_x = res_pma_r | res_pma_r1 | (res_pma_r2 | res_pma_r3) | (res_pma_r4 | res_pma_r5 | (
    res_pma_r6 | res_pma_r7)) ? _res_pma_T_13_cfg_x : _res_pma_T_29_cfg_x; // @[ParallelMux.scala 90:77]
  wire  res_pma_cfg_w = res_pma_r | res_pma_r1 | (res_pma_r2 | res_pma_r3) | (res_pma_r4 | res_pma_r5 | (
    res_pma_r6 | res_pma_r7)) ? _res_pma_T_13_cfg_w : _res_pma_T_29_cfg_w; // @[ParallelMux.scala 90:77]
  wire  res_pma_cfg_r = res_pma_r | res_pma_r1 | (res_pma_r2 | res_pma_r3) | (res_pma_r4 | res_pma_r5 | (
    res_pma_r6 | res_pma_r7)) ? _res_pma_T_13_cfg_r : _res_pma_T_29_cfg_r; // @[ParallelMux.scala 90:77]
  assign io_resp_c = res_pma_r | res_pma_r1 | (res_pma_r2 | res_pma_r3) | (res_pma_r4 | res_pma_r5 | (res_pma_r6
     | res_pma_r7)) ? _res_pma_T_13_cfg_c : _res_pma_T_29_cfg_c; // @[ParallelMux.scala 90:77]
  assign io_resp_atomic = res_pma_r | res_pma_r1 | (res_pma_r2 | res_pma_r3) | (res_pma_r4 | res_pma_r5 | (
    res_pma_r6 | res_pma_r7)) ? _res_pma_T_13_cfg_atomic : _res_pma_T_29_cfg_atomic; // @[ParallelMux.scala 90:77]
  assign io_resp_x = res_pmp_cfg_x & res_pma_cfg_x; // @[PMP.scala 580:28]
  assign io_resp_w = res_pmp_cfg_w & res_pma_cfg_w; // @[PMP.scala 579:28]
  assign io_resp_r = res_pmp_cfg_r & res_pma_cfg_r; // @[PMP.scala 578:28]
  always @(posedge clock) begin
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pmp_r17_0_cfg_x <= res_pmp_cur_cfg_x; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pmp_r17_0_cfg_w <= res_pmp_cur_cfg_w; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pmp_r17_0_cfg_r <= res_pmp_cur_cfg_r; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pmp_r17_1_cfg_x <= res_pmp_cur_1_cfg_x; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pmp_r17_1_cfg_w <= res_pmp_cur_1_cfg_w; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pmp_r17_1_cfg_r <= res_pmp_cur_1_cfg_r; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pmp_r17_2_cfg_x <= res_pmp_cur_2_cfg_x; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pmp_r17_2_cfg_w <= res_pmp_cur_2_cfg_w; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pmp_r17_2_cfg_r <= res_pmp_cur_2_cfg_r; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pmp_r17_3_cfg_x <= res_pmp_cur_3_cfg_x; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pmp_r17_3_cfg_w <= res_pmp_cur_3_cfg_w; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pmp_r17_3_cfg_r <= res_pmp_cur_3_cfg_r; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pmp_r17_4_cfg_x <= res_pmp_cur_4_cfg_x; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pmp_r17_4_cfg_w <= res_pmp_cur_4_cfg_w; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pmp_r17_4_cfg_r <= res_pmp_cur_4_cfg_r; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pmp_r17_5_cfg_x <= res_pmp_cur_5_cfg_x; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pmp_r17_5_cfg_w <= res_pmp_cur_5_cfg_w; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pmp_r17_5_cfg_r <= res_pmp_cur_5_cfg_r; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pmp_r17_6_cfg_x <= res_pmp_cur_6_cfg_x; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pmp_r17_6_cfg_w <= res_pmp_cur_6_cfg_w; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pmp_r17_6_cfg_r <= res_pmp_cur_6_cfg_r; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pmp_r17_7_cfg_x <= res_pmp_cur_7_cfg_x; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pmp_r17_7_cfg_w <= res_pmp_cur_7_cfg_w; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pmp_r17_7_cfg_r <= res_pmp_cur_7_cfg_r; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pmp_r17_8_cfg_x <= res_pmp_cur_8_cfg_x; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pmp_r17_8_cfg_w <= res_pmp_cur_8_cfg_w; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pmp_r17_8_cfg_r <= res_pmp_cur_8_cfg_r; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pmp_r17_9_cfg_x <= res_pmp_cur_9_cfg_x; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pmp_r17_9_cfg_w <= res_pmp_cur_9_cfg_w; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pmp_r17_9_cfg_r <= res_pmp_cur_9_cfg_r; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pmp_r17_10_cfg_x <= res_pmp_cur_10_cfg_x; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pmp_r17_10_cfg_w <= res_pmp_cur_10_cfg_w; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pmp_r17_10_cfg_r <= res_pmp_cur_10_cfg_r; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pmp_r17_11_cfg_x <= res_pmp_cur_11_cfg_x; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pmp_r17_11_cfg_w <= res_pmp_cur_11_cfg_w; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pmp_r17_11_cfg_r <= res_pmp_cur_11_cfg_r; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pmp_r17_12_cfg_x <= res_pmp_cur_12_cfg_x; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pmp_r17_12_cfg_w <= res_pmp_cur_12_cfg_w; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pmp_r17_12_cfg_r <= res_pmp_cur_12_cfg_r; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pmp_r17_13_cfg_x <= res_pmp_cur_13_cfg_x; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pmp_r17_13_cfg_w <= res_pmp_cur_13_cfg_w; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pmp_r17_13_cfg_r <= res_pmp_cur_13_cfg_r; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pmp_r17_14_cfg_x <= res_pmp_cur_14_cfg_x; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pmp_r17_14_cfg_w <= res_pmp_cur_14_cfg_w; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pmp_r17_14_cfg_r <= res_pmp_cur_14_cfg_r; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pmp_r17_15_cfg_x <= res_pmp_cur_15_cfg_x; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pmp_r17_15_cfg_w <= res_pmp_cur_15_cfg_w; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pmp_r17_15_cfg_r <= res_pmp_cur_15_cfg_r; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pmp_r17_16_cfg_x <= res_pmp_passThrough; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pmp_r17_16_cfg_w <= res_pmp_passThrough; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pmp_r17_16_cfg_r <= res_pmp_passThrough; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pma_r17_0_cfg_c <= io_check_env_pma_0_cfg_c; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pma_r17_0_cfg_atomic <= io_check_env_pma_0_cfg_atomic; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pma_r17_0_cfg_x <= io_check_env_pma_0_cfg_x; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pma_r17_0_cfg_w <= io_check_env_pma_0_cfg_w; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pma_r17_0_cfg_r <= io_check_env_pma_0_cfg_r; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pma_r17_1_cfg_c <= io_check_env_pma_1_cfg_c; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pma_r17_1_cfg_atomic <= io_check_env_pma_1_cfg_atomic; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pma_r17_1_cfg_x <= io_check_env_pma_1_cfg_x; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pma_r17_1_cfg_w <= io_check_env_pma_1_cfg_w; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pma_r17_1_cfg_r <= io_check_env_pma_1_cfg_r; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pma_r17_2_cfg_c <= io_check_env_pma_2_cfg_c; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pma_r17_2_cfg_atomic <= io_check_env_pma_2_cfg_atomic; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pma_r17_2_cfg_x <= io_check_env_pma_2_cfg_x; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pma_r17_2_cfg_w <= io_check_env_pma_2_cfg_w; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pma_r17_2_cfg_r <= io_check_env_pma_2_cfg_r; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pma_r17_3_cfg_c <= io_check_env_pma_3_cfg_c; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pma_r17_3_cfg_atomic <= io_check_env_pma_3_cfg_atomic; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pma_r17_3_cfg_x <= io_check_env_pma_3_cfg_x; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pma_r17_3_cfg_w <= io_check_env_pma_3_cfg_w; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pma_r17_3_cfg_r <= io_check_env_pma_3_cfg_r; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pma_r17_4_cfg_c <= io_check_env_pma_4_cfg_c; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pma_r17_4_cfg_atomic <= io_check_env_pma_4_cfg_atomic; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pma_r17_4_cfg_x <= io_check_env_pma_4_cfg_x; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pma_r17_4_cfg_w <= io_check_env_pma_4_cfg_w; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pma_r17_4_cfg_r <= io_check_env_pma_4_cfg_r; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pma_r17_5_cfg_c <= io_check_env_pma_5_cfg_c; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pma_r17_5_cfg_atomic <= io_check_env_pma_5_cfg_atomic; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pma_r17_5_cfg_x <= io_check_env_pma_5_cfg_x; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pma_r17_5_cfg_w <= io_check_env_pma_5_cfg_w; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pma_r17_5_cfg_r <= io_check_env_pma_5_cfg_r; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pma_r17_6_cfg_c <= io_check_env_pma_6_cfg_c; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pma_r17_6_cfg_atomic <= io_check_env_pma_6_cfg_atomic; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pma_r17_6_cfg_x <= io_check_env_pma_6_cfg_x; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pma_r17_6_cfg_w <= io_check_env_pma_6_cfg_w; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pma_r17_6_cfg_r <= io_check_env_pma_6_cfg_r; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pma_r17_7_cfg_c <= io_check_env_pma_7_cfg_c; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pma_r17_7_cfg_atomic <= io_check_env_pma_7_cfg_atomic; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pma_r17_7_cfg_x <= io_check_env_pma_7_cfg_x; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pma_r17_7_cfg_w <= io_check_env_pma_7_cfg_w; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pma_r17_7_cfg_r <= io_check_env_pma_7_cfg_r; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pma_r17_8_cfg_c <= io_check_env_pma_8_cfg_c; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pma_r17_8_cfg_atomic <= io_check_env_pma_8_cfg_atomic; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pma_r17_8_cfg_x <= io_check_env_pma_8_cfg_x; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pma_r17_8_cfg_w <= io_check_env_pma_8_cfg_w; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pma_r17_8_cfg_r <= io_check_env_pma_8_cfg_r; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pma_r17_9_cfg_c <= io_check_env_pma_9_cfg_c; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pma_r17_9_cfg_atomic <= io_check_env_pma_9_cfg_atomic; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pma_r17_9_cfg_x <= io_check_env_pma_9_cfg_x; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pma_r17_9_cfg_w <= io_check_env_pma_9_cfg_w; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pma_r17_9_cfg_r <= io_check_env_pma_9_cfg_r; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pma_r17_10_cfg_c <= io_check_env_pma_10_cfg_c; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pma_r17_10_cfg_atomic <= io_check_env_pma_10_cfg_atomic; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pma_r17_10_cfg_x <= io_check_env_pma_10_cfg_x; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pma_r17_10_cfg_w <= io_check_env_pma_10_cfg_w; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pma_r17_10_cfg_r <= io_check_env_pma_10_cfg_r; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pma_r17_11_cfg_c <= io_check_env_pma_11_cfg_c; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pma_r17_11_cfg_atomic <= io_check_env_pma_11_cfg_atomic; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pma_r17_11_cfg_x <= io_check_env_pma_11_cfg_x; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pma_r17_11_cfg_w <= io_check_env_pma_11_cfg_w; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pma_r17_11_cfg_r <= io_check_env_pma_11_cfg_r; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pma_r17_12_cfg_c <= io_check_env_pma_12_cfg_c; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pma_r17_12_cfg_atomic <= io_check_env_pma_12_cfg_atomic; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pma_r17_12_cfg_x <= io_check_env_pma_12_cfg_x; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pma_r17_12_cfg_w <= io_check_env_pma_12_cfg_w; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pma_r17_12_cfg_r <= io_check_env_pma_12_cfg_r; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pma_r17_13_cfg_c <= io_check_env_pma_13_cfg_c; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pma_r17_13_cfg_atomic <= io_check_env_pma_13_cfg_atomic; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pma_r17_13_cfg_x <= io_check_env_pma_13_cfg_x; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pma_r17_13_cfg_w <= io_check_env_pma_13_cfg_w; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pma_r17_13_cfg_r <= io_check_env_pma_13_cfg_r; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pma_r17_14_cfg_c <= io_check_env_pma_14_cfg_c; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pma_r17_14_cfg_atomic <= io_check_env_pma_14_cfg_atomic; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pma_r17_14_cfg_x <= io_check_env_pma_14_cfg_x; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pma_r17_14_cfg_w <= io_check_env_pma_14_cfg_w; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pma_r17_14_cfg_r <= io_check_env_pma_14_cfg_r; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pma_r17_15_cfg_c <= io_check_env_pma_15_cfg_c; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pma_r17_15_cfg_atomic <= io_check_env_pma_15_cfg_atomic; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pma_r17_15_cfg_x <= io_check_env_pma_15_cfg_x; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pma_r17_15_cfg_w <= io_check_env_pma_15_cfg_w; // @[Reg.scala 17:22]
    end
    if (io_req_valid) begin // @[Reg.scala 17:18]
      res_pma_r17_15_cfg_r <= io_check_env_pma_15_cfg_r; // @[Reg.scala 17:22]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      res_pmp_r <= 1'h0; // @[PMP.scala 199:8]
    end else if (io_req_valid) begin // @[Reg.scala 28:20]
      if (io_check_env_pmp_0_cfg_a[1]) begin
        res_pmp_r <= _res_pmp_is_match_T_8;
      end else begin
        res_pmp_r <= _res_pmp_is_match_T_20;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      res_pmp_r1 <= 1'h0; // @[PMP.scala 199:8]
    end else if (io_req_valid) begin // @[Reg.scala 28:20]
      if (io_check_env_pmp_1_cfg_a[1]) begin
        res_pmp_r1 <= _res_pmp_is_match_T_29;
      end else begin
        res_pmp_r1 <= _res_pmp_is_match_T_41;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      res_pmp_r2 <= 1'h0; // @[PMP.scala 199:8]
    end else if (io_req_valid) begin // @[Reg.scala 28:20]
      if (io_check_env_pmp_2_cfg_a[1]) begin
        res_pmp_r2 <= _res_pmp_is_match_T_50;
      end else begin
        res_pmp_r2 <= _res_pmp_is_match_T_62;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      res_pmp_r3 <= 1'h0; // @[PMP.scala 199:8]
    end else if (io_req_valid) begin // @[Reg.scala 28:20]
      if (io_check_env_pmp_3_cfg_a[1]) begin
        res_pmp_r3 <= _res_pmp_is_match_T_71;
      end else begin
        res_pmp_r3 <= _res_pmp_is_match_T_83;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      res_pmp_r4 <= 1'h0; // @[PMP.scala 199:8]
    end else if (io_req_valid) begin // @[Reg.scala 28:20]
      if (io_check_env_pmp_4_cfg_a[1]) begin
        res_pmp_r4 <= _res_pmp_is_match_T_92;
      end else begin
        res_pmp_r4 <= _res_pmp_is_match_T_104;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      res_pmp_r5 <= 1'h0; // @[PMP.scala 199:8]
    end else if (io_req_valid) begin // @[Reg.scala 28:20]
      if (io_check_env_pmp_5_cfg_a[1]) begin
        res_pmp_r5 <= _res_pmp_is_match_T_113;
      end else begin
        res_pmp_r5 <= _res_pmp_is_match_T_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      res_pmp_r6 <= 1'h0; // @[PMP.scala 199:8]
    end else if (io_req_valid) begin // @[Reg.scala 28:20]
      if (io_check_env_pmp_6_cfg_a[1]) begin
        res_pmp_r6 <= _res_pmp_is_match_T_134;
      end else begin
        res_pmp_r6 <= _res_pmp_is_match_T_146;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      res_pmp_r7 <= 1'h0; // @[PMP.scala 199:8]
    end else if (io_req_valid) begin // @[Reg.scala 28:20]
      if (io_check_env_pmp_7_cfg_a[1]) begin
        res_pmp_r7 <= _res_pmp_is_match_T_155;
      end else begin
        res_pmp_r7 <= _res_pmp_is_match_T_167;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      res_pmp_r8 <= 1'h0; // @[PMP.scala 199:8]
    end else if (io_req_valid) begin // @[Reg.scala 28:20]
      if (io_check_env_pmp_8_cfg_a[1]) begin
        res_pmp_r8 <= _res_pmp_is_match_T_176;
      end else begin
        res_pmp_r8 <= _res_pmp_is_match_T_188;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      res_pmp_r9 <= 1'h0; // @[PMP.scala 199:8]
    end else if (io_req_valid) begin // @[Reg.scala 28:20]
      if (io_check_env_pmp_9_cfg_a[1]) begin
        res_pmp_r9 <= _res_pmp_is_match_T_197;
      end else begin
        res_pmp_r9 <= _res_pmp_is_match_T_209;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      res_pmp_r10 <= 1'h0; // @[PMP.scala 199:8]
    end else if (io_req_valid) begin // @[Reg.scala 28:20]
      if (io_check_env_pmp_10_cfg_a[1]) begin
        res_pmp_r10 <= _res_pmp_is_match_T_218;
      end else begin
        res_pmp_r10 <= _res_pmp_is_match_T_230;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      res_pmp_r11 <= 1'h0; // @[PMP.scala 199:8]
    end else if (io_req_valid) begin // @[Reg.scala 28:20]
      if (io_check_env_pmp_11_cfg_a[1]) begin
        res_pmp_r11 <= _res_pmp_is_match_T_239;
      end else begin
        res_pmp_r11 <= _res_pmp_is_match_T_251;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      res_pmp_r12 <= 1'h0; // @[PMP.scala 199:8]
    end else if (io_req_valid) begin // @[Reg.scala 28:20]
      if (io_check_env_pmp_12_cfg_a[1]) begin
        res_pmp_r12 <= _res_pmp_is_match_T_260;
      end else begin
        res_pmp_r12 <= _res_pmp_is_match_T_272;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      res_pmp_r13 <= 1'h0; // @[PMP.scala 199:8]
    end else if (io_req_valid) begin // @[Reg.scala 28:20]
      if (io_check_env_pmp_13_cfg_a[1]) begin
        res_pmp_r13 <= _res_pmp_is_match_T_281;
      end else begin
        res_pmp_r13 <= _res_pmp_is_match_T_293;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      res_pmp_r14 <= 1'h0; // @[PMP.scala 199:8]
    end else if (io_req_valid) begin // @[Reg.scala 28:20]
      if (io_check_env_pmp_14_cfg_a[1]) begin
        res_pmp_r14 <= _res_pmp_is_match_T_302;
      end else begin
        res_pmp_r14 <= _res_pmp_is_match_T_314;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      res_pmp_r15 <= 1'h0; // @[PMP.scala 199:8]
    end else if (io_req_valid) begin // @[Reg.scala 28:20]
      if (io_check_env_pmp_15_cfg_a[1]) begin
        res_pmp_r15 <= _res_pmp_is_match_T_323;
      end else begin
        res_pmp_r15 <= _res_pmp_is_match_T_335;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      res_pma_r <= 1'h0; // @[PMP.scala 199:8]
    end else if (io_req_valid) begin // @[Reg.scala 28:20]
      if (io_check_env_pma_0_cfg_a[1]) begin
        res_pma_r <= _res_pma_is_match_T_8;
      end else begin
        res_pma_r <= _res_pma_is_match_T_20;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      res_pma_r1 <= 1'h0; // @[PMP.scala 199:8]
    end else if (io_req_valid) begin // @[Reg.scala 28:20]
      if (io_check_env_pma_1_cfg_a[1]) begin
        res_pma_r1 <= _res_pma_is_match_T_29;
      end else begin
        res_pma_r1 <= _res_pma_is_match_T_41;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      res_pma_r2 <= 1'h0; // @[PMP.scala 199:8]
    end else if (io_req_valid) begin // @[Reg.scala 28:20]
      if (io_check_env_pma_2_cfg_a[1]) begin
        res_pma_r2 <= _res_pma_is_match_T_50;
      end else begin
        res_pma_r2 <= _res_pma_is_match_T_62;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      res_pma_r3 <= 1'h0; // @[PMP.scala 199:8]
    end else if (io_req_valid) begin // @[Reg.scala 28:20]
      if (io_check_env_pma_3_cfg_a[1]) begin
        res_pma_r3 <= _res_pma_is_match_T_71;
      end else begin
        res_pma_r3 <= _res_pma_is_match_T_83;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      res_pma_r4 <= 1'h0; // @[PMP.scala 199:8]
    end else if (io_req_valid) begin // @[Reg.scala 28:20]
      if (io_check_env_pma_4_cfg_a[1]) begin
        res_pma_r4 <= _res_pma_is_match_T_92;
      end else begin
        res_pma_r4 <= _res_pma_is_match_T_104;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      res_pma_r5 <= 1'h0; // @[PMP.scala 199:8]
    end else if (io_req_valid) begin // @[Reg.scala 28:20]
      if (io_check_env_pma_5_cfg_a[1]) begin
        res_pma_r5 <= _res_pma_is_match_T_113;
      end else begin
        res_pma_r5 <= _res_pma_is_match_T_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      res_pma_r6 <= 1'h0; // @[PMP.scala 199:8]
    end else if (io_req_valid) begin // @[Reg.scala 28:20]
      if (io_check_env_pma_6_cfg_a[1]) begin
        res_pma_r6 <= _res_pma_is_match_T_134;
      end else begin
        res_pma_r6 <= _res_pma_is_match_T_146;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      res_pma_r7 <= 1'h0; // @[PMP.scala 199:8]
    end else if (io_req_valid) begin // @[Reg.scala 28:20]
      if (io_check_env_pma_7_cfg_a[1]) begin
        res_pma_r7 <= _res_pma_is_match_T_155;
      end else begin
        res_pma_r7 <= _res_pma_is_match_T_167;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      res_pma_r8 <= 1'h0; // @[PMP.scala 199:8]
    end else if (io_req_valid) begin // @[Reg.scala 28:20]
      if (io_check_env_pma_8_cfg_a[1]) begin
        res_pma_r8 <= _res_pma_is_match_T_176;
      end else begin
        res_pma_r8 <= _res_pma_is_match_T_188;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      res_pma_r9 <= 1'h0; // @[PMP.scala 199:8]
    end else if (io_req_valid) begin // @[Reg.scala 28:20]
      if (io_check_env_pma_9_cfg_a[1]) begin
        res_pma_r9 <= _res_pma_is_match_T_197;
      end else begin
        res_pma_r9 <= _res_pma_is_match_T_209;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      res_pma_r10 <= 1'h0; // @[PMP.scala 199:8]
    end else if (io_req_valid) begin // @[Reg.scala 28:20]
      if (io_check_env_pma_10_cfg_a[1]) begin
        res_pma_r10 <= _res_pma_is_match_T_218;
      end else begin
        res_pma_r10 <= _res_pma_is_match_T_230;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      res_pma_r11 <= 1'h0; // @[PMP.scala 199:8]
    end else if (io_req_valid) begin // @[Reg.scala 28:20]
      if (io_check_env_pma_11_cfg_a[1]) begin
        res_pma_r11 <= _res_pma_is_match_T_239;
      end else begin
        res_pma_r11 <= _res_pma_is_match_T_251;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      res_pma_r12 <= 1'h0; // @[PMP.scala 199:8]
    end else if (io_req_valid) begin // @[Reg.scala 28:20]
      if (io_check_env_pma_12_cfg_a[1]) begin
        res_pma_r12 <= _res_pma_is_match_T_260;
      end else begin
        res_pma_r12 <= _res_pma_is_match_T_272;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      res_pma_r13 <= 1'h0; // @[PMP.scala 199:8]
    end else if (io_req_valid) begin // @[Reg.scala 28:20]
      if (io_check_env_pma_13_cfg_a[1]) begin
        res_pma_r13 <= _res_pma_is_match_T_281;
      end else begin
        res_pma_r13 <= _res_pma_is_match_T_293;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      res_pma_r14 <= 1'h0; // @[PMP.scala 199:8]
    end else if (io_req_valid) begin // @[Reg.scala 28:20]
      if (io_check_env_pma_14_cfg_a[1]) begin
        res_pma_r14 <= _res_pma_is_match_T_302;
      end else begin
        res_pma_r14 <= _res_pma_is_match_T_314;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      res_pma_r15 <= 1'h0; // @[PMP.scala 199:8]
    end else if (io_req_valid) begin // @[Reg.scala 28:20]
      if (io_check_env_pma_15_cfg_a[1]) begin
        res_pma_r15 <= _res_pma_is_match_T_323;
      end else begin
        res_pma_r15 <= _res_pma_is_match_T_335;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  res_pmp_r = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  res_pmp_r1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  res_pmp_r2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  res_pmp_r3 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  res_pmp_r4 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  res_pmp_r5 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  res_pmp_r6 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  res_pmp_r7 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  res_pmp_r8 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  res_pmp_r9 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  res_pmp_r10 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  res_pmp_r11 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  res_pmp_r12 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  res_pmp_r13 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  res_pmp_r14 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  res_pmp_r15 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  res_pmp_r17_0_cfg_x = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  res_pmp_r17_0_cfg_w = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  res_pmp_r17_0_cfg_r = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  res_pmp_r17_1_cfg_x = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  res_pmp_r17_1_cfg_w = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  res_pmp_r17_1_cfg_r = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  res_pmp_r17_2_cfg_x = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  res_pmp_r17_2_cfg_w = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  res_pmp_r17_2_cfg_r = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  res_pmp_r17_3_cfg_x = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  res_pmp_r17_3_cfg_w = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  res_pmp_r17_3_cfg_r = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  res_pmp_r17_4_cfg_x = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  res_pmp_r17_4_cfg_w = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  res_pmp_r17_4_cfg_r = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  res_pmp_r17_5_cfg_x = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  res_pmp_r17_5_cfg_w = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  res_pmp_r17_5_cfg_r = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  res_pmp_r17_6_cfg_x = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  res_pmp_r17_6_cfg_w = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  res_pmp_r17_6_cfg_r = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  res_pmp_r17_7_cfg_x = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  res_pmp_r17_7_cfg_w = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  res_pmp_r17_7_cfg_r = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  res_pmp_r17_8_cfg_x = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  res_pmp_r17_8_cfg_w = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  res_pmp_r17_8_cfg_r = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  res_pmp_r17_9_cfg_x = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  res_pmp_r17_9_cfg_w = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  res_pmp_r17_9_cfg_r = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  res_pmp_r17_10_cfg_x = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  res_pmp_r17_10_cfg_w = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  res_pmp_r17_10_cfg_r = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  res_pmp_r17_11_cfg_x = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  res_pmp_r17_11_cfg_w = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  res_pmp_r17_11_cfg_r = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  res_pmp_r17_12_cfg_x = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  res_pmp_r17_12_cfg_w = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  res_pmp_r17_12_cfg_r = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  res_pmp_r17_13_cfg_x = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  res_pmp_r17_13_cfg_w = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  res_pmp_r17_13_cfg_r = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  res_pmp_r17_14_cfg_x = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  res_pmp_r17_14_cfg_w = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  res_pmp_r17_14_cfg_r = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  res_pmp_r17_15_cfg_x = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  res_pmp_r17_15_cfg_w = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  res_pmp_r17_15_cfg_r = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  res_pmp_r17_16_cfg_x = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  res_pmp_r17_16_cfg_w = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  res_pmp_r17_16_cfg_r = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  res_pma_r = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  res_pma_r1 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  res_pma_r2 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  res_pma_r3 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  res_pma_r4 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  res_pma_r5 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  res_pma_r6 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  res_pma_r7 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  res_pma_r8 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  res_pma_r9 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  res_pma_r10 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  res_pma_r11 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  res_pma_r12 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  res_pma_r13 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  res_pma_r14 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  res_pma_r15 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  res_pma_r17_0_cfg_c = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  res_pma_r17_0_cfg_atomic = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  res_pma_r17_0_cfg_x = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  res_pma_r17_0_cfg_w = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  res_pma_r17_0_cfg_r = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  res_pma_r17_1_cfg_c = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  res_pma_r17_1_cfg_atomic = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  res_pma_r17_1_cfg_x = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  res_pma_r17_1_cfg_w = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  res_pma_r17_1_cfg_r = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  res_pma_r17_2_cfg_c = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  res_pma_r17_2_cfg_atomic = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  res_pma_r17_2_cfg_x = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  res_pma_r17_2_cfg_w = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  res_pma_r17_2_cfg_r = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  res_pma_r17_3_cfg_c = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  res_pma_r17_3_cfg_atomic = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  res_pma_r17_3_cfg_x = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  res_pma_r17_3_cfg_w = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  res_pma_r17_3_cfg_r = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  res_pma_r17_4_cfg_c = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  res_pma_r17_4_cfg_atomic = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  res_pma_r17_4_cfg_x = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  res_pma_r17_4_cfg_w = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  res_pma_r17_4_cfg_r = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  res_pma_r17_5_cfg_c = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  res_pma_r17_5_cfg_atomic = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  res_pma_r17_5_cfg_x = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  res_pma_r17_5_cfg_w = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  res_pma_r17_5_cfg_r = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  res_pma_r17_6_cfg_c = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  res_pma_r17_6_cfg_atomic = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  res_pma_r17_6_cfg_x = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  res_pma_r17_6_cfg_w = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  res_pma_r17_6_cfg_r = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  res_pma_r17_7_cfg_c = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  res_pma_r17_7_cfg_atomic = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  res_pma_r17_7_cfg_x = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  res_pma_r17_7_cfg_w = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  res_pma_r17_7_cfg_r = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  res_pma_r17_8_cfg_c = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  res_pma_r17_8_cfg_atomic = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  res_pma_r17_8_cfg_x = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  res_pma_r17_8_cfg_w = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  res_pma_r17_8_cfg_r = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  res_pma_r17_9_cfg_c = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  res_pma_r17_9_cfg_atomic = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  res_pma_r17_9_cfg_x = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  res_pma_r17_9_cfg_w = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  res_pma_r17_9_cfg_r = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  res_pma_r17_10_cfg_c = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  res_pma_r17_10_cfg_atomic = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  res_pma_r17_10_cfg_x = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  res_pma_r17_10_cfg_w = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  res_pma_r17_10_cfg_r = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  res_pma_r17_11_cfg_c = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  res_pma_r17_11_cfg_atomic = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  res_pma_r17_11_cfg_x = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  res_pma_r17_11_cfg_w = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  res_pma_r17_11_cfg_r = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  res_pma_r17_12_cfg_c = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  res_pma_r17_12_cfg_atomic = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  res_pma_r17_12_cfg_x = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  res_pma_r17_12_cfg_w = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  res_pma_r17_12_cfg_r = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  res_pma_r17_13_cfg_c = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  res_pma_r17_13_cfg_atomic = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  res_pma_r17_13_cfg_x = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  res_pma_r17_13_cfg_w = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  res_pma_r17_13_cfg_r = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  res_pma_r17_14_cfg_c = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  res_pma_r17_14_cfg_atomic = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  res_pma_r17_14_cfg_x = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  res_pma_r17_14_cfg_w = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  res_pma_r17_14_cfg_r = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  res_pma_r17_15_cfg_c = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  res_pma_r17_15_cfg_atomic = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  res_pma_r17_15_cfg_x = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  res_pma_r17_15_cfg_w = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  res_pma_r17_15_cfg_r = _RAND_162[0:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    res_pmp_r = 1'h0;
  end
  if (reset) begin
    res_pmp_r1 = 1'h0;
  end
  if (reset) begin
    res_pmp_r2 = 1'h0;
  end
  if (reset) begin
    res_pmp_r3 = 1'h0;
  end
  if (reset) begin
    res_pmp_r4 = 1'h0;
  end
  if (reset) begin
    res_pmp_r5 = 1'h0;
  end
  if (reset) begin
    res_pmp_r6 = 1'h0;
  end
  if (reset) begin
    res_pmp_r7 = 1'h0;
  end
  if (reset) begin
    res_pmp_r8 = 1'h0;
  end
  if (reset) begin
    res_pmp_r9 = 1'h0;
  end
  if (reset) begin
    res_pmp_r10 = 1'h0;
  end
  if (reset) begin
    res_pmp_r11 = 1'h0;
  end
  if (reset) begin
    res_pmp_r12 = 1'h0;
  end
  if (reset) begin
    res_pmp_r13 = 1'h0;
  end
  if (reset) begin
    res_pmp_r14 = 1'h0;
  end
  if (reset) begin
    res_pmp_r15 = 1'h0;
  end
  if (reset) begin
    res_pma_r = 1'h0;
  end
  if (reset) begin
    res_pma_r1 = 1'h0;
  end
  if (reset) begin
    res_pma_r2 = 1'h0;
  end
  if (reset) begin
    res_pma_r3 = 1'h0;
  end
  if (reset) begin
    res_pma_r4 = 1'h0;
  end
  if (reset) begin
    res_pma_r5 = 1'h0;
  end
  if (reset) begin
    res_pma_r6 = 1'h0;
  end
  if (reset) begin
    res_pma_r7 = 1'h0;
  end
  if (reset) begin
    res_pma_r8 = 1'h0;
  end
  if (reset) begin
    res_pma_r9 = 1'h0;
  end
  if (reset) begin
    res_pma_r10 = 1'h0;
  end
  if (reset) begin
    res_pma_r11 = 1'h0;
  end
  if (reset) begin
    res_pma_r12 = 1'h0;
  end
  if (reset) begin
    res_pma_r13 = 1'h0;
  end
  if (reset) begin
    res_pma_r14 = 1'h0;
  end
  if (reset) begin
    res_pma_r15 = 1'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule

