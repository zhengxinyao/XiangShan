module PayloadArray_2(
  input         clock,
  input  [7:0]  io_read_0_addr,
  output        io_read_0_data_cf_pd_isRVC,
  output [1:0]  io_read_0_data_cf_pd_brType,
  output        io_read_0_data_cf_pd_isCall,
  output        io_read_0_data_cf_pd_isRet,
  output        io_read_0_data_cf_pred_taken,
  output        io_read_0_data_cf_ftqPtr_flag,
  output [2:0]  io_read_0_data_cf_ftqPtr_value,
  output [2:0]  io_read_0_data_cf_ftqOffset,
  output [3:0]  io_read_0_data_ctrl_fuType,
  output [6:0]  io_read_0_data_ctrl_fuOpType,
  output        io_read_0_data_ctrl_rfWen,
  output        io_read_0_data_ctrl_fpWen,
  output [19:0] io_read_0_data_ctrl_imm,
  output        io_read_0_data_ctrl_fpu_isAddSub,
  output        io_read_0_data_ctrl_fpu_typeTagIn,
  output        io_read_0_data_ctrl_fpu_typeTagOut,
  output        io_read_0_data_ctrl_fpu_fromInt,
  output        io_read_0_data_ctrl_fpu_wflags,
  output        io_read_0_data_ctrl_fpu_fpWen,
  output [1:0]  io_read_0_data_ctrl_fpu_fmaCmd,
  output        io_read_0_data_ctrl_fpu_div,
  output        io_read_0_data_ctrl_fpu_sqrt,
  output        io_read_0_data_ctrl_fpu_fcvt,
  output [1:0]  io_read_0_data_ctrl_fpu_typ,
  output [1:0]  io_read_0_data_ctrl_fpu_fmt,
  output        io_read_0_data_ctrl_fpu_ren3,
  output [2:0]  io_read_0_data_ctrl_fpu_rm,
  output [5:0]  io_read_0_data_pdest,
  output        io_read_0_data_robIdx_flag,
  output [4:0]  io_read_0_data_robIdx_value,
  input  [7:0]  io_read_1_addr,
  output        io_read_1_data_cf_pd_isRVC,
  output [1:0]  io_read_1_data_cf_pd_brType,
  output        io_read_1_data_cf_pd_isCall,
  output        io_read_1_data_cf_pd_isRet,
  output        io_read_1_data_cf_pred_taken,
  output        io_read_1_data_cf_ftqPtr_flag,
  output [2:0]  io_read_1_data_cf_ftqPtr_value,
  output [2:0]  io_read_1_data_cf_ftqOffset,
  output [3:0]  io_read_1_data_ctrl_fuType,
  output [6:0]  io_read_1_data_ctrl_fuOpType,
  output        io_read_1_data_ctrl_rfWen,
  output        io_read_1_data_ctrl_fpWen,
  output [19:0] io_read_1_data_ctrl_imm,
  output        io_read_1_data_ctrl_fpu_isAddSub,
  output        io_read_1_data_ctrl_fpu_typeTagIn,
  output        io_read_1_data_ctrl_fpu_typeTagOut,
  output        io_read_1_data_ctrl_fpu_fromInt,
  output        io_read_1_data_ctrl_fpu_wflags,
  output        io_read_1_data_ctrl_fpu_fpWen,
  output [1:0]  io_read_1_data_ctrl_fpu_fmaCmd,
  output        io_read_1_data_ctrl_fpu_div,
  output        io_read_1_data_ctrl_fpu_sqrt,
  output        io_read_1_data_ctrl_fpu_fcvt,
  output [1:0]  io_read_1_data_ctrl_fpu_typ,
  output [1:0]  io_read_1_data_ctrl_fpu_fmt,
  output        io_read_1_data_ctrl_fpu_ren3,
  output [2:0]  io_read_1_data_ctrl_fpu_rm,
  output [5:0]  io_read_1_data_pdest,
  output        io_read_1_data_robIdx_flag,
  output [4:0]  io_read_1_data_robIdx_value,
  input         io_write_0_enable,
  input  [7:0]  io_write_0_addr,
  input         io_write_0_data_cf_pd_isRVC,
  input  [1:0]  io_write_0_data_cf_pd_brType,
  input         io_write_0_data_cf_pd_isCall,
  input         io_write_0_data_cf_pd_isRet,
  input         io_write_0_data_cf_pred_taken,
  input         io_write_0_data_cf_ftqPtr_flag,
  input  [2:0]  io_write_0_data_cf_ftqPtr_value,
  input  [2:0]  io_write_0_data_cf_ftqOffset,
  input  [3:0]  io_write_0_data_ctrl_fuType,
  input  [6:0]  io_write_0_data_ctrl_fuOpType,
  input         io_write_0_data_ctrl_rfWen,
  input         io_write_0_data_ctrl_fpWen,
  input  [19:0] io_write_0_data_ctrl_imm,
  input         io_write_0_data_ctrl_fpu_isAddSub,
  input         io_write_0_data_ctrl_fpu_typeTagIn,
  input         io_write_0_data_ctrl_fpu_typeTagOut,
  input         io_write_0_data_ctrl_fpu_fromInt,
  input         io_write_0_data_ctrl_fpu_wflags,
  input         io_write_0_data_ctrl_fpu_fpWen,
  input  [1:0]  io_write_0_data_ctrl_fpu_fmaCmd,
  input         io_write_0_data_ctrl_fpu_div,
  input         io_write_0_data_ctrl_fpu_sqrt,
  input         io_write_0_data_ctrl_fpu_fcvt,
  input  [1:0]  io_write_0_data_ctrl_fpu_typ,
  input  [1:0]  io_write_0_data_ctrl_fpu_fmt,
  input         io_write_0_data_ctrl_fpu_ren3,
  input  [2:0]  io_write_0_data_ctrl_fpu_rm,
  input  [5:0]  io_write_0_data_pdest,
  input         io_write_0_data_robIdx_flag,
  input  [4:0]  io_write_0_data_robIdx_value
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
`endif // RANDOMIZE_REG_INIT
  reg  payload_0_cf_pd_isRVC; // @[PayloadArray.scala 45:20]
  reg [1:0] payload_0_cf_pd_brType; // @[PayloadArray.scala 45:20]
  reg  payload_0_cf_pd_isCall; // @[PayloadArray.scala 45:20]
  reg  payload_0_cf_pd_isRet; // @[PayloadArray.scala 45:20]
  reg  payload_0_cf_pred_taken; // @[PayloadArray.scala 45:20]
  reg  payload_0_cf_ftqPtr_flag; // @[PayloadArray.scala 45:20]
  reg [2:0] payload_0_cf_ftqPtr_value; // @[PayloadArray.scala 45:20]
  reg [2:0] payload_0_cf_ftqOffset; // @[PayloadArray.scala 45:20]
  reg [3:0] payload_0_ctrl_fuType; // @[PayloadArray.scala 45:20]
  reg [6:0] payload_0_ctrl_fuOpType; // @[PayloadArray.scala 45:20]
  reg  payload_0_ctrl_rfWen; // @[PayloadArray.scala 45:20]
  reg  payload_0_ctrl_fpWen; // @[PayloadArray.scala 45:20]
  reg [19:0] payload_0_ctrl_imm; // @[PayloadArray.scala 45:20]
  reg  payload_0_ctrl_fpu_isAddSub; // @[PayloadArray.scala 45:20]
  reg  payload_0_ctrl_fpu_typeTagIn; // @[PayloadArray.scala 45:20]
  reg  payload_0_ctrl_fpu_typeTagOut; // @[PayloadArray.scala 45:20]
  reg  payload_0_ctrl_fpu_fromInt; // @[PayloadArray.scala 45:20]
  reg  payload_0_ctrl_fpu_wflags; // @[PayloadArray.scala 45:20]
  reg  payload_0_ctrl_fpu_fpWen; // @[PayloadArray.scala 45:20]
  reg [1:0] payload_0_ctrl_fpu_fmaCmd; // @[PayloadArray.scala 45:20]
  reg  payload_0_ctrl_fpu_div; // @[PayloadArray.scala 45:20]
  reg  payload_0_ctrl_fpu_sqrt; // @[PayloadArray.scala 45:20]
  reg  payload_0_ctrl_fpu_fcvt; // @[PayloadArray.scala 45:20]
  reg [1:0] payload_0_ctrl_fpu_typ; // @[PayloadArray.scala 45:20]
  reg [1:0] payload_0_ctrl_fpu_fmt; // @[PayloadArray.scala 45:20]
  reg  payload_0_ctrl_fpu_ren3; // @[PayloadArray.scala 45:20]
  reg [2:0] payload_0_ctrl_fpu_rm; // @[PayloadArray.scala 45:20]
  reg [5:0] payload_0_pdest; // @[PayloadArray.scala 45:20]
  reg  payload_0_robIdx_flag; // @[PayloadArray.scala 45:20]
  reg [4:0] payload_0_robIdx_value; // @[PayloadArray.scala 45:20]
  reg  payload_1_cf_pd_isRVC; // @[PayloadArray.scala 45:20]
  reg [1:0] payload_1_cf_pd_brType; // @[PayloadArray.scala 45:20]
  reg  payload_1_cf_pd_isCall; // @[PayloadArray.scala 45:20]
  reg  payload_1_cf_pd_isRet; // @[PayloadArray.scala 45:20]
  reg  payload_1_cf_pred_taken; // @[PayloadArray.scala 45:20]
  reg  payload_1_cf_ftqPtr_flag; // @[PayloadArray.scala 45:20]
  reg [2:0] payload_1_cf_ftqPtr_value; // @[PayloadArray.scala 45:20]
  reg [2:0] payload_1_cf_ftqOffset; // @[PayloadArray.scala 45:20]
  reg [3:0] payload_1_ctrl_fuType; // @[PayloadArray.scala 45:20]
  reg [6:0] payload_1_ctrl_fuOpType; // @[PayloadArray.scala 45:20]
  reg  payload_1_ctrl_rfWen; // @[PayloadArray.scala 45:20]
  reg  payload_1_ctrl_fpWen; // @[PayloadArray.scala 45:20]
  reg [19:0] payload_1_ctrl_imm; // @[PayloadArray.scala 45:20]
  reg  payload_1_ctrl_fpu_isAddSub; // @[PayloadArray.scala 45:20]
  reg  payload_1_ctrl_fpu_typeTagIn; // @[PayloadArray.scala 45:20]
  reg  payload_1_ctrl_fpu_typeTagOut; // @[PayloadArray.scala 45:20]
  reg  payload_1_ctrl_fpu_fromInt; // @[PayloadArray.scala 45:20]
  reg  payload_1_ctrl_fpu_wflags; // @[PayloadArray.scala 45:20]
  reg  payload_1_ctrl_fpu_fpWen; // @[PayloadArray.scala 45:20]
  reg [1:0] payload_1_ctrl_fpu_fmaCmd; // @[PayloadArray.scala 45:20]
  reg  payload_1_ctrl_fpu_div; // @[PayloadArray.scala 45:20]
  reg  payload_1_ctrl_fpu_sqrt; // @[PayloadArray.scala 45:20]
  reg  payload_1_ctrl_fpu_fcvt; // @[PayloadArray.scala 45:20]
  reg [1:0] payload_1_ctrl_fpu_typ; // @[PayloadArray.scala 45:20]
  reg [1:0] payload_1_ctrl_fpu_fmt; // @[PayloadArray.scala 45:20]
  reg  payload_1_ctrl_fpu_ren3; // @[PayloadArray.scala 45:20]
  reg [2:0] payload_1_ctrl_fpu_rm; // @[PayloadArray.scala 45:20]
  reg [5:0] payload_1_pdest; // @[PayloadArray.scala 45:20]
  reg  payload_1_robIdx_flag; // @[PayloadArray.scala 45:20]
  reg [4:0] payload_1_robIdx_value; // @[PayloadArray.scala 45:20]
  reg  payload_2_cf_pd_isRVC; // @[PayloadArray.scala 45:20]
  reg [1:0] payload_2_cf_pd_brType; // @[PayloadArray.scala 45:20]
  reg  payload_2_cf_pd_isCall; // @[PayloadArray.scala 45:20]
  reg  payload_2_cf_pd_isRet; // @[PayloadArray.scala 45:20]
  reg  payload_2_cf_pred_taken; // @[PayloadArray.scala 45:20]
  reg  payload_2_cf_ftqPtr_flag; // @[PayloadArray.scala 45:20]
  reg [2:0] payload_2_cf_ftqPtr_value; // @[PayloadArray.scala 45:20]
  reg [2:0] payload_2_cf_ftqOffset; // @[PayloadArray.scala 45:20]
  reg [3:0] payload_2_ctrl_fuType; // @[PayloadArray.scala 45:20]
  reg [6:0] payload_2_ctrl_fuOpType; // @[PayloadArray.scala 45:20]
  reg  payload_2_ctrl_rfWen; // @[PayloadArray.scala 45:20]
  reg  payload_2_ctrl_fpWen; // @[PayloadArray.scala 45:20]
  reg [19:0] payload_2_ctrl_imm; // @[PayloadArray.scala 45:20]
  reg  payload_2_ctrl_fpu_isAddSub; // @[PayloadArray.scala 45:20]
  reg  payload_2_ctrl_fpu_typeTagIn; // @[PayloadArray.scala 45:20]
  reg  payload_2_ctrl_fpu_typeTagOut; // @[PayloadArray.scala 45:20]
  reg  payload_2_ctrl_fpu_fromInt; // @[PayloadArray.scala 45:20]
  reg  payload_2_ctrl_fpu_wflags; // @[PayloadArray.scala 45:20]
  reg  payload_2_ctrl_fpu_fpWen; // @[PayloadArray.scala 45:20]
  reg [1:0] payload_2_ctrl_fpu_fmaCmd; // @[PayloadArray.scala 45:20]
  reg  payload_2_ctrl_fpu_div; // @[PayloadArray.scala 45:20]
  reg  payload_2_ctrl_fpu_sqrt; // @[PayloadArray.scala 45:20]
  reg  payload_2_ctrl_fpu_fcvt; // @[PayloadArray.scala 45:20]
  reg [1:0] payload_2_ctrl_fpu_typ; // @[PayloadArray.scala 45:20]
  reg [1:0] payload_2_ctrl_fpu_fmt; // @[PayloadArray.scala 45:20]
  reg  payload_2_ctrl_fpu_ren3; // @[PayloadArray.scala 45:20]
  reg [2:0] payload_2_ctrl_fpu_rm; // @[PayloadArray.scala 45:20]
  reg [5:0] payload_2_pdest; // @[PayloadArray.scala 45:20]
  reg  payload_2_robIdx_flag; // @[PayloadArray.scala 45:20]
  reg [4:0] payload_2_robIdx_value; // @[PayloadArray.scala 45:20]
  reg  payload_3_cf_pd_isRVC; // @[PayloadArray.scala 45:20]
  reg [1:0] payload_3_cf_pd_brType; // @[PayloadArray.scala 45:20]
  reg  payload_3_cf_pd_isCall; // @[PayloadArray.scala 45:20]
  reg  payload_3_cf_pd_isRet; // @[PayloadArray.scala 45:20]
  reg  payload_3_cf_pred_taken; // @[PayloadArray.scala 45:20]
  reg  payload_3_cf_ftqPtr_flag; // @[PayloadArray.scala 45:20]
  reg [2:0] payload_3_cf_ftqPtr_value; // @[PayloadArray.scala 45:20]
  reg [2:0] payload_3_cf_ftqOffset; // @[PayloadArray.scala 45:20]
  reg [3:0] payload_3_ctrl_fuType; // @[PayloadArray.scala 45:20]
  reg [6:0] payload_3_ctrl_fuOpType; // @[PayloadArray.scala 45:20]
  reg  payload_3_ctrl_rfWen; // @[PayloadArray.scala 45:20]
  reg  payload_3_ctrl_fpWen; // @[PayloadArray.scala 45:20]
  reg [19:0] payload_3_ctrl_imm; // @[PayloadArray.scala 45:20]
  reg  payload_3_ctrl_fpu_isAddSub; // @[PayloadArray.scala 45:20]
  reg  payload_3_ctrl_fpu_typeTagIn; // @[PayloadArray.scala 45:20]
  reg  payload_3_ctrl_fpu_typeTagOut; // @[PayloadArray.scala 45:20]
  reg  payload_3_ctrl_fpu_fromInt; // @[PayloadArray.scala 45:20]
  reg  payload_3_ctrl_fpu_wflags; // @[PayloadArray.scala 45:20]
  reg  payload_3_ctrl_fpu_fpWen; // @[PayloadArray.scala 45:20]
  reg [1:0] payload_3_ctrl_fpu_fmaCmd; // @[PayloadArray.scala 45:20]
  reg  payload_3_ctrl_fpu_div; // @[PayloadArray.scala 45:20]
  reg  payload_3_ctrl_fpu_sqrt; // @[PayloadArray.scala 45:20]
  reg  payload_3_ctrl_fpu_fcvt; // @[PayloadArray.scala 45:20]
  reg [1:0] payload_3_ctrl_fpu_typ; // @[PayloadArray.scala 45:20]
  reg [1:0] payload_3_ctrl_fpu_fmt; // @[PayloadArray.scala 45:20]
  reg  payload_3_ctrl_fpu_ren3; // @[PayloadArray.scala 45:20]
  reg [2:0] payload_3_ctrl_fpu_rm; // @[PayloadArray.scala 45:20]
  reg [5:0] payload_3_pdest; // @[PayloadArray.scala 45:20]
  reg  payload_3_robIdx_flag; // @[PayloadArray.scala 45:20]
  reg [4:0] payload_3_robIdx_value; // @[PayloadArray.scala 45:20]
  reg  payload_4_cf_pd_isRVC; // @[PayloadArray.scala 45:20]
  reg [1:0] payload_4_cf_pd_brType; // @[PayloadArray.scala 45:20]
  reg  payload_4_cf_pd_isCall; // @[PayloadArray.scala 45:20]
  reg  payload_4_cf_pd_isRet; // @[PayloadArray.scala 45:20]
  reg  payload_4_cf_pred_taken; // @[PayloadArray.scala 45:20]
  reg  payload_4_cf_ftqPtr_flag; // @[PayloadArray.scala 45:20]
  reg [2:0] payload_4_cf_ftqPtr_value; // @[PayloadArray.scala 45:20]
  reg [2:0] payload_4_cf_ftqOffset; // @[PayloadArray.scala 45:20]
  reg [3:0] payload_4_ctrl_fuType; // @[PayloadArray.scala 45:20]
  reg [6:0] payload_4_ctrl_fuOpType; // @[PayloadArray.scala 45:20]
  reg  payload_4_ctrl_rfWen; // @[PayloadArray.scala 45:20]
  reg  payload_4_ctrl_fpWen; // @[PayloadArray.scala 45:20]
  reg [19:0] payload_4_ctrl_imm; // @[PayloadArray.scala 45:20]
  reg  payload_4_ctrl_fpu_isAddSub; // @[PayloadArray.scala 45:20]
  reg  payload_4_ctrl_fpu_typeTagIn; // @[PayloadArray.scala 45:20]
  reg  payload_4_ctrl_fpu_typeTagOut; // @[PayloadArray.scala 45:20]
  reg  payload_4_ctrl_fpu_fromInt; // @[PayloadArray.scala 45:20]
  reg  payload_4_ctrl_fpu_wflags; // @[PayloadArray.scala 45:20]
  reg  payload_4_ctrl_fpu_fpWen; // @[PayloadArray.scala 45:20]
  reg [1:0] payload_4_ctrl_fpu_fmaCmd; // @[PayloadArray.scala 45:20]
  reg  payload_4_ctrl_fpu_div; // @[PayloadArray.scala 45:20]
  reg  payload_4_ctrl_fpu_sqrt; // @[PayloadArray.scala 45:20]
  reg  payload_4_ctrl_fpu_fcvt; // @[PayloadArray.scala 45:20]
  reg [1:0] payload_4_ctrl_fpu_typ; // @[PayloadArray.scala 45:20]
  reg [1:0] payload_4_ctrl_fpu_fmt; // @[PayloadArray.scala 45:20]
  reg  payload_4_ctrl_fpu_ren3; // @[PayloadArray.scala 45:20]
  reg [2:0] payload_4_ctrl_fpu_rm; // @[PayloadArray.scala 45:20]
  reg [5:0] payload_4_pdest; // @[PayloadArray.scala 45:20]
  reg  payload_4_robIdx_flag; // @[PayloadArray.scala 45:20]
  reg [4:0] payload_4_robIdx_value; // @[PayloadArray.scala 45:20]
  reg  payload_5_cf_pd_isRVC; // @[PayloadArray.scala 45:20]
  reg [1:0] payload_5_cf_pd_brType; // @[PayloadArray.scala 45:20]
  reg  payload_5_cf_pd_isCall; // @[PayloadArray.scala 45:20]
  reg  payload_5_cf_pd_isRet; // @[PayloadArray.scala 45:20]
  reg  payload_5_cf_pred_taken; // @[PayloadArray.scala 45:20]
  reg  payload_5_cf_ftqPtr_flag; // @[PayloadArray.scala 45:20]
  reg [2:0] payload_5_cf_ftqPtr_value; // @[PayloadArray.scala 45:20]
  reg [2:0] payload_5_cf_ftqOffset; // @[PayloadArray.scala 45:20]
  reg [3:0] payload_5_ctrl_fuType; // @[PayloadArray.scala 45:20]
  reg [6:0] payload_5_ctrl_fuOpType; // @[PayloadArray.scala 45:20]
  reg  payload_5_ctrl_rfWen; // @[PayloadArray.scala 45:20]
  reg  payload_5_ctrl_fpWen; // @[PayloadArray.scala 45:20]
  reg [19:0] payload_5_ctrl_imm; // @[PayloadArray.scala 45:20]
  reg  payload_5_ctrl_fpu_isAddSub; // @[PayloadArray.scala 45:20]
  reg  payload_5_ctrl_fpu_typeTagIn; // @[PayloadArray.scala 45:20]
  reg  payload_5_ctrl_fpu_typeTagOut; // @[PayloadArray.scala 45:20]
  reg  payload_5_ctrl_fpu_fromInt; // @[PayloadArray.scala 45:20]
  reg  payload_5_ctrl_fpu_wflags; // @[PayloadArray.scala 45:20]
  reg  payload_5_ctrl_fpu_fpWen; // @[PayloadArray.scala 45:20]
  reg [1:0] payload_5_ctrl_fpu_fmaCmd; // @[PayloadArray.scala 45:20]
  reg  payload_5_ctrl_fpu_div; // @[PayloadArray.scala 45:20]
  reg  payload_5_ctrl_fpu_sqrt; // @[PayloadArray.scala 45:20]
  reg  payload_5_ctrl_fpu_fcvt; // @[PayloadArray.scala 45:20]
  reg [1:0] payload_5_ctrl_fpu_typ; // @[PayloadArray.scala 45:20]
  reg [1:0] payload_5_ctrl_fpu_fmt; // @[PayloadArray.scala 45:20]
  reg  payload_5_ctrl_fpu_ren3; // @[PayloadArray.scala 45:20]
  reg [2:0] payload_5_ctrl_fpu_rm; // @[PayloadArray.scala 45:20]
  reg [5:0] payload_5_pdest; // @[PayloadArray.scala 45:20]
  reg  payload_5_robIdx_flag; // @[PayloadArray.scala 45:20]
  reg [4:0] payload_5_robIdx_value; // @[PayloadArray.scala 45:20]
  reg  payload_6_cf_pd_isRVC; // @[PayloadArray.scala 45:20]
  reg [1:0] payload_6_cf_pd_brType; // @[PayloadArray.scala 45:20]
  reg  payload_6_cf_pd_isCall; // @[PayloadArray.scala 45:20]
  reg  payload_6_cf_pd_isRet; // @[PayloadArray.scala 45:20]
  reg  payload_6_cf_pred_taken; // @[PayloadArray.scala 45:20]
  reg  payload_6_cf_ftqPtr_flag; // @[PayloadArray.scala 45:20]
  reg [2:0] payload_6_cf_ftqPtr_value; // @[PayloadArray.scala 45:20]
  reg [2:0] payload_6_cf_ftqOffset; // @[PayloadArray.scala 45:20]
  reg [3:0] payload_6_ctrl_fuType; // @[PayloadArray.scala 45:20]
  reg [6:0] payload_6_ctrl_fuOpType; // @[PayloadArray.scala 45:20]
  reg  payload_6_ctrl_rfWen; // @[PayloadArray.scala 45:20]
  reg  payload_6_ctrl_fpWen; // @[PayloadArray.scala 45:20]
  reg [19:0] payload_6_ctrl_imm; // @[PayloadArray.scala 45:20]
  reg  payload_6_ctrl_fpu_isAddSub; // @[PayloadArray.scala 45:20]
  reg  payload_6_ctrl_fpu_typeTagIn; // @[PayloadArray.scala 45:20]
  reg  payload_6_ctrl_fpu_typeTagOut; // @[PayloadArray.scala 45:20]
  reg  payload_6_ctrl_fpu_fromInt; // @[PayloadArray.scala 45:20]
  reg  payload_6_ctrl_fpu_wflags; // @[PayloadArray.scala 45:20]
  reg  payload_6_ctrl_fpu_fpWen; // @[PayloadArray.scala 45:20]
  reg [1:0] payload_6_ctrl_fpu_fmaCmd; // @[PayloadArray.scala 45:20]
  reg  payload_6_ctrl_fpu_div; // @[PayloadArray.scala 45:20]
  reg  payload_6_ctrl_fpu_sqrt; // @[PayloadArray.scala 45:20]
  reg  payload_6_ctrl_fpu_fcvt; // @[PayloadArray.scala 45:20]
  reg [1:0] payload_6_ctrl_fpu_typ; // @[PayloadArray.scala 45:20]
  reg [1:0] payload_6_ctrl_fpu_fmt; // @[PayloadArray.scala 45:20]
  reg  payload_6_ctrl_fpu_ren3; // @[PayloadArray.scala 45:20]
  reg [2:0] payload_6_ctrl_fpu_rm; // @[PayloadArray.scala 45:20]
  reg [5:0] payload_6_pdest; // @[PayloadArray.scala 45:20]
  reg  payload_6_robIdx_flag; // @[PayloadArray.scala 45:20]
  reg [4:0] payload_6_robIdx_value; // @[PayloadArray.scala 45:20]
  reg  payload_7_cf_pd_isRVC; // @[PayloadArray.scala 45:20]
  reg [1:0] payload_7_cf_pd_brType; // @[PayloadArray.scala 45:20]
  reg  payload_7_cf_pd_isCall; // @[PayloadArray.scala 45:20]
  reg  payload_7_cf_pd_isRet; // @[PayloadArray.scala 45:20]
  reg  payload_7_cf_pred_taken; // @[PayloadArray.scala 45:20]
  reg  payload_7_cf_ftqPtr_flag; // @[PayloadArray.scala 45:20]
  reg [2:0] payload_7_cf_ftqPtr_value; // @[PayloadArray.scala 45:20]
  reg [2:0] payload_7_cf_ftqOffset; // @[PayloadArray.scala 45:20]
  reg [3:0] payload_7_ctrl_fuType; // @[PayloadArray.scala 45:20]
  reg [6:0] payload_7_ctrl_fuOpType; // @[PayloadArray.scala 45:20]
  reg  payload_7_ctrl_rfWen; // @[PayloadArray.scala 45:20]
  reg  payload_7_ctrl_fpWen; // @[PayloadArray.scala 45:20]
  reg [19:0] payload_7_ctrl_imm; // @[PayloadArray.scala 45:20]
  reg  payload_7_ctrl_fpu_isAddSub; // @[PayloadArray.scala 45:20]
  reg  payload_7_ctrl_fpu_typeTagIn; // @[PayloadArray.scala 45:20]
  reg  payload_7_ctrl_fpu_typeTagOut; // @[PayloadArray.scala 45:20]
  reg  payload_7_ctrl_fpu_fromInt; // @[PayloadArray.scala 45:20]
  reg  payload_7_ctrl_fpu_wflags; // @[PayloadArray.scala 45:20]
  reg  payload_7_ctrl_fpu_fpWen; // @[PayloadArray.scala 45:20]
  reg [1:0] payload_7_ctrl_fpu_fmaCmd; // @[PayloadArray.scala 45:20]
  reg  payload_7_ctrl_fpu_div; // @[PayloadArray.scala 45:20]
  reg  payload_7_ctrl_fpu_sqrt; // @[PayloadArray.scala 45:20]
  reg  payload_7_ctrl_fpu_fcvt; // @[PayloadArray.scala 45:20]
  reg [1:0] payload_7_ctrl_fpu_typ; // @[PayloadArray.scala 45:20]
  reg [1:0] payload_7_ctrl_fpu_fmt; // @[PayloadArray.scala 45:20]
  reg  payload_7_ctrl_fpu_ren3; // @[PayloadArray.scala 45:20]
  reg [2:0] payload_7_ctrl_fpu_rm; // @[PayloadArray.scala 45:20]
  reg [5:0] payload_7_pdest; // @[PayloadArray.scala 45:20]
  reg  payload_7_robIdx_flag; // @[PayloadArray.scala 45:20]
  reg [4:0] payload_7_robIdx_value; // @[PayloadArray.scala 45:20]
  wire [4:0] _io_read_0_data_T_233 = io_read_0_addr[0] ? payload_0_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_234 = io_read_0_addr[1] ? payload_1_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_235 = io_read_0_addr[2] ? payload_2_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_236 = io_read_0_addr[3] ? payload_3_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_237 = io_read_0_addr[4] ? payload_4_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_238 = io_read_0_addr[5] ? payload_5_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_239 = io_read_0_addr[6] ? payload_6_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_240 = io_read_0_addr[7] ? payload_7_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_241 = _io_read_0_data_T_233 | _io_read_0_data_T_234; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_242 = _io_read_0_data_T_241 | _io_read_0_data_T_235; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_243 = _io_read_0_data_T_242 | _io_read_0_data_T_236; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_244 = _io_read_0_data_T_243 | _io_read_0_data_T_237; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_245 = _io_read_0_data_T_244 | _io_read_0_data_T_238; // @[Mux.scala 27:73]
  wire [4:0] _io_read_0_data_T_246 = _io_read_0_data_T_245 | _io_read_0_data_T_239; // @[Mux.scala 27:73]
  wire [5:0] _io_read_0_data_T_278 = io_read_0_addr[0] ? payload_0_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] _io_read_0_data_T_279 = io_read_0_addr[1] ? payload_1_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] _io_read_0_data_T_280 = io_read_0_addr[2] ? payload_2_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] _io_read_0_data_T_281 = io_read_0_addr[3] ? payload_3_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] _io_read_0_data_T_282 = io_read_0_addr[4] ? payload_4_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] _io_read_0_data_T_283 = io_read_0_addr[5] ? payload_5_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] _io_read_0_data_T_284 = io_read_0_addr[6] ? payload_6_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] _io_read_0_data_T_285 = io_read_0_addr[7] ? payload_7_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] _io_read_0_data_T_286 = _io_read_0_data_T_278 | _io_read_0_data_T_279; // @[Mux.scala 27:73]
  wire [5:0] _io_read_0_data_T_287 = _io_read_0_data_T_286 | _io_read_0_data_T_280; // @[Mux.scala 27:73]
  wire [5:0] _io_read_0_data_T_288 = _io_read_0_data_T_287 | _io_read_0_data_T_281; // @[Mux.scala 27:73]
  wire [5:0] _io_read_0_data_T_289 = _io_read_0_data_T_288 | _io_read_0_data_T_282; // @[Mux.scala 27:73]
  wire [5:0] _io_read_0_data_T_290 = _io_read_0_data_T_289 | _io_read_0_data_T_283; // @[Mux.scala 27:73]
  wire [5:0] _io_read_0_data_T_291 = _io_read_0_data_T_290 | _io_read_0_data_T_284; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_428 = io_read_0_addr[0] ? payload_0_ctrl_fpu_rm : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_429 = io_read_0_addr[1] ? payload_1_ctrl_fpu_rm : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_430 = io_read_0_addr[2] ? payload_2_ctrl_fpu_rm : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_431 = io_read_0_addr[3] ? payload_3_ctrl_fpu_rm : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_432 = io_read_0_addr[4] ? payload_4_ctrl_fpu_rm : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_433 = io_read_0_addr[5] ? payload_5_ctrl_fpu_rm : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_434 = io_read_0_addr[6] ? payload_6_ctrl_fpu_rm : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_435 = io_read_0_addr[7] ? payload_7_ctrl_fpu_rm : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_436 = _io_read_0_data_T_428 | _io_read_0_data_T_429; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_437 = _io_read_0_data_T_436 | _io_read_0_data_T_430; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_438 = _io_read_0_data_T_437 | _io_read_0_data_T_431; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_439 = _io_read_0_data_T_438 | _io_read_0_data_T_432; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_440 = _io_read_0_data_T_439 | _io_read_0_data_T_433; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_441 = _io_read_0_data_T_440 | _io_read_0_data_T_434; // @[Mux.scala 27:73]
  wire [1:0] _io_read_0_data_T_458 = io_read_0_addr[0] ? payload_0_ctrl_fpu_fmt : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_0_data_T_459 = io_read_0_addr[1] ? payload_1_ctrl_fpu_fmt : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_0_data_T_460 = io_read_0_addr[2] ? payload_2_ctrl_fpu_fmt : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_0_data_T_461 = io_read_0_addr[3] ? payload_3_ctrl_fpu_fmt : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_0_data_T_462 = io_read_0_addr[4] ? payload_4_ctrl_fpu_fmt : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_0_data_T_463 = io_read_0_addr[5] ? payload_5_ctrl_fpu_fmt : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_0_data_T_464 = io_read_0_addr[6] ? payload_6_ctrl_fpu_fmt : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_0_data_T_465 = io_read_0_addr[7] ? payload_7_ctrl_fpu_fmt : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_0_data_T_466 = _io_read_0_data_T_458 | _io_read_0_data_T_459; // @[Mux.scala 27:73]
  wire [1:0] _io_read_0_data_T_467 = _io_read_0_data_T_466 | _io_read_0_data_T_460; // @[Mux.scala 27:73]
  wire [1:0] _io_read_0_data_T_468 = _io_read_0_data_T_467 | _io_read_0_data_T_461; // @[Mux.scala 27:73]
  wire [1:0] _io_read_0_data_T_469 = _io_read_0_data_T_468 | _io_read_0_data_T_462; // @[Mux.scala 27:73]
  wire [1:0] _io_read_0_data_T_470 = _io_read_0_data_T_469 | _io_read_0_data_T_463; // @[Mux.scala 27:73]
  wire [1:0] _io_read_0_data_T_471 = _io_read_0_data_T_470 | _io_read_0_data_T_464; // @[Mux.scala 27:73]
  wire [1:0] _io_read_0_data_T_473 = io_read_0_addr[0] ? payload_0_ctrl_fpu_typ : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_0_data_T_474 = io_read_0_addr[1] ? payload_1_ctrl_fpu_typ : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_0_data_T_475 = io_read_0_addr[2] ? payload_2_ctrl_fpu_typ : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_0_data_T_476 = io_read_0_addr[3] ? payload_3_ctrl_fpu_typ : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_0_data_T_477 = io_read_0_addr[4] ? payload_4_ctrl_fpu_typ : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_0_data_T_478 = io_read_0_addr[5] ? payload_5_ctrl_fpu_typ : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_0_data_T_479 = io_read_0_addr[6] ? payload_6_ctrl_fpu_typ : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_0_data_T_480 = io_read_0_addr[7] ? payload_7_ctrl_fpu_typ : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_0_data_T_481 = _io_read_0_data_T_473 | _io_read_0_data_T_474; // @[Mux.scala 27:73]
  wire [1:0] _io_read_0_data_T_482 = _io_read_0_data_T_481 | _io_read_0_data_T_475; // @[Mux.scala 27:73]
  wire [1:0] _io_read_0_data_T_483 = _io_read_0_data_T_482 | _io_read_0_data_T_476; // @[Mux.scala 27:73]
  wire [1:0] _io_read_0_data_T_484 = _io_read_0_data_T_483 | _io_read_0_data_T_477; // @[Mux.scala 27:73]
  wire [1:0] _io_read_0_data_T_485 = _io_read_0_data_T_484 | _io_read_0_data_T_478; // @[Mux.scala 27:73]
  wire [1:0] _io_read_0_data_T_486 = _io_read_0_data_T_485 | _io_read_0_data_T_479; // @[Mux.scala 27:73]
  wire [1:0] _io_read_0_data_T_533 = io_read_0_addr[0] ? payload_0_ctrl_fpu_fmaCmd : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_0_data_T_534 = io_read_0_addr[1] ? payload_1_ctrl_fpu_fmaCmd : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_0_data_T_535 = io_read_0_addr[2] ? payload_2_ctrl_fpu_fmaCmd : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_0_data_T_536 = io_read_0_addr[3] ? payload_3_ctrl_fpu_fmaCmd : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_0_data_T_537 = io_read_0_addr[4] ? payload_4_ctrl_fpu_fmaCmd : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_0_data_T_538 = io_read_0_addr[5] ? payload_5_ctrl_fpu_fmaCmd : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_0_data_T_539 = io_read_0_addr[6] ? payload_6_ctrl_fpu_fmaCmd : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_0_data_T_540 = io_read_0_addr[7] ? payload_7_ctrl_fpu_fmaCmd : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_0_data_T_541 = _io_read_0_data_T_533 | _io_read_0_data_T_534; // @[Mux.scala 27:73]
  wire [1:0] _io_read_0_data_T_542 = _io_read_0_data_T_541 | _io_read_0_data_T_535; // @[Mux.scala 27:73]
  wire [1:0] _io_read_0_data_T_543 = _io_read_0_data_T_542 | _io_read_0_data_T_536; // @[Mux.scala 27:73]
  wire [1:0] _io_read_0_data_T_544 = _io_read_0_data_T_543 | _io_read_0_data_T_537; // @[Mux.scala 27:73]
  wire [1:0] _io_read_0_data_T_545 = _io_read_0_data_T_544 | _io_read_0_data_T_538; // @[Mux.scala 27:73]
  wire [1:0] _io_read_0_data_T_546 = _io_read_0_data_T_545 | _io_read_0_data_T_539; // @[Mux.scala 27:73]
  wire [19:0] _io_read_0_data_T_653 = io_read_0_addr[0] ? payload_0_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _io_read_0_data_T_654 = io_read_0_addr[1] ? payload_1_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _io_read_0_data_T_655 = io_read_0_addr[2] ? payload_2_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _io_read_0_data_T_656 = io_read_0_addr[3] ? payload_3_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _io_read_0_data_T_657 = io_read_0_addr[4] ? payload_4_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _io_read_0_data_T_658 = io_read_0_addr[5] ? payload_5_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _io_read_0_data_T_659 = io_read_0_addr[6] ? payload_6_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _io_read_0_data_T_660 = io_read_0_addr[7] ? payload_7_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _io_read_0_data_T_661 = _io_read_0_data_T_653 | _io_read_0_data_T_654; // @[Mux.scala 27:73]
  wire [19:0] _io_read_0_data_T_662 = _io_read_0_data_T_661 | _io_read_0_data_T_655; // @[Mux.scala 27:73]
  wire [19:0] _io_read_0_data_T_663 = _io_read_0_data_T_662 | _io_read_0_data_T_656; // @[Mux.scala 27:73]
  wire [19:0] _io_read_0_data_T_664 = _io_read_0_data_T_663 | _io_read_0_data_T_657; // @[Mux.scala 27:73]
  wire [19:0] _io_read_0_data_T_665 = _io_read_0_data_T_664 | _io_read_0_data_T_658; // @[Mux.scala 27:73]
  wire [19:0] _io_read_0_data_T_666 = _io_read_0_data_T_665 | _io_read_0_data_T_659; // @[Mux.scala 27:73]
  wire [6:0] _io_read_0_data_T_773 = io_read_0_addr[0] ? payload_0_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _io_read_0_data_T_774 = io_read_0_addr[1] ? payload_1_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _io_read_0_data_T_775 = io_read_0_addr[2] ? payload_2_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _io_read_0_data_T_776 = io_read_0_addr[3] ? payload_3_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _io_read_0_data_T_777 = io_read_0_addr[4] ? payload_4_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _io_read_0_data_T_778 = io_read_0_addr[5] ? payload_5_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _io_read_0_data_T_779 = io_read_0_addr[6] ? payload_6_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _io_read_0_data_T_780 = io_read_0_addr[7] ? payload_7_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _io_read_0_data_T_781 = _io_read_0_data_T_773 | _io_read_0_data_T_774; // @[Mux.scala 27:73]
  wire [6:0] _io_read_0_data_T_782 = _io_read_0_data_T_781 | _io_read_0_data_T_775; // @[Mux.scala 27:73]
  wire [6:0] _io_read_0_data_T_783 = _io_read_0_data_T_782 | _io_read_0_data_T_776; // @[Mux.scala 27:73]
  wire [6:0] _io_read_0_data_T_784 = _io_read_0_data_T_783 | _io_read_0_data_T_777; // @[Mux.scala 27:73]
  wire [6:0] _io_read_0_data_T_785 = _io_read_0_data_T_784 | _io_read_0_data_T_778; // @[Mux.scala 27:73]
  wire [6:0] _io_read_0_data_T_786 = _io_read_0_data_T_785 | _io_read_0_data_T_779; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_788 = io_read_0_addr[0] ? payload_0_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_789 = io_read_0_addr[1] ? payload_1_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_790 = io_read_0_addr[2] ? payload_2_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_791 = io_read_0_addr[3] ? payload_3_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_792 = io_read_0_addr[4] ? payload_4_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_793 = io_read_0_addr[5] ? payload_5_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_794 = io_read_0_addr[6] ? payload_6_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_795 = io_read_0_addr[7] ? payload_7_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_796 = _io_read_0_data_T_788 | _io_read_0_data_T_789; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_797 = _io_read_0_data_T_796 | _io_read_0_data_T_790; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_798 = _io_read_0_data_T_797 | _io_read_0_data_T_791; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_799 = _io_read_0_data_T_798 | _io_read_0_data_T_792; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_800 = _io_read_0_data_T_799 | _io_read_0_data_T_793; // @[Mux.scala 27:73]
  wire [3:0] _io_read_0_data_T_801 = _io_read_0_data_T_800 | _io_read_0_data_T_794; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_923 = io_read_0_addr[0] ? payload_0_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_924 = io_read_0_addr[1] ? payload_1_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_925 = io_read_0_addr[2] ? payload_2_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_926 = io_read_0_addr[3] ? payload_3_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_927 = io_read_0_addr[4] ? payload_4_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_928 = io_read_0_addr[5] ? payload_5_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_929 = io_read_0_addr[6] ? payload_6_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_930 = io_read_0_addr[7] ? payload_7_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_931 = _io_read_0_data_T_923 | _io_read_0_data_T_924; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_932 = _io_read_0_data_T_931 | _io_read_0_data_T_925; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_933 = _io_read_0_data_T_932 | _io_read_0_data_T_926; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_934 = _io_read_0_data_T_933 | _io_read_0_data_T_927; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_935 = _io_read_0_data_T_934 | _io_read_0_data_T_928; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_936 = _io_read_0_data_T_935 | _io_read_0_data_T_929; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_938 = io_read_0_addr[0] ? payload_0_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_939 = io_read_0_addr[1] ? payload_1_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_940 = io_read_0_addr[2] ? payload_2_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_941 = io_read_0_addr[3] ? payload_3_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_942 = io_read_0_addr[4] ? payload_4_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_943 = io_read_0_addr[5] ? payload_5_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_944 = io_read_0_addr[6] ? payload_6_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_945 = io_read_0_addr[7] ? payload_7_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_946 = _io_read_0_data_T_938 | _io_read_0_data_T_939; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_947 = _io_read_0_data_T_946 | _io_read_0_data_T_940; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_948 = _io_read_0_data_T_947 | _io_read_0_data_T_941; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_949 = _io_read_0_data_T_948 | _io_read_0_data_T_942; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_950 = _io_read_0_data_T_949 | _io_read_0_data_T_943; // @[Mux.scala 27:73]
  wire [2:0] _io_read_0_data_T_951 = _io_read_0_data_T_950 | _io_read_0_data_T_944; // @[Mux.scala 27:73]
  wire [1:0] _io_read_0_data_T_1118 = io_read_0_addr[0] ? payload_0_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_0_data_T_1119 = io_read_0_addr[1] ? payload_1_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_0_data_T_1120 = io_read_0_addr[2] ? payload_2_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_0_data_T_1121 = io_read_0_addr[3] ? payload_3_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_0_data_T_1122 = io_read_0_addr[4] ? payload_4_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_0_data_T_1123 = io_read_0_addr[5] ? payload_5_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_0_data_T_1124 = io_read_0_addr[6] ? payload_6_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_0_data_T_1125 = io_read_0_addr[7] ? payload_7_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_0_data_T_1126 = _io_read_0_data_T_1118 | _io_read_0_data_T_1119; // @[Mux.scala 27:73]
  wire [1:0] _io_read_0_data_T_1127 = _io_read_0_data_T_1126 | _io_read_0_data_T_1120; // @[Mux.scala 27:73]
  wire [1:0] _io_read_0_data_T_1128 = _io_read_0_data_T_1127 | _io_read_0_data_T_1121; // @[Mux.scala 27:73]
  wire [1:0] _io_read_0_data_T_1129 = _io_read_0_data_T_1128 | _io_read_0_data_T_1122; // @[Mux.scala 27:73]
  wire [1:0] _io_read_0_data_T_1130 = _io_read_0_data_T_1129 | _io_read_0_data_T_1123; // @[Mux.scala 27:73]
  wire [1:0] _io_read_0_data_T_1131 = _io_read_0_data_T_1130 | _io_read_0_data_T_1124; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_233 = io_read_1_addr[0] ? payload_0_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_234 = io_read_1_addr[1] ? payload_1_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_235 = io_read_1_addr[2] ? payload_2_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_236 = io_read_1_addr[3] ? payload_3_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_237 = io_read_1_addr[4] ? payload_4_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_238 = io_read_1_addr[5] ? payload_5_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_239 = io_read_1_addr[6] ? payload_6_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_240 = io_read_1_addr[7] ? payload_7_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_241 = _io_read_1_data_T_233 | _io_read_1_data_T_234; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_242 = _io_read_1_data_T_241 | _io_read_1_data_T_235; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_243 = _io_read_1_data_T_242 | _io_read_1_data_T_236; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_244 = _io_read_1_data_T_243 | _io_read_1_data_T_237; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_245 = _io_read_1_data_T_244 | _io_read_1_data_T_238; // @[Mux.scala 27:73]
  wire [4:0] _io_read_1_data_T_246 = _io_read_1_data_T_245 | _io_read_1_data_T_239; // @[Mux.scala 27:73]
  wire [5:0] _io_read_1_data_T_278 = io_read_1_addr[0] ? payload_0_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] _io_read_1_data_T_279 = io_read_1_addr[1] ? payload_1_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] _io_read_1_data_T_280 = io_read_1_addr[2] ? payload_2_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] _io_read_1_data_T_281 = io_read_1_addr[3] ? payload_3_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] _io_read_1_data_T_282 = io_read_1_addr[4] ? payload_4_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] _io_read_1_data_T_283 = io_read_1_addr[5] ? payload_5_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] _io_read_1_data_T_284 = io_read_1_addr[6] ? payload_6_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] _io_read_1_data_T_285 = io_read_1_addr[7] ? payload_7_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] _io_read_1_data_T_286 = _io_read_1_data_T_278 | _io_read_1_data_T_279; // @[Mux.scala 27:73]
  wire [5:0] _io_read_1_data_T_287 = _io_read_1_data_T_286 | _io_read_1_data_T_280; // @[Mux.scala 27:73]
  wire [5:0] _io_read_1_data_T_288 = _io_read_1_data_T_287 | _io_read_1_data_T_281; // @[Mux.scala 27:73]
  wire [5:0] _io_read_1_data_T_289 = _io_read_1_data_T_288 | _io_read_1_data_T_282; // @[Mux.scala 27:73]
  wire [5:0] _io_read_1_data_T_290 = _io_read_1_data_T_289 | _io_read_1_data_T_283; // @[Mux.scala 27:73]
  wire [5:0] _io_read_1_data_T_291 = _io_read_1_data_T_290 | _io_read_1_data_T_284; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_428 = io_read_1_addr[0] ? payload_0_ctrl_fpu_rm : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_429 = io_read_1_addr[1] ? payload_1_ctrl_fpu_rm : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_430 = io_read_1_addr[2] ? payload_2_ctrl_fpu_rm : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_431 = io_read_1_addr[3] ? payload_3_ctrl_fpu_rm : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_432 = io_read_1_addr[4] ? payload_4_ctrl_fpu_rm : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_433 = io_read_1_addr[5] ? payload_5_ctrl_fpu_rm : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_434 = io_read_1_addr[6] ? payload_6_ctrl_fpu_rm : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_435 = io_read_1_addr[7] ? payload_7_ctrl_fpu_rm : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_436 = _io_read_1_data_T_428 | _io_read_1_data_T_429; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_437 = _io_read_1_data_T_436 | _io_read_1_data_T_430; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_438 = _io_read_1_data_T_437 | _io_read_1_data_T_431; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_439 = _io_read_1_data_T_438 | _io_read_1_data_T_432; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_440 = _io_read_1_data_T_439 | _io_read_1_data_T_433; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_441 = _io_read_1_data_T_440 | _io_read_1_data_T_434; // @[Mux.scala 27:73]
  wire [1:0] _io_read_1_data_T_458 = io_read_1_addr[0] ? payload_0_ctrl_fpu_fmt : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_1_data_T_459 = io_read_1_addr[1] ? payload_1_ctrl_fpu_fmt : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_1_data_T_460 = io_read_1_addr[2] ? payload_2_ctrl_fpu_fmt : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_1_data_T_461 = io_read_1_addr[3] ? payload_3_ctrl_fpu_fmt : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_1_data_T_462 = io_read_1_addr[4] ? payload_4_ctrl_fpu_fmt : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_1_data_T_463 = io_read_1_addr[5] ? payload_5_ctrl_fpu_fmt : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_1_data_T_464 = io_read_1_addr[6] ? payload_6_ctrl_fpu_fmt : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_1_data_T_465 = io_read_1_addr[7] ? payload_7_ctrl_fpu_fmt : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_1_data_T_466 = _io_read_1_data_T_458 | _io_read_1_data_T_459; // @[Mux.scala 27:73]
  wire [1:0] _io_read_1_data_T_467 = _io_read_1_data_T_466 | _io_read_1_data_T_460; // @[Mux.scala 27:73]
  wire [1:0] _io_read_1_data_T_468 = _io_read_1_data_T_467 | _io_read_1_data_T_461; // @[Mux.scala 27:73]
  wire [1:0] _io_read_1_data_T_469 = _io_read_1_data_T_468 | _io_read_1_data_T_462; // @[Mux.scala 27:73]
  wire [1:0] _io_read_1_data_T_470 = _io_read_1_data_T_469 | _io_read_1_data_T_463; // @[Mux.scala 27:73]
  wire [1:0] _io_read_1_data_T_471 = _io_read_1_data_T_470 | _io_read_1_data_T_464; // @[Mux.scala 27:73]
  wire [1:0] _io_read_1_data_T_473 = io_read_1_addr[0] ? payload_0_ctrl_fpu_typ : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_1_data_T_474 = io_read_1_addr[1] ? payload_1_ctrl_fpu_typ : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_1_data_T_475 = io_read_1_addr[2] ? payload_2_ctrl_fpu_typ : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_1_data_T_476 = io_read_1_addr[3] ? payload_3_ctrl_fpu_typ : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_1_data_T_477 = io_read_1_addr[4] ? payload_4_ctrl_fpu_typ : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_1_data_T_478 = io_read_1_addr[5] ? payload_5_ctrl_fpu_typ : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_1_data_T_479 = io_read_1_addr[6] ? payload_6_ctrl_fpu_typ : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_1_data_T_480 = io_read_1_addr[7] ? payload_7_ctrl_fpu_typ : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_1_data_T_481 = _io_read_1_data_T_473 | _io_read_1_data_T_474; // @[Mux.scala 27:73]
  wire [1:0] _io_read_1_data_T_482 = _io_read_1_data_T_481 | _io_read_1_data_T_475; // @[Mux.scala 27:73]
  wire [1:0] _io_read_1_data_T_483 = _io_read_1_data_T_482 | _io_read_1_data_T_476; // @[Mux.scala 27:73]
  wire [1:0] _io_read_1_data_T_484 = _io_read_1_data_T_483 | _io_read_1_data_T_477; // @[Mux.scala 27:73]
  wire [1:0] _io_read_1_data_T_485 = _io_read_1_data_T_484 | _io_read_1_data_T_478; // @[Mux.scala 27:73]
  wire [1:0] _io_read_1_data_T_486 = _io_read_1_data_T_485 | _io_read_1_data_T_479; // @[Mux.scala 27:73]
  wire [1:0] _io_read_1_data_T_533 = io_read_1_addr[0] ? payload_0_ctrl_fpu_fmaCmd : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_1_data_T_534 = io_read_1_addr[1] ? payload_1_ctrl_fpu_fmaCmd : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_1_data_T_535 = io_read_1_addr[2] ? payload_2_ctrl_fpu_fmaCmd : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_1_data_T_536 = io_read_1_addr[3] ? payload_3_ctrl_fpu_fmaCmd : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_1_data_T_537 = io_read_1_addr[4] ? payload_4_ctrl_fpu_fmaCmd : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_1_data_T_538 = io_read_1_addr[5] ? payload_5_ctrl_fpu_fmaCmd : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_1_data_T_539 = io_read_1_addr[6] ? payload_6_ctrl_fpu_fmaCmd : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_1_data_T_540 = io_read_1_addr[7] ? payload_7_ctrl_fpu_fmaCmd : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_1_data_T_541 = _io_read_1_data_T_533 | _io_read_1_data_T_534; // @[Mux.scala 27:73]
  wire [1:0] _io_read_1_data_T_542 = _io_read_1_data_T_541 | _io_read_1_data_T_535; // @[Mux.scala 27:73]
  wire [1:0] _io_read_1_data_T_543 = _io_read_1_data_T_542 | _io_read_1_data_T_536; // @[Mux.scala 27:73]
  wire [1:0] _io_read_1_data_T_544 = _io_read_1_data_T_543 | _io_read_1_data_T_537; // @[Mux.scala 27:73]
  wire [1:0] _io_read_1_data_T_545 = _io_read_1_data_T_544 | _io_read_1_data_T_538; // @[Mux.scala 27:73]
  wire [1:0] _io_read_1_data_T_546 = _io_read_1_data_T_545 | _io_read_1_data_T_539; // @[Mux.scala 27:73]
  wire [19:0] _io_read_1_data_T_653 = io_read_1_addr[0] ? payload_0_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _io_read_1_data_T_654 = io_read_1_addr[1] ? payload_1_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _io_read_1_data_T_655 = io_read_1_addr[2] ? payload_2_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _io_read_1_data_T_656 = io_read_1_addr[3] ? payload_3_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _io_read_1_data_T_657 = io_read_1_addr[4] ? payload_4_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _io_read_1_data_T_658 = io_read_1_addr[5] ? payload_5_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _io_read_1_data_T_659 = io_read_1_addr[6] ? payload_6_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _io_read_1_data_T_660 = io_read_1_addr[7] ? payload_7_ctrl_imm : 20'h0; // @[Mux.scala 27:73]
  wire [19:0] _io_read_1_data_T_661 = _io_read_1_data_T_653 | _io_read_1_data_T_654; // @[Mux.scala 27:73]
  wire [19:0] _io_read_1_data_T_662 = _io_read_1_data_T_661 | _io_read_1_data_T_655; // @[Mux.scala 27:73]
  wire [19:0] _io_read_1_data_T_663 = _io_read_1_data_T_662 | _io_read_1_data_T_656; // @[Mux.scala 27:73]
  wire [19:0] _io_read_1_data_T_664 = _io_read_1_data_T_663 | _io_read_1_data_T_657; // @[Mux.scala 27:73]
  wire [19:0] _io_read_1_data_T_665 = _io_read_1_data_T_664 | _io_read_1_data_T_658; // @[Mux.scala 27:73]
  wire [19:0] _io_read_1_data_T_666 = _io_read_1_data_T_665 | _io_read_1_data_T_659; // @[Mux.scala 27:73]
  wire [6:0] _io_read_1_data_T_773 = io_read_1_addr[0] ? payload_0_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _io_read_1_data_T_774 = io_read_1_addr[1] ? payload_1_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _io_read_1_data_T_775 = io_read_1_addr[2] ? payload_2_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _io_read_1_data_T_776 = io_read_1_addr[3] ? payload_3_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _io_read_1_data_T_777 = io_read_1_addr[4] ? payload_4_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _io_read_1_data_T_778 = io_read_1_addr[5] ? payload_5_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _io_read_1_data_T_779 = io_read_1_addr[6] ? payload_6_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _io_read_1_data_T_780 = io_read_1_addr[7] ? payload_7_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _io_read_1_data_T_781 = _io_read_1_data_T_773 | _io_read_1_data_T_774; // @[Mux.scala 27:73]
  wire [6:0] _io_read_1_data_T_782 = _io_read_1_data_T_781 | _io_read_1_data_T_775; // @[Mux.scala 27:73]
  wire [6:0] _io_read_1_data_T_783 = _io_read_1_data_T_782 | _io_read_1_data_T_776; // @[Mux.scala 27:73]
  wire [6:0] _io_read_1_data_T_784 = _io_read_1_data_T_783 | _io_read_1_data_T_777; // @[Mux.scala 27:73]
  wire [6:0] _io_read_1_data_T_785 = _io_read_1_data_T_784 | _io_read_1_data_T_778; // @[Mux.scala 27:73]
  wire [6:0] _io_read_1_data_T_786 = _io_read_1_data_T_785 | _io_read_1_data_T_779; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_788 = io_read_1_addr[0] ? payload_0_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_789 = io_read_1_addr[1] ? payload_1_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_790 = io_read_1_addr[2] ? payload_2_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_791 = io_read_1_addr[3] ? payload_3_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_792 = io_read_1_addr[4] ? payload_4_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_793 = io_read_1_addr[5] ? payload_5_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_794 = io_read_1_addr[6] ? payload_6_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_795 = io_read_1_addr[7] ? payload_7_ctrl_fuType : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_796 = _io_read_1_data_T_788 | _io_read_1_data_T_789; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_797 = _io_read_1_data_T_796 | _io_read_1_data_T_790; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_798 = _io_read_1_data_T_797 | _io_read_1_data_T_791; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_799 = _io_read_1_data_T_798 | _io_read_1_data_T_792; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_800 = _io_read_1_data_T_799 | _io_read_1_data_T_793; // @[Mux.scala 27:73]
  wire [3:0] _io_read_1_data_T_801 = _io_read_1_data_T_800 | _io_read_1_data_T_794; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_923 = io_read_1_addr[0] ? payload_0_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_924 = io_read_1_addr[1] ? payload_1_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_925 = io_read_1_addr[2] ? payload_2_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_926 = io_read_1_addr[3] ? payload_3_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_927 = io_read_1_addr[4] ? payload_4_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_928 = io_read_1_addr[5] ? payload_5_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_929 = io_read_1_addr[6] ? payload_6_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_930 = io_read_1_addr[7] ? payload_7_cf_ftqOffset : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_931 = _io_read_1_data_T_923 | _io_read_1_data_T_924; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_932 = _io_read_1_data_T_931 | _io_read_1_data_T_925; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_933 = _io_read_1_data_T_932 | _io_read_1_data_T_926; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_934 = _io_read_1_data_T_933 | _io_read_1_data_T_927; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_935 = _io_read_1_data_T_934 | _io_read_1_data_T_928; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_936 = _io_read_1_data_T_935 | _io_read_1_data_T_929; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_938 = io_read_1_addr[0] ? payload_0_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_939 = io_read_1_addr[1] ? payload_1_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_940 = io_read_1_addr[2] ? payload_2_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_941 = io_read_1_addr[3] ? payload_3_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_942 = io_read_1_addr[4] ? payload_4_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_943 = io_read_1_addr[5] ? payload_5_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_944 = io_read_1_addr[6] ? payload_6_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_945 = io_read_1_addr[7] ? payload_7_cf_ftqPtr_value : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_946 = _io_read_1_data_T_938 | _io_read_1_data_T_939; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_947 = _io_read_1_data_T_946 | _io_read_1_data_T_940; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_948 = _io_read_1_data_T_947 | _io_read_1_data_T_941; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_949 = _io_read_1_data_T_948 | _io_read_1_data_T_942; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_950 = _io_read_1_data_T_949 | _io_read_1_data_T_943; // @[Mux.scala 27:73]
  wire [2:0] _io_read_1_data_T_951 = _io_read_1_data_T_950 | _io_read_1_data_T_944; // @[Mux.scala 27:73]
  wire [1:0] _io_read_1_data_T_1118 = io_read_1_addr[0] ? payload_0_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_1_data_T_1119 = io_read_1_addr[1] ? payload_1_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_1_data_T_1120 = io_read_1_addr[2] ? payload_2_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_1_data_T_1121 = io_read_1_addr[3] ? payload_3_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_1_data_T_1122 = io_read_1_addr[4] ? payload_4_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_1_data_T_1123 = io_read_1_addr[5] ? payload_5_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_1_data_T_1124 = io_read_1_addr[6] ? payload_6_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_1_data_T_1125 = io_read_1_addr[7] ? payload_7_cf_pd_brType : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_read_1_data_T_1126 = _io_read_1_data_T_1118 | _io_read_1_data_T_1119; // @[Mux.scala 27:73]
  wire [1:0] _io_read_1_data_T_1127 = _io_read_1_data_T_1126 | _io_read_1_data_T_1120; // @[Mux.scala 27:73]
  wire [1:0] _io_read_1_data_T_1128 = _io_read_1_data_T_1127 | _io_read_1_data_T_1121; // @[Mux.scala 27:73]
  wire [1:0] _io_read_1_data_T_1129 = _io_read_1_data_T_1128 | _io_read_1_data_T_1122; // @[Mux.scala 27:73]
  wire [1:0] _io_read_1_data_T_1130 = _io_read_1_data_T_1129 | _io_read_1_data_T_1123; // @[Mux.scala 27:73]
  wire [1:0] _io_read_1_data_T_1131 = _io_read_1_data_T_1130 | _io_read_1_data_T_1124; // @[Mux.scala 27:73]
  wire  wenVec_0 = io_write_0_enable & io_write_0_addr[0]; // @[PayloadArray.scala 55:53]
  wire  wen = |wenVec_0; // @[PayloadArray.scala 56:29]
  wire  wenVec_1_0 = io_write_0_enable & io_write_0_addr[1]; // @[PayloadArray.scala 55:53]
  wire  wen_1 = |wenVec_1_0; // @[PayloadArray.scala 56:29]
  wire  wenVec_2_0 = io_write_0_enable & io_write_0_addr[2]; // @[PayloadArray.scala 55:53]
  wire  wen_2 = |wenVec_2_0; // @[PayloadArray.scala 56:29]
  wire  wenVec_3_0 = io_write_0_enable & io_write_0_addr[3]; // @[PayloadArray.scala 55:53]
  wire  wen_3 = |wenVec_3_0; // @[PayloadArray.scala 56:29]
  wire  wenVec_4_0 = io_write_0_enable & io_write_0_addr[4]; // @[PayloadArray.scala 55:53]
  wire  wen_4 = |wenVec_4_0; // @[PayloadArray.scala 56:29]
  wire  wenVec_5_0 = io_write_0_enable & io_write_0_addr[5]; // @[PayloadArray.scala 55:53]
  wire  wen_5 = |wenVec_5_0; // @[PayloadArray.scala 56:29]
  wire  wenVec_6_0 = io_write_0_enable & io_write_0_addr[6]; // @[PayloadArray.scala 55:53]
  wire  wen_6 = |wenVec_6_0; // @[PayloadArray.scala 56:29]
  wire  wenVec_7_0 = io_write_0_enable & io_write_0_addr[7]; // @[PayloadArray.scala 55:53]
  wire  wen_7 = |wenVec_7_0; // @[PayloadArray.scala 56:29]
  assign io_read_0_data_cf_pd_isRVC = io_read_0_addr[0] & payload_0_cf_pd_isRVC | io_read_0_addr[1] &
    payload_1_cf_pd_isRVC | io_read_0_addr[2] & payload_2_cf_pd_isRVC | io_read_0_addr[3] & payload_3_cf_pd_isRVC |
    io_read_0_addr[4] & payload_4_cf_pd_isRVC | io_read_0_addr[5] & payload_5_cf_pd_isRVC | io_read_0_addr[6] &
    payload_6_cf_pd_isRVC | io_read_0_addr[7] & payload_7_cf_pd_isRVC; // @[Mux.scala 27:73]
  assign io_read_0_data_cf_pd_brType = _io_read_0_data_T_1131 | _io_read_0_data_T_1125; // @[Mux.scala 27:73]
  assign io_read_0_data_cf_pd_isCall = io_read_0_addr[0] & payload_0_cf_pd_isCall | io_read_0_addr[1] &
    payload_1_cf_pd_isCall | io_read_0_addr[2] & payload_2_cf_pd_isCall | io_read_0_addr[3] & payload_3_cf_pd_isCall |
    io_read_0_addr[4] & payload_4_cf_pd_isCall | io_read_0_addr[5] & payload_5_cf_pd_isCall | io_read_0_addr[6] &
    payload_6_cf_pd_isCall | io_read_0_addr[7] & payload_7_cf_pd_isCall; // @[Mux.scala 27:73]
  assign io_read_0_data_cf_pd_isRet = io_read_0_addr[0] & payload_0_cf_pd_isRet | io_read_0_addr[1] &
    payload_1_cf_pd_isRet | io_read_0_addr[2] & payload_2_cf_pd_isRet | io_read_0_addr[3] & payload_3_cf_pd_isRet |
    io_read_0_addr[4] & payload_4_cf_pd_isRet | io_read_0_addr[5] & payload_5_cf_pd_isRet | io_read_0_addr[6] &
    payload_6_cf_pd_isRet | io_read_0_addr[7] & payload_7_cf_pd_isRet; // @[Mux.scala 27:73]
  assign io_read_0_data_cf_pred_taken = io_read_0_addr[0] & payload_0_cf_pred_taken | io_read_0_addr[1] &
    payload_1_cf_pred_taken | io_read_0_addr[2] & payload_2_cf_pred_taken | io_read_0_addr[3] & payload_3_cf_pred_taken
     | io_read_0_addr[4] & payload_4_cf_pred_taken | io_read_0_addr[5] & payload_5_cf_pred_taken | io_read_0_addr[6] &
    payload_6_cf_pred_taken | io_read_0_addr[7] & payload_7_cf_pred_taken; // @[Mux.scala 27:73]
  assign io_read_0_data_cf_ftqPtr_flag = io_read_0_addr[0] & payload_0_cf_ftqPtr_flag | io_read_0_addr[1] &
    payload_1_cf_ftqPtr_flag | io_read_0_addr[2] & payload_2_cf_ftqPtr_flag | io_read_0_addr[3] &
    payload_3_cf_ftqPtr_flag | io_read_0_addr[4] & payload_4_cf_ftqPtr_flag | io_read_0_addr[5] &
    payload_5_cf_ftqPtr_flag | io_read_0_addr[6] & payload_6_cf_ftqPtr_flag | io_read_0_addr[7] &
    payload_7_cf_ftqPtr_flag; // @[Mux.scala 27:73]
  assign io_read_0_data_cf_ftqPtr_value = _io_read_0_data_T_951 | _io_read_0_data_T_945; // @[Mux.scala 27:73]
  assign io_read_0_data_cf_ftqOffset = _io_read_0_data_T_936 | _io_read_0_data_T_930; // @[Mux.scala 27:73]
  assign io_read_0_data_ctrl_fuType = _io_read_0_data_T_801 | _io_read_0_data_T_795; // @[Mux.scala 27:73]
  assign io_read_0_data_ctrl_fuOpType = _io_read_0_data_T_786 | _io_read_0_data_T_780; // @[Mux.scala 27:73]
  assign io_read_0_data_ctrl_rfWen = io_read_0_addr[0] & payload_0_ctrl_rfWen | io_read_0_addr[1] & payload_1_ctrl_rfWen
     | io_read_0_addr[2] & payload_2_ctrl_rfWen | io_read_0_addr[3] & payload_3_ctrl_rfWen | io_read_0_addr[4] &
    payload_4_ctrl_rfWen | io_read_0_addr[5] & payload_5_ctrl_rfWen | io_read_0_addr[6] & payload_6_ctrl_rfWen |
    io_read_0_addr[7] & payload_7_ctrl_rfWen; // @[Mux.scala 27:73]
  assign io_read_0_data_ctrl_fpWen = io_read_0_addr[0] & payload_0_ctrl_fpWen | io_read_0_addr[1] & payload_1_ctrl_fpWen
     | io_read_0_addr[2] & payload_2_ctrl_fpWen | io_read_0_addr[3] & payload_3_ctrl_fpWen | io_read_0_addr[4] &
    payload_4_ctrl_fpWen | io_read_0_addr[5] & payload_5_ctrl_fpWen | io_read_0_addr[6] & payload_6_ctrl_fpWen |
    io_read_0_addr[7] & payload_7_ctrl_fpWen; // @[Mux.scala 27:73]
  assign io_read_0_data_ctrl_imm = _io_read_0_data_T_666 | _io_read_0_data_T_660; // @[Mux.scala 27:73]
  assign io_read_0_data_ctrl_fpu_isAddSub = io_read_0_addr[0] & payload_0_ctrl_fpu_isAddSub | io_read_0_addr[1] &
    payload_1_ctrl_fpu_isAddSub | io_read_0_addr[2] & payload_2_ctrl_fpu_isAddSub | io_read_0_addr[3] &
    payload_3_ctrl_fpu_isAddSub | io_read_0_addr[4] & payload_4_ctrl_fpu_isAddSub | io_read_0_addr[5] &
    payload_5_ctrl_fpu_isAddSub | io_read_0_addr[6] & payload_6_ctrl_fpu_isAddSub | io_read_0_addr[7] &
    payload_7_ctrl_fpu_isAddSub; // @[Mux.scala 27:73]
  assign io_read_0_data_ctrl_fpu_typeTagIn = io_read_0_addr[0] & payload_0_ctrl_fpu_typeTagIn | io_read_0_addr[1] &
    payload_1_ctrl_fpu_typeTagIn | io_read_0_addr[2] & payload_2_ctrl_fpu_typeTagIn | io_read_0_addr[3] &
    payload_3_ctrl_fpu_typeTagIn | io_read_0_addr[4] & payload_4_ctrl_fpu_typeTagIn | io_read_0_addr[5] &
    payload_5_ctrl_fpu_typeTagIn | io_read_0_addr[6] & payload_6_ctrl_fpu_typeTagIn | io_read_0_addr[7] &
    payload_7_ctrl_fpu_typeTagIn; // @[Mux.scala 27:73]
  assign io_read_0_data_ctrl_fpu_typeTagOut = io_read_0_addr[0] & payload_0_ctrl_fpu_typeTagOut | io_read_0_addr[1] &
    payload_1_ctrl_fpu_typeTagOut | io_read_0_addr[2] & payload_2_ctrl_fpu_typeTagOut | io_read_0_addr[3] &
    payload_3_ctrl_fpu_typeTagOut | io_read_0_addr[4] & payload_4_ctrl_fpu_typeTagOut | io_read_0_addr[5] &
    payload_5_ctrl_fpu_typeTagOut | io_read_0_addr[6] & payload_6_ctrl_fpu_typeTagOut | io_read_0_addr[7] &
    payload_7_ctrl_fpu_typeTagOut; // @[Mux.scala 27:73]
  assign io_read_0_data_ctrl_fpu_fromInt = io_read_0_addr[0] & payload_0_ctrl_fpu_fromInt | io_read_0_addr[1] &
    payload_1_ctrl_fpu_fromInt | io_read_0_addr[2] & payload_2_ctrl_fpu_fromInt | io_read_0_addr[3] &
    payload_3_ctrl_fpu_fromInt | io_read_0_addr[4] & payload_4_ctrl_fpu_fromInt | io_read_0_addr[5] &
    payload_5_ctrl_fpu_fromInt | io_read_0_addr[6] & payload_6_ctrl_fpu_fromInt | io_read_0_addr[7] &
    payload_7_ctrl_fpu_fromInt; // @[Mux.scala 27:73]
  assign io_read_0_data_ctrl_fpu_wflags = io_read_0_addr[0] & payload_0_ctrl_fpu_wflags | io_read_0_addr[1] &
    payload_1_ctrl_fpu_wflags | io_read_0_addr[2] & payload_2_ctrl_fpu_wflags | io_read_0_addr[3] &
    payload_3_ctrl_fpu_wflags | io_read_0_addr[4] & payload_4_ctrl_fpu_wflags | io_read_0_addr[5] &
    payload_5_ctrl_fpu_wflags | io_read_0_addr[6] & payload_6_ctrl_fpu_wflags | io_read_0_addr[7] &
    payload_7_ctrl_fpu_wflags; // @[Mux.scala 27:73]
  assign io_read_0_data_ctrl_fpu_fpWen = io_read_0_addr[0] & payload_0_ctrl_fpu_fpWen | io_read_0_addr[1] &
    payload_1_ctrl_fpu_fpWen | io_read_0_addr[2] & payload_2_ctrl_fpu_fpWen | io_read_0_addr[3] &
    payload_3_ctrl_fpu_fpWen | io_read_0_addr[4] & payload_4_ctrl_fpu_fpWen | io_read_0_addr[5] &
    payload_5_ctrl_fpu_fpWen | io_read_0_addr[6] & payload_6_ctrl_fpu_fpWen | io_read_0_addr[7] &
    payload_7_ctrl_fpu_fpWen; // @[Mux.scala 27:73]
  assign io_read_0_data_ctrl_fpu_fmaCmd = _io_read_0_data_T_546 | _io_read_0_data_T_540; // @[Mux.scala 27:73]
  assign io_read_0_data_ctrl_fpu_div = io_read_0_addr[0] & payload_0_ctrl_fpu_div | io_read_0_addr[1] &
    payload_1_ctrl_fpu_div | io_read_0_addr[2] & payload_2_ctrl_fpu_div | io_read_0_addr[3] & payload_3_ctrl_fpu_div |
    io_read_0_addr[4] & payload_4_ctrl_fpu_div | io_read_0_addr[5] & payload_5_ctrl_fpu_div | io_read_0_addr[6] &
    payload_6_ctrl_fpu_div | io_read_0_addr[7] & payload_7_ctrl_fpu_div; // @[Mux.scala 27:73]
  assign io_read_0_data_ctrl_fpu_sqrt = io_read_0_addr[0] & payload_0_ctrl_fpu_sqrt | io_read_0_addr[1] &
    payload_1_ctrl_fpu_sqrt | io_read_0_addr[2] & payload_2_ctrl_fpu_sqrt | io_read_0_addr[3] & payload_3_ctrl_fpu_sqrt
     | io_read_0_addr[4] & payload_4_ctrl_fpu_sqrt | io_read_0_addr[5] & payload_5_ctrl_fpu_sqrt | io_read_0_addr[6] &
    payload_6_ctrl_fpu_sqrt | io_read_0_addr[7] & payload_7_ctrl_fpu_sqrt; // @[Mux.scala 27:73]
  assign io_read_0_data_ctrl_fpu_fcvt = io_read_0_addr[0] & payload_0_ctrl_fpu_fcvt | io_read_0_addr[1] &
    payload_1_ctrl_fpu_fcvt | io_read_0_addr[2] & payload_2_ctrl_fpu_fcvt | io_read_0_addr[3] & payload_3_ctrl_fpu_fcvt
     | io_read_0_addr[4] & payload_4_ctrl_fpu_fcvt | io_read_0_addr[5] & payload_5_ctrl_fpu_fcvt | io_read_0_addr[6] &
    payload_6_ctrl_fpu_fcvt | io_read_0_addr[7] & payload_7_ctrl_fpu_fcvt; // @[Mux.scala 27:73]
  assign io_read_0_data_ctrl_fpu_typ = _io_read_0_data_T_486 | _io_read_0_data_T_480; // @[Mux.scala 27:73]
  assign io_read_0_data_ctrl_fpu_fmt = _io_read_0_data_T_471 | _io_read_0_data_T_465; // @[Mux.scala 27:73]
  assign io_read_0_data_ctrl_fpu_ren3 = io_read_0_addr[0] & payload_0_ctrl_fpu_ren3 | io_read_0_addr[1] &
    payload_1_ctrl_fpu_ren3 | io_read_0_addr[2] & payload_2_ctrl_fpu_ren3 | io_read_0_addr[3] & payload_3_ctrl_fpu_ren3
     | io_read_0_addr[4] & payload_4_ctrl_fpu_ren3 | io_read_0_addr[5] & payload_5_ctrl_fpu_ren3 | io_read_0_addr[6] &
    payload_6_ctrl_fpu_ren3 | io_read_0_addr[7] & payload_7_ctrl_fpu_ren3; // @[Mux.scala 27:73]
  assign io_read_0_data_ctrl_fpu_rm = _io_read_0_data_T_441 | _io_read_0_data_T_435; // @[Mux.scala 27:73]
  assign io_read_0_data_pdest = _io_read_0_data_T_291 | _io_read_0_data_T_285; // @[Mux.scala 27:73]
  assign io_read_0_data_robIdx_flag = io_read_0_addr[0] & payload_0_robIdx_flag | io_read_0_addr[1] &
    payload_1_robIdx_flag | io_read_0_addr[2] & payload_2_robIdx_flag | io_read_0_addr[3] & payload_3_robIdx_flag |
    io_read_0_addr[4] & payload_4_robIdx_flag | io_read_0_addr[5] & payload_5_robIdx_flag | io_read_0_addr[6] &
    payload_6_robIdx_flag | io_read_0_addr[7] & payload_7_robIdx_flag; // @[Mux.scala 27:73]
  assign io_read_0_data_robIdx_value = _io_read_0_data_T_246 | _io_read_0_data_T_240; // @[Mux.scala 27:73]
  assign io_read_1_data_cf_pd_isRVC = io_read_1_addr[0] & payload_0_cf_pd_isRVC | io_read_1_addr[1] &
    payload_1_cf_pd_isRVC | io_read_1_addr[2] & payload_2_cf_pd_isRVC | io_read_1_addr[3] & payload_3_cf_pd_isRVC |
    io_read_1_addr[4] & payload_4_cf_pd_isRVC | io_read_1_addr[5] & payload_5_cf_pd_isRVC | io_read_1_addr[6] &
    payload_6_cf_pd_isRVC | io_read_1_addr[7] & payload_7_cf_pd_isRVC; // @[Mux.scala 27:73]
  assign io_read_1_data_cf_pd_brType = _io_read_1_data_T_1131 | _io_read_1_data_T_1125; // @[Mux.scala 27:73]
  assign io_read_1_data_cf_pd_isCall = io_read_1_addr[0] & payload_0_cf_pd_isCall | io_read_1_addr[1] &
    payload_1_cf_pd_isCall | io_read_1_addr[2] & payload_2_cf_pd_isCall | io_read_1_addr[3] & payload_3_cf_pd_isCall |
    io_read_1_addr[4] & payload_4_cf_pd_isCall | io_read_1_addr[5] & payload_5_cf_pd_isCall | io_read_1_addr[6] &
    payload_6_cf_pd_isCall | io_read_1_addr[7] & payload_7_cf_pd_isCall; // @[Mux.scala 27:73]
  assign io_read_1_data_cf_pd_isRet = io_read_1_addr[0] & payload_0_cf_pd_isRet | io_read_1_addr[1] &
    payload_1_cf_pd_isRet | io_read_1_addr[2] & payload_2_cf_pd_isRet | io_read_1_addr[3] & payload_3_cf_pd_isRet |
    io_read_1_addr[4] & payload_4_cf_pd_isRet | io_read_1_addr[5] & payload_5_cf_pd_isRet | io_read_1_addr[6] &
    payload_6_cf_pd_isRet | io_read_1_addr[7] & payload_7_cf_pd_isRet; // @[Mux.scala 27:73]
  assign io_read_1_data_cf_pred_taken = io_read_1_addr[0] & payload_0_cf_pred_taken | io_read_1_addr[1] &
    payload_1_cf_pred_taken | io_read_1_addr[2] & payload_2_cf_pred_taken | io_read_1_addr[3] & payload_3_cf_pred_taken
     | io_read_1_addr[4] & payload_4_cf_pred_taken | io_read_1_addr[5] & payload_5_cf_pred_taken | io_read_1_addr[6] &
    payload_6_cf_pred_taken | io_read_1_addr[7] & payload_7_cf_pred_taken; // @[Mux.scala 27:73]
  assign io_read_1_data_cf_ftqPtr_flag = io_read_1_addr[0] & payload_0_cf_ftqPtr_flag | io_read_1_addr[1] &
    payload_1_cf_ftqPtr_flag | io_read_1_addr[2] & payload_2_cf_ftqPtr_flag | io_read_1_addr[3] &
    payload_3_cf_ftqPtr_flag | io_read_1_addr[4] & payload_4_cf_ftqPtr_flag | io_read_1_addr[5] &
    payload_5_cf_ftqPtr_flag | io_read_1_addr[6] & payload_6_cf_ftqPtr_flag | io_read_1_addr[7] &
    payload_7_cf_ftqPtr_flag; // @[Mux.scala 27:73]
  assign io_read_1_data_cf_ftqPtr_value = _io_read_1_data_T_951 | _io_read_1_data_T_945; // @[Mux.scala 27:73]
  assign io_read_1_data_cf_ftqOffset = _io_read_1_data_T_936 | _io_read_1_data_T_930; // @[Mux.scala 27:73]
  assign io_read_1_data_ctrl_fuType = _io_read_1_data_T_801 | _io_read_1_data_T_795; // @[Mux.scala 27:73]
  assign io_read_1_data_ctrl_fuOpType = _io_read_1_data_T_786 | _io_read_1_data_T_780; // @[Mux.scala 27:73]
  assign io_read_1_data_ctrl_rfWen = io_read_1_addr[0] & payload_0_ctrl_rfWen | io_read_1_addr[1] & payload_1_ctrl_rfWen
     | io_read_1_addr[2] & payload_2_ctrl_rfWen | io_read_1_addr[3] & payload_3_ctrl_rfWen | io_read_1_addr[4] &
    payload_4_ctrl_rfWen | io_read_1_addr[5] & payload_5_ctrl_rfWen | io_read_1_addr[6] & payload_6_ctrl_rfWen |
    io_read_1_addr[7] & payload_7_ctrl_rfWen; // @[Mux.scala 27:73]
  assign io_read_1_data_ctrl_fpWen = io_read_1_addr[0] & payload_0_ctrl_fpWen | io_read_1_addr[1] & payload_1_ctrl_fpWen
     | io_read_1_addr[2] & payload_2_ctrl_fpWen | io_read_1_addr[3] & payload_3_ctrl_fpWen | io_read_1_addr[4] &
    payload_4_ctrl_fpWen | io_read_1_addr[5] & payload_5_ctrl_fpWen | io_read_1_addr[6] & payload_6_ctrl_fpWen |
    io_read_1_addr[7] & payload_7_ctrl_fpWen; // @[Mux.scala 27:73]
  assign io_read_1_data_ctrl_imm = _io_read_1_data_T_666 | _io_read_1_data_T_660; // @[Mux.scala 27:73]
  assign io_read_1_data_ctrl_fpu_isAddSub = io_read_1_addr[0] & payload_0_ctrl_fpu_isAddSub | io_read_1_addr[1] &
    payload_1_ctrl_fpu_isAddSub | io_read_1_addr[2] & payload_2_ctrl_fpu_isAddSub | io_read_1_addr[3] &
    payload_3_ctrl_fpu_isAddSub | io_read_1_addr[4] & payload_4_ctrl_fpu_isAddSub | io_read_1_addr[5] &
    payload_5_ctrl_fpu_isAddSub | io_read_1_addr[6] & payload_6_ctrl_fpu_isAddSub | io_read_1_addr[7] &
    payload_7_ctrl_fpu_isAddSub; // @[Mux.scala 27:73]
  assign io_read_1_data_ctrl_fpu_typeTagIn = io_read_1_addr[0] & payload_0_ctrl_fpu_typeTagIn | io_read_1_addr[1] &
    payload_1_ctrl_fpu_typeTagIn | io_read_1_addr[2] & payload_2_ctrl_fpu_typeTagIn | io_read_1_addr[3] &
    payload_3_ctrl_fpu_typeTagIn | io_read_1_addr[4] & payload_4_ctrl_fpu_typeTagIn | io_read_1_addr[5] &
    payload_5_ctrl_fpu_typeTagIn | io_read_1_addr[6] & payload_6_ctrl_fpu_typeTagIn | io_read_1_addr[7] &
    payload_7_ctrl_fpu_typeTagIn; // @[Mux.scala 27:73]
  assign io_read_1_data_ctrl_fpu_typeTagOut = io_read_1_addr[0] & payload_0_ctrl_fpu_typeTagOut | io_read_1_addr[1] &
    payload_1_ctrl_fpu_typeTagOut | io_read_1_addr[2] & payload_2_ctrl_fpu_typeTagOut | io_read_1_addr[3] &
    payload_3_ctrl_fpu_typeTagOut | io_read_1_addr[4] & payload_4_ctrl_fpu_typeTagOut | io_read_1_addr[5] &
    payload_5_ctrl_fpu_typeTagOut | io_read_1_addr[6] & payload_6_ctrl_fpu_typeTagOut | io_read_1_addr[7] &
    payload_7_ctrl_fpu_typeTagOut; // @[Mux.scala 27:73]
  assign io_read_1_data_ctrl_fpu_fromInt = io_read_1_addr[0] & payload_0_ctrl_fpu_fromInt | io_read_1_addr[1] &
    payload_1_ctrl_fpu_fromInt | io_read_1_addr[2] & payload_2_ctrl_fpu_fromInt | io_read_1_addr[3] &
    payload_3_ctrl_fpu_fromInt | io_read_1_addr[4] & payload_4_ctrl_fpu_fromInt | io_read_1_addr[5] &
    payload_5_ctrl_fpu_fromInt | io_read_1_addr[6] & payload_6_ctrl_fpu_fromInt | io_read_1_addr[7] &
    payload_7_ctrl_fpu_fromInt; // @[Mux.scala 27:73]
  assign io_read_1_data_ctrl_fpu_wflags = io_read_1_addr[0] & payload_0_ctrl_fpu_wflags | io_read_1_addr[1] &
    payload_1_ctrl_fpu_wflags | io_read_1_addr[2] & payload_2_ctrl_fpu_wflags | io_read_1_addr[3] &
    payload_3_ctrl_fpu_wflags | io_read_1_addr[4] & payload_4_ctrl_fpu_wflags | io_read_1_addr[5] &
    payload_5_ctrl_fpu_wflags | io_read_1_addr[6] & payload_6_ctrl_fpu_wflags | io_read_1_addr[7] &
    payload_7_ctrl_fpu_wflags; // @[Mux.scala 27:73]
  assign io_read_1_data_ctrl_fpu_fpWen = io_read_1_addr[0] & payload_0_ctrl_fpu_fpWen | io_read_1_addr[1] &
    payload_1_ctrl_fpu_fpWen | io_read_1_addr[2] & payload_2_ctrl_fpu_fpWen | io_read_1_addr[3] &
    payload_3_ctrl_fpu_fpWen | io_read_1_addr[4] & payload_4_ctrl_fpu_fpWen | io_read_1_addr[5] &
    payload_5_ctrl_fpu_fpWen | io_read_1_addr[6] & payload_6_ctrl_fpu_fpWen | io_read_1_addr[7] &
    payload_7_ctrl_fpu_fpWen; // @[Mux.scala 27:73]
  assign io_read_1_data_ctrl_fpu_fmaCmd = _io_read_1_data_T_546 | _io_read_1_data_T_540; // @[Mux.scala 27:73]
  assign io_read_1_data_ctrl_fpu_div = io_read_1_addr[0] & payload_0_ctrl_fpu_div | io_read_1_addr[1] &
    payload_1_ctrl_fpu_div | io_read_1_addr[2] & payload_2_ctrl_fpu_div | io_read_1_addr[3] & payload_3_ctrl_fpu_div |
    io_read_1_addr[4] & payload_4_ctrl_fpu_div | io_read_1_addr[5] & payload_5_ctrl_fpu_div | io_read_1_addr[6] &
    payload_6_ctrl_fpu_div | io_read_1_addr[7] & payload_7_ctrl_fpu_div; // @[Mux.scala 27:73]
  assign io_read_1_data_ctrl_fpu_sqrt = io_read_1_addr[0] & payload_0_ctrl_fpu_sqrt | io_read_1_addr[1] &
    payload_1_ctrl_fpu_sqrt | io_read_1_addr[2] & payload_2_ctrl_fpu_sqrt | io_read_1_addr[3] & payload_3_ctrl_fpu_sqrt
     | io_read_1_addr[4] & payload_4_ctrl_fpu_sqrt | io_read_1_addr[5] & payload_5_ctrl_fpu_sqrt | io_read_1_addr[6] &
    payload_6_ctrl_fpu_sqrt | io_read_1_addr[7] & payload_7_ctrl_fpu_sqrt; // @[Mux.scala 27:73]
  assign io_read_1_data_ctrl_fpu_fcvt = io_read_1_addr[0] & payload_0_ctrl_fpu_fcvt | io_read_1_addr[1] &
    payload_1_ctrl_fpu_fcvt | io_read_1_addr[2] & payload_2_ctrl_fpu_fcvt | io_read_1_addr[3] & payload_3_ctrl_fpu_fcvt
     | io_read_1_addr[4] & payload_4_ctrl_fpu_fcvt | io_read_1_addr[5] & payload_5_ctrl_fpu_fcvt | io_read_1_addr[6] &
    payload_6_ctrl_fpu_fcvt | io_read_1_addr[7] & payload_7_ctrl_fpu_fcvt; // @[Mux.scala 27:73]
  assign io_read_1_data_ctrl_fpu_typ = _io_read_1_data_T_486 | _io_read_1_data_T_480; // @[Mux.scala 27:73]
  assign io_read_1_data_ctrl_fpu_fmt = _io_read_1_data_T_471 | _io_read_1_data_T_465; // @[Mux.scala 27:73]
  assign io_read_1_data_ctrl_fpu_ren3 = io_read_1_addr[0] & payload_0_ctrl_fpu_ren3 | io_read_1_addr[1] &
    payload_1_ctrl_fpu_ren3 | io_read_1_addr[2] & payload_2_ctrl_fpu_ren3 | io_read_1_addr[3] & payload_3_ctrl_fpu_ren3
     | io_read_1_addr[4] & payload_4_ctrl_fpu_ren3 | io_read_1_addr[5] & payload_5_ctrl_fpu_ren3 | io_read_1_addr[6] &
    payload_6_ctrl_fpu_ren3 | io_read_1_addr[7] & payload_7_ctrl_fpu_ren3; // @[Mux.scala 27:73]
  assign io_read_1_data_ctrl_fpu_rm = _io_read_1_data_T_441 | _io_read_1_data_T_435; // @[Mux.scala 27:73]
  assign io_read_1_data_pdest = _io_read_1_data_T_291 | _io_read_1_data_T_285; // @[Mux.scala 27:73]
  assign io_read_1_data_robIdx_flag = io_read_1_addr[0] & payload_0_robIdx_flag | io_read_1_addr[1] &
    payload_1_robIdx_flag | io_read_1_addr[2] & payload_2_robIdx_flag | io_read_1_addr[3] & payload_3_robIdx_flag |
    io_read_1_addr[4] & payload_4_robIdx_flag | io_read_1_addr[5] & payload_5_robIdx_flag | io_read_1_addr[6] &
    payload_6_robIdx_flag | io_read_1_addr[7] & payload_7_robIdx_flag; // @[Mux.scala 27:73]
  assign io_read_1_data_robIdx_value = _io_read_1_data_T_246 | _io_read_1_data_T_240; // @[Mux.scala 27:73]
  always @(posedge clock) begin
    if (wen) begin // @[PayloadArray.scala 58:16]
      payload_0_cf_pd_isRVC <= io_write_0_data_cf_pd_isRVC; // @[PayloadArray.scala 59:18]
    end
    if (wen) begin // @[PayloadArray.scala 58:16]
      payload_0_cf_pd_brType <= io_write_0_data_cf_pd_brType; // @[PayloadArray.scala 59:18]
    end
    if (wen) begin // @[PayloadArray.scala 58:16]
      payload_0_cf_pd_isCall <= io_write_0_data_cf_pd_isCall; // @[PayloadArray.scala 59:18]
    end
    if (wen) begin // @[PayloadArray.scala 58:16]
      payload_0_cf_pd_isRet <= io_write_0_data_cf_pd_isRet; // @[PayloadArray.scala 59:18]
    end
    if (wen) begin // @[PayloadArray.scala 58:16]
      payload_0_cf_pred_taken <= io_write_0_data_cf_pred_taken; // @[PayloadArray.scala 59:18]
    end
    if (wen) begin // @[PayloadArray.scala 58:16]
      payload_0_cf_ftqPtr_flag <= io_write_0_data_cf_ftqPtr_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen) begin // @[PayloadArray.scala 58:16]
      payload_0_cf_ftqPtr_value <= io_write_0_data_cf_ftqPtr_value; // @[PayloadArray.scala 59:18]
    end
    if (wen) begin // @[PayloadArray.scala 58:16]
      payload_0_cf_ftqOffset <= io_write_0_data_cf_ftqOffset; // @[PayloadArray.scala 59:18]
    end
    if (wen) begin // @[PayloadArray.scala 58:16]
      payload_0_ctrl_fuType <= io_write_0_data_ctrl_fuType; // @[PayloadArray.scala 59:18]
    end
    if (wen) begin // @[PayloadArray.scala 58:16]
      payload_0_ctrl_fuOpType <= io_write_0_data_ctrl_fuOpType; // @[PayloadArray.scala 59:18]
    end
    if (wen) begin // @[PayloadArray.scala 58:16]
      payload_0_ctrl_rfWen <= io_write_0_data_ctrl_rfWen; // @[PayloadArray.scala 59:18]
    end
    if (wen) begin // @[PayloadArray.scala 58:16]
      payload_0_ctrl_fpWen <= io_write_0_data_ctrl_fpWen; // @[PayloadArray.scala 59:18]
    end
    if (wen) begin // @[PayloadArray.scala 58:16]
      payload_0_ctrl_imm <= io_write_0_data_ctrl_imm; // @[PayloadArray.scala 59:18]
    end
    if (wen) begin // @[PayloadArray.scala 58:16]
      payload_0_ctrl_fpu_isAddSub <= io_write_0_data_ctrl_fpu_isAddSub; // @[PayloadArray.scala 59:18]
    end
    if (wen) begin // @[PayloadArray.scala 58:16]
      payload_0_ctrl_fpu_typeTagIn <= io_write_0_data_ctrl_fpu_typeTagIn; // @[PayloadArray.scala 59:18]
    end
    if (wen) begin // @[PayloadArray.scala 58:16]
      payload_0_ctrl_fpu_typeTagOut <= io_write_0_data_ctrl_fpu_typeTagOut; // @[PayloadArray.scala 59:18]
    end
    if (wen) begin // @[PayloadArray.scala 58:16]
      payload_0_ctrl_fpu_fromInt <= io_write_0_data_ctrl_fpu_fromInt; // @[PayloadArray.scala 59:18]
    end
    if (wen) begin // @[PayloadArray.scala 58:16]
      payload_0_ctrl_fpu_wflags <= io_write_0_data_ctrl_fpu_wflags; // @[PayloadArray.scala 59:18]
    end
    if (wen) begin // @[PayloadArray.scala 58:16]
      payload_0_ctrl_fpu_fpWen <= io_write_0_data_ctrl_fpu_fpWen; // @[PayloadArray.scala 59:18]
    end
    if (wen) begin // @[PayloadArray.scala 58:16]
      payload_0_ctrl_fpu_fmaCmd <= io_write_0_data_ctrl_fpu_fmaCmd; // @[PayloadArray.scala 59:18]
    end
    if (wen) begin // @[PayloadArray.scala 58:16]
      payload_0_ctrl_fpu_div <= io_write_0_data_ctrl_fpu_div; // @[PayloadArray.scala 59:18]
    end
    if (wen) begin // @[PayloadArray.scala 58:16]
      payload_0_ctrl_fpu_sqrt <= io_write_0_data_ctrl_fpu_sqrt; // @[PayloadArray.scala 59:18]
    end
    if (wen) begin // @[PayloadArray.scala 58:16]
      payload_0_ctrl_fpu_fcvt <= io_write_0_data_ctrl_fpu_fcvt; // @[PayloadArray.scala 59:18]
    end
    if (wen) begin // @[PayloadArray.scala 58:16]
      payload_0_ctrl_fpu_typ <= io_write_0_data_ctrl_fpu_typ; // @[PayloadArray.scala 59:18]
    end
    if (wen) begin // @[PayloadArray.scala 58:16]
      payload_0_ctrl_fpu_fmt <= io_write_0_data_ctrl_fpu_fmt; // @[PayloadArray.scala 59:18]
    end
    if (wen) begin // @[PayloadArray.scala 58:16]
      payload_0_ctrl_fpu_ren3 <= io_write_0_data_ctrl_fpu_ren3; // @[PayloadArray.scala 59:18]
    end
    if (wen) begin // @[PayloadArray.scala 58:16]
      payload_0_ctrl_fpu_rm <= io_write_0_data_ctrl_fpu_rm; // @[PayloadArray.scala 59:18]
    end
    if (wen) begin // @[PayloadArray.scala 58:16]
      payload_0_pdest <= io_write_0_data_pdest; // @[PayloadArray.scala 59:18]
    end
    if (wen) begin // @[PayloadArray.scala 58:16]
      payload_0_robIdx_flag <= io_write_0_data_robIdx_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen) begin // @[PayloadArray.scala 58:16]
      payload_0_robIdx_value <= io_write_0_data_robIdx_value; // @[PayloadArray.scala 59:18]
    end
    if (wen_1) begin // @[PayloadArray.scala 58:16]
      payload_1_cf_pd_isRVC <= io_write_0_data_cf_pd_isRVC; // @[PayloadArray.scala 59:18]
    end
    if (wen_1) begin // @[PayloadArray.scala 58:16]
      payload_1_cf_pd_brType <= io_write_0_data_cf_pd_brType; // @[PayloadArray.scala 59:18]
    end
    if (wen_1) begin // @[PayloadArray.scala 58:16]
      payload_1_cf_pd_isCall <= io_write_0_data_cf_pd_isCall; // @[PayloadArray.scala 59:18]
    end
    if (wen_1) begin // @[PayloadArray.scala 58:16]
      payload_1_cf_pd_isRet <= io_write_0_data_cf_pd_isRet; // @[PayloadArray.scala 59:18]
    end
    if (wen_1) begin // @[PayloadArray.scala 58:16]
      payload_1_cf_pred_taken <= io_write_0_data_cf_pred_taken; // @[PayloadArray.scala 59:18]
    end
    if (wen_1) begin // @[PayloadArray.scala 58:16]
      payload_1_cf_ftqPtr_flag <= io_write_0_data_cf_ftqPtr_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen_1) begin // @[PayloadArray.scala 58:16]
      payload_1_cf_ftqPtr_value <= io_write_0_data_cf_ftqPtr_value; // @[PayloadArray.scala 59:18]
    end
    if (wen_1) begin // @[PayloadArray.scala 58:16]
      payload_1_cf_ftqOffset <= io_write_0_data_cf_ftqOffset; // @[PayloadArray.scala 59:18]
    end
    if (wen_1) begin // @[PayloadArray.scala 58:16]
      payload_1_ctrl_fuType <= io_write_0_data_ctrl_fuType; // @[PayloadArray.scala 59:18]
    end
    if (wen_1) begin // @[PayloadArray.scala 58:16]
      payload_1_ctrl_fuOpType <= io_write_0_data_ctrl_fuOpType; // @[PayloadArray.scala 59:18]
    end
    if (wen_1) begin // @[PayloadArray.scala 58:16]
      payload_1_ctrl_rfWen <= io_write_0_data_ctrl_rfWen; // @[PayloadArray.scala 59:18]
    end
    if (wen_1) begin // @[PayloadArray.scala 58:16]
      payload_1_ctrl_fpWen <= io_write_0_data_ctrl_fpWen; // @[PayloadArray.scala 59:18]
    end
    if (wen_1) begin // @[PayloadArray.scala 58:16]
      payload_1_ctrl_imm <= io_write_0_data_ctrl_imm; // @[PayloadArray.scala 59:18]
    end
    if (wen_1) begin // @[PayloadArray.scala 58:16]
      payload_1_ctrl_fpu_isAddSub <= io_write_0_data_ctrl_fpu_isAddSub; // @[PayloadArray.scala 59:18]
    end
    if (wen_1) begin // @[PayloadArray.scala 58:16]
      payload_1_ctrl_fpu_typeTagIn <= io_write_0_data_ctrl_fpu_typeTagIn; // @[PayloadArray.scala 59:18]
    end
    if (wen_1) begin // @[PayloadArray.scala 58:16]
      payload_1_ctrl_fpu_typeTagOut <= io_write_0_data_ctrl_fpu_typeTagOut; // @[PayloadArray.scala 59:18]
    end
    if (wen_1) begin // @[PayloadArray.scala 58:16]
      payload_1_ctrl_fpu_fromInt <= io_write_0_data_ctrl_fpu_fromInt; // @[PayloadArray.scala 59:18]
    end
    if (wen_1) begin // @[PayloadArray.scala 58:16]
      payload_1_ctrl_fpu_wflags <= io_write_0_data_ctrl_fpu_wflags; // @[PayloadArray.scala 59:18]
    end
    if (wen_1) begin // @[PayloadArray.scala 58:16]
      payload_1_ctrl_fpu_fpWen <= io_write_0_data_ctrl_fpu_fpWen; // @[PayloadArray.scala 59:18]
    end
    if (wen_1) begin // @[PayloadArray.scala 58:16]
      payload_1_ctrl_fpu_fmaCmd <= io_write_0_data_ctrl_fpu_fmaCmd; // @[PayloadArray.scala 59:18]
    end
    if (wen_1) begin // @[PayloadArray.scala 58:16]
      payload_1_ctrl_fpu_div <= io_write_0_data_ctrl_fpu_div; // @[PayloadArray.scala 59:18]
    end
    if (wen_1) begin // @[PayloadArray.scala 58:16]
      payload_1_ctrl_fpu_sqrt <= io_write_0_data_ctrl_fpu_sqrt; // @[PayloadArray.scala 59:18]
    end
    if (wen_1) begin // @[PayloadArray.scala 58:16]
      payload_1_ctrl_fpu_fcvt <= io_write_0_data_ctrl_fpu_fcvt; // @[PayloadArray.scala 59:18]
    end
    if (wen_1) begin // @[PayloadArray.scala 58:16]
      payload_1_ctrl_fpu_typ <= io_write_0_data_ctrl_fpu_typ; // @[PayloadArray.scala 59:18]
    end
    if (wen_1) begin // @[PayloadArray.scala 58:16]
      payload_1_ctrl_fpu_fmt <= io_write_0_data_ctrl_fpu_fmt; // @[PayloadArray.scala 59:18]
    end
    if (wen_1) begin // @[PayloadArray.scala 58:16]
      payload_1_ctrl_fpu_ren3 <= io_write_0_data_ctrl_fpu_ren3; // @[PayloadArray.scala 59:18]
    end
    if (wen_1) begin // @[PayloadArray.scala 58:16]
      payload_1_ctrl_fpu_rm <= io_write_0_data_ctrl_fpu_rm; // @[PayloadArray.scala 59:18]
    end
    if (wen_1) begin // @[PayloadArray.scala 58:16]
      payload_1_pdest <= io_write_0_data_pdest; // @[PayloadArray.scala 59:18]
    end
    if (wen_1) begin // @[PayloadArray.scala 58:16]
      payload_1_robIdx_flag <= io_write_0_data_robIdx_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen_1) begin // @[PayloadArray.scala 58:16]
      payload_1_robIdx_value <= io_write_0_data_robIdx_value; // @[PayloadArray.scala 59:18]
    end
    if (wen_2) begin // @[PayloadArray.scala 58:16]
      payload_2_cf_pd_isRVC <= io_write_0_data_cf_pd_isRVC; // @[PayloadArray.scala 59:18]
    end
    if (wen_2) begin // @[PayloadArray.scala 58:16]
      payload_2_cf_pd_brType <= io_write_0_data_cf_pd_brType; // @[PayloadArray.scala 59:18]
    end
    if (wen_2) begin // @[PayloadArray.scala 58:16]
      payload_2_cf_pd_isCall <= io_write_0_data_cf_pd_isCall; // @[PayloadArray.scala 59:18]
    end
    if (wen_2) begin // @[PayloadArray.scala 58:16]
      payload_2_cf_pd_isRet <= io_write_0_data_cf_pd_isRet; // @[PayloadArray.scala 59:18]
    end
    if (wen_2) begin // @[PayloadArray.scala 58:16]
      payload_2_cf_pred_taken <= io_write_0_data_cf_pred_taken; // @[PayloadArray.scala 59:18]
    end
    if (wen_2) begin // @[PayloadArray.scala 58:16]
      payload_2_cf_ftqPtr_flag <= io_write_0_data_cf_ftqPtr_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen_2) begin // @[PayloadArray.scala 58:16]
      payload_2_cf_ftqPtr_value <= io_write_0_data_cf_ftqPtr_value; // @[PayloadArray.scala 59:18]
    end
    if (wen_2) begin // @[PayloadArray.scala 58:16]
      payload_2_cf_ftqOffset <= io_write_0_data_cf_ftqOffset; // @[PayloadArray.scala 59:18]
    end
    if (wen_2) begin // @[PayloadArray.scala 58:16]
      payload_2_ctrl_fuType <= io_write_0_data_ctrl_fuType; // @[PayloadArray.scala 59:18]
    end
    if (wen_2) begin // @[PayloadArray.scala 58:16]
      payload_2_ctrl_fuOpType <= io_write_0_data_ctrl_fuOpType; // @[PayloadArray.scala 59:18]
    end
    if (wen_2) begin // @[PayloadArray.scala 58:16]
      payload_2_ctrl_rfWen <= io_write_0_data_ctrl_rfWen; // @[PayloadArray.scala 59:18]
    end
    if (wen_2) begin // @[PayloadArray.scala 58:16]
      payload_2_ctrl_fpWen <= io_write_0_data_ctrl_fpWen; // @[PayloadArray.scala 59:18]
    end
    if (wen_2) begin // @[PayloadArray.scala 58:16]
      payload_2_ctrl_imm <= io_write_0_data_ctrl_imm; // @[PayloadArray.scala 59:18]
    end
    if (wen_2) begin // @[PayloadArray.scala 58:16]
      payload_2_ctrl_fpu_isAddSub <= io_write_0_data_ctrl_fpu_isAddSub; // @[PayloadArray.scala 59:18]
    end
    if (wen_2) begin // @[PayloadArray.scala 58:16]
      payload_2_ctrl_fpu_typeTagIn <= io_write_0_data_ctrl_fpu_typeTagIn; // @[PayloadArray.scala 59:18]
    end
    if (wen_2) begin // @[PayloadArray.scala 58:16]
      payload_2_ctrl_fpu_typeTagOut <= io_write_0_data_ctrl_fpu_typeTagOut; // @[PayloadArray.scala 59:18]
    end
    if (wen_2) begin // @[PayloadArray.scala 58:16]
      payload_2_ctrl_fpu_fromInt <= io_write_0_data_ctrl_fpu_fromInt; // @[PayloadArray.scala 59:18]
    end
    if (wen_2) begin // @[PayloadArray.scala 58:16]
      payload_2_ctrl_fpu_wflags <= io_write_0_data_ctrl_fpu_wflags; // @[PayloadArray.scala 59:18]
    end
    if (wen_2) begin // @[PayloadArray.scala 58:16]
      payload_2_ctrl_fpu_fpWen <= io_write_0_data_ctrl_fpu_fpWen; // @[PayloadArray.scala 59:18]
    end
    if (wen_2) begin // @[PayloadArray.scala 58:16]
      payload_2_ctrl_fpu_fmaCmd <= io_write_0_data_ctrl_fpu_fmaCmd; // @[PayloadArray.scala 59:18]
    end
    if (wen_2) begin // @[PayloadArray.scala 58:16]
      payload_2_ctrl_fpu_div <= io_write_0_data_ctrl_fpu_div; // @[PayloadArray.scala 59:18]
    end
    if (wen_2) begin // @[PayloadArray.scala 58:16]
      payload_2_ctrl_fpu_sqrt <= io_write_0_data_ctrl_fpu_sqrt; // @[PayloadArray.scala 59:18]
    end
    if (wen_2) begin // @[PayloadArray.scala 58:16]
      payload_2_ctrl_fpu_fcvt <= io_write_0_data_ctrl_fpu_fcvt; // @[PayloadArray.scala 59:18]
    end
    if (wen_2) begin // @[PayloadArray.scala 58:16]
      payload_2_ctrl_fpu_typ <= io_write_0_data_ctrl_fpu_typ; // @[PayloadArray.scala 59:18]
    end
    if (wen_2) begin // @[PayloadArray.scala 58:16]
      payload_2_ctrl_fpu_fmt <= io_write_0_data_ctrl_fpu_fmt; // @[PayloadArray.scala 59:18]
    end
    if (wen_2) begin // @[PayloadArray.scala 58:16]
      payload_2_ctrl_fpu_ren3 <= io_write_0_data_ctrl_fpu_ren3; // @[PayloadArray.scala 59:18]
    end
    if (wen_2) begin // @[PayloadArray.scala 58:16]
      payload_2_ctrl_fpu_rm <= io_write_0_data_ctrl_fpu_rm; // @[PayloadArray.scala 59:18]
    end
    if (wen_2) begin // @[PayloadArray.scala 58:16]
      payload_2_pdest <= io_write_0_data_pdest; // @[PayloadArray.scala 59:18]
    end
    if (wen_2) begin // @[PayloadArray.scala 58:16]
      payload_2_robIdx_flag <= io_write_0_data_robIdx_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen_2) begin // @[PayloadArray.scala 58:16]
      payload_2_robIdx_value <= io_write_0_data_robIdx_value; // @[PayloadArray.scala 59:18]
    end
    if (wen_3) begin // @[PayloadArray.scala 58:16]
      payload_3_cf_pd_isRVC <= io_write_0_data_cf_pd_isRVC; // @[PayloadArray.scala 59:18]
    end
    if (wen_3) begin // @[PayloadArray.scala 58:16]
      payload_3_cf_pd_brType <= io_write_0_data_cf_pd_brType; // @[PayloadArray.scala 59:18]
    end
    if (wen_3) begin // @[PayloadArray.scala 58:16]
      payload_3_cf_pd_isCall <= io_write_0_data_cf_pd_isCall; // @[PayloadArray.scala 59:18]
    end
    if (wen_3) begin // @[PayloadArray.scala 58:16]
      payload_3_cf_pd_isRet <= io_write_0_data_cf_pd_isRet; // @[PayloadArray.scala 59:18]
    end
    if (wen_3) begin // @[PayloadArray.scala 58:16]
      payload_3_cf_pred_taken <= io_write_0_data_cf_pred_taken; // @[PayloadArray.scala 59:18]
    end
    if (wen_3) begin // @[PayloadArray.scala 58:16]
      payload_3_cf_ftqPtr_flag <= io_write_0_data_cf_ftqPtr_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen_3) begin // @[PayloadArray.scala 58:16]
      payload_3_cf_ftqPtr_value <= io_write_0_data_cf_ftqPtr_value; // @[PayloadArray.scala 59:18]
    end
    if (wen_3) begin // @[PayloadArray.scala 58:16]
      payload_3_cf_ftqOffset <= io_write_0_data_cf_ftqOffset; // @[PayloadArray.scala 59:18]
    end
    if (wen_3) begin // @[PayloadArray.scala 58:16]
      payload_3_ctrl_fuType <= io_write_0_data_ctrl_fuType; // @[PayloadArray.scala 59:18]
    end
    if (wen_3) begin // @[PayloadArray.scala 58:16]
      payload_3_ctrl_fuOpType <= io_write_0_data_ctrl_fuOpType; // @[PayloadArray.scala 59:18]
    end
    if (wen_3) begin // @[PayloadArray.scala 58:16]
      payload_3_ctrl_rfWen <= io_write_0_data_ctrl_rfWen; // @[PayloadArray.scala 59:18]
    end
    if (wen_3) begin // @[PayloadArray.scala 58:16]
      payload_3_ctrl_fpWen <= io_write_0_data_ctrl_fpWen; // @[PayloadArray.scala 59:18]
    end
    if (wen_3) begin // @[PayloadArray.scala 58:16]
      payload_3_ctrl_imm <= io_write_0_data_ctrl_imm; // @[PayloadArray.scala 59:18]
    end
    if (wen_3) begin // @[PayloadArray.scala 58:16]
      payload_3_ctrl_fpu_isAddSub <= io_write_0_data_ctrl_fpu_isAddSub; // @[PayloadArray.scala 59:18]
    end
    if (wen_3) begin // @[PayloadArray.scala 58:16]
      payload_3_ctrl_fpu_typeTagIn <= io_write_0_data_ctrl_fpu_typeTagIn; // @[PayloadArray.scala 59:18]
    end
    if (wen_3) begin // @[PayloadArray.scala 58:16]
      payload_3_ctrl_fpu_typeTagOut <= io_write_0_data_ctrl_fpu_typeTagOut; // @[PayloadArray.scala 59:18]
    end
    if (wen_3) begin // @[PayloadArray.scala 58:16]
      payload_3_ctrl_fpu_fromInt <= io_write_0_data_ctrl_fpu_fromInt; // @[PayloadArray.scala 59:18]
    end
    if (wen_3) begin // @[PayloadArray.scala 58:16]
      payload_3_ctrl_fpu_wflags <= io_write_0_data_ctrl_fpu_wflags; // @[PayloadArray.scala 59:18]
    end
    if (wen_3) begin // @[PayloadArray.scala 58:16]
      payload_3_ctrl_fpu_fpWen <= io_write_0_data_ctrl_fpu_fpWen; // @[PayloadArray.scala 59:18]
    end
    if (wen_3) begin // @[PayloadArray.scala 58:16]
      payload_3_ctrl_fpu_fmaCmd <= io_write_0_data_ctrl_fpu_fmaCmd; // @[PayloadArray.scala 59:18]
    end
    if (wen_3) begin // @[PayloadArray.scala 58:16]
      payload_3_ctrl_fpu_div <= io_write_0_data_ctrl_fpu_div; // @[PayloadArray.scala 59:18]
    end
    if (wen_3) begin // @[PayloadArray.scala 58:16]
      payload_3_ctrl_fpu_sqrt <= io_write_0_data_ctrl_fpu_sqrt; // @[PayloadArray.scala 59:18]
    end
    if (wen_3) begin // @[PayloadArray.scala 58:16]
      payload_3_ctrl_fpu_fcvt <= io_write_0_data_ctrl_fpu_fcvt; // @[PayloadArray.scala 59:18]
    end
    if (wen_3) begin // @[PayloadArray.scala 58:16]
      payload_3_ctrl_fpu_typ <= io_write_0_data_ctrl_fpu_typ; // @[PayloadArray.scala 59:18]
    end
    if (wen_3) begin // @[PayloadArray.scala 58:16]
      payload_3_ctrl_fpu_fmt <= io_write_0_data_ctrl_fpu_fmt; // @[PayloadArray.scala 59:18]
    end
    if (wen_3) begin // @[PayloadArray.scala 58:16]
      payload_3_ctrl_fpu_ren3 <= io_write_0_data_ctrl_fpu_ren3; // @[PayloadArray.scala 59:18]
    end
    if (wen_3) begin // @[PayloadArray.scala 58:16]
      payload_3_ctrl_fpu_rm <= io_write_0_data_ctrl_fpu_rm; // @[PayloadArray.scala 59:18]
    end
    if (wen_3) begin // @[PayloadArray.scala 58:16]
      payload_3_pdest <= io_write_0_data_pdest; // @[PayloadArray.scala 59:18]
    end
    if (wen_3) begin // @[PayloadArray.scala 58:16]
      payload_3_robIdx_flag <= io_write_0_data_robIdx_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen_3) begin // @[PayloadArray.scala 58:16]
      payload_3_robIdx_value <= io_write_0_data_robIdx_value; // @[PayloadArray.scala 59:18]
    end
    if (wen_4) begin // @[PayloadArray.scala 58:16]
      payload_4_cf_pd_isRVC <= io_write_0_data_cf_pd_isRVC; // @[PayloadArray.scala 59:18]
    end
    if (wen_4) begin // @[PayloadArray.scala 58:16]
      payload_4_cf_pd_brType <= io_write_0_data_cf_pd_brType; // @[PayloadArray.scala 59:18]
    end
    if (wen_4) begin // @[PayloadArray.scala 58:16]
      payload_4_cf_pd_isCall <= io_write_0_data_cf_pd_isCall; // @[PayloadArray.scala 59:18]
    end
    if (wen_4) begin // @[PayloadArray.scala 58:16]
      payload_4_cf_pd_isRet <= io_write_0_data_cf_pd_isRet; // @[PayloadArray.scala 59:18]
    end
    if (wen_4) begin // @[PayloadArray.scala 58:16]
      payload_4_cf_pred_taken <= io_write_0_data_cf_pred_taken; // @[PayloadArray.scala 59:18]
    end
    if (wen_4) begin // @[PayloadArray.scala 58:16]
      payload_4_cf_ftqPtr_flag <= io_write_0_data_cf_ftqPtr_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen_4) begin // @[PayloadArray.scala 58:16]
      payload_4_cf_ftqPtr_value <= io_write_0_data_cf_ftqPtr_value; // @[PayloadArray.scala 59:18]
    end
    if (wen_4) begin // @[PayloadArray.scala 58:16]
      payload_4_cf_ftqOffset <= io_write_0_data_cf_ftqOffset; // @[PayloadArray.scala 59:18]
    end
    if (wen_4) begin // @[PayloadArray.scala 58:16]
      payload_4_ctrl_fuType <= io_write_0_data_ctrl_fuType; // @[PayloadArray.scala 59:18]
    end
    if (wen_4) begin // @[PayloadArray.scala 58:16]
      payload_4_ctrl_fuOpType <= io_write_0_data_ctrl_fuOpType; // @[PayloadArray.scala 59:18]
    end
    if (wen_4) begin // @[PayloadArray.scala 58:16]
      payload_4_ctrl_rfWen <= io_write_0_data_ctrl_rfWen; // @[PayloadArray.scala 59:18]
    end
    if (wen_4) begin // @[PayloadArray.scala 58:16]
      payload_4_ctrl_fpWen <= io_write_0_data_ctrl_fpWen; // @[PayloadArray.scala 59:18]
    end
    if (wen_4) begin // @[PayloadArray.scala 58:16]
      payload_4_ctrl_imm <= io_write_0_data_ctrl_imm; // @[PayloadArray.scala 59:18]
    end
    if (wen_4) begin // @[PayloadArray.scala 58:16]
      payload_4_ctrl_fpu_isAddSub <= io_write_0_data_ctrl_fpu_isAddSub; // @[PayloadArray.scala 59:18]
    end
    if (wen_4) begin // @[PayloadArray.scala 58:16]
      payload_4_ctrl_fpu_typeTagIn <= io_write_0_data_ctrl_fpu_typeTagIn; // @[PayloadArray.scala 59:18]
    end
    if (wen_4) begin // @[PayloadArray.scala 58:16]
      payload_4_ctrl_fpu_typeTagOut <= io_write_0_data_ctrl_fpu_typeTagOut; // @[PayloadArray.scala 59:18]
    end
    if (wen_4) begin // @[PayloadArray.scala 58:16]
      payload_4_ctrl_fpu_fromInt <= io_write_0_data_ctrl_fpu_fromInt; // @[PayloadArray.scala 59:18]
    end
    if (wen_4) begin // @[PayloadArray.scala 58:16]
      payload_4_ctrl_fpu_wflags <= io_write_0_data_ctrl_fpu_wflags; // @[PayloadArray.scala 59:18]
    end
    if (wen_4) begin // @[PayloadArray.scala 58:16]
      payload_4_ctrl_fpu_fpWen <= io_write_0_data_ctrl_fpu_fpWen; // @[PayloadArray.scala 59:18]
    end
    if (wen_4) begin // @[PayloadArray.scala 58:16]
      payload_4_ctrl_fpu_fmaCmd <= io_write_0_data_ctrl_fpu_fmaCmd; // @[PayloadArray.scala 59:18]
    end
    if (wen_4) begin // @[PayloadArray.scala 58:16]
      payload_4_ctrl_fpu_div <= io_write_0_data_ctrl_fpu_div; // @[PayloadArray.scala 59:18]
    end
    if (wen_4) begin // @[PayloadArray.scala 58:16]
      payload_4_ctrl_fpu_sqrt <= io_write_0_data_ctrl_fpu_sqrt; // @[PayloadArray.scala 59:18]
    end
    if (wen_4) begin // @[PayloadArray.scala 58:16]
      payload_4_ctrl_fpu_fcvt <= io_write_0_data_ctrl_fpu_fcvt; // @[PayloadArray.scala 59:18]
    end
    if (wen_4) begin // @[PayloadArray.scala 58:16]
      payload_4_ctrl_fpu_typ <= io_write_0_data_ctrl_fpu_typ; // @[PayloadArray.scala 59:18]
    end
    if (wen_4) begin // @[PayloadArray.scala 58:16]
      payload_4_ctrl_fpu_fmt <= io_write_0_data_ctrl_fpu_fmt; // @[PayloadArray.scala 59:18]
    end
    if (wen_4) begin // @[PayloadArray.scala 58:16]
      payload_4_ctrl_fpu_ren3 <= io_write_0_data_ctrl_fpu_ren3; // @[PayloadArray.scala 59:18]
    end
    if (wen_4) begin // @[PayloadArray.scala 58:16]
      payload_4_ctrl_fpu_rm <= io_write_0_data_ctrl_fpu_rm; // @[PayloadArray.scala 59:18]
    end
    if (wen_4) begin // @[PayloadArray.scala 58:16]
      payload_4_pdest <= io_write_0_data_pdest; // @[PayloadArray.scala 59:18]
    end
    if (wen_4) begin // @[PayloadArray.scala 58:16]
      payload_4_robIdx_flag <= io_write_0_data_robIdx_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen_4) begin // @[PayloadArray.scala 58:16]
      payload_4_robIdx_value <= io_write_0_data_robIdx_value; // @[PayloadArray.scala 59:18]
    end
    if (wen_5) begin // @[PayloadArray.scala 58:16]
      payload_5_cf_pd_isRVC <= io_write_0_data_cf_pd_isRVC; // @[PayloadArray.scala 59:18]
    end
    if (wen_5) begin // @[PayloadArray.scala 58:16]
      payload_5_cf_pd_brType <= io_write_0_data_cf_pd_brType; // @[PayloadArray.scala 59:18]
    end
    if (wen_5) begin // @[PayloadArray.scala 58:16]
      payload_5_cf_pd_isCall <= io_write_0_data_cf_pd_isCall; // @[PayloadArray.scala 59:18]
    end
    if (wen_5) begin // @[PayloadArray.scala 58:16]
      payload_5_cf_pd_isRet <= io_write_0_data_cf_pd_isRet; // @[PayloadArray.scala 59:18]
    end
    if (wen_5) begin // @[PayloadArray.scala 58:16]
      payload_5_cf_pred_taken <= io_write_0_data_cf_pred_taken; // @[PayloadArray.scala 59:18]
    end
    if (wen_5) begin // @[PayloadArray.scala 58:16]
      payload_5_cf_ftqPtr_flag <= io_write_0_data_cf_ftqPtr_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen_5) begin // @[PayloadArray.scala 58:16]
      payload_5_cf_ftqPtr_value <= io_write_0_data_cf_ftqPtr_value; // @[PayloadArray.scala 59:18]
    end
    if (wen_5) begin // @[PayloadArray.scala 58:16]
      payload_5_cf_ftqOffset <= io_write_0_data_cf_ftqOffset; // @[PayloadArray.scala 59:18]
    end
    if (wen_5) begin // @[PayloadArray.scala 58:16]
      payload_5_ctrl_fuType <= io_write_0_data_ctrl_fuType; // @[PayloadArray.scala 59:18]
    end
    if (wen_5) begin // @[PayloadArray.scala 58:16]
      payload_5_ctrl_fuOpType <= io_write_0_data_ctrl_fuOpType; // @[PayloadArray.scala 59:18]
    end
    if (wen_5) begin // @[PayloadArray.scala 58:16]
      payload_5_ctrl_rfWen <= io_write_0_data_ctrl_rfWen; // @[PayloadArray.scala 59:18]
    end
    if (wen_5) begin // @[PayloadArray.scala 58:16]
      payload_5_ctrl_fpWen <= io_write_0_data_ctrl_fpWen; // @[PayloadArray.scala 59:18]
    end
    if (wen_5) begin // @[PayloadArray.scala 58:16]
      payload_5_ctrl_imm <= io_write_0_data_ctrl_imm; // @[PayloadArray.scala 59:18]
    end
    if (wen_5) begin // @[PayloadArray.scala 58:16]
      payload_5_ctrl_fpu_isAddSub <= io_write_0_data_ctrl_fpu_isAddSub; // @[PayloadArray.scala 59:18]
    end
    if (wen_5) begin // @[PayloadArray.scala 58:16]
      payload_5_ctrl_fpu_typeTagIn <= io_write_0_data_ctrl_fpu_typeTagIn; // @[PayloadArray.scala 59:18]
    end
    if (wen_5) begin // @[PayloadArray.scala 58:16]
      payload_5_ctrl_fpu_typeTagOut <= io_write_0_data_ctrl_fpu_typeTagOut; // @[PayloadArray.scala 59:18]
    end
    if (wen_5) begin // @[PayloadArray.scala 58:16]
      payload_5_ctrl_fpu_fromInt <= io_write_0_data_ctrl_fpu_fromInt; // @[PayloadArray.scala 59:18]
    end
    if (wen_5) begin // @[PayloadArray.scala 58:16]
      payload_5_ctrl_fpu_wflags <= io_write_0_data_ctrl_fpu_wflags; // @[PayloadArray.scala 59:18]
    end
    if (wen_5) begin // @[PayloadArray.scala 58:16]
      payload_5_ctrl_fpu_fpWen <= io_write_0_data_ctrl_fpu_fpWen; // @[PayloadArray.scala 59:18]
    end
    if (wen_5) begin // @[PayloadArray.scala 58:16]
      payload_5_ctrl_fpu_fmaCmd <= io_write_0_data_ctrl_fpu_fmaCmd; // @[PayloadArray.scala 59:18]
    end
    if (wen_5) begin // @[PayloadArray.scala 58:16]
      payload_5_ctrl_fpu_div <= io_write_0_data_ctrl_fpu_div; // @[PayloadArray.scala 59:18]
    end
    if (wen_5) begin // @[PayloadArray.scala 58:16]
      payload_5_ctrl_fpu_sqrt <= io_write_0_data_ctrl_fpu_sqrt; // @[PayloadArray.scala 59:18]
    end
    if (wen_5) begin // @[PayloadArray.scala 58:16]
      payload_5_ctrl_fpu_fcvt <= io_write_0_data_ctrl_fpu_fcvt; // @[PayloadArray.scala 59:18]
    end
    if (wen_5) begin // @[PayloadArray.scala 58:16]
      payload_5_ctrl_fpu_typ <= io_write_0_data_ctrl_fpu_typ; // @[PayloadArray.scala 59:18]
    end
    if (wen_5) begin // @[PayloadArray.scala 58:16]
      payload_5_ctrl_fpu_fmt <= io_write_0_data_ctrl_fpu_fmt; // @[PayloadArray.scala 59:18]
    end
    if (wen_5) begin // @[PayloadArray.scala 58:16]
      payload_5_ctrl_fpu_ren3 <= io_write_0_data_ctrl_fpu_ren3; // @[PayloadArray.scala 59:18]
    end
    if (wen_5) begin // @[PayloadArray.scala 58:16]
      payload_5_ctrl_fpu_rm <= io_write_0_data_ctrl_fpu_rm; // @[PayloadArray.scala 59:18]
    end
    if (wen_5) begin // @[PayloadArray.scala 58:16]
      payload_5_pdest <= io_write_0_data_pdest; // @[PayloadArray.scala 59:18]
    end
    if (wen_5) begin // @[PayloadArray.scala 58:16]
      payload_5_robIdx_flag <= io_write_0_data_robIdx_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen_5) begin // @[PayloadArray.scala 58:16]
      payload_5_robIdx_value <= io_write_0_data_robIdx_value; // @[PayloadArray.scala 59:18]
    end
    if (wen_6) begin // @[PayloadArray.scala 58:16]
      payload_6_cf_pd_isRVC <= io_write_0_data_cf_pd_isRVC; // @[PayloadArray.scala 59:18]
    end
    if (wen_6) begin // @[PayloadArray.scala 58:16]
      payload_6_cf_pd_brType <= io_write_0_data_cf_pd_brType; // @[PayloadArray.scala 59:18]
    end
    if (wen_6) begin // @[PayloadArray.scala 58:16]
      payload_6_cf_pd_isCall <= io_write_0_data_cf_pd_isCall; // @[PayloadArray.scala 59:18]
    end
    if (wen_6) begin // @[PayloadArray.scala 58:16]
      payload_6_cf_pd_isRet <= io_write_0_data_cf_pd_isRet; // @[PayloadArray.scala 59:18]
    end
    if (wen_6) begin // @[PayloadArray.scala 58:16]
      payload_6_cf_pred_taken <= io_write_0_data_cf_pred_taken; // @[PayloadArray.scala 59:18]
    end
    if (wen_6) begin // @[PayloadArray.scala 58:16]
      payload_6_cf_ftqPtr_flag <= io_write_0_data_cf_ftqPtr_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen_6) begin // @[PayloadArray.scala 58:16]
      payload_6_cf_ftqPtr_value <= io_write_0_data_cf_ftqPtr_value; // @[PayloadArray.scala 59:18]
    end
    if (wen_6) begin // @[PayloadArray.scala 58:16]
      payload_6_cf_ftqOffset <= io_write_0_data_cf_ftqOffset; // @[PayloadArray.scala 59:18]
    end
    if (wen_6) begin // @[PayloadArray.scala 58:16]
      payload_6_ctrl_fuType <= io_write_0_data_ctrl_fuType; // @[PayloadArray.scala 59:18]
    end
    if (wen_6) begin // @[PayloadArray.scala 58:16]
      payload_6_ctrl_fuOpType <= io_write_0_data_ctrl_fuOpType; // @[PayloadArray.scala 59:18]
    end
    if (wen_6) begin // @[PayloadArray.scala 58:16]
      payload_6_ctrl_rfWen <= io_write_0_data_ctrl_rfWen; // @[PayloadArray.scala 59:18]
    end
    if (wen_6) begin // @[PayloadArray.scala 58:16]
      payload_6_ctrl_fpWen <= io_write_0_data_ctrl_fpWen; // @[PayloadArray.scala 59:18]
    end
    if (wen_6) begin // @[PayloadArray.scala 58:16]
      payload_6_ctrl_imm <= io_write_0_data_ctrl_imm; // @[PayloadArray.scala 59:18]
    end
    if (wen_6) begin // @[PayloadArray.scala 58:16]
      payload_6_ctrl_fpu_isAddSub <= io_write_0_data_ctrl_fpu_isAddSub; // @[PayloadArray.scala 59:18]
    end
    if (wen_6) begin // @[PayloadArray.scala 58:16]
      payload_6_ctrl_fpu_typeTagIn <= io_write_0_data_ctrl_fpu_typeTagIn; // @[PayloadArray.scala 59:18]
    end
    if (wen_6) begin // @[PayloadArray.scala 58:16]
      payload_6_ctrl_fpu_typeTagOut <= io_write_0_data_ctrl_fpu_typeTagOut; // @[PayloadArray.scala 59:18]
    end
    if (wen_6) begin // @[PayloadArray.scala 58:16]
      payload_6_ctrl_fpu_fromInt <= io_write_0_data_ctrl_fpu_fromInt; // @[PayloadArray.scala 59:18]
    end
    if (wen_6) begin // @[PayloadArray.scala 58:16]
      payload_6_ctrl_fpu_wflags <= io_write_0_data_ctrl_fpu_wflags; // @[PayloadArray.scala 59:18]
    end
    if (wen_6) begin // @[PayloadArray.scala 58:16]
      payload_6_ctrl_fpu_fpWen <= io_write_0_data_ctrl_fpu_fpWen; // @[PayloadArray.scala 59:18]
    end
    if (wen_6) begin // @[PayloadArray.scala 58:16]
      payload_6_ctrl_fpu_fmaCmd <= io_write_0_data_ctrl_fpu_fmaCmd; // @[PayloadArray.scala 59:18]
    end
    if (wen_6) begin // @[PayloadArray.scala 58:16]
      payload_6_ctrl_fpu_div <= io_write_0_data_ctrl_fpu_div; // @[PayloadArray.scala 59:18]
    end
    if (wen_6) begin // @[PayloadArray.scala 58:16]
      payload_6_ctrl_fpu_sqrt <= io_write_0_data_ctrl_fpu_sqrt; // @[PayloadArray.scala 59:18]
    end
    if (wen_6) begin // @[PayloadArray.scala 58:16]
      payload_6_ctrl_fpu_fcvt <= io_write_0_data_ctrl_fpu_fcvt; // @[PayloadArray.scala 59:18]
    end
    if (wen_6) begin // @[PayloadArray.scala 58:16]
      payload_6_ctrl_fpu_typ <= io_write_0_data_ctrl_fpu_typ; // @[PayloadArray.scala 59:18]
    end
    if (wen_6) begin // @[PayloadArray.scala 58:16]
      payload_6_ctrl_fpu_fmt <= io_write_0_data_ctrl_fpu_fmt; // @[PayloadArray.scala 59:18]
    end
    if (wen_6) begin // @[PayloadArray.scala 58:16]
      payload_6_ctrl_fpu_ren3 <= io_write_0_data_ctrl_fpu_ren3; // @[PayloadArray.scala 59:18]
    end
    if (wen_6) begin // @[PayloadArray.scala 58:16]
      payload_6_ctrl_fpu_rm <= io_write_0_data_ctrl_fpu_rm; // @[PayloadArray.scala 59:18]
    end
    if (wen_6) begin // @[PayloadArray.scala 58:16]
      payload_6_pdest <= io_write_0_data_pdest; // @[PayloadArray.scala 59:18]
    end
    if (wen_6) begin // @[PayloadArray.scala 58:16]
      payload_6_robIdx_flag <= io_write_0_data_robIdx_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen_6) begin // @[PayloadArray.scala 58:16]
      payload_6_robIdx_value <= io_write_0_data_robIdx_value; // @[PayloadArray.scala 59:18]
    end
    if (wen_7) begin // @[PayloadArray.scala 58:16]
      payload_7_cf_pd_isRVC <= io_write_0_data_cf_pd_isRVC; // @[PayloadArray.scala 59:18]
    end
    if (wen_7) begin // @[PayloadArray.scala 58:16]
      payload_7_cf_pd_brType <= io_write_0_data_cf_pd_brType; // @[PayloadArray.scala 59:18]
    end
    if (wen_7) begin // @[PayloadArray.scala 58:16]
      payload_7_cf_pd_isCall <= io_write_0_data_cf_pd_isCall; // @[PayloadArray.scala 59:18]
    end
    if (wen_7) begin // @[PayloadArray.scala 58:16]
      payload_7_cf_pd_isRet <= io_write_0_data_cf_pd_isRet; // @[PayloadArray.scala 59:18]
    end
    if (wen_7) begin // @[PayloadArray.scala 58:16]
      payload_7_cf_pred_taken <= io_write_0_data_cf_pred_taken; // @[PayloadArray.scala 59:18]
    end
    if (wen_7) begin // @[PayloadArray.scala 58:16]
      payload_7_cf_ftqPtr_flag <= io_write_0_data_cf_ftqPtr_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen_7) begin // @[PayloadArray.scala 58:16]
      payload_7_cf_ftqPtr_value <= io_write_0_data_cf_ftqPtr_value; // @[PayloadArray.scala 59:18]
    end
    if (wen_7) begin // @[PayloadArray.scala 58:16]
      payload_7_cf_ftqOffset <= io_write_0_data_cf_ftqOffset; // @[PayloadArray.scala 59:18]
    end
    if (wen_7) begin // @[PayloadArray.scala 58:16]
      payload_7_ctrl_fuType <= io_write_0_data_ctrl_fuType; // @[PayloadArray.scala 59:18]
    end
    if (wen_7) begin // @[PayloadArray.scala 58:16]
      payload_7_ctrl_fuOpType <= io_write_0_data_ctrl_fuOpType; // @[PayloadArray.scala 59:18]
    end
    if (wen_7) begin // @[PayloadArray.scala 58:16]
      payload_7_ctrl_rfWen <= io_write_0_data_ctrl_rfWen; // @[PayloadArray.scala 59:18]
    end
    if (wen_7) begin // @[PayloadArray.scala 58:16]
      payload_7_ctrl_fpWen <= io_write_0_data_ctrl_fpWen; // @[PayloadArray.scala 59:18]
    end
    if (wen_7) begin // @[PayloadArray.scala 58:16]
      payload_7_ctrl_imm <= io_write_0_data_ctrl_imm; // @[PayloadArray.scala 59:18]
    end
    if (wen_7) begin // @[PayloadArray.scala 58:16]
      payload_7_ctrl_fpu_isAddSub <= io_write_0_data_ctrl_fpu_isAddSub; // @[PayloadArray.scala 59:18]
    end
    if (wen_7) begin // @[PayloadArray.scala 58:16]
      payload_7_ctrl_fpu_typeTagIn <= io_write_0_data_ctrl_fpu_typeTagIn; // @[PayloadArray.scala 59:18]
    end
    if (wen_7) begin // @[PayloadArray.scala 58:16]
      payload_7_ctrl_fpu_typeTagOut <= io_write_0_data_ctrl_fpu_typeTagOut; // @[PayloadArray.scala 59:18]
    end
    if (wen_7) begin // @[PayloadArray.scala 58:16]
      payload_7_ctrl_fpu_fromInt <= io_write_0_data_ctrl_fpu_fromInt; // @[PayloadArray.scala 59:18]
    end
    if (wen_7) begin // @[PayloadArray.scala 58:16]
      payload_7_ctrl_fpu_wflags <= io_write_0_data_ctrl_fpu_wflags; // @[PayloadArray.scala 59:18]
    end
    if (wen_7) begin // @[PayloadArray.scala 58:16]
      payload_7_ctrl_fpu_fpWen <= io_write_0_data_ctrl_fpu_fpWen; // @[PayloadArray.scala 59:18]
    end
    if (wen_7) begin // @[PayloadArray.scala 58:16]
      payload_7_ctrl_fpu_fmaCmd <= io_write_0_data_ctrl_fpu_fmaCmd; // @[PayloadArray.scala 59:18]
    end
    if (wen_7) begin // @[PayloadArray.scala 58:16]
      payload_7_ctrl_fpu_div <= io_write_0_data_ctrl_fpu_div; // @[PayloadArray.scala 59:18]
    end
    if (wen_7) begin // @[PayloadArray.scala 58:16]
      payload_7_ctrl_fpu_sqrt <= io_write_0_data_ctrl_fpu_sqrt; // @[PayloadArray.scala 59:18]
    end
    if (wen_7) begin // @[PayloadArray.scala 58:16]
      payload_7_ctrl_fpu_fcvt <= io_write_0_data_ctrl_fpu_fcvt; // @[PayloadArray.scala 59:18]
    end
    if (wen_7) begin // @[PayloadArray.scala 58:16]
      payload_7_ctrl_fpu_typ <= io_write_0_data_ctrl_fpu_typ; // @[PayloadArray.scala 59:18]
    end
    if (wen_7) begin // @[PayloadArray.scala 58:16]
      payload_7_ctrl_fpu_fmt <= io_write_0_data_ctrl_fpu_fmt; // @[PayloadArray.scala 59:18]
    end
    if (wen_7) begin // @[PayloadArray.scala 58:16]
      payload_7_ctrl_fpu_ren3 <= io_write_0_data_ctrl_fpu_ren3; // @[PayloadArray.scala 59:18]
    end
    if (wen_7) begin // @[PayloadArray.scala 58:16]
      payload_7_ctrl_fpu_rm <= io_write_0_data_ctrl_fpu_rm; // @[PayloadArray.scala 59:18]
    end
    if (wen_7) begin // @[PayloadArray.scala 58:16]
      payload_7_pdest <= io_write_0_data_pdest; // @[PayloadArray.scala 59:18]
    end
    if (wen_7) begin // @[PayloadArray.scala 58:16]
      payload_7_robIdx_flag <= io_write_0_data_robIdx_flag; // @[PayloadArray.scala 59:18]
    end
    if (wen_7) begin // @[PayloadArray.scala 58:16]
      payload_7_robIdx_value <= io_write_0_data_robIdx_value; // @[PayloadArray.scala 59:18]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  payload_0_cf_pd_isRVC = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  payload_0_cf_pd_brType = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  payload_0_cf_pd_isCall = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  payload_0_cf_pd_isRet = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  payload_0_cf_pred_taken = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  payload_0_cf_ftqPtr_flag = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  payload_0_cf_ftqPtr_value = _RAND_6[2:0];
  _RAND_7 = {1{`RANDOM}};
  payload_0_cf_ftqOffset = _RAND_7[2:0];
  _RAND_8 = {1{`RANDOM}};
  payload_0_ctrl_fuType = _RAND_8[3:0];
  _RAND_9 = {1{`RANDOM}};
  payload_0_ctrl_fuOpType = _RAND_9[6:0];
  _RAND_10 = {1{`RANDOM}};
  payload_0_ctrl_rfWen = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  payload_0_ctrl_fpWen = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  payload_0_ctrl_imm = _RAND_12[19:0];
  _RAND_13 = {1{`RANDOM}};
  payload_0_ctrl_fpu_isAddSub = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  payload_0_ctrl_fpu_typeTagIn = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  payload_0_ctrl_fpu_typeTagOut = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  payload_0_ctrl_fpu_fromInt = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  payload_0_ctrl_fpu_wflags = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  payload_0_ctrl_fpu_fpWen = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  payload_0_ctrl_fpu_fmaCmd = _RAND_19[1:0];
  _RAND_20 = {1{`RANDOM}};
  payload_0_ctrl_fpu_div = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  payload_0_ctrl_fpu_sqrt = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  payload_0_ctrl_fpu_fcvt = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  payload_0_ctrl_fpu_typ = _RAND_23[1:0];
  _RAND_24 = {1{`RANDOM}};
  payload_0_ctrl_fpu_fmt = _RAND_24[1:0];
  _RAND_25 = {1{`RANDOM}};
  payload_0_ctrl_fpu_ren3 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  payload_0_ctrl_fpu_rm = _RAND_26[2:0];
  _RAND_27 = {1{`RANDOM}};
  payload_0_pdest = _RAND_27[5:0];
  _RAND_28 = {1{`RANDOM}};
  payload_0_robIdx_flag = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  payload_0_robIdx_value = _RAND_29[4:0];
  _RAND_30 = {1{`RANDOM}};
  payload_1_cf_pd_isRVC = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  payload_1_cf_pd_brType = _RAND_31[1:0];
  _RAND_32 = {1{`RANDOM}};
  payload_1_cf_pd_isCall = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  payload_1_cf_pd_isRet = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  payload_1_cf_pred_taken = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  payload_1_cf_ftqPtr_flag = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  payload_1_cf_ftqPtr_value = _RAND_36[2:0];
  _RAND_37 = {1{`RANDOM}};
  payload_1_cf_ftqOffset = _RAND_37[2:0];
  _RAND_38 = {1{`RANDOM}};
  payload_1_ctrl_fuType = _RAND_38[3:0];
  _RAND_39 = {1{`RANDOM}};
  payload_1_ctrl_fuOpType = _RAND_39[6:0];
  _RAND_40 = {1{`RANDOM}};
  payload_1_ctrl_rfWen = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  payload_1_ctrl_fpWen = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  payload_1_ctrl_imm = _RAND_42[19:0];
  _RAND_43 = {1{`RANDOM}};
  payload_1_ctrl_fpu_isAddSub = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  payload_1_ctrl_fpu_typeTagIn = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  payload_1_ctrl_fpu_typeTagOut = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  payload_1_ctrl_fpu_fromInt = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  payload_1_ctrl_fpu_wflags = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  payload_1_ctrl_fpu_fpWen = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  payload_1_ctrl_fpu_fmaCmd = _RAND_49[1:0];
  _RAND_50 = {1{`RANDOM}};
  payload_1_ctrl_fpu_div = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  payload_1_ctrl_fpu_sqrt = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  payload_1_ctrl_fpu_fcvt = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  payload_1_ctrl_fpu_typ = _RAND_53[1:0];
  _RAND_54 = {1{`RANDOM}};
  payload_1_ctrl_fpu_fmt = _RAND_54[1:0];
  _RAND_55 = {1{`RANDOM}};
  payload_1_ctrl_fpu_ren3 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  payload_1_ctrl_fpu_rm = _RAND_56[2:0];
  _RAND_57 = {1{`RANDOM}};
  payload_1_pdest = _RAND_57[5:0];
  _RAND_58 = {1{`RANDOM}};
  payload_1_robIdx_flag = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  payload_1_robIdx_value = _RAND_59[4:0];
  _RAND_60 = {1{`RANDOM}};
  payload_2_cf_pd_isRVC = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  payload_2_cf_pd_brType = _RAND_61[1:0];
  _RAND_62 = {1{`RANDOM}};
  payload_2_cf_pd_isCall = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  payload_2_cf_pd_isRet = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  payload_2_cf_pred_taken = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  payload_2_cf_ftqPtr_flag = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  payload_2_cf_ftqPtr_value = _RAND_66[2:0];
  _RAND_67 = {1{`RANDOM}};
  payload_2_cf_ftqOffset = _RAND_67[2:0];
  _RAND_68 = {1{`RANDOM}};
  payload_2_ctrl_fuType = _RAND_68[3:0];
  _RAND_69 = {1{`RANDOM}};
  payload_2_ctrl_fuOpType = _RAND_69[6:0];
  _RAND_70 = {1{`RANDOM}};
  payload_2_ctrl_rfWen = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  payload_2_ctrl_fpWen = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  payload_2_ctrl_imm = _RAND_72[19:0];
  _RAND_73 = {1{`RANDOM}};
  payload_2_ctrl_fpu_isAddSub = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  payload_2_ctrl_fpu_typeTagIn = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  payload_2_ctrl_fpu_typeTagOut = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  payload_2_ctrl_fpu_fromInt = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  payload_2_ctrl_fpu_wflags = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  payload_2_ctrl_fpu_fpWen = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  payload_2_ctrl_fpu_fmaCmd = _RAND_79[1:0];
  _RAND_80 = {1{`RANDOM}};
  payload_2_ctrl_fpu_div = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  payload_2_ctrl_fpu_sqrt = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  payload_2_ctrl_fpu_fcvt = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  payload_2_ctrl_fpu_typ = _RAND_83[1:0];
  _RAND_84 = {1{`RANDOM}};
  payload_2_ctrl_fpu_fmt = _RAND_84[1:0];
  _RAND_85 = {1{`RANDOM}};
  payload_2_ctrl_fpu_ren3 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  payload_2_ctrl_fpu_rm = _RAND_86[2:0];
  _RAND_87 = {1{`RANDOM}};
  payload_2_pdest = _RAND_87[5:0];
  _RAND_88 = {1{`RANDOM}};
  payload_2_robIdx_flag = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  payload_2_robIdx_value = _RAND_89[4:0];
  _RAND_90 = {1{`RANDOM}};
  payload_3_cf_pd_isRVC = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  payload_3_cf_pd_brType = _RAND_91[1:0];
  _RAND_92 = {1{`RANDOM}};
  payload_3_cf_pd_isCall = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  payload_3_cf_pd_isRet = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  payload_3_cf_pred_taken = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  payload_3_cf_ftqPtr_flag = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  payload_3_cf_ftqPtr_value = _RAND_96[2:0];
  _RAND_97 = {1{`RANDOM}};
  payload_3_cf_ftqOffset = _RAND_97[2:0];
  _RAND_98 = {1{`RANDOM}};
  payload_3_ctrl_fuType = _RAND_98[3:0];
  _RAND_99 = {1{`RANDOM}};
  payload_3_ctrl_fuOpType = _RAND_99[6:0];
  _RAND_100 = {1{`RANDOM}};
  payload_3_ctrl_rfWen = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  payload_3_ctrl_fpWen = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  payload_3_ctrl_imm = _RAND_102[19:0];
  _RAND_103 = {1{`RANDOM}};
  payload_3_ctrl_fpu_isAddSub = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  payload_3_ctrl_fpu_typeTagIn = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  payload_3_ctrl_fpu_typeTagOut = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  payload_3_ctrl_fpu_fromInt = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  payload_3_ctrl_fpu_wflags = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  payload_3_ctrl_fpu_fpWen = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  payload_3_ctrl_fpu_fmaCmd = _RAND_109[1:0];
  _RAND_110 = {1{`RANDOM}};
  payload_3_ctrl_fpu_div = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  payload_3_ctrl_fpu_sqrt = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  payload_3_ctrl_fpu_fcvt = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  payload_3_ctrl_fpu_typ = _RAND_113[1:0];
  _RAND_114 = {1{`RANDOM}};
  payload_3_ctrl_fpu_fmt = _RAND_114[1:0];
  _RAND_115 = {1{`RANDOM}};
  payload_3_ctrl_fpu_ren3 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  payload_3_ctrl_fpu_rm = _RAND_116[2:0];
  _RAND_117 = {1{`RANDOM}};
  payload_3_pdest = _RAND_117[5:0];
  _RAND_118 = {1{`RANDOM}};
  payload_3_robIdx_flag = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  payload_3_robIdx_value = _RAND_119[4:0];
  _RAND_120 = {1{`RANDOM}};
  payload_4_cf_pd_isRVC = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  payload_4_cf_pd_brType = _RAND_121[1:0];
  _RAND_122 = {1{`RANDOM}};
  payload_4_cf_pd_isCall = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  payload_4_cf_pd_isRet = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  payload_4_cf_pred_taken = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  payload_4_cf_ftqPtr_flag = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  payload_4_cf_ftqPtr_value = _RAND_126[2:0];
  _RAND_127 = {1{`RANDOM}};
  payload_4_cf_ftqOffset = _RAND_127[2:0];
  _RAND_128 = {1{`RANDOM}};
  payload_4_ctrl_fuType = _RAND_128[3:0];
  _RAND_129 = {1{`RANDOM}};
  payload_4_ctrl_fuOpType = _RAND_129[6:0];
  _RAND_130 = {1{`RANDOM}};
  payload_4_ctrl_rfWen = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  payload_4_ctrl_fpWen = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  payload_4_ctrl_imm = _RAND_132[19:0];
  _RAND_133 = {1{`RANDOM}};
  payload_4_ctrl_fpu_isAddSub = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  payload_4_ctrl_fpu_typeTagIn = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  payload_4_ctrl_fpu_typeTagOut = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  payload_4_ctrl_fpu_fromInt = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  payload_4_ctrl_fpu_wflags = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  payload_4_ctrl_fpu_fpWen = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  payload_4_ctrl_fpu_fmaCmd = _RAND_139[1:0];
  _RAND_140 = {1{`RANDOM}};
  payload_4_ctrl_fpu_div = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  payload_4_ctrl_fpu_sqrt = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  payload_4_ctrl_fpu_fcvt = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  payload_4_ctrl_fpu_typ = _RAND_143[1:0];
  _RAND_144 = {1{`RANDOM}};
  payload_4_ctrl_fpu_fmt = _RAND_144[1:0];
  _RAND_145 = {1{`RANDOM}};
  payload_4_ctrl_fpu_ren3 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  payload_4_ctrl_fpu_rm = _RAND_146[2:0];
  _RAND_147 = {1{`RANDOM}};
  payload_4_pdest = _RAND_147[5:0];
  _RAND_148 = {1{`RANDOM}};
  payload_4_robIdx_flag = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  payload_4_robIdx_value = _RAND_149[4:0];
  _RAND_150 = {1{`RANDOM}};
  payload_5_cf_pd_isRVC = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  payload_5_cf_pd_brType = _RAND_151[1:0];
  _RAND_152 = {1{`RANDOM}};
  payload_5_cf_pd_isCall = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  payload_5_cf_pd_isRet = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  payload_5_cf_pred_taken = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  payload_5_cf_ftqPtr_flag = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  payload_5_cf_ftqPtr_value = _RAND_156[2:0];
  _RAND_157 = {1{`RANDOM}};
  payload_5_cf_ftqOffset = _RAND_157[2:0];
  _RAND_158 = {1{`RANDOM}};
  payload_5_ctrl_fuType = _RAND_158[3:0];
  _RAND_159 = {1{`RANDOM}};
  payload_5_ctrl_fuOpType = _RAND_159[6:0];
  _RAND_160 = {1{`RANDOM}};
  payload_5_ctrl_rfWen = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  payload_5_ctrl_fpWen = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  payload_5_ctrl_imm = _RAND_162[19:0];
  _RAND_163 = {1{`RANDOM}};
  payload_5_ctrl_fpu_isAddSub = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  payload_5_ctrl_fpu_typeTagIn = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  payload_5_ctrl_fpu_typeTagOut = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  payload_5_ctrl_fpu_fromInt = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  payload_5_ctrl_fpu_wflags = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  payload_5_ctrl_fpu_fpWen = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  payload_5_ctrl_fpu_fmaCmd = _RAND_169[1:0];
  _RAND_170 = {1{`RANDOM}};
  payload_5_ctrl_fpu_div = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  payload_5_ctrl_fpu_sqrt = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  payload_5_ctrl_fpu_fcvt = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  payload_5_ctrl_fpu_typ = _RAND_173[1:0];
  _RAND_174 = {1{`RANDOM}};
  payload_5_ctrl_fpu_fmt = _RAND_174[1:0];
  _RAND_175 = {1{`RANDOM}};
  payload_5_ctrl_fpu_ren3 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  payload_5_ctrl_fpu_rm = _RAND_176[2:0];
  _RAND_177 = {1{`RANDOM}};
  payload_5_pdest = _RAND_177[5:0];
  _RAND_178 = {1{`RANDOM}};
  payload_5_robIdx_flag = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  payload_5_robIdx_value = _RAND_179[4:0];
  _RAND_180 = {1{`RANDOM}};
  payload_6_cf_pd_isRVC = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  payload_6_cf_pd_brType = _RAND_181[1:0];
  _RAND_182 = {1{`RANDOM}};
  payload_6_cf_pd_isCall = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  payload_6_cf_pd_isRet = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  payload_6_cf_pred_taken = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  payload_6_cf_ftqPtr_flag = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  payload_6_cf_ftqPtr_value = _RAND_186[2:0];
  _RAND_187 = {1{`RANDOM}};
  payload_6_cf_ftqOffset = _RAND_187[2:0];
  _RAND_188 = {1{`RANDOM}};
  payload_6_ctrl_fuType = _RAND_188[3:0];
  _RAND_189 = {1{`RANDOM}};
  payload_6_ctrl_fuOpType = _RAND_189[6:0];
  _RAND_190 = {1{`RANDOM}};
  payload_6_ctrl_rfWen = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  payload_6_ctrl_fpWen = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  payload_6_ctrl_imm = _RAND_192[19:0];
  _RAND_193 = {1{`RANDOM}};
  payload_6_ctrl_fpu_isAddSub = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  payload_6_ctrl_fpu_typeTagIn = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  payload_6_ctrl_fpu_typeTagOut = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  payload_6_ctrl_fpu_fromInt = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  payload_6_ctrl_fpu_wflags = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  payload_6_ctrl_fpu_fpWen = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  payload_6_ctrl_fpu_fmaCmd = _RAND_199[1:0];
  _RAND_200 = {1{`RANDOM}};
  payload_6_ctrl_fpu_div = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  payload_6_ctrl_fpu_sqrt = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  payload_6_ctrl_fpu_fcvt = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  payload_6_ctrl_fpu_typ = _RAND_203[1:0];
  _RAND_204 = {1{`RANDOM}};
  payload_6_ctrl_fpu_fmt = _RAND_204[1:0];
  _RAND_205 = {1{`RANDOM}};
  payload_6_ctrl_fpu_ren3 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  payload_6_ctrl_fpu_rm = _RAND_206[2:0];
  _RAND_207 = {1{`RANDOM}};
  payload_6_pdest = _RAND_207[5:0];
  _RAND_208 = {1{`RANDOM}};
  payload_6_robIdx_flag = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  payload_6_robIdx_value = _RAND_209[4:0];
  _RAND_210 = {1{`RANDOM}};
  payload_7_cf_pd_isRVC = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  payload_7_cf_pd_brType = _RAND_211[1:0];
  _RAND_212 = {1{`RANDOM}};
  payload_7_cf_pd_isCall = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  payload_7_cf_pd_isRet = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  payload_7_cf_pred_taken = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  payload_7_cf_ftqPtr_flag = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  payload_7_cf_ftqPtr_value = _RAND_216[2:0];
  _RAND_217 = {1{`RANDOM}};
  payload_7_cf_ftqOffset = _RAND_217[2:0];
  _RAND_218 = {1{`RANDOM}};
  payload_7_ctrl_fuType = _RAND_218[3:0];
  _RAND_219 = {1{`RANDOM}};
  payload_7_ctrl_fuOpType = _RAND_219[6:0];
  _RAND_220 = {1{`RANDOM}};
  payload_7_ctrl_rfWen = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  payload_7_ctrl_fpWen = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  payload_7_ctrl_imm = _RAND_222[19:0];
  _RAND_223 = {1{`RANDOM}};
  payload_7_ctrl_fpu_isAddSub = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  payload_7_ctrl_fpu_typeTagIn = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  payload_7_ctrl_fpu_typeTagOut = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  payload_7_ctrl_fpu_fromInt = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  payload_7_ctrl_fpu_wflags = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  payload_7_ctrl_fpu_fpWen = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  payload_7_ctrl_fpu_fmaCmd = _RAND_229[1:0];
  _RAND_230 = {1{`RANDOM}};
  payload_7_ctrl_fpu_div = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  payload_7_ctrl_fpu_sqrt = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  payload_7_ctrl_fpu_fcvt = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  payload_7_ctrl_fpu_typ = _RAND_233[1:0];
  _RAND_234 = {1{`RANDOM}};
  payload_7_ctrl_fpu_fmt = _RAND_234[1:0];
  _RAND_235 = {1{`RANDOM}};
  payload_7_ctrl_fpu_ren3 = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  payload_7_ctrl_fpu_rm = _RAND_236[2:0];
  _RAND_237 = {1{`RANDOM}};
  payload_7_pdest = _RAND_237[5:0];
  _RAND_238 = {1{`RANDOM}};
  payload_7_robIdx_flag = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  payload_7_robIdx_value = _RAND_239[4:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule

