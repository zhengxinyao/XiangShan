module BankedAsyncDataModuleTemplateWithDup(
  input         clock,
  input  [3:0]  io_raddr_0,
  input  [3:0]  io_raddr_1,
  output [26:0] io_rdata_0_0_tag,
  output [15:0] io_rdata_0_0_asid,
  output [23:0] io_rdata_0_0_ppn,
  output        io_rdata_0_0_perm_pf,
  output        io_rdata_0_0_perm_af,
  output        io_rdata_0_0_perm_d,
  output        io_rdata_0_0_perm_a,
  output        io_rdata_0_0_perm_u,
  output        io_rdata_0_0_perm_x,
  output        io_rdata_0_0_perm_w,
  output        io_rdata_0_0_perm_r,
  output        io_rdata_0_0_perm_pm_r,
  output        io_rdata_0_0_perm_pm_w,
  output        io_rdata_0_0_perm_pm_c,
  output [23:0] io_rdata_0_1_ppn,
  output [26:0] io_rdata_1_0_tag,
  output [15:0] io_rdata_1_0_asid,
  output [23:0] io_rdata_1_0_ppn,
  output        io_rdata_1_0_perm_pf,
  output        io_rdata_1_0_perm_af,
  output        io_rdata_1_0_perm_a,
  output        io_rdata_1_0_perm_u,
  output        io_rdata_1_0_perm_x,
  output        io_rdata_1_0_perm_r,
  output        io_rdata_1_0_perm_pm_r,
  output        io_rdata_1_0_perm_pm_c,
  output [23:0] io_rdata_1_1_ppn,
  input         io_wen,
  input  [3:0]  io_waddr,
  input  [26:0] io_wdata_tag,
  input  [15:0] io_wdata_asid,
  input  [23:0] io_wdata_ppn,
  input         io_wdata_perm_pf,
  input         io_wdata_perm_af,
  input         io_wdata_perm_d,
  input         io_wdata_perm_a,
  input         io_wdata_perm_u,
  input         io_wdata_perm_x,
  input         io_wdata_perm_w,
  input         io_wdata_perm_r,
  input         io_wdata_perm_pm_r,
  input         io_wdata_perm_pm_w,
  input         io_wdata_perm_pm_c
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
`endif // RANDOMIZE_REG_INIT
  reg [26:0] dataBanks_0_tag [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_tag_data_read_0_0_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_tag_data_read_0_0_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire [26:0] dataBanks_0_tag_data_read_0_0_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_tag_data_read_1_0_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_tag_data_read_1_0_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire [26:0] dataBanks_0_tag_data_read_1_0_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_tag_data_read_0_0_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_tag_data_read_0_0_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire [26:0] dataBanks_0_tag_data_read_0_0_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_tag_data_read_1_0_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_tag_data_read_1_0_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire [26:0] dataBanks_0_tag_data_read_1_0_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire [26:0] dataBanks_0_tag_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_tag_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_tag_MPORT_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_tag_MPORT_en; // @[TLBStorage.scala 58:8]
  reg [15:0] dataBanks_0_asid [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_asid_data_read_0_0_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_asid_data_read_0_0_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire [15:0] dataBanks_0_asid_data_read_0_0_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_asid_data_read_1_0_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_asid_data_read_1_0_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire [15:0] dataBanks_0_asid_data_read_1_0_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_asid_data_read_0_0_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_asid_data_read_0_0_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire [15:0] dataBanks_0_asid_data_read_0_0_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_asid_data_read_1_0_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_asid_data_read_1_0_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire [15:0] dataBanks_0_asid_data_read_1_0_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire [15:0] dataBanks_0_asid_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_asid_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_asid_MPORT_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_asid_MPORT_en; // @[TLBStorage.scala 58:8]
  reg [23:0] dataBanks_0_ppn [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_ppn_data_read_0_0_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_ppn_data_read_0_0_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire [23:0] dataBanks_0_ppn_data_read_0_0_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_ppn_data_read_1_0_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_ppn_data_read_1_0_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire [23:0] dataBanks_0_ppn_data_read_1_0_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_ppn_data_read_0_0_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_ppn_data_read_0_0_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire [23:0] dataBanks_0_ppn_data_read_0_0_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_ppn_data_read_1_0_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_ppn_data_read_1_0_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire [23:0] dataBanks_0_ppn_data_read_1_0_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire [23:0] dataBanks_0_ppn_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_ppn_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_ppn_MPORT_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_ppn_MPORT_en; // @[TLBStorage.scala 58:8]
  reg  dataBanks_0_perm_pf [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_pf_data_read_0_0_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_pf_data_read_0_0_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_pf_data_read_0_0_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_pf_data_read_1_0_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_pf_data_read_1_0_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_pf_data_read_1_0_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_pf_data_read_0_0_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_pf_data_read_0_0_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_pf_data_read_0_0_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_pf_data_read_1_0_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_pf_data_read_1_0_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_pf_data_read_1_0_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_pf_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_pf_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_pf_MPORT_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_pf_MPORT_en; // @[TLBStorage.scala 58:8]
  reg  dataBanks_0_perm_af [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_af_data_read_0_0_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_af_data_read_0_0_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_af_data_read_0_0_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_af_data_read_1_0_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_af_data_read_1_0_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_af_data_read_1_0_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_af_data_read_0_0_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_af_data_read_0_0_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_af_data_read_0_0_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_af_data_read_1_0_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_af_data_read_1_0_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_af_data_read_1_0_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_af_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_af_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_af_MPORT_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_af_MPORT_en; // @[TLBStorage.scala 58:8]
  reg  dataBanks_0_perm_d [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_d_data_read_0_0_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_d_data_read_0_0_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_d_data_read_0_0_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_d_data_read_1_0_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_d_data_read_1_0_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_d_data_read_1_0_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_d_data_read_0_0_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_d_data_read_0_0_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_d_data_read_0_0_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_d_data_read_1_0_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_d_data_read_1_0_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_d_data_read_1_0_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_d_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_d_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_d_MPORT_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_d_MPORT_en; // @[TLBStorage.scala 58:8]
  reg  dataBanks_0_perm_a [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_a_data_read_0_0_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_a_data_read_0_0_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_a_data_read_0_0_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_a_data_read_1_0_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_a_data_read_1_0_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_a_data_read_1_0_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_a_data_read_0_0_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_a_data_read_0_0_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_a_data_read_0_0_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_a_data_read_1_0_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_a_data_read_1_0_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_a_data_read_1_0_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_a_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_a_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_a_MPORT_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_a_MPORT_en; // @[TLBStorage.scala 58:8]
  reg  dataBanks_0_perm_u [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_u_data_read_0_0_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_u_data_read_0_0_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_u_data_read_0_0_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_u_data_read_1_0_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_u_data_read_1_0_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_u_data_read_1_0_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_u_data_read_0_0_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_u_data_read_0_0_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_u_data_read_0_0_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_u_data_read_1_0_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_u_data_read_1_0_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_u_data_read_1_0_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_u_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_u_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_u_MPORT_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_u_MPORT_en; // @[TLBStorage.scala 58:8]
  reg  dataBanks_0_perm_x [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_x_data_read_0_0_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_x_data_read_0_0_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_x_data_read_0_0_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_x_data_read_1_0_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_x_data_read_1_0_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_x_data_read_1_0_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_x_data_read_0_0_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_x_data_read_0_0_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_x_data_read_0_0_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_x_data_read_1_0_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_x_data_read_1_0_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_x_data_read_1_0_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_x_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_x_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_x_MPORT_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_x_MPORT_en; // @[TLBStorage.scala 58:8]
  reg  dataBanks_0_perm_w [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_wdata_read_0_0_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_wdata_read_0_0_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_wdata_read_0_0_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_wdata_read_1_0_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_wdata_read_1_0_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_wdata_read_1_0_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_wdata_read_0_0_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_wdata_read_0_0_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_wdata_read_0_0_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_wdata_read_1_0_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_wdata_read_1_0_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_wdata_read_1_0_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_wMPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_wMPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_wMPORT_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_wMPORT_en; // @[TLBStorage.scala 58:8]
  reg  dataBanks_0_perm_r [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_rdata_read_0_0_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_rdata_read_0_0_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_rdata_read_0_0_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_rdata_read_1_0_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_rdata_read_1_0_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_rdata_read_1_0_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_rdata_read_0_0_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_rdata_read_0_0_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_rdata_read_0_0_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_rdata_read_1_0_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_rdata_read_1_0_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_rdata_read_1_0_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_rMPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_rMPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_rMPORT_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_rMPORT_en; // @[TLBStorage.scala 58:8]
  reg  dataBanks_0_perm_pm_r [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_pm_rdata_read_0_0_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_pm_rdata_read_0_0_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_pm_rdata_read_0_0_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_pm_rdata_read_1_0_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_pm_rdata_read_1_0_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_pm_rdata_read_1_0_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_pm_rdata_read_0_0_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_pm_rdata_read_0_0_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_pm_rdata_read_0_0_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_pm_rdata_read_1_0_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_pm_rdata_read_1_0_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_pm_rdata_read_1_0_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_pm_rMPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_pm_rMPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_pm_rMPORT_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_pm_rMPORT_en; // @[TLBStorage.scala 58:8]
  reg  dataBanks_0_perm_pm_w [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_pm_wdata_read_0_0_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_pm_wdata_read_0_0_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_pm_wdata_read_0_0_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_pm_wdata_read_1_0_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_pm_wdata_read_1_0_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_pm_wdata_read_1_0_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_pm_wdata_read_0_0_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_pm_wdata_read_0_0_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_pm_wdata_read_0_0_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_pm_wdata_read_1_0_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_pm_wdata_read_1_0_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_pm_wdata_read_1_0_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_pm_wMPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_pm_wMPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_pm_wMPORT_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_pm_wMPORT_en; // @[TLBStorage.scala 58:8]
  reg  dataBanks_0_perm_pm_c [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_pm_c_data_read_0_0_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_pm_c_data_read_0_0_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_pm_c_data_read_0_0_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_pm_c_data_read_1_0_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_pm_c_data_read_1_0_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_pm_c_data_read_1_0_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_pm_c_data_read_0_0_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_pm_c_data_read_0_0_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_pm_c_data_read_0_0_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_pm_c_data_read_1_0_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_pm_c_data_read_1_0_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_pm_c_data_read_1_0_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_pm_c_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_pm_c_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_pm_c_MPORT_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_0_perm_pm_c_MPORT_en; // @[TLBStorage.scala 58:8]
  reg [26:0] dataBanks_1_tag [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_tag_data_read_0_1_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_tag_data_read_0_1_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire [26:0] dataBanks_1_tag_data_read_0_1_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_tag_data_read_1_1_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_tag_data_read_1_1_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire [26:0] dataBanks_1_tag_data_read_1_1_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_tag_data_read_0_1_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_tag_data_read_0_1_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire [26:0] dataBanks_1_tag_data_read_0_1_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_tag_data_read_1_1_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_tag_data_read_1_1_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire [26:0] dataBanks_1_tag_data_read_1_1_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire [26:0] dataBanks_1_tag_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_tag_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_tag_MPORT_1_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_tag_MPORT_1_en; // @[TLBStorage.scala 58:8]
  reg [15:0] dataBanks_1_asid [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_asid_data_read_0_1_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_asid_data_read_0_1_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire [15:0] dataBanks_1_asid_data_read_0_1_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_asid_data_read_1_1_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_asid_data_read_1_1_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire [15:0] dataBanks_1_asid_data_read_1_1_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_asid_data_read_0_1_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_asid_data_read_0_1_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire [15:0] dataBanks_1_asid_data_read_0_1_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_asid_data_read_1_1_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_asid_data_read_1_1_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire [15:0] dataBanks_1_asid_data_read_1_1_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire [15:0] dataBanks_1_asid_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_asid_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_asid_MPORT_1_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_asid_MPORT_1_en; // @[TLBStorage.scala 58:8]
  reg [23:0] dataBanks_1_ppn [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_ppn_data_read_0_1_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_ppn_data_read_0_1_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire [23:0] dataBanks_1_ppn_data_read_0_1_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_ppn_data_read_1_1_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_ppn_data_read_1_1_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire [23:0] dataBanks_1_ppn_data_read_1_1_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_ppn_data_read_0_1_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_ppn_data_read_0_1_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire [23:0] dataBanks_1_ppn_data_read_0_1_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_ppn_data_read_1_1_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_ppn_data_read_1_1_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire [23:0] dataBanks_1_ppn_data_read_1_1_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire [23:0] dataBanks_1_ppn_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_ppn_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_ppn_MPORT_1_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_ppn_MPORT_1_en; // @[TLBStorage.scala 58:8]
  reg  dataBanks_1_perm_pf [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_pf_data_read_0_1_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_pf_data_read_0_1_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_pf_data_read_0_1_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_pf_data_read_1_1_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_pf_data_read_1_1_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_pf_data_read_1_1_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_pf_data_read_0_1_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_pf_data_read_0_1_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_pf_data_read_0_1_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_pf_data_read_1_1_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_pf_data_read_1_1_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_pf_data_read_1_1_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_pf_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_pf_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_pf_MPORT_1_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_pf_MPORT_1_en; // @[TLBStorage.scala 58:8]
  reg  dataBanks_1_perm_af [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_af_data_read_0_1_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_af_data_read_0_1_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_af_data_read_0_1_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_af_data_read_1_1_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_af_data_read_1_1_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_af_data_read_1_1_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_af_data_read_0_1_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_af_data_read_0_1_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_af_data_read_0_1_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_af_data_read_1_1_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_af_data_read_1_1_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_af_data_read_1_1_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_af_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_af_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_af_MPORT_1_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_af_MPORT_1_en; // @[TLBStorage.scala 58:8]
  reg  dataBanks_1_perm_d [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_d_data_read_0_1_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_d_data_read_0_1_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_d_data_read_0_1_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_d_data_read_1_1_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_d_data_read_1_1_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_d_data_read_1_1_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_d_data_read_0_1_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_d_data_read_0_1_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_d_data_read_0_1_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_d_data_read_1_1_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_d_data_read_1_1_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_d_data_read_1_1_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_d_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_d_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_d_MPORT_1_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_d_MPORT_1_en; // @[TLBStorage.scala 58:8]
  reg  dataBanks_1_perm_a [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_a_data_read_0_1_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_a_data_read_0_1_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_a_data_read_0_1_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_a_data_read_1_1_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_a_data_read_1_1_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_a_data_read_1_1_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_a_data_read_0_1_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_a_data_read_0_1_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_a_data_read_0_1_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_a_data_read_1_1_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_a_data_read_1_1_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_a_data_read_1_1_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_a_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_a_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_a_MPORT_1_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_a_MPORT_1_en; // @[TLBStorage.scala 58:8]
  reg  dataBanks_1_perm_u [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_u_data_read_0_1_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_u_data_read_0_1_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_u_data_read_0_1_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_u_data_read_1_1_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_u_data_read_1_1_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_u_data_read_1_1_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_u_data_read_0_1_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_u_data_read_0_1_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_u_data_read_0_1_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_u_data_read_1_1_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_u_data_read_1_1_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_u_data_read_1_1_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_u_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_u_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_u_MPORT_1_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_u_MPORT_1_en; // @[TLBStorage.scala 58:8]
  reg  dataBanks_1_perm_x [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_x_data_read_0_1_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_x_data_read_0_1_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_x_data_read_0_1_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_x_data_read_1_1_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_x_data_read_1_1_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_x_data_read_1_1_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_x_data_read_0_1_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_x_data_read_0_1_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_x_data_read_0_1_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_x_data_read_1_1_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_x_data_read_1_1_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_x_data_read_1_1_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_x_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_x_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_x_MPORT_1_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_x_MPORT_1_en; // @[TLBStorage.scala 58:8]
  reg  dataBanks_1_perm_w [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_wdata_read_0_1_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_wdata_read_0_1_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_wdata_read_0_1_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_wdata_read_1_1_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_wdata_read_1_1_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_wdata_read_1_1_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_wdata_read_0_1_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_wdata_read_0_1_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_wdata_read_0_1_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_wdata_read_1_1_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_wdata_read_1_1_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_wdata_read_1_1_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_wMPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_wMPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_wMPORT_1_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_wMPORT_1_en; // @[TLBStorage.scala 58:8]
  reg  dataBanks_1_perm_r [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_rdata_read_0_1_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_rdata_read_0_1_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_rdata_read_0_1_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_rdata_read_1_1_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_rdata_read_1_1_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_rdata_read_1_1_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_rdata_read_0_1_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_rdata_read_0_1_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_rdata_read_0_1_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_rdata_read_1_1_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_rdata_read_1_1_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_rdata_read_1_1_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_rMPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_rMPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_rMPORT_1_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_rMPORT_1_en; // @[TLBStorage.scala 58:8]
  reg  dataBanks_1_perm_pm_r [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_pm_rdata_read_0_1_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_pm_rdata_read_0_1_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_pm_rdata_read_0_1_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_pm_rdata_read_1_1_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_pm_rdata_read_1_1_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_pm_rdata_read_1_1_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_pm_rdata_read_0_1_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_pm_rdata_read_0_1_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_pm_rdata_read_0_1_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_pm_rdata_read_1_1_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_pm_rdata_read_1_1_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_pm_rdata_read_1_1_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_pm_rMPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_pm_rMPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_pm_rMPORT_1_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_pm_rMPORT_1_en; // @[TLBStorage.scala 58:8]
  reg  dataBanks_1_perm_pm_w [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_pm_wdata_read_0_1_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_pm_wdata_read_0_1_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_pm_wdata_read_0_1_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_pm_wdata_read_1_1_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_pm_wdata_read_1_1_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_pm_wdata_read_1_1_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_pm_wdata_read_0_1_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_pm_wdata_read_0_1_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_pm_wdata_read_0_1_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_pm_wdata_read_1_1_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_pm_wdata_read_1_1_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_pm_wdata_read_1_1_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_pm_wMPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_pm_wMPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_pm_wMPORT_1_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_pm_wMPORT_1_en; // @[TLBStorage.scala 58:8]
  reg  dataBanks_1_perm_pm_c [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_pm_c_data_read_0_1_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_pm_c_data_read_0_1_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_pm_c_data_read_0_1_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_pm_c_data_read_1_1_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_pm_c_data_read_1_1_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_pm_c_data_read_1_1_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_pm_c_data_read_0_1_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_pm_c_data_read_0_1_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_pm_c_data_read_0_1_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_pm_c_data_read_1_1_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_pm_c_data_read_1_1_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_pm_c_data_read_1_1_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_pm_c_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_pm_c_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_pm_c_MPORT_1_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_1_perm_pm_c_MPORT_1_en; // @[TLBStorage.scala 58:8]
  reg [26:0] dataBanks_2_tag [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_tag_data_read_0_2_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_tag_data_read_0_2_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire [26:0] dataBanks_2_tag_data_read_0_2_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_tag_data_read_1_2_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_tag_data_read_1_2_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire [26:0] dataBanks_2_tag_data_read_1_2_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_tag_data_read_0_2_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_tag_data_read_0_2_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire [26:0] dataBanks_2_tag_data_read_0_2_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_tag_data_read_1_2_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_tag_data_read_1_2_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire [26:0] dataBanks_2_tag_data_read_1_2_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire [26:0] dataBanks_2_tag_MPORT_2_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_tag_MPORT_2_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_tag_MPORT_2_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_tag_MPORT_2_en; // @[TLBStorage.scala 58:8]
  reg [15:0] dataBanks_2_asid [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_asid_data_read_0_2_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_asid_data_read_0_2_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire [15:0] dataBanks_2_asid_data_read_0_2_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_asid_data_read_1_2_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_asid_data_read_1_2_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire [15:0] dataBanks_2_asid_data_read_1_2_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_asid_data_read_0_2_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_asid_data_read_0_2_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire [15:0] dataBanks_2_asid_data_read_0_2_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_asid_data_read_1_2_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_asid_data_read_1_2_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire [15:0] dataBanks_2_asid_data_read_1_2_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire [15:0] dataBanks_2_asid_MPORT_2_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_asid_MPORT_2_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_asid_MPORT_2_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_asid_MPORT_2_en; // @[TLBStorage.scala 58:8]
  reg [23:0] dataBanks_2_ppn [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_ppn_data_read_0_2_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_ppn_data_read_0_2_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire [23:0] dataBanks_2_ppn_data_read_0_2_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_ppn_data_read_1_2_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_ppn_data_read_1_2_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire [23:0] dataBanks_2_ppn_data_read_1_2_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_ppn_data_read_0_2_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_ppn_data_read_0_2_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire [23:0] dataBanks_2_ppn_data_read_0_2_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_ppn_data_read_1_2_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_ppn_data_read_1_2_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire [23:0] dataBanks_2_ppn_data_read_1_2_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire [23:0] dataBanks_2_ppn_MPORT_2_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_ppn_MPORT_2_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_ppn_MPORT_2_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_ppn_MPORT_2_en; // @[TLBStorage.scala 58:8]
  reg  dataBanks_2_perm_pf [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_pf_data_read_0_2_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_pf_data_read_0_2_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_pf_data_read_0_2_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_pf_data_read_1_2_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_pf_data_read_1_2_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_pf_data_read_1_2_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_pf_data_read_0_2_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_pf_data_read_0_2_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_pf_data_read_0_2_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_pf_data_read_1_2_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_pf_data_read_1_2_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_pf_data_read_1_2_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_pf_MPORT_2_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_pf_MPORT_2_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_pf_MPORT_2_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_pf_MPORT_2_en; // @[TLBStorage.scala 58:8]
  reg  dataBanks_2_perm_af [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_af_data_read_0_2_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_af_data_read_0_2_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_af_data_read_0_2_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_af_data_read_1_2_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_af_data_read_1_2_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_af_data_read_1_2_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_af_data_read_0_2_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_af_data_read_0_2_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_af_data_read_0_2_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_af_data_read_1_2_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_af_data_read_1_2_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_af_data_read_1_2_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_af_MPORT_2_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_af_MPORT_2_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_af_MPORT_2_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_af_MPORT_2_en; // @[TLBStorage.scala 58:8]
  reg  dataBanks_2_perm_d [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_d_data_read_0_2_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_d_data_read_0_2_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_d_data_read_0_2_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_d_data_read_1_2_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_d_data_read_1_2_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_d_data_read_1_2_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_d_data_read_0_2_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_d_data_read_0_2_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_d_data_read_0_2_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_d_data_read_1_2_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_d_data_read_1_2_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_d_data_read_1_2_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_d_MPORT_2_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_d_MPORT_2_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_d_MPORT_2_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_d_MPORT_2_en; // @[TLBStorage.scala 58:8]
  reg  dataBanks_2_perm_a [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_a_data_read_0_2_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_a_data_read_0_2_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_a_data_read_0_2_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_a_data_read_1_2_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_a_data_read_1_2_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_a_data_read_1_2_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_a_data_read_0_2_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_a_data_read_0_2_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_a_data_read_0_2_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_a_data_read_1_2_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_a_data_read_1_2_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_a_data_read_1_2_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_a_MPORT_2_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_a_MPORT_2_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_a_MPORT_2_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_a_MPORT_2_en; // @[TLBStorage.scala 58:8]
  reg  dataBanks_2_perm_u [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_u_data_read_0_2_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_u_data_read_0_2_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_u_data_read_0_2_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_u_data_read_1_2_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_u_data_read_1_2_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_u_data_read_1_2_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_u_data_read_0_2_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_u_data_read_0_2_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_u_data_read_0_2_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_u_data_read_1_2_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_u_data_read_1_2_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_u_data_read_1_2_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_u_MPORT_2_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_u_MPORT_2_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_u_MPORT_2_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_u_MPORT_2_en; // @[TLBStorage.scala 58:8]
  reg  dataBanks_2_perm_x [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_x_data_read_0_2_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_x_data_read_0_2_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_x_data_read_0_2_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_x_data_read_1_2_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_x_data_read_1_2_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_x_data_read_1_2_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_x_data_read_0_2_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_x_data_read_0_2_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_x_data_read_0_2_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_x_data_read_1_2_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_x_data_read_1_2_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_x_data_read_1_2_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_x_MPORT_2_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_x_MPORT_2_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_x_MPORT_2_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_x_MPORT_2_en; // @[TLBStorage.scala 58:8]
  reg  dataBanks_2_perm_w [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_wdata_read_0_2_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_wdata_read_0_2_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_wdata_read_0_2_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_wdata_read_1_2_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_wdata_read_1_2_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_wdata_read_1_2_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_wdata_read_0_2_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_wdata_read_0_2_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_wdata_read_0_2_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_wdata_read_1_2_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_wdata_read_1_2_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_wdata_read_1_2_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_wMPORT_2_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_wMPORT_2_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_wMPORT_2_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_wMPORT_2_en; // @[TLBStorage.scala 58:8]
  reg  dataBanks_2_perm_r [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_rdata_read_0_2_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_rdata_read_0_2_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_rdata_read_0_2_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_rdata_read_1_2_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_rdata_read_1_2_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_rdata_read_1_2_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_rdata_read_0_2_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_rdata_read_0_2_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_rdata_read_0_2_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_rdata_read_1_2_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_rdata_read_1_2_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_rdata_read_1_2_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_rMPORT_2_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_rMPORT_2_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_rMPORT_2_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_rMPORT_2_en; // @[TLBStorage.scala 58:8]
  reg  dataBanks_2_perm_pm_r [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_pm_rdata_read_0_2_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_pm_rdata_read_0_2_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_pm_rdata_read_0_2_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_pm_rdata_read_1_2_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_pm_rdata_read_1_2_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_pm_rdata_read_1_2_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_pm_rdata_read_0_2_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_pm_rdata_read_0_2_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_pm_rdata_read_0_2_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_pm_rdata_read_1_2_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_pm_rdata_read_1_2_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_pm_rdata_read_1_2_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_pm_rMPORT_2_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_pm_rMPORT_2_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_pm_rMPORT_2_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_pm_rMPORT_2_en; // @[TLBStorage.scala 58:8]
  reg  dataBanks_2_perm_pm_w [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_pm_wdata_read_0_2_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_pm_wdata_read_0_2_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_pm_wdata_read_0_2_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_pm_wdata_read_1_2_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_pm_wdata_read_1_2_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_pm_wdata_read_1_2_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_pm_wdata_read_0_2_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_pm_wdata_read_0_2_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_pm_wdata_read_0_2_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_pm_wdata_read_1_2_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_pm_wdata_read_1_2_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_pm_wdata_read_1_2_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_pm_wMPORT_2_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_pm_wMPORT_2_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_pm_wMPORT_2_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_pm_wMPORT_2_en; // @[TLBStorage.scala 58:8]
  reg  dataBanks_2_perm_pm_c [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_pm_c_data_read_0_2_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_pm_c_data_read_0_2_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_pm_c_data_read_0_2_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_pm_c_data_read_1_2_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_pm_c_data_read_1_2_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_pm_c_data_read_1_2_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_pm_c_data_read_0_2_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_pm_c_data_read_0_2_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_pm_c_data_read_0_2_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_pm_c_data_read_1_2_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_pm_c_data_read_1_2_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_pm_c_data_read_1_2_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_pm_c_MPORT_2_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_pm_c_MPORT_2_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_pm_c_MPORT_2_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_2_perm_pm_c_MPORT_2_en; // @[TLBStorage.scala 58:8]
  reg [26:0] dataBanks_3_tag [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_tag_data_read_0_3_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_tag_data_read_0_3_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire [26:0] dataBanks_3_tag_data_read_0_3_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_tag_data_read_1_3_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_tag_data_read_1_3_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire [26:0] dataBanks_3_tag_data_read_1_3_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_tag_data_read_0_3_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_tag_data_read_0_3_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire [26:0] dataBanks_3_tag_data_read_0_3_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_tag_data_read_1_3_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_tag_data_read_1_3_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire [26:0] dataBanks_3_tag_data_read_1_3_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire [26:0] dataBanks_3_tag_MPORT_3_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_tag_MPORT_3_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_tag_MPORT_3_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_tag_MPORT_3_en; // @[TLBStorage.scala 58:8]
  reg [15:0] dataBanks_3_asid [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_asid_data_read_0_3_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_asid_data_read_0_3_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire [15:0] dataBanks_3_asid_data_read_0_3_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_asid_data_read_1_3_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_asid_data_read_1_3_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire [15:0] dataBanks_3_asid_data_read_1_3_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_asid_data_read_0_3_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_asid_data_read_0_3_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire [15:0] dataBanks_3_asid_data_read_0_3_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_asid_data_read_1_3_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_asid_data_read_1_3_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire [15:0] dataBanks_3_asid_data_read_1_3_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire [15:0] dataBanks_3_asid_MPORT_3_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_asid_MPORT_3_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_asid_MPORT_3_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_asid_MPORT_3_en; // @[TLBStorage.scala 58:8]
  reg [23:0] dataBanks_3_ppn [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_ppn_data_read_0_3_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_ppn_data_read_0_3_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire [23:0] dataBanks_3_ppn_data_read_0_3_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_ppn_data_read_1_3_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_ppn_data_read_1_3_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire [23:0] dataBanks_3_ppn_data_read_1_3_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_ppn_data_read_0_3_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_ppn_data_read_0_3_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire [23:0] dataBanks_3_ppn_data_read_0_3_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_ppn_data_read_1_3_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_ppn_data_read_1_3_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire [23:0] dataBanks_3_ppn_data_read_1_3_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire [23:0] dataBanks_3_ppn_MPORT_3_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_ppn_MPORT_3_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_ppn_MPORT_3_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_ppn_MPORT_3_en; // @[TLBStorage.scala 58:8]
  reg  dataBanks_3_perm_pf [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_pf_data_read_0_3_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_pf_data_read_0_3_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_pf_data_read_0_3_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_pf_data_read_1_3_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_pf_data_read_1_3_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_pf_data_read_1_3_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_pf_data_read_0_3_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_pf_data_read_0_3_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_pf_data_read_0_3_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_pf_data_read_1_3_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_pf_data_read_1_3_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_pf_data_read_1_3_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_pf_MPORT_3_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_pf_MPORT_3_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_pf_MPORT_3_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_pf_MPORT_3_en; // @[TLBStorage.scala 58:8]
  reg  dataBanks_3_perm_af [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_af_data_read_0_3_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_af_data_read_0_3_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_af_data_read_0_3_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_af_data_read_1_3_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_af_data_read_1_3_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_af_data_read_1_3_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_af_data_read_0_3_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_af_data_read_0_3_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_af_data_read_0_3_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_af_data_read_1_3_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_af_data_read_1_3_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_af_data_read_1_3_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_af_MPORT_3_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_af_MPORT_3_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_af_MPORT_3_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_af_MPORT_3_en; // @[TLBStorage.scala 58:8]
  reg  dataBanks_3_perm_d [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_d_data_read_0_3_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_d_data_read_0_3_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_d_data_read_0_3_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_d_data_read_1_3_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_d_data_read_1_3_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_d_data_read_1_3_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_d_data_read_0_3_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_d_data_read_0_3_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_d_data_read_0_3_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_d_data_read_1_3_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_d_data_read_1_3_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_d_data_read_1_3_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_d_MPORT_3_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_d_MPORT_3_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_d_MPORT_3_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_d_MPORT_3_en; // @[TLBStorage.scala 58:8]
  reg  dataBanks_3_perm_a [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_a_data_read_0_3_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_a_data_read_0_3_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_a_data_read_0_3_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_a_data_read_1_3_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_a_data_read_1_3_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_a_data_read_1_3_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_a_data_read_0_3_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_a_data_read_0_3_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_a_data_read_0_3_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_a_data_read_1_3_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_a_data_read_1_3_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_a_data_read_1_3_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_a_MPORT_3_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_a_MPORT_3_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_a_MPORT_3_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_a_MPORT_3_en; // @[TLBStorage.scala 58:8]
  reg  dataBanks_3_perm_u [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_u_data_read_0_3_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_u_data_read_0_3_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_u_data_read_0_3_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_u_data_read_1_3_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_u_data_read_1_3_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_u_data_read_1_3_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_u_data_read_0_3_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_u_data_read_0_3_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_u_data_read_0_3_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_u_data_read_1_3_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_u_data_read_1_3_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_u_data_read_1_3_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_u_MPORT_3_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_u_MPORT_3_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_u_MPORT_3_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_u_MPORT_3_en; // @[TLBStorage.scala 58:8]
  reg  dataBanks_3_perm_x [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_x_data_read_0_3_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_x_data_read_0_3_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_x_data_read_0_3_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_x_data_read_1_3_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_x_data_read_1_3_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_x_data_read_1_3_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_x_data_read_0_3_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_x_data_read_0_3_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_x_data_read_0_3_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_x_data_read_1_3_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_x_data_read_1_3_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_x_data_read_1_3_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_x_MPORT_3_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_x_MPORT_3_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_x_MPORT_3_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_x_MPORT_3_en; // @[TLBStorage.scala 58:8]
  reg  dataBanks_3_perm_w [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_wdata_read_0_3_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_wdata_read_0_3_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_wdata_read_0_3_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_wdata_read_1_3_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_wdata_read_1_3_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_wdata_read_1_3_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_wdata_read_0_3_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_wdata_read_0_3_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_wdata_read_0_3_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_wdata_read_1_3_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_wdata_read_1_3_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_wdata_read_1_3_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_wMPORT_3_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_wMPORT_3_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_wMPORT_3_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_wMPORT_3_en; // @[TLBStorage.scala 58:8]
  reg  dataBanks_3_perm_r [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_rdata_read_0_3_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_rdata_read_0_3_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_rdata_read_0_3_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_rdata_read_1_3_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_rdata_read_1_3_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_rdata_read_1_3_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_rdata_read_0_3_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_rdata_read_0_3_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_rdata_read_0_3_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_rdata_read_1_3_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_rdata_read_1_3_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_rdata_read_1_3_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_rMPORT_3_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_rMPORT_3_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_rMPORT_3_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_rMPORT_3_en; // @[TLBStorage.scala 58:8]
  reg  dataBanks_3_perm_pm_r [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_pm_rdata_read_0_3_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_pm_rdata_read_0_3_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_pm_rdata_read_0_3_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_pm_rdata_read_1_3_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_pm_rdata_read_1_3_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_pm_rdata_read_1_3_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_pm_rdata_read_0_3_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_pm_rdata_read_0_3_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_pm_rdata_read_0_3_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_pm_rdata_read_1_3_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_pm_rdata_read_1_3_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_pm_rdata_read_1_3_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_pm_rMPORT_3_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_pm_rMPORT_3_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_pm_rMPORT_3_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_pm_rMPORT_3_en; // @[TLBStorage.scala 58:8]
  reg  dataBanks_3_perm_pm_w [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_pm_wdata_read_0_3_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_pm_wdata_read_0_3_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_pm_wdata_read_0_3_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_pm_wdata_read_1_3_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_pm_wdata_read_1_3_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_pm_wdata_read_1_3_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_pm_wdata_read_0_3_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_pm_wdata_read_0_3_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_pm_wdata_read_0_3_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_pm_wdata_read_1_3_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_pm_wdata_read_1_3_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_pm_wdata_read_1_3_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_pm_wMPORT_3_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_pm_wMPORT_3_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_pm_wMPORT_3_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_pm_wMPORT_3_en; // @[TLBStorage.scala 58:8]
  reg  dataBanks_3_perm_pm_c [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_pm_c_data_read_0_3_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_pm_c_data_read_0_3_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_pm_c_data_read_0_3_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_pm_c_data_read_1_3_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_pm_c_data_read_1_3_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_pm_c_data_read_1_3_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_pm_c_data_read_0_3_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_pm_c_data_read_0_3_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_pm_c_data_read_0_3_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_pm_c_data_read_1_3_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_pm_c_data_read_1_3_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_pm_c_data_read_1_3_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_pm_c_MPORT_3_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_pm_c_MPORT_3_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_pm_c_MPORT_3_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_3_perm_pm_c_MPORT_3_en; // @[TLBStorage.scala 58:8]
  reg [26:0] dataBanks_4_tag [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_tag_data_read_0_4_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_tag_data_read_0_4_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire [26:0] dataBanks_4_tag_data_read_0_4_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_tag_data_read_1_4_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_tag_data_read_1_4_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire [26:0] dataBanks_4_tag_data_read_1_4_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_tag_data_read_0_4_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_tag_data_read_0_4_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire [26:0] dataBanks_4_tag_data_read_0_4_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_tag_data_read_1_4_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_tag_data_read_1_4_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire [26:0] dataBanks_4_tag_data_read_1_4_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire [26:0] dataBanks_4_tag_MPORT_4_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_tag_MPORT_4_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_tag_MPORT_4_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_tag_MPORT_4_en; // @[TLBStorage.scala 58:8]
  reg [15:0] dataBanks_4_asid [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_asid_data_read_0_4_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_asid_data_read_0_4_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire [15:0] dataBanks_4_asid_data_read_0_4_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_asid_data_read_1_4_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_asid_data_read_1_4_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire [15:0] dataBanks_4_asid_data_read_1_4_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_asid_data_read_0_4_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_asid_data_read_0_4_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire [15:0] dataBanks_4_asid_data_read_0_4_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_asid_data_read_1_4_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_asid_data_read_1_4_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire [15:0] dataBanks_4_asid_data_read_1_4_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire [15:0] dataBanks_4_asid_MPORT_4_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_asid_MPORT_4_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_asid_MPORT_4_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_asid_MPORT_4_en; // @[TLBStorage.scala 58:8]
  reg [23:0] dataBanks_4_ppn [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_ppn_data_read_0_4_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_ppn_data_read_0_4_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire [23:0] dataBanks_4_ppn_data_read_0_4_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_ppn_data_read_1_4_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_ppn_data_read_1_4_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire [23:0] dataBanks_4_ppn_data_read_1_4_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_ppn_data_read_0_4_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_ppn_data_read_0_4_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire [23:0] dataBanks_4_ppn_data_read_0_4_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_ppn_data_read_1_4_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_ppn_data_read_1_4_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire [23:0] dataBanks_4_ppn_data_read_1_4_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire [23:0] dataBanks_4_ppn_MPORT_4_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_ppn_MPORT_4_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_ppn_MPORT_4_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_ppn_MPORT_4_en; // @[TLBStorage.scala 58:8]
  reg  dataBanks_4_perm_pf [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_pf_data_read_0_4_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_pf_data_read_0_4_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_pf_data_read_0_4_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_pf_data_read_1_4_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_pf_data_read_1_4_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_pf_data_read_1_4_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_pf_data_read_0_4_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_pf_data_read_0_4_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_pf_data_read_0_4_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_pf_data_read_1_4_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_pf_data_read_1_4_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_pf_data_read_1_4_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_pf_MPORT_4_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_pf_MPORT_4_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_pf_MPORT_4_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_pf_MPORT_4_en; // @[TLBStorage.scala 58:8]
  reg  dataBanks_4_perm_af [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_af_data_read_0_4_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_af_data_read_0_4_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_af_data_read_0_4_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_af_data_read_1_4_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_af_data_read_1_4_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_af_data_read_1_4_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_af_data_read_0_4_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_af_data_read_0_4_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_af_data_read_0_4_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_af_data_read_1_4_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_af_data_read_1_4_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_af_data_read_1_4_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_af_MPORT_4_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_af_MPORT_4_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_af_MPORT_4_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_af_MPORT_4_en; // @[TLBStorage.scala 58:8]
  reg  dataBanks_4_perm_d [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_d_data_read_0_4_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_d_data_read_0_4_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_d_data_read_0_4_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_d_data_read_1_4_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_d_data_read_1_4_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_d_data_read_1_4_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_d_data_read_0_4_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_d_data_read_0_4_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_d_data_read_0_4_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_d_data_read_1_4_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_d_data_read_1_4_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_d_data_read_1_4_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_d_MPORT_4_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_d_MPORT_4_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_d_MPORT_4_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_d_MPORT_4_en; // @[TLBStorage.scala 58:8]
  reg  dataBanks_4_perm_a [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_a_data_read_0_4_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_a_data_read_0_4_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_a_data_read_0_4_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_a_data_read_1_4_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_a_data_read_1_4_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_a_data_read_1_4_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_a_data_read_0_4_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_a_data_read_0_4_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_a_data_read_0_4_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_a_data_read_1_4_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_a_data_read_1_4_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_a_data_read_1_4_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_a_MPORT_4_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_a_MPORT_4_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_a_MPORT_4_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_a_MPORT_4_en; // @[TLBStorage.scala 58:8]
  reg  dataBanks_4_perm_u [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_u_data_read_0_4_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_u_data_read_0_4_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_u_data_read_0_4_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_u_data_read_1_4_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_u_data_read_1_4_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_u_data_read_1_4_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_u_data_read_0_4_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_u_data_read_0_4_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_u_data_read_0_4_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_u_data_read_1_4_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_u_data_read_1_4_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_u_data_read_1_4_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_u_MPORT_4_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_u_MPORT_4_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_u_MPORT_4_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_u_MPORT_4_en; // @[TLBStorage.scala 58:8]
  reg  dataBanks_4_perm_x [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_x_data_read_0_4_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_x_data_read_0_4_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_x_data_read_0_4_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_x_data_read_1_4_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_x_data_read_1_4_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_x_data_read_1_4_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_x_data_read_0_4_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_x_data_read_0_4_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_x_data_read_0_4_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_x_data_read_1_4_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_x_data_read_1_4_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_x_data_read_1_4_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_x_MPORT_4_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_x_MPORT_4_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_x_MPORT_4_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_x_MPORT_4_en; // @[TLBStorage.scala 58:8]
  reg  dataBanks_4_perm_w [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_wdata_read_0_4_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_wdata_read_0_4_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_wdata_read_0_4_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_wdata_read_1_4_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_wdata_read_1_4_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_wdata_read_1_4_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_wdata_read_0_4_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_wdata_read_0_4_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_wdata_read_0_4_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_wdata_read_1_4_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_wdata_read_1_4_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_wdata_read_1_4_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_wMPORT_4_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_wMPORT_4_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_wMPORT_4_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_wMPORT_4_en; // @[TLBStorage.scala 58:8]
  reg  dataBanks_4_perm_r [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_rdata_read_0_4_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_rdata_read_0_4_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_rdata_read_0_4_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_rdata_read_1_4_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_rdata_read_1_4_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_rdata_read_1_4_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_rdata_read_0_4_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_rdata_read_0_4_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_rdata_read_0_4_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_rdata_read_1_4_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_rdata_read_1_4_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_rdata_read_1_4_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_rMPORT_4_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_rMPORT_4_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_rMPORT_4_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_rMPORT_4_en; // @[TLBStorage.scala 58:8]
  reg  dataBanks_4_perm_pm_r [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_pm_rdata_read_0_4_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_pm_rdata_read_0_4_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_pm_rdata_read_0_4_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_pm_rdata_read_1_4_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_pm_rdata_read_1_4_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_pm_rdata_read_1_4_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_pm_rdata_read_0_4_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_pm_rdata_read_0_4_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_pm_rdata_read_0_4_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_pm_rdata_read_1_4_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_pm_rdata_read_1_4_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_pm_rdata_read_1_4_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_pm_rMPORT_4_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_pm_rMPORT_4_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_pm_rMPORT_4_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_pm_rMPORT_4_en; // @[TLBStorage.scala 58:8]
  reg  dataBanks_4_perm_pm_w [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_pm_wdata_read_0_4_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_pm_wdata_read_0_4_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_pm_wdata_read_0_4_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_pm_wdata_read_1_4_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_pm_wdata_read_1_4_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_pm_wdata_read_1_4_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_pm_wdata_read_0_4_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_pm_wdata_read_0_4_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_pm_wdata_read_0_4_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_pm_wdata_read_1_4_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_pm_wdata_read_1_4_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_pm_wdata_read_1_4_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_pm_wMPORT_4_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_pm_wMPORT_4_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_pm_wMPORT_4_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_pm_wMPORT_4_en; // @[TLBStorage.scala 58:8]
  reg  dataBanks_4_perm_pm_c [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_pm_c_data_read_0_4_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_pm_c_data_read_0_4_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_pm_c_data_read_0_4_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_pm_c_data_read_1_4_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_pm_c_data_read_1_4_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_pm_c_data_read_1_4_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_pm_c_data_read_0_4_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_pm_c_data_read_0_4_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_pm_c_data_read_0_4_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_pm_c_data_read_1_4_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_pm_c_data_read_1_4_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_pm_c_data_read_1_4_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_pm_c_MPORT_4_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_pm_c_MPORT_4_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_pm_c_MPORT_4_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_4_perm_pm_c_MPORT_4_en; // @[TLBStorage.scala 58:8]
  reg [26:0] dataBanks_5_tag [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_tag_data_read_0_5_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_tag_data_read_0_5_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire [26:0] dataBanks_5_tag_data_read_0_5_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_tag_data_read_1_5_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_tag_data_read_1_5_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire [26:0] dataBanks_5_tag_data_read_1_5_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_tag_data_read_0_5_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_tag_data_read_0_5_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire [26:0] dataBanks_5_tag_data_read_0_5_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_tag_data_read_1_5_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_tag_data_read_1_5_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire [26:0] dataBanks_5_tag_data_read_1_5_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire [26:0] dataBanks_5_tag_MPORT_5_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_tag_MPORT_5_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_tag_MPORT_5_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_tag_MPORT_5_en; // @[TLBStorage.scala 58:8]
  reg [15:0] dataBanks_5_asid [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_asid_data_read_0_5_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_asid_data_read_0_5_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire [15:0] dataBanks_5_asid_data_read_0_5_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_asid_data_read_1_5_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_asid_data_read_1_5_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire [15:0] dataBanks_5_asid_data_read_1_5_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_asid_data_read_0_5_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_asid_data_read_0_5_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire [15:0] dataBanks_5_asid_data_read_0_5_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_asid_data_read_1_5_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_asid_data_read_1_5_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire [15:0] dataBanks_5_asid_data_read_1_5_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire [15:0] dataBanks_5_asid_MPORT_5_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_asid_MPORT_5_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_asid_MPORT_5_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_asid_MPORT_5_en; // @[TLBStorage.scala 58:8]
  reg [23:0] dataBanks_5_ppn [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_ppn_data_read_0_5_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_ppn_data_read_0_5_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire [23:0] dataBanks_5_ppn_data_read_0_5_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_ppn_data_read_1_5_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_ppn_data_read_1_5_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire [23:0] dataBanks_5_ppn_data_read_1_5_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_ppn_data_read_0_5_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_ppn_data_read_0_5_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire [23:0] dataBanks_5_ppn_data_read_0_5_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_ppn_data_read_1_5_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_ppn_data_read_1_5_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire [23:0] dataBanks_5_ppn_data_read_1_5_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire [23:0] dataBanks_5_ppn_MPORT_5_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_ppn_MPORT_5_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_ppn_MPORT_5_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_ppn_MPORT_5_en; // @[TLBStorage.scala 58:8]
  reg  dataBanks_5_perm_pf [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_pf_data_read_0_5_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_pf_data_read_0_5_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_pf_data_read_0_5_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_pf_data_read_1_5_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_pf_data_read_1_5_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_pf_data_read_1_5_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_pf_data_read_0_5_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_pf_data_read_0_5_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_pf_data_read_0_5_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_pf_data_read_1_5_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_pf_data_read_1_5_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_pf_data_read_1_5_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_pf_MPORT_5_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_pf_MPORT_5_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_pf_MPORT_5_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_pf_MPORT_5_en; // @[TLBStorage.scala 58:8]
  reg  dataBanks_5_perm_af [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_af_data_read_0_5_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_af_data_read_0_5_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_af_data_read_0_5_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_af_data_read_1_5_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_af_data_read_1_5_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_af_data_read_1_5_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_af_data_read_0_5_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_af_data_read_0_5_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_af_data_read_0_5_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_af_data_read_1_5_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_af_data_read_1_5_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_af_data_read_1_5_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_af_MPORT_5_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_af_MPORT_5_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_af_MPORT_5_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_af_MPORT_5_en; // @[TLBStorage.scala 58:8]
  reg  dataBanks_5_perm_d [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_d_data_read_0_5_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_d_data_read_0_5_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_d_data_read_0_5_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_d_data_read_1_5_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_d_data_read_1_5_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_d_data_read_1_5_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_d_data_read_0_5_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_d_data_read_0_5_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_d_data_read_0_5_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_d_data_read_1_5_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_d_data_read_1_5_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_d_data_read_1_5_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_d_MPORT_5_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_d_MPORT_5_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_d_MPORT_5_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_d_MPORT_5_en; // @[TLBStorage.scala 58:8]
  reg  dataBanks_5_perm_a [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_a_data_read_0_5_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_a_data_read_0_5_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_a_data_read_0_5_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_a_data_read_1_5_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_a_data_read_1_5_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_a_data_read_1_5_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_a_data_read_0_5_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_a_data_read_0_5_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_a_data_read_0_5_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_a_data_read_1_5_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_a_data_read_1_5_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_a_data_read_1_5_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_a_MPORT_5_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_a_MPORT_5_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_a_MPORT_5_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_a_MPORT_5_en; // @[TLBStorage.scala 58:8]
  reg  dataBanks_5_perm_u [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_u_data_read_0_5_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_u_data_read_0_5_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_u_data_read_0_5_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_u_data_read_1_5_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_u_data_read_1_5_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_u_data_read_1_5_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_u_data_read_0_5_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_u_data_read_0_5_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_u_data_read_0_5_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_u_data_read_1_5_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_u_data_read_1_5_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_u_data_read_1_5_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_u_MPORT_5_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_u_MPORT_5_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_u_MPORT_5_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_u_MPORT_5_en; // @[TLBStorage.scala 58:8]
  reg  dataBanks_5_perm_x [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_x_data_read_0_5_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_x_data_read_0_5_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_x_data_read_0_5_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_x_data_read_1_5_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_x_data_read_1_5_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_x_data_read_1_5_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_x_data_read_0_5_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_x_data_read_0_5_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_x_data_read_0_5_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_x_data_read_1_5_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_x_data_read_1_5_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_x_data_read_1_5_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_x_MPORT_5_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_x_MPORT_5_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_x_MPORT_5_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_x_MPORT_5_en; // @[TLBStorage.scala 58:8]
  reg  dataBanks_5_perm_w [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_wdata_read_0_5_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_wdata_read_0_5_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_wdata_read_0_5_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_wdata_read_1_5_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_wdata_read_1_5_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_wdata_read_1_5_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_wdata_read_0_5_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_wdata_read_0_5_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_wdata_read_0_5_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_wdata_read_1_5_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_wdata_read_1_5_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_wdata_read_1_5_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_wMPORT_5_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_wMPORT_5_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_wMPORT_5_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_wMPORT_5_en; // @[TLBStorage.scala 58:8]
  reg  dataBanks_5_perm_r [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_rdata_read_0_5_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_rdata_read_0_5_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_rdata_read_0_5_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_rdata_read_1_5_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_rdata_read_1_5_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_rdata_read_1_5_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_rdata_read_0_5_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_rdata_read_0_5_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_rdata_read_0_5_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_rdata_read_1_5_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_rdata_read_1_5_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_rdata_read_1_5_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_rMPORT_5_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_rMPORT_5_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_rMPORT_5_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_rMPORT_5_en; // @[TLBStorage.scala 58:8]
  reg  dataBanks_5_perm_pm_r [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_pm_rdata_read_0_5_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_pm_rdata_read_0_5_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_pm_rdata_read_0_5_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_pm_rdata_read_1_5_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_pm_rdata_read_1_5_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_pm_rdata_read_1_5_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_pm_rdata_read_0_5_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_pm_rdata_read_0_5_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_pm_rdata_read_0_5_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_pm_rdata_read_1_5_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_pm_rdata_read_1_5_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_pm_rdata_read_1_5_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_pm_rMPORT_5_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_pm_rMPORT_5_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_pm_rMPORT_5_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_pm_rMPORT_5_en; // @[TLBStorage.scala 58:8]
  reg  dataBanks_5_perm_pm_w [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_pm_wdata_read_0_5_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_pm_wdata_read_0_5_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_pm_wdata_read_0_5_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_pm_wdata_read_1_5_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_pm_wdata_read_1_5_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_pm_wdata_read_1_5_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_pm_wdata_read_0_5_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_pm_wdata_read_0_5_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_pm_wdata_read_0_5_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_pm_wdata_read_1_5_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_pm_wdata_read_1_5_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_pm_wdata_read_1_5_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_pm_wMPORT_5_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_pm_wMPORT_5_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_pm_wMPORT_5_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_pm_wMPORT_5_en; // @[TLBStorage.scala 58:8]
  reg  dataBanks_5_perm_pm_c [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_pm_c_data_read_0_5_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_pm_c_data_read_0_5_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_pm_c_data_read_0_5_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_pm_c_data_read_1_5_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_pm_c_data_read_1_5_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_pm_c_data_read_1_5_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_pm_c_data_read_0_5_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_pm_c_data_read_0_5_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_pm_c_data_read_0_5_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_pm_c_data_read_1_5_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_pm_c_data_read_1_5_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_pm_c_data_read_1_5_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_pm_c_MPORT_5_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_pm_c_MPORT_5_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_pm_c_MPORT_5_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_5_perm_pm_c_MPORT_5_en; // @[TLBStorage.scala 58:8]
  reg [26:0] dataBanks_6_tag [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_tag_data_read_0_6_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_tag_data_read_0_6_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire [26:0] dataBanks_6_tag_data_read_0_6_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_tag_data_read_1_6_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_tag_data_read_1_6_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire [26:0] dataBanks_6_tag_data_read_1_6_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_tag_data_read_0_6_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_tag_data_read_0_6_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire [26:0] dataBanks_6_tag_data_read_0_6_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_tag_data_read_1_6_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_tag_data_read_1_6_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire [26:0] dataBanks_6_tag_data_read_1_6_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire [26:0] dataBanks_6_tag_MPORT_6_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_tag_MPORT_6_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_tag_MPORT_6_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_tag_MPORT_6_en; // @[TLBStorage.scala 58:8]
  reg [15:0] dataBanks_6_asid [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_asid_data_read_0_6_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_asid_data_read_0_6_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire [15:0] dataBanks_6_asid_data_read_0_6_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_asid_data_read_1_6_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_asid_data_read_1_6_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire [15:0] dataBanks_6_asid_data_read_1_6_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_asid_data_read_0_6_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_asid_data_read_0_6_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire [15:0] dataBanks_6_asid_data_read_0_6_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_asid_data_read_1_6_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_asid_data_read_1_6_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire [15:0] dataBanks_6_asid_data_read_1_6_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire [15:0] dataBanks_6_asid_MPORT_6_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_asid_MPORT_6_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_asid_MPORT_6_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_asid_MPORT_6_en; // @[TLBStorage.scala 58:8]
  reg [23:0] dataBanks_6_ppn [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_ppn_data_read_0_6_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_ppn_data_read_0_6_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire [23:0] dataBanks_6_ppn_data_read_0_6_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_ppn_data_read_1_6_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_ppn_data_read_1_6_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire [23:0] dataBanks_6_ppn_data_read_1_6_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_ppn_data_read_0_6_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_ppn_data_read_0_6_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire [23:0] dataBanks_6_ppn_data_read_0_6_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_ppn_data_read_1_6_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_ppn_data_read_1_6_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire [23:0] dataBanks_6_ppn_data_read_1_6_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire [23:0] dataBanks_6_ppn_MPORT_6_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_ppn_MPORT_6_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_ppn_MPORT_6_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_ppn_MPORT_6_en; // @[TLBStorage.scala 58:8]
  reg  dataBanks_6_perm_pf [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_pf_data_read_0_6_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_pf_data_read_0_6_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_pf_data_read_0_6_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_pf_data_read_1_6_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_pf_data_read_1_6_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_pf_data_read_1_6_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_pf_data_read_0_6_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_pf_data_read_0_6_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_pf_data_read_0_6_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_pf_data_read_1_6_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_pf_data_read_1_6_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_pf_data_read_1_6_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_pf_MPORT_6_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_pf_MPORT_6_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_pf_MPORT_6_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_pf_MPORT_6_en; // @[TLBStorage.scala 58:8]
  reg  dataBanks_6_perm_af [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_af_data_read_0_6_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_af_data_read_0_6_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_af_data_read_0_6_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_af_data_read_1_6_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_af_data_read_1_6_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_af_data_read_1_6_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_af_data_read_0_6_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_af_data_read_0_6_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_af_data_read_0_6_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_af_data_read_1_6_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_af_data_read_1_6_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_af_data_read_1_6_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_af_MPORT_6_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_af_MPORT_6_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_af_MPORT_6_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_af_MPORT_6_en; // @[TLBStorage.scala 58:8]
  reg  dataBanks_6_perm_d [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_d_data_read_0_6_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_d_data_read_0_6_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_d_data_read_0_6_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_d_data_read_1_6_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_d_data_read_1_6_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_d_data_read_1_6_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_d_data_read_0_6_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_d_data_read_0_6_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_d_data_read_0_6_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_d_data_read_1_6_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_d_data_read_1_6_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_d_data_read_1_6_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_d_MPORT_6_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_d_MPORT_6_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_d_MPORT_6_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_d_MPORT_6_en; // @[TLBStorage.scala 58:8]
  reg  dataBanks_6_perm_a [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_a_data_read_0_6_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_a_data_read_0_6_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_a_data_read_0_6_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_a_data_read_1_6_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_a_data_read_1_6_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_a_data_read_1_6_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_a_data_read_0_6_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_a_data_read_0_6_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_a_data_read_0_6_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_a_data_read_1_6_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_a_data_read_1_6_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_a_data_read_1_6_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_a_MPORT_6_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_a_MPORT_6_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_a_MPORT_6_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_a_MPORT_6_en; // @[TLBStorage.scala 58:8]
  reg  dataBanks_6_perm_u [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_u_data_read_0_6_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_u_data_read_0_6_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_u_data_read_0_6_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_u_data_read_1_6_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_u_data_read_1_6_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_u_data_read_1_6_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_u_data_read_0_6_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_u_data_read_0_6_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_u_data_read_0_6_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_u_data_read_1_6_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_u_data_read_1_6_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_u_data_read_1_6_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_u_MPORT_6_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_u_MPORT_6_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_u_MPORT_6_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_u_MPORT_6_en; // @[TLBStorage.scala 58:8]
  reg  dataBanks_6_perm_x [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_x_data_read_0_6_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_x_data_read_0_6_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_x_data_read_0_6_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_x_data_read_1_6_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_x_data_read_1_6_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_x_data_read_1_6_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_x_data_read_0_6_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_x_data_read_0_6_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_x_data_read_0_6_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_x_data_read_1_6_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_x_data_read_1_6_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_x_data_read_1_6_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_x_MPORT_6_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_x_MPORT_6_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_x_MPORT_6_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_x_MPORT_6_en; // @[TLBStorage.scala 58:8]
  reg  dataBanks_6_perm_w [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_wdata_read_0_6_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_wdata_read_0_6_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_wdata_read_0_6_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_wdata_read_1_6_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_wdata_read_1_6_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_wdata_read_1_6_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_wdata_read_0_6_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_wdata_read_0_6_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_wdata_read_0_6_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_wdata_read_1_6_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_wdata_read_1_6_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_wdata_read_1_6_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_wMPORT_6_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_wMPORT_6_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_wMPORT_6_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_wMPORT_6_en; // @[TLBStorage.scala 58:8]
  reg  dataBanks_6_perm_r [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_rdata_read_0_6_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_rdata_read_0_6_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_rdata_read_0_6_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_rdata_read_1_6_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_rdata_read_1_6_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_rdata_read_1_6_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_rdata_read_0_6_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_rdata_read_0_6_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_rdata_read_0_6_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_rdata_read_1_6_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_rdata_read_1_6_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_rdata_read_1_6_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_rMPORT_6_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_rMPORT_6_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_rMPORT_6_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_rMPORT_6_en; // @[TLBStorage.scala 58:8]
  reg  dataBanks_6_perm_pm_r [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_pm_rdata_read_0_6_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_pm_rdata_read_0_6_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_pm_rdata_read_0_6_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_pm_rdata_read_1_6_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_pm_rdata_read_1_6_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_pm_rdata_read_1_6_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_pm_rdata_read_0_6_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_pm_rdata_read_0_6_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_pm_rdata_read_0_6_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_pm_rdata_read_1_6_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_pm_rdata_read_1_6_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_pm_rdata_read_1_6_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_pm_rMPORT_6_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_pm_rMPORT_6_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_pm_rMPORT_6_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_pm_rMPORT_6_en; // @[TLBStorage.scala 58:8]
  reg  dataBanks_6_perm_pm_w [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_pm_wdata_read_0_6_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_pm_wdata_read_0_6_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_pm_wdata_read_0_6_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_pm_wdata_read_1_6_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_pm_wdata_read_1_6_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_pm_wdata_read_1_6_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_pm_wdata_read_0_6_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_pm_wdata_read_0_6_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_pm_wdata_read_0_6_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_pm_wdata_read_1_6_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_pm_wdata_read_1_6_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_pm_wdata_read_1_6_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_pm_wMPORT_6_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_pm_wMPORT_6_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_pm_wMPORT_6_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_pm_wMPORT_6_en; // @[TLBStorage.scala 58:8]
  reg  dataBanks_6_perm_pm_c [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_pm_c_data_read_0_6_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_pm_c_data_read_0_6_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_pm_c_data_read_0_6_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_pm_c_data_read_1_6_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_pm_c_data_read_1_6_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_pm_c_data_read_1_6_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_pm_c_data_read_0_6_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_pm_c_data_read_0_6_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_pm_c_data_read_0_6_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_pm_c_data_read_1_6_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_pm_c_data_read_1_6_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_pm_c_data_read_1_6_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_pm_c_MPORT_6_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_pm_c_MPORT_6_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_pm_c_MPORT_6_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_6_perm_pm_c_MPORT_6_en; // @[TLBStorage.scala 58:8]
  reg [26:0] dataBanks_7_tag [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_tag_data_read_0_7_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_tag_data_read_0_7_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire [26:0] dataBanks_7_tag_data_read_0_7_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_tag_data_read_1_7_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_tag_data_read_1_7_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire [26:0] dataBanks_7_tag_data_read_1_7_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_tag_data_read_0_7_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_tag_data_read_0_7_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire [26:0] dataBanks_7_tag_data_read_0_7_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_tag_data_read_1_7_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_tag_data_read_1_7_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire [26:0] dataBanks_7_tag_data_read_1_7_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire [26:0] dataBanks_7_tag_MPORT_7_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_tag_MPORT_7_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_tag_MPORT_7_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_tag_MPORT_7_en; // @[TLBStorage.scala 58:8]
  reg [15:0] dataBanks_7_asid [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_asid_data_read_0_7_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_asid_data_read_0_7_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire [15:0] dataBanks_7_asid_data_read_0_7_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_asid_data_read_1_7_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_asid_data_read_1_7_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire [15:0] dataBanks_7_asid_data_read_1_7_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_asid_data_read_0_7_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_asid_data_read_0_7_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire [15:0] dataBanks_7_asid_data_read_0_7_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_asid_data_read_1_7_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_asid_data_read_1_7_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire [15:0] dataBanks_7_asid_data_read_1_7_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire [15:0] dataBanks_7_asid_MPORT_7_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_asid_MPORT_7_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_asid_MPORT_7_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_asid_MPORT_7_en; // @[TLBStorage.scala 58:8]
  reg [23:0] dataBanks_7_ppn [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_ppn_data_read_0_7_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_ppn_data_read_0_7_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire [23:0] dataBanks_7_ppn_data_read_0_7_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_ppn_data_read_1_7_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_ppn_data_read_1_7_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire [23:0] dataBanks_7_ppn_data_read_1_7_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_ppn_data_read_0_7_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_ppn_data_read_0_7_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire [23:0] dataBanks_7_ppn_data_read_0_7_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_ppn_data_read_1_7_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_ppn_data_read_1_7_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire [23:0] dataBanks_7_ppn_data_read_1_7_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire [23:0] dataBanks_7_ppn_MPORT_7_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_ppn_MPORT_7_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_ppn_MPORT_7_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_ppn_MPORT_7_en; // @[TLBStorage.scala 58:8]
  reg  dataBanks_7_perm_pf [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_pf_data_read_0_7_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_pf_data_read_0_7_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_pf_data_read_0_7_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_pf_data_read_1_7_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_pf_data_read_1_7_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_pf_data_read_1_7_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_pf_data_read_0_7_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_pf_data_read_0_7_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_pf_data_read_0_7_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_pf_data_read_1_7_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_pf_data_read_1_7_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_pf_data_read_1_7_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_pf_MPORT_7_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_pf_MPORT_7_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_pf_MPORT_7_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_pf_MPORT_7_en; // @[TLBStorage.scala 58:8]
  reg  dataBanks_7_perm_af [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_af_data_read_0_7_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_af_data_read_0_7_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_af_data_read_0_7_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_af_data_read_1_7_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_af_data_read_1_7_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_af_data_read_1_7_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_af_data_read_0_7_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_af_data_read_0_7_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_af_data_read_0_7_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_af_data_read_1_7_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_af_data_read_1_7_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_af_data_read_1_7_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_af_MPORT_7_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_af_MPORT_7_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_af_MPORT_7_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_af_MPORT_7_en; // @[TLBStorage.scala 58:8]
  reg  dataBanks_7_perm_d [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_d_data_read_0_7_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_d_data_read_0_7_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_d_data_read_0_7_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_d_data_read_1_7_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_d_data_read_1_7_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_d_data_read_1_7_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_d_data_read_0_7_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_d_data_read_0_7_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_d_data_read_0_7_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_d_data_read_1_7_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_d_data_read_1_7_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_d_data_read_1_7_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_d_MPORT_7_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_d_MPORT_7_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_d_MPORT_7_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_d_MPORT_7_en; // @[TLBStorage.scala 58:8]
  reg  dataBanks_7_perm_a [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_a_data_read_0_7_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_a_data_read_0_7_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_a_data_read_0_7_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_a_data_read_1_7_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_a_data_read_1_7_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_a_data_read_1_7_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_a_data_read_0_7_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_a_data_read_0_7_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_a_data_read_0_7_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_a_data_read_1_7_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_a_data_read_1_7_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_a_data_read_1_7_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_a_MPORT_7_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_a_MPORT_7_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_a_MPORT_7_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_a_MPORT_7_en; // @[TLBStorage.scala 58:8]
  reg  dataBanks_7_perm_u [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_u_data_read_0_7_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_u_data_read_0_7_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_u_data_read_0_7_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_u_data_read_1_7_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_u_data_read_1_7_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_u_data_read_1_7_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_u_data_read_0_7_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_u_data_read_0_7_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_u_data_read_0_7_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_u_data_read_1_7_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_u_data_read_1_7_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_u_data_read_1_7_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_u_MPORT_7_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_u_MPORT_7_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_u_MPORT_7_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_u_MPORT_7_en; // @[TLBStorage.scala 58:8]
  reg  dataBanks_7_perm_x [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_x_data_read_0_7_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_x_data_read_0_7_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_x_data_read_0_7_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_x_data_read_1_7_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_x_data_read_1_7_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_x_data_read_1_7_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_x_data_read_0_7_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_x_data_read_0_7_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_x_data_read_0_7_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_x_data_read_1_7_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_x_data_read_1_7_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_x_data_read_1_7_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_x_MPORT_7_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_x_MPORT_7_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_x_MPORT_7_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_x_MPORT_7_en; // @[TLBStorage.scala 58:8]
  reg  dataBanks_7_perm_w [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_wdata_read_0_7_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_wdata_read_0_7_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_wdata_read_0_7_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_wdata_read_1_7_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_wdata_read_1_7_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_wdata_read_1_7_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_wdata_read_0_7_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_wdata_read_0_7_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_wdata_read_0_7_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_wdata_read_1_7_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_wdata_read_1_7_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_wdata_read_1_7_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_wMPORT_7_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_wMPORT_7_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_wMPORT_7_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_wMPORT_7_en; // @[TLBStorage.scala 58:8]
  reg  dataBanks_7_perm_r [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_rdata_read_0_7_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_rdata_read_0_7_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_rdata_read_0_7_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_rdata_read_1_7_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_rdata_read_1_7_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_rdata_read_1_7_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_rdata_read_0_7_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_rdata_read_0_7_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_rdata_read_0_7_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_rdata_read_1_7_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_rdata_read_1_7_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_rdata_read_1_7_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_rMPORT_7_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_rMPORT_7_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_rMPORT_7_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_rMPORT_7_en; // @[TLBStorage.scala 58:8]
  reg  dataBanks_7_perm_pm_r [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_pm_rdata_read_0_7_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_pm_rdata_read_0_7_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_pm_rdata_read_0_7_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_pm_rdata_read_1_7_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_pm_rdata_read_1_7_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_pm_rdata_read_1_7_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_pm_rdata_read_0_7_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_pm_rdata_read_0_7_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_pm_rdata_read_0_7_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_pm_rdata_read_1_7_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_pm_rdata_read_1_7_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_pm_rdata_read_1_7_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_pm_rMPORT_7_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_pm_rMPORT_7_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_pm_rMPORT_7_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_pm_rMPORT_7_en; // @[TLBStorage.scala 58:8]
  reg  dataBanks_7_perm_pm_w [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_pm_wdata_read_0_7_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_pm_wdata_read_0_7_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_pm_wdata_read_0_7_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_pm_wdata_read_1_7_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_pm_wdata_read_1_7_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_pm_wdata_read_1_7_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_pm_wdata_read_0_7_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_pm_wdata_read_0_7_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_pm_wdata_read_0_7_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_pm_wdata_read_1_7_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_pm_wdata_read_1_7_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_pm_wdata_read_1_7_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_pm_wMPORT_7_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_pm_wMPORT_7_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_pm_wMPORT_7_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_pm_wMPORT_7_en; // @[TLBStorage.scala 58:8]
  reg  dataBanks_7_perm_pm_c [0:1]; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_pm_c_data_read_0_7_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_pm_c_data_read_0_7_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_pm_c_data_read_0_7_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_pm_c_data_read_1_7_MPORT_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_pm_c_data_read_1_7_MPORT_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_pm_c_data_read_1_7_MPORT_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_pm_c_data_read_0_7_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_pm_c_data_read_0_7_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_pm_c_data_read_0_7_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_pm_c_data_read_1_7_MPORT_1_en; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_pm_c_data_read_1_7_MPORT_1_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_pm_c_data_read_1_7_MPORT_1_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_pm_c_MPORT_7_data; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_pm_c_MPORT_7_addr; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_pm_c_MPORT_7_mask; // @[TLBStorage.scala 58:8]
  wire  dataBanks_7_perm_pm_c_MPORT_7_en; // @[TLBStorage.scala 58:8]
  reg [26:0] data_read__0_0_tag; // @[TLBStorage.scala 63:24]
  reg [15:0] data_read__0_0_asid; // @[TLBStorage.scala 63:24]
  reg [23:0] data_read__0_0_ppn; // @[TLBStorage.scala 63:24]
  reg  data_read__0_0_perm_pf; // @[TLBStorage.scala 63:24]
  reg  data_read__0_0_perm_af; // @[TLBStorage.scala 63:24]
  reg  data_read__0_0_perm_d; // @[TLBStorage.scala 63:24]
  reg  data_read__0_0_perm_a; // @[TLBStorage.scala 63:24]
  reg  data_read__0_0_perm_u; // @[TLBStorage.scala 63:24]
  reg  data_read__0_0_perm_x; // @[TLBStorage.scala 63:24]
  reg  data_read__0_0_perm_w; // @[TLBStorage.scala 63:24]
  reg  data_read__0_0_perm_r; // @[TLBStorage.scala 63:24]
  reg  data_read__0_0_perm_pm_r; // @[TLBStorage.scala 63:24]
  reg  data_read__0_0_perm_pm_w; // @[TLBStorage.scala 63:24]
  reg  data_read__0_0_perm_pm_c; // @[TLBStorage.scala 63:24]
  reg [26:0] data_read__0_1_tag; // @[TLBStorage.scala 63:24]
  reg [15:0] data_read__0_1_asid; // @[TLBStorage.scala 63:24]
  reg [23:0] data_read__0_1_ppn; // @[TLBStorage.scala 63:24]
  reg  data_read__0_1_perm_pf; // @[TLBStorage.scala 63:24]
  reg  data_read__0_1_perm_af; // @[TLBStorage.scala 63:24]
  reg  data_read__0_1_perm_d; // @[TLBStorage.scala 63:24]
  reg  data_read__0_1_perm_a; // @[TLBStorage.scala 63:24]
  reg  data_read__0_1_perm_u; // @[TLBStorage.scala 63:24]
  reg  data_read__0_1_perm_x; // @[TLBStorage.scala 63:24]
  reg  data_read__0_1_perm_w; // @[TLBStorage.scala 63:24]
  reg  data_read__0_1_perm_r; // @[TLBStorage.scala 63:24]
  reg  data_read__0_1_perm_pm_r; // @[TLBStorage.scala 63:24]
  reg  data_read__0_1_perm_pm_w; // @[TLBStorage.scala 63:24]
  reg  data_read__0_1_perm_pm_c; // @[TLBStorage.scala 63:24]
  reg [26:0] data_read__0_2_tag; // @[TLBStorage.scala 63:24]
  reg [15:0] data_read__0_2_asid; // @[TLBStorage.scala 63:24]
  reg [23:0] data_read__0_2_ppn; // @[TLBStorage.scala 63:24]
  reg  data_read__0_2_perm_pf; // @[TLBStorage.scala 63:24]
  reg  data_read__0_2_perm_af; // @[TLBStorage.scala 63:24]
  reg  data_read__0_2_perm_d; // @[TLBStorage.scala 63:24]
  reg  data_read__0_2_perm_a; // @[TLBStorage.scala 63:24]
  reg  data_read__0_2_perm_u; // @[TLBStorage.scala 63:24]
  reg  data_read__0_2_perm_x; // @[TLBStorage.scala 63:24]
  reg  data_read__0_2_perm_w; // @[TLBStorage.scala 63:24]
  reg  data_read__0_2_perm_r; // @[TLBStorage.scala 63:24]
  reg  data_read__0_2_perm_pm_r; // @[TLBStorage.scala 63:24]
  reg  data_read__0_2_perm_pm_w; // @[TLBStorage.scala 63:24]
  reg  data_read__0_2_perm_pm_c; // @[TLBStorage.scala 63:24]
  reg [26:0] data_read__0_3_tag; // @[TLBStorage.scala 63:24]
  reg [15:0] data_read__0_3_asid; // @[TLBStorage.scala 63:24]
  reg [23:0] data_read__0_3_ppn; // @[TLBStorage.scala 63:24]
  reg  data_read__0_3_perm_pf; // @[TLBStorage.scala 63:24]
  reg  data_read__0_3_perm_af; // @[TLBStorage.scala 63:24]
  reg  data_read__0_3_perm_d; // @[TLBStorage.scala 63:24]
  reg  data_read__0_3_perm_a; // @[TLBStorage.scala 63:24]
  reg  data_read__0_3_perm_u; // @[TLBStorage.scala 63:24]
  reg  data_read__0_3_perm_x; // @[TLBStorage.scala 63:24]
  reg  data_read__0_3_perm_w; // @[TLBStorage.scala 63:24]
  reg  data_read__0_3_perm_r; // @[TLBStorage.scala 63:24]
  reg  data_read__0_3_perm_pm_r; // @[TLBStorage.scala 63:24]
  reg  data_read__0_3_perm_pm_w; // @[TLBStorage.scala 63:24]
  reg  data_read__0_3_perm_pm_c; // @[TLBStorage.scala 63:24]
  reg [26:0] data_read__0_4_tag; // @[TLBStorage.scala 63:24]
  reg [15:0] data_read__0_4_asid; // @[TLBStorage.scala 63:24]
  reg [23:0] data_read__0_4_ppn; // @[TLBStorage.scala 63:24]
  reg  data_read__0_4_perm_pf; // @[TLBStorage.scala 63:24]
  reg  data_read__0_4_perm_af; // @[TLBStorage.scala 63:24]
  reg  data_read__0_4_perm_d; // @[TLBStorage.scala 63:24]
  reg  data_read__0_4_perm_a; // @[TLBStorage.scala 63:24]
  reg  data_read__0_4_perm_u; // @[TLBStorage.scala 63:24]
  reg  data_read__0_4_perm_x; // @[TLBStorage.scala 63:24]
  reg  data_read__0_4_perm_w; // @[TLBStorage.scala 63:24]
  reg  data_read__0_4_perm_r; // @[TLBStorage.scala 63:24]
  reg  data_read__0_4_perm_pm_r; // @[TLBStorage.scala 63:24]
  reg  data_read__0_4_perm_pm_w; // @[TLBStorage.scala 63:24]
  reg  data_read__0_4_perm_pm_c; // @[TLBStorage.scala 63:24]
  reg [26:0] data_read__0_5_tag; // @[TLBStorage.scala 63:24]
  reg [15:0] data_read__0_5_asid; // @[TLBStorage.scala 63:24]
  reg [23:0] data_read__0_5_ppn; // @[TLBStorage.scala 63:24]
  reg  data_read__0_5_perm_pf; // @[TLBStorage.scala 63:24]
  reg  data_read__0_5_perm_af; // @[TLBStorage.scala 63:24]
  reg  data_read__0_5_perm_d; // @[TLBStorage.scala 63:24]
  reg  data_read__0_5_perm_a; // @[TLBStorage.scala 63:24]
  reg  data_read__0_5_perm_u; // @[TLBStorage.scala 63:24]
  reg  data_read__0_5_perm_x; // @[TLBStorage.scala 63:24]
  reg  data_read__0_5_perm_w; // @[TLBStorage.scala 63:24]
  reg  data_read__0_5_perm_r; // @[TLBStorage.scala 63:24]
  reg  data_read__0_5_perm_pm_r; // @[TLBStorage.scala 63:24]
  reg  data_read__0_5_perm_pm_w; // @[TLBStorage.scala 63:24]
  reg  data_read__0_5_perm_pm_c; // @[TLBStorage.scala 63:24]
  reg [26:0] data_read__0_6_tag; // @[TLBStorage.scala 63:24]
  reg [15:0] data_read__0_6_asid; // @[TLBStorage.scala 63:24]
  reg [23:0] data_read__0_6_ppn; // @[TLBStorage.scala 63:24]
  reg  data_read__0_6_perm_pf; // @[TLBStorage.scala 63:24]
  reg  data_read__0_6_perm_af; // @[TLBStorage.scala 63:24]
  reg  data_read__0_6_perm_d; // @[TLBStorage.scala 63:24]
  reg  data_read__0_6_perm_a; // @[TLBStorage.scala 63:24]
  reg  data_read__0_6_perm_u; // @[TLBStorage.scala 63:24]
  reg  data_read__0_6_perm_x; // @[TLBStorage.scala 63:24]
  reg  data_read__0_6_perm_w; // @[TLBStorage.scala 63:24]
  reg  data_read__0_6_perm_r; // @[TLBStorage.scala 63:24]
  reg  data_read__0_6_perm_pm_r; // @[TLBStorage.scala 63:24]
  reg  data_read__0_6_perm_pm_w; // @[TLBStorage.scala 63:24]
  reg  data_read__0_6_perm_pm_c; // @[TLBStorage.scala 63:24]
  reg [26:0] data_read__0_7_tag; // @[TLBStorage.scala 63:24]
  reg [15:0] data_read__0_7_asid; // @[TLBStorage.scala 63:24]
  reg [23:0] data_read__0_7_ppn; // @[TLBStorage.scala 63:24]
  reg  data_read__0_7_perm_pf; // @[TLBStorage.scala 63:24]
  reg  data_read__0_7_perm_af; // @[TLBStorage.scala 63:24]
  reg  data_read__0_7_perm_d; // @[TLBStorage.scala 63:24]
  reg  data_read__0_7_perm_a; // @[TLBStorage.scala 63:24]
  reg  data_read__0_7_perm_u; // @[TLBStorage.scala 63:24]
  reg  data_read__0_7_perm_x; // @[TLBStorage.scala 63:24]
  reg  data_read__0_7_perm_w; // @[TLBStorage.scala 63:24]
  reg  data_read__0_7_perm_r; // @[TLBStorage.scala 63:24]
  reg  data_read__0_7_perm_pm_r; // @[TLBStorage.scala 63:24]
  reg  data_read__0_7_perm_pm_w; // @[TLBStorage.scala 63:24]
  reg  data_read__0_7_perm_pm_c; // @[TLBStorage.scala 63:24]
  reg [23:0] data_read__1_0_ppn; // @[TLBStorage.scala 63:24]
  reg [23:0] data_read__1_1_ppn; // @[TLBStorage.scala 63:24]
  reg [23:0] data_read__1_2_ppn; // @[TLBStorage.scala 63:24]
  reg [23:0] data_read__1_3_ppn; // @[TLBStorage.scala 63:24]
  reg [23:0] data_read__1_4_ppn; // @[TLBStorage.scala 63:24]
  reg [23:0] data_read__1_5_ppn; // @[TLBStorage.scala 63:24]
  reg [23:0] data_read__1_6_ppn; // @[TLBStorage.scala 63:24]
  reg [23:0] data_read__1_7_ppn; // @[TLBStorage.scala 63:24]
  reg [7:0] bank_index__0; // @[TLBStorage.scala 64:25]
  reg [7:0] bank_index__1; // @[TLBStorage.scala 64:25]
  wire [23:0] _io_rdata_0_0_T_218 = bank_index__0[0] ? data_read__0_0_ppn : 24'h0; // @[Mux.scala 27:73]
  wire [23:0] _io_rdata_0_0_T_219 = bank_index__0[1] ? data_read__0_1_ppn : 24'h0; // @[Mux.scala 27:73]
  wire [23:0] _io_rdata_0_0_T_220 = bank_index__0[2] ? data_read__0_2_ppn : 24'h0; // @[Mux.scala 27:73]
  wire [23:0] _io_rdata_0_0_T_221 = bank_index__0[3] ? data_read__0_3_ppn : 24'h0; // @[Mux.scala 27:73]
  wire [23:0] _io_rdata_0_0_T_222 = bank_index__0[4] ? data_read__0_4_ppn : 24'h0; // @[Mux.scala 27:73]
  wire [23:0] _io_rdata_0_0_T_223 = bank_index__0[5] ? data_read__0_5_ppn : 24'h0; // @[Mux.scala 27:73]
  wire [23:0] _io_rdata_0_0_T_224 = bank_index__0[6] ? data_read__0_6_ppn : 24'h0; // @[Mux.scala 27:73]
  wire [23:0] _io_rdata_0_0_T_225 = bank_index__0[7] ? data_read__0_7_ppn : 24'h0; // @[Mux.scala 27:73]
  wire [23:0] _io_rdata_0_0_T_226 = _io_rdata_0_0_T_218 | _io_rdata_0_0_T_219; // @[Mux.scala 27:73]
  wire [23:0] _io_rdata_0_0_T_227 = _io_rdata_0_0_T_226 | _io_rdata_0_0_T_220; // @[Mux.scala 27:73]
  wire [23:0] _io_rdata_0_0_T_228 = _io_rdata_0_0_T_227 | _io_rdata_0_0_T_221; // @[Mux.scala 27:73]
  wire [23:0] _io_rdata_0_0_T_229 = _io_rdata_0_0_T_228 | _io_rdata_0_0_T_222; // @[Mux.scala 27:73]
  wire [23:0] _io_rdata_0_0_T_230 = _io_rdata_0_0_T_229 | _io_rdata_0_0_T_223; // @[Mux.scala 27:73]
  wire [23:0] _io_rdata_0_0_T_231 = _io_rdata_0_0_T_230 | _io_rdata_0_0_T_224; // @[Mux.scala 27:73]
  wire [15:0] _io_rdata_0_0_T_233 = bank_index__0[0] ? data_read__0_0_asid : 16'h0; // @[Mux.scala 27:73]
  wire [15:0] _io_rdata_0_0_T_234 = bank_index__0[1] ? data_read__0_1_asid : 16'h0; // @[Mux.scala 27:73]
  wire [15:0] _io_rdata_0_0_T_235 = bank_index__0[2] ? data_read__0_2_asid : 16'h0; // @[Mux.scala 27:73]
  wire [15:0] _io_rdata_0_0_T_236 = bank_index__0[3] ? data_read__0_3_asid : 16'h0; // @[Mux.scala 27:73]
  wire [15:0] _io_rdata_0_0_T_237 = bank_index__0[4] ? data_read__0_4_asid : 16'h0; // @[Mux.scala 27:73]
  wire [15:0] _io_rdata_0_0_T_238 = bank_index__0[5] ? data_read__0_5_asid : 16'h0; // @[Mux.scala 27:73]
  wire [15:0] _io_rdata_0_0_T_239 = bank_index__0[6] ? data_read__0_6_asid : 16'h0; // @[Mux.scala 27:73]
  wire [15:0] _io_rdata_0_0_T_240 = bank_index__0[7] ? data_read__0_7_asid : 16'h0; // @[Mux.scala 27:73]
  wire [15:0] _io_rdata_0_0_T_241 = _io_rdata_0_0_T_233 | _io_rdata_0_0_T_234; // @[Mux.scala 27:73]
  wire [15:0] _io_rdata_0_0_T_242 = _io_rdata_0_0_T_241 | _io_rdata_0_0_T_235; // @[Mux.scala 27:73]
  wire [15:0] _io_rdata_0_0_T_243 = _io_rdata_0_0_T_242 | _io_rdata_0_0_T_236; // @[Mux.scala 27:73]
  wire [15:0] _io_rdata_0_0_T_244 = _io_rdata_0_0_T_243 | _io_rdata_0_0_T_237; // @[Mux.scala 27:73]
  wire [15:0] _io_rdata_0_0_T_245 = _io_rdata_0_0_T_244 | _io_rdata_0_0_T_238; // @[Mux.scala 27:73]
  wire [15:0] _io_rdata_0_0_T_246 = _io_rdata_0_0_T_245 | _io_rdata_0_0_T_239; // @[Mux.scala 27:73]
  wire [26:0] _io_rdata_0_0_T_248 = bank_index__0[0] ? data_read__0_0_tag : 27'h0; // @[Mux.scala 27:73]
  wire [26:0] _io_rdata_0_0_T_249 = bank_index__0[1] ? data_read__0_1_tag : 27'h0; // @[Mux.scala 27:73]
  wire [26:0] _io_rdata_0_0_T_250 = bank_index__0[2] ? data_read__0_2_tag : 27'h0; // @[Mux.scala 27:73]
  wire [26:0] _io_rdata_0_0_T_251 = bank_index__0[3] ? data_read__0_3_tag : 27'h0; // @[Mux.scala 27:73]
  wire [26:0] _io_rdata_0_0_T_252 = bank_index__0[4] ? data_read__0_4_tag : 27'h0; // @[Mux.scala 27:73]
  wire [26:0] _io_rdata_0_0_T_253 = bank_index__0[5] ? data_read__0_5_tag : 27'h0; // @[Mux.scala 27:73]
  wire [26:0] _io_rdata_0_0_T_254 = bank_index__0[6] ? data_read__0_6_tag : 27'h0; // @[Mux.scala 27:73]
  wire [26:0] _io_rdata_0_0_T_255 = bank_index__0[7] ? data_read__0_7_tag : 27'h0; // @[Mux.scala 27:73]
  wire [26:0] _io_rdata_0_0_T_256 = _io_rdata_0_0_T_248 | _io_rdata_0_0_T_249; // @[Mux.scala 27:73]
  wire [26:0] _io_rdata_0_0_T_257 = _io_rdata_0_0_T_256 | _io_rdata_0_0_T_250; // @[Mux.scala 27:73]
  wire [26:0] _io_rdata_0_0_T_258 = _io_rdata_0_0_T_257 | _io_rdata_0_0_T_251; // @[Mux.scala 27:73]
  wire [26:0] _io_rdata_0_0_T_259 = _io_rdata_0_0_T_258 | _io_rdata_0_0_T_252; // @[Mux.scala 27:73]
  wire [26:0] _io_rdata_0_0_T_260 = _io_rdata_0_0_T_259 | _io_rdata_0_0_T_253; // @[Mux.scala 27:73]
  wire [26:0] _io_rdata_0_0_T_261 = _io_rdata_0_0_T_260 | _io_rdata_0_0_T_254; // @[Mux.scala 27:73]
  wire [23:0] _io_rdata_0_1_T_218 = bank_index__1[0] ? data_read__1_0_ppn : 24'h0; // @[Mux.scala 27:73]
  wire [23:0] _io_rdata_0_1_T_219 = bank_index__1[1] ? data_read__1_1_ppn : 24'h0; // @[Mux.scala 27:73]
  wire [23:0] _io_rdata_0_1_T_220 = bank_index__1[2] ? data_read__1_2_ppn : 24'h0; // @[Mux.scala 27:73]
  wire [23:0] _io_rdata_0_1_T_221 = bank_index__1[3] ? data_read__1_3_ppn : 24'h0; // @[Mux.scala 27:73]
  wire [23:0] _io_rdata_0_1_T_222 = bank_index__1[4] ? data_read__1_4_ppn : 24'h0; // @[Mux.scala 27:73]
  wire [23:0] _io_rdata_0_1_T_223 = bank_index__1[5] ? data_read__1_5_ppn : 24'h0; // @[Mux.scala 27:73]
  wire [23:0] _io_rdata_0_1_T_224 = bank_index__1[6] ? data_read__1_6_ppn : 24'h0; // @[Mux.scala 27:73]
  wire [23:0] _io_rdata_0_1_T_225 = bank_index__1[7] ? data_read__1_7_ppn : 24'h0; // @[Mux.scala 27:73]
  wire [23:0] _io_rdata_0_1_T_226 = _io_rdata_0_1_T_218 | _io_rdata_0_1_T_219; // @[Mux.scala 27:73]
  wire [23:0] _io_rdata_0_1_T_227 = _io_rdata_0_1_T_226 | _io_rdata_0_1_T_220; // @[Mux.scala 27:73]
  wire [23:0] _io_rdata_0_1_T_228 = _io_rdata_0_1_T_227 | _io_rdata_0_1_T_221; // @[Mux.scala 27:73]
  wire [23:0] _io_rdata_0_1_T_229 = _io_rdata_0_1_T_228 | _io_rdata_0_1_T_222; // @[Mux.scala 27:73]
  wire [23:0] _io_rdata_0_1_T_230 = _io_rdata_0_1_T_229 | _io_rdata_0_1_T_223; // @[Mux.scala 27:73]
  wire [23:0] _io_rdata_0_1_T_231 = _io_rdata_0_1_T_230 | _io_rdata_0_1_T_224; // @[Mux.scala 27:73]
  reg [26:0] data_read_1_0_0_tag; // @[TLBStorage.scala 63:24]
  reg [15:0] data_read_1_0_0_asid; // @[TLBStorage.scala 63:24]
  reg [23:0] data_read_1_0_0_ppn; // @[TLBStorage.scala 63:24]
  reg  data_read_1_0_0_perm_pf; // @[TLBStorage.scala 63:24]
  reg  data_read_1_0_0_perm_af; // @[TLBStorage.scala 63:24]
  reg  data_read_1_0_0_perm_a; // @[TLBStorage.scala 63:24]
  reg  data_read_1_0_0_perm_u; // @[TLBStorage.scala 63:24]
  reg  data_read_1_0_0_perm_x; // @[TLBStorage.scala 63:24]
  reg  data_read_1_0_0_perm_r; // @[TLBStorage.scala 63:24]
  reg  data_read_1_0_0_perm_pm_r; // @[TLBStorage.scala 63:24]
  reg  data_read_1_0_0_perm_pm_c; // @[TLBStorage.scala 63:24]
  reg [26:0] data_read_1_0_1_tag; // @[TLBStorage.scala 63:24]
  reg [15:0] data_read_1_0_1_asid; // @[TLBStorage.scala 63:24]
  reg [23:0] data_read_1_0_1_ppn; // @[TLBStorage.scala 63:24]
  reg  data_read_1_0_1_perm_pf; // @[TLBStorage.scala 63:24]
  reg  data_read_1_0_1_perm_af; // @[TLBStorage.scala 63:24]
  reg  data_read_1_0_1_perm_a; // @[TLBStorage.scala 63:24]
  reg  data_read_1_0_1_perm_u; // @[TLBStorage.scala 63:24]
  reg  data_read_1_0_1_perm_x; // @[TLBStorage.scala 63:24]
  reg  data_read_1_0_1_perm_r; // @[TLBStorage.scala 63:24]
  reg  data_read_1_0_1_perm_pm_r; // @[TLBStorage.scala 63:24]
  reg  data_read_1_0_1_perm_pm_c; // @[TLBStorage.scala 63:24]
  reg [26:0] data_read_1_0_2_tag; // @[TLBStorage.scala 63:24]
  reg [15:0] data_read_1_0_2_asid; // @[TLBStorage.scala 63:24]
  reg [23:0] data_read_1_0_2_ppn; // @[TLBStorage.scala 63:24]
  reg  data_read_1_0_2_perm_pf; // @[TLBStorage.scala 63:24]
  reg  data_read_1_0_2_perm_af; // @[TLBStorage.scala 63:24]
  reg  data_read_1_0_2_perm_a; // @[TLBStorage.scala 63:24]
  reg  data_read_1_0_2_perm_u; // @[TLBStorage.scala 63:24]
  reg  data_read_1_0_2_perm_x; // @[TLBStorage.scala 63:24]
  reg  data_read_1_0_2_perm_r; // @[TLBStorage.scala 63:24]
  reg  data_read_1_0_2_perm_pm_r; // @[TLBStorage.scala 63:24]
  reg  data_read_1_0_2_perm_pm_c; // @[TLBStorage.scala 63:24]
  reg [26:0] data_read_1_0_3_tag; // @[TLBStorage.scala 63:24]
  reg [15:0] data_read_1_0_3_asid; // @[TLBStorage.scala 63:24]
  reg [23:0] data_read_1_0_3_ppn; // @[TLBStorage.scala 63:24]
  reg  data_read_1_0_3_perm_pf; // @[TLBStorage.scala 63:24]
  reg  data_read_1_0_3_perm_af; // @[TLBStorage.scala 63:24]
  reg  data_read_1_0_3_perm_a; // @[TLBStorage.scala 63:24]
  reg  data_read_1_0_3_perm_u; // @[TLBStorage.scala 63:24]
  reg  data_read_1_0_3_perm_x; // @[TLBStorage.scala 63:24]
  reg  data_read_1_0_3_perm_r; // @[TLBStorage.scala 63:24]
  reg  data_read_1_0_3_perm_pm_r; // @[TLBStorage.scala 63:24]
  reg  data_read_1_0_3_perm_pm_c; // @[TLBStorage.scala 63:24]
  reg [26:0] data_read_1_0_4_tag; // @[TLBStorage.scala 63:24]
  reg [15:0] data_read_1_0_4_asid; // @[TLBStorage.scala 63:24]
  reg [23:0] data_read_1_0_4_ppn; // @[TLBStorage.scala 63:24]
  reg  data_read_1_0_4_perm_pf; // @[TLBStorage.scala 63:24]
  reg  data_read_1_0_4_perm_af; // @[TLBStorage.scala 63:24]
  reg  data_read_1_0_4_perm_a; // @[TLBStorage.scala 63:24]
  reg  data_read_1_0_4_perm_u; // @[TLBStorage.scala 63:24]
  reg  data_read_1_0_4_perm_x; // @[TLBStorage.scala 63:24]
  reg  data_read_1_0_4_perm_r; // @[TLBStorage.scala 63:24]
  reg  data_read_1_0_4_perm_pm_r; // @[TLBStorage.scala 63:24]
  reg  data_read_1_0_4_perm_pm_c; // @[TLBStorage.scala 63:24]
  reg [26:0] data_read_1_0_5_tag; // @[TLBStorage.scala 63:24]
  reg [15:0] data_read_1_0_5_asid; // @[TLBStorage.scala 63:24]
  reg [23:0] data_read_1_0_5_ppn; // @[TLBStorage.scala 63:24]
  reg  data_read_1_0_5_perm_pf; // @[TLBStorage.scala 63:24]
  reg  data_read_1_0_5_perm_af; // @[TLBStorage.scala 63:24]
  reg  data_read_1_0_5_perm_a; // @[TLBStorage.scala 63:24]
  reg  data_read_1_0_5_perm_u; // @[TLBStorage.scala 63:24]
  reg  data_read_1_0_5_perm_x; // @[TLBStorage.scala 63:24]
  reg  data_read_1_0_5_perm_r; // @[TLBStorage.scala 63:24]
  reg  data_read_1_0_5_perm_pm_r; // @[TLBStorage.scala 63:24]
  reg  data_read_1_0_5_perm_pm_c; // @[TLBStorage.scala 63:24]
  reg [26:0] data_read_1_0_6_tag; // @[TLBStorage.scala 63:24]
  reg [15:0] data_read_1_0_6_asid; // @[TLBStorage.scala 63:24]
  reg [23:0] data_read_1_0_6_ppn; // @[TLBStorage.scala 63:24]
  reg  data_read_1_0_6_perm_pf; // @[TLBStorage.scala 63:24]
  reg  data_read_1_0_6_perm_af; // @[TLBStorage.scala 63:24]
  reg  data_read_1_0_6_perm_a; // @[TLBStorage.scala 63:24]
  reg  data_read_1_0_6_perm_u; // @[TLBStorage.scala 63:24]
  reg  data_read_1_0_6_perm_x; // @[TLBStorage.scala 63:24]
  reg  data_read_1_0_6_perm_r; // @[TLBStorage.scala 63:24]
  reg  data_read_1_0_6_perm_pm_r; // @[TLBStorage.scala 63:24]
  reg  data_read_1_0_6_perm_pm_c; // @[TLBStorage.scala 63:24]
  reg [26:0] data_read_1_0_7_tag; // @[TLBStorage.scala 63:24]
  reg [15:0] data_read_1_0_7_asid; // @[TLBStorage.scala 63:24]
  reg [23:0] data_read_1_0_7_ppn; // @[TLBStorage.scala 63:24]
  reg  data_read_1_0_7_perm_pf; // @[TLBStorage.scala 63:24]
  reg  data_read_1_0_7_perm_af; // @[TLBStorage.scala 63:24]
  reg  data_read_1_0_7_perm_a; // @[TLBStorage.scala 63:24]
  reg  data_read_1_0_7_perm_u; // @[TLBStorage.scala 63:24]
  reg  data_read_1_0_7_perm_x; // @[TLBStorage.scala 63:24]
  reg  data_read_1_0_7_perm_r; // @[TLBStorage.scala 63:24]
  reg  data_read_1_0_7_perm_pm_r; // @[TLBStorage.scala 63:24]
  reg  data_read_1_0_7_perm_pm_c; // @[TLBStorage.scala 63:24]
  reg [23:0] data_read_1_1_0_ppn; // @[TLBStorage.scala 63:24]
  reg [23:0] data_read_1_1_1_ppn; // @[TLBStorage.scala 63:24]
  reg [23:0] data_read_1_1_2_ppn; // @[TLBStorage.scala 63:24]
  reg [23:0] data_read_1_1_3_ppn; // @[TLBStorage.scala 63:24]
  reg [23:0] data_read_1_1_4_ppn; // @[TLBStorage.scala 63:24]
  reg [23:0] data_read_1_1_5_ppn; // @[TLBStorage.scala 63:24]
  reg [23:0] data_read_1_1_6_ppn; // @[TLBStorage.scala 63:24]
  reg [23:0] data_read_1_1_7_ppn; // @[TLBStorage.scala 63:24]
  reg [7:0] bank_index_1_0; // @[TLBStorage.scala 64:25]
  reg [7:0] bank_index_1_1; // @[TLBStorage.scala 64:25]
  wire [23:0] _io_rdata_1_0_T_218 = bank_index_1_0[0] ? data_read_1_0_0_ppn : 24'h0; // @[Mux.scala 27:73]
  wire [23:0] _io_rdata_1_0_T_219 = bank_index_1_0[1] ? data_read_1_0_1_ppn : 24'h0; // @[Mux.scala 27:73]
  wire [23:0] _io_rdata_1_0_T_220 = bank_index_1_0[2] ? data_read_1_0_2_ppn : 24'h0; // @[Mux.scala 27:73]
  wire [23:0] _io_rdata_1_0_T_221 = bank_index_1_0[3] ? data_read_1_0_3_ppn : 24'h0; // @[Mux.scala 27:73]
  wire [23:0] _io_rdata_1_0_T_222 = bank_index_1_0[4] ? data_read_1_0_4_ppn : 24'h0; // @[Mux.scala 27:73]
  wire [23:0] _io_rdata_1_0_T_223 = bank_index_1_0[5] ? data_read_1_0_5_ppn : 24'h0; // @[Mux.scala 27:73]
  wire [23:0] _io_rdata_1_0_T_224 = bank_index_1_0[6] ? data_read_1_0_6_ppn : 24'h0; // @[Mux.scala 27:73]
  wire [23:0] _io_rdata_1_0_T_225 = bank_index_1_0[7] ? data_read_1_0_7_ppn : 24'h0; // @[Mux.scala 27:73]
  wire [23:0] _io_rdata_1_0_T_226 = _io_rdata_1_0_T_218 | _io_rdata_1_0_T_219; // @[Mux.scala 27:73]
  wire [23:0] _io_rdata_1_0_T_227 = _io_rdata_1_0_T_226 | _io_rdata_1_0_T_220; // @[Mux.scala 27:73]
  wire [23:0] _io_rdata_1_0_T_228 = _io_rdata_1_0_T_227 | _io_rdata_1_0_T_221; // @[Mux.scala 27:73]
  wire [23:0] _io_rdata_1_0_T_229 = _io_rdata_1_0_T_228 | _io_rdata_1_0_T_222; // @[Mux.scala 27:73]
  wire [23:0] _io_rdata_1_0_T_230 = _io_rdata_1_0_T_229 | _io_rdata_1_0_T_223; // @[Mux.scala 27:73]
  wire [23:0] _io_rdata_1_0_T_231 = _io_rdata_1_0_T_230 | _io_rdata_1_0_T_224; // @[Mux.scala 27:73]
  wire [15:0] _io_rdata_1_0_T_233 = bank_index_1_0[0] ? data_read_1_0_0_asid : 16'h0; // @[Mux.scala 27:73]
  wire [15:0] _io_rdata_1_0_T_234 = bank_index_1_0[1] ? data_read_1_0_1_asid : 16'h0; // @[Mux.scala 27:73]
  wire [15:0] _io_rdata_1_0_T_235 = bank_index_1_0[2] ? data_read_1_0_2_asid : 16'h0; // @[Mux.scala 27:73]
  wire [15:0] _io_rdata_1_0_T_236 = bank_index_1_0[3] ? data_read_1_0_3_asid : 16'h0; // @[Mux.scala 27:73]
  wire [15:0] _io_rdata_1_0_T_237 = bank_index_1_0[4] ? data_read_1_0_4_asid : 16'h0; // @[Mux.scala 27:73]
  wire [15:0] _io_rdata_1_0_T_238 = bank_index_1_0[5] ? data_read_1_0_5_asid : 16'h0; // @[Mux.scala 27:73]
  wire [15:0] _io_rdata_1_0_T_239 = bank_index_1_0[6] ? data_read_1_0_6_asid : 16'h0; // @[Mux.scala 27:73]
  wire [15:0] _io_rdata_1_0_T_240 = bank_index_1_0[7] ? data_read_1_0_7_asid : 16'h0; // @[Mux.scala 27:73]
  wire [15:0] _io_rdata_1_0_T_241 = _io_rdata_1_0_T_233 | _io_rdata_1_0_T_234; // @[Mux.scala 27:73]
  wire [15:0] _io_rdata_1_0_T_242 = _io_rdata_1_0_T_241 | _io_rdata_1_0_T_235; // @[Mux.scala 27:73]
  wire [15:0] _io_rdata_1_0_T_243 = _io_rdata_1_0_T_242 | _io_rdata_1_0_T_236; // @[Mux.scala 27:73]
  wire [15:0] _io_rdata_1_0_T_244 = _io_rdata_1_0_T_243 | _io_rdata_1_0_T_237; // @[Mux.scala 27:73]
  wire [15:0] _io_rdata_1_0_T_245 = _io_rdata_1_0_T_244 | _io_rdata_1_0_T_238; // @[Mux.scala 27:73]
  wire [15:0] _io_rdata_1_0_T_246 = _io_rdata_1_0_T_245 | _io_rdata_1_0_T_239; // @[Mux.scala 27:73]
  wire [26:0] _io_rdata_1_0_T_248 = bank_index_1_0[0] ? data_read_1_0_0_tag : 27'h0; // @[Mux.scala 27:73]
  wire [26:0] _io_rdata_1_0_T_249 = bank_index_1_0[1] ? data_read_1_0_1_tag : 27'h0; // @[Mux.scala 27:73]
  wire [26:0] _io_rdata_1_0_T_250 = bank_index_1_0[2] ? data_read_1_0_2_tag : 27'h0; // @[Mux.scala 27:73]
  wire [26:0] _io_rdata_1_0_T_251 = bank_index_1_0[3] ? data_read_1_0_3_tag : 27'h0; // @[Mux.scala 27:73]
  wire [26:0] _io_rdata_1_0_T_252 = bank_index_1_0[4] ? data_read_1_0_4_tag : 27'h0; // @[Mux.scala 27:73]
  wire [26:0] _io_rdata_1_0_T_253 = bank_index_1_0[5] ? data_read_1_0_5_tag : 27'h0; // @[Mux.scala 27:73]
  wire [26:0] _io_rdata_1_0_T_254 = bank_index_1_0[6] ? data_read_1_0_6_tag : 27'h0; // @[Mux.scala 27:73]
  wire [26:0] _io_rdata_1_0_T_255 = bank_index_1_0[7] ? data_read_1_0_7_tag : 27'h0; // @[Mux.scala 27:73]
  wire [26:0] _io_rdata_1_0_T_256 = _io_rdata_1_0_T_248 | _io_rdata_1_0_T_249; // @[Mux.scala 27:73]
  wire [26:0] _io_rdata_1_0_T_257 = _io_rdata_1_0_T_256 | _io_rdata_1_0_T_250; // @[Mux.scala 27:73]
  wire [26:0] _io_rdata_1_0_T_258 = _io_rdata_1_0_T_257 | _io_rdata_1_0_T_251; // @[Mux.scala 27:73]
  wire [26:0] _io_rdata_1_0_T_259 = _io_rdata_1_0_T_258 | _io_rdata_1_0_T_252; // @[Mux.scala 27:73]
  wire [26:0] _io_rdata_1_0_T_260 = _io_rdata_1_0_T_259 | _io_rdata_1_0_T_253; // @[Mux.scala 27:73]
  wire [26:0] _io_rdata_1_0_T_261 = _io_rdata_1_0_T_260 | _io_rdata_1_0_T_254; // @[Mux.scala 27:73]
  wire [23:0] _io_rdata_1_1_T_218 = bank_index_1_1[0] ? data_read_1_1_0_ppn : 24'h0; // @[Mux.scala 27:73]
  wire [23:0] _io_rdata_1_1_T_219 = bank_index_1_1[1] ? data_read_1_1_1_ppn : 24'h0; // @[Mux.scala 27:73]
  wire [23:0] _io_rdata_1_1_T_220 = bank_index_1_1[2] ? data_read_1_1_2_ppn : 24'h0; // @[Mux.scala 27:73]
  wire [23:0] _io_rdata_1_1_T_221 = bank_index_1_1[3] ? data_read_1_1_3_ppn : 24'h0; // @[Mux.scala 27:73]
  wire [23:0] _io_rdata_1_1_T_222 = bank_index_1_1[4] ? data_read_1_1_4_ppn : 24'h0; // @[Mux.scala 27:73]
  wire [23:0] _io_rdata_1_1_T_223 = bank_index_1_1[5] ? data_read_1_1_5_ppn : 24'h0; // @[Mux.scala 27:73]
  wire [23:0] _io_rdata_1_1_T_224 = bank_index_1_1[6] ? data_read_1_1_6_ppn : 24'h0; // @[Mux.scala 27:73]
  wire [23:0] _io_rdata_1_1_T_225 = bank_index_1_1[7] ? data_read_1_1_7_ppn : 24'h0; // @[Mux.scala 27:73]
  wire [23:0] _io_rdata_1_1_T_226 = _io_rdata_1_1_T_218 | _io_rdata_1_1_T_219; // @[Mux.scala 27:73]
  wire [23:0] _io_rdata_1_1_T_227 = _io_rdata_1_1_T_226 | _io_rdata_1_1_T_220; // @[Mux.scala 27:73]
  wire [23:0] _io_rdata_1_1_T_228 = _io_rdata_1_1_T_227 | _io_rdata_1_1_T_221; // @[Mux.scala 27:73]
  wire [23:0] _io_rdata_1_1_T_229 = _io_rdata_1_1_T_228 | _io_rdata_1_1_T_222; // @[Mux.scala 27:73]
  wire [23:0] _io_rdata_1_1_T_230 = _io_rdata_1_1_T_229 | _io_rdata_1_1_T_223; // @[Mux.scala 27:73]
  wire [23:0] _io_rdata_1_1_T_231 = _io_rdata_1_1_T_230 | _io_rdata_1_1_T_224; // @[Mux.scala 27:73]
  wire  _T_1 = io_waddr[3:1] == 3'h0; // @[TLBStorage.scala 80:42]
  wire  _T_5 = io_waddr[3:1] == 3'h1; // @[TLBStorage.scala 80:42]
  wire  _T_9 = io_waddr[3:1] == 3'h2; // @[TLBStorage.scala 80:42]
  wire  _T_13 = io_waddr[3:1] == 3'h3; // @[TLBStorage.scala 80:42]
  wire  _T_17 = io_waddr[3:1] == 3'h4; // @[TLBStorage.scala 80:42]
  wire  _T_21 = io_waddr[3:1] == 3'h5; // @[TLBStorage.scala 80:42]
  wire  _T_25 = io_waddr[3:1] == 3'h6; // @[TLBStorage.scala 80:42]
  wire  _T_29 = io_waddr[3:1] == 3'h7; // @[TLBStorage.scala 80:42]
  assign dataBanks_0_tag_data_read_0_0_MPORT_en = 1'h1;
  assign dataBanks_0_tag_data_read_0_0_MPORT_addr = io_raddr_0[0];
  assign dataBanks_0_tag_data_read_0_0_MPORT_data = dataBanks_0_tag[dataBanks_0_tag_data_read_0_0_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_0_tag_data_read_1_0_MPORT_en = 1'h1;
  assign dataBanks_0_tag_data_read_1_0_MPORT_addr = io_raddr_0[0];
  assign dataBanks_0_tag_data_read_1_0_MPORT_data = dataBanks_0_tag[dataBanks_0_tag_data_read_1_0_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_0_tag_data_read_0_0_MPORT_1_en = 1'h1;
  assign dataBanks_0_tag_data_read_0_0_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_0_tag_data_read_0_0_MPORT_1_data = dataBanks_0_tag[dataBanks_0_tag_data_read_0_0_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_0_tag_data_read_1_0_MPORT_1_en = 1'h1;
  assign dataBanks_0_tag_data_read_1_0_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_0_tag_data_read_1_0_MPORT_1_data = dataBanks_0_tag[dataBanks_0_tag_data_read_1_0_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_0_tag_MPORT_data = io_wdata_tag;
  assign dataBanks_0_tag_MPORT_addr = io_waddr[0];
  assign dataBanks_0_tag_MPORT_mask = 1'h1;
  assign dataBanks_0_tag_MPORT_en = io_wen & _T_1;
  assign dataBanks_0_asid_data_read_0_0_MPORT_en = 1'h1;
  assign dataBanks_0_asid_data_read_0_0_MPORT_addr = io_raddr_0[0];
  assign dataBanks_0_asid_data_read_0_0_MPORT_data = dataBanks_0_asid[dataBanks_0_asid_data_read_0_0_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_0_asid_data_read_1_0_MPORT_en = 1'h1;
  assign dataBanks_0_asid_data_read_1_0_MPORT_addr = io_raddr_0[0];
  assign dataBanks_0_asid_data_read_1_0_MPORT_data = dataBanks_0_asid[dataBanks_0_asid_data_read_1_0_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_0_asid_data_read_0_0_MPORT_1_en = 1'h1;
  assign dataBanks_0_asid_data_read_0_0_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_0_asid_data_read_0_0_MPORT_1_data = dataBanks_0_asid[dataBanks_0_asid_data_read_0_0_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_0_asid_data_read_1_0_MPORT_1_en = 1'h1;
  assign dataBanks_0_asid_data_read_1_0_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_0_asid_data_read_1_0_MPORT_1_data = dataBanks_0_asid[dataBanks_0_asid_data_read_1_0_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_0_asid_MPORT_data = io_wdata_asid;
  assign dataBanks_0_asid_MPORT_addr = io_waddr[0];
  assign dataBanks_0_asid_MPORT_mask = 1'h1;
  assign dataBanks_0_asid_MPORT_en = io_wen & _T_1;
  assign dataBanks_0_ppn_data_read_0_0_MPORT_en = 1'h1;
  assign dataBanks_0_ppn_data_read_0_0_MPORT_addr = io_raddr_0[0];
  assign dataBanks_0_ppn_data_read_0_0_MPORT_data = dataBanks_0_ppn[dataBanks_0_ppn_data_read_0_0_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_0_ppn_data_read_1_0_MPORT_en = 1'h1;
  assign dataBanks_0_ppn_data_read_1_0_MPORT_addr = io_raddr_0[0];
  assign dataBanks_0_ppn_data_read_1_0_MPORT_data = dataBanks_0_ppn[dataBanks_0_ppn_data_read_1_0_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_0_ppn_data_read_0_0_MPORT_1_en = 1'h1;
  assign dataBanks_0_ppn_data_read_0_0_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_0_ppn_data_read_0_0_MPORT_1_data = dataBanks_0_ppn[dataBanks_0_ppn_data_read_0_0_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_0_ppn_data_read_1_0_MPORT_1_en = 1'h1;
  assign dataBanks_0_ppn_data_read_1_0_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_0_ppn_data_read_1_0_MPORT_1_data = dataBanks_0_ppn[dataBanks_0_ppn_data_read_1_0_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_0_ppn_MPORT_data = io_wdata_ppn;
  assign dataBanks_0_ppn_MPORT_addr = io_waddr[0];
  assign dataBanks_0_ppn_MPORT_mask = 1'h1;
  assign dataBanks_0_ppn_MPORT_en = io_wen & _T_1;
  assign dataBanks_0_perm_pf_data_read_0_0_MPORT_en = 1'h1;
  assign dataBanks_0_perm_pf_data_read_0_0_MPORT_addr = io_raddr_0[0];
  assign dataBanks_0_perm_pf_data_read_0_0_MPORT_data =
    dataBanks_0_perm_pf[dataBanks_0_perm_pf_data_read_0_0_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_0_perm_pf_data_read_1_0_MPORT_en = 1'h1;
  assign dataBanks_0_perm_pf_data_read_1_0_MPORT_addr = io_raddr_0[0];
  assign dataBanks_0_perm_pf_data_read_1_0_MPORT_data =
    dataBanks_0_perm_pf[dataBanks_0_perm_pf_data_read_1_0_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_0_perm_pf_data_read_0_0_MPORT_1_en = 1'h1;
  assign dataBanks_0_perm_pf_data_read_0_0_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_0_perm_pf_data_read_0_0_MPORT_1_data =
    dataBanks_0_perm_pf[dataBanks_0_perm_pf_data_read_0_0_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_0_perm_pf_data_read_1_0_MPORT_1_en = 1'h1;
  assign dataBanks_0_perm_pf_data_read_1_0_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_0_perm_pf_data_read_1_0_MPORT_1_data =
    dataBanks_0_perm_pf[dataBanks_0_perm_pf_data_read_1_0_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_0_perm_pf_MPORT_data = io_wdata_perm_pf;
  assign dataBanks_0_perm_pf_MPORT_addr = io_waddr[0];
  assign dataBanks_0_perm_pf_MPORT_mask = 1'h1;
  assign dataBanks_0_perm_pf_MPORT_en = io_wen & _T_1;
  assign dataBanks_0_perm_af_data_read_0_0_MPORT_en = 1'h1;
  assign dataBanks_0_perm_af_data_read_0_0_MPORT_addr = io_raddr_0[0];
  assign dataBanks_0_perm_af_data_read_0_0_MPORT_data =
    dataBanks_0_perm_af[dataBanks_0_perm_af_data_read_0_0_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_0_perm_af_data_read_1_0_MPORT_en = 1'h1;
  assign dataBanks_0_perm_af_data_read_1_0_MPORT_addr = io_raddr_0[0];
  assign dataBanks_0_perm_af_data_read_1_0_MPORT_data =
    dataBanks_0_perm_af[dataBanks_0_perm_af_data_read_1_0_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_0_perm_af_data_read_0_0_MPORT_1_en = 1'h1;
  assign dataBanks_0_perm_af_data_read_0_0_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_0_perm_af_data_read_0_0_MPORT_1_data =
    dataBanks_0_perm_af[dataBanks_0_perm_af_data_read_0_0_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_0_perm_af_data_read_1_0_MPORT_1_en = 1'h1;
  assign dataBanks_0_perm_af_data_read_1_0_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_0_perm_af_data_read_1_0_MPORT_1_data =
    dataBanks_0_perm_af[dataBanks_0_perm_af_data_read_1_0_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_0_perm_af_MPORT_data = io_wdata_perm_af;
  assign dataBanks_0_perm_af_MPORT_addr = io_waddr[0];
  assign dataBanks_0_perm_af_MPORT_mask = 1'h1;
  assign dataBanks_0_perm_af_MPORT_en = io_wen & _T_1;
  assign dataBanks_0_perm_d_data_read_0_0_MPORT_en = 1'h1;
  assign dataBanks_0_perm_d_data_read_0_0_MPORT_addr = io_raddr_0[0];
  assign dataBanks_0_perm_d_data_read_0_0_MPORT_data = dataBanks_0_perm_d[dataBanks_0_perm_d_data_read_0_0_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_0_perm_d_data_read_1_0_MPORT_en = 1'h1;
  assign dataBanks_0_perm_d_data_read_1_0_MPORT_addr = io_raddr_0[0];
  assign dataBanks_0_perm_d_data_read_1_0_MPORT_data = dataBanks_0_perm_d[dataBanks_0_perm_d_data_read_1_0_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_0_perm_d_data_read_0_0_MPORT_1_en = 1'h1;
  assign dataBanks_0_perm_d_data_read_0_0_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_0_perm_d_data_read_0_0_MPORT_1_data =
    dataBanks_0_perm_d[dataBanks_0_perm_d_data_read_0_0_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_0_perm_d_data_read_1_0_MPORT_1_en = 1'h1;
  assign dataBanks_0_perm_d_data_read_1_0_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_0_perm_d_data_read_1_0_MPORT_1_data =
    dataBanks_0_perm_d[dataBanks_0_perm_d_data_read_1_0_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_0_perm_d_MPORT_data = io_wdata_perm_d;
  assign dataBanks_0_perm_d_MPORT_addr = io_waddr[0];
  assign dataBanks_0_perm_d_MPORT_mask = 1'h1;
  assign dataBanks_0_perm_d_MPORT_en = io_wen & _T_1;
  assign dataBanks_0_perm_a_data_read_0_0_MPORT_en = 1'h1;
  assign dataBanks_0_perm_a_data_read_0_0_MPORT_addr = io_raddr_0[0];
  assign dataBanks_0_perm_a_data_read_0_0_MPORT_data = dataBanks_0_perm_a[dataBanks_0_perm_a_data_read_0_0_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_0_perm_a_data_read_1_0_MPORT_en = 1'h1;
  assign dataBanks_0_perm_a_data_read_1_0_MPORT_addr = io_raddr_0[0];
  assign dataBanks_0_perm_a_data_read_1_0_MPORT_data = dataBanks_0_perm_a[dataBanks_0_perm_a_data_read_1_0_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_0_perm_a_data_read_0_0_MPORT_1_en = 1'h1;
  assign dataBanks_0_perm_a_data_read_0_0_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_0_perm_a_data_read_0_0_MPORT_1_data =
    dataBanks_0_perm_a[dataBanks_0_perm_a_data_read_0_0_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_0_perm_a_data_read_1_0_MPORT_1_en = 1'h1;
  assign dataBanks_0_perm_a_data_read_1_0_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_0_perm_a_data_read_1_0_MPORT_1_data =
    dataBanks_0_perm_a[dataBanks_0_perm_a_data_read_1_0_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_0_perm_a_MPORT_data = io_wdata_perm_a;
  assign dataBanks_0_perm_a_MPORT_addr = io_waddr[0];
  assign dataBanks_0_perm_a_MPORT_mask = 1'h1;
  assign dataBanks_0_perm_a_MPORT_en = io_wen & _T_1;
  assign dataBanks_0_perm_u_data_read_0_0_MPORT_en = 1'h1;
  assign dataBanks_0_perm_u_data_read_0_0_MPORT_addr = io_raddr_0[0];
  assign dataBanks_0_perm_u_data_read_0_0_MPORT_data = dataBanks_0_perm_u[dataBanks_0_perm_u_data_read_0_0_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_0_perm_u_data_read_1_0_MPORT_en = 1'h1;
  assign dataBanks_0_perm_u_data_read_1_0_MPORT_addr = io_raddr_0[0];
  assign dataBanks_0_perm_u_data_read_1_0_MPORT_data = dataBanks_0_perm_u[dataBanks_0_perm_u_data_read_1_0_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_0_perm_u_data_read_0_0_MPORT_1_en = 1'h1;
  assign dataBanks_0_perm_u_data_read_0_0_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_0_perm_u_data_read_0_0_MPORT_1_data =
    dataBanks_0_perm_u[dataBanks_0_perm_u_data_read_0_0_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_0_perm_u_data_read_1_0_MPORT_1_en = 1'h1;
  assign dataBanks_0_perm_u_data_read_1_0_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_0_perm_u_data_read_1_0_MPORT_1_data =
    dataBanks_0_perm_u[dataBanks_0_perm_u_data_read_1_0_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_0_perm_u_MPORT_data = io_wdata_perm_u;
  assign dataBanks_0_perm_u_MPORT_addr = io_waddr[0];
  assign dataBanks_0_perm_u_MPORT_mask = 1'h1;
  assign dataBanks_0_perm_u_MPORT_en = io_wen & _T_1;
  assign dataBanks_0_perm_x_data_read_0_0_MPORT_en = 1'h1;
  assign dataBanks_0_perm_x_data_read_0_0_MPORT_addr = io_raddr_0[0];
  assign dataBanks_0_perm_x_data_read_0_0_MPORT_data = dataBanks_0_perm_x[dataBanks_0_perm_x_data_read_0_0_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_0_perm_x_data_read_1_0_MPORT_en = 1'h1;
  assign dataBanks_0_perm_x_data_read_1_0_MPORT_addr = io_raddr_0[0];
  assign dataBanks_0_perm_x_data_read_1_0_MPORT_data = dataBanks_0_perm_x[dataBanks_0_perm_x_data_read_1_0_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_0_perm_x_data_read_0_0_MPORT_1_en = 1'h1;
  assign dataBanks_0_perm_x_data_read_0_0_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_0_perm_x_data_read_0_0_MPORT_1_data =
    dataBanks_0_perm_x[dataBanks_0_perm_x_data_read_0_0_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_0_perm_x_data_read_1_0_MPORT_1_en = 1'h1;
  assign dataBanks_0_perm_x_data_read_1_0_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_0_perm_x_data_read_1_0_MPORT_1_data =
    dataBanks_0_perm_x[dataBanks_0_perm_x_data_read_1_0_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_0_perm_x_MPORT_data = io_wdata_perm_x;
  assign dataBanks_0_perm_x_MPORT_addr = io_waddr[0];
  assign dataBanks_0_perm_x_MPORT_mask = 1'h1;
  assign dataBanks_0_perm_x_MPORT_en = io_wen & _T_1;
  assign dataBanks_0_perm_wdata_read_0_0_MPORT_en = 1'h1;
  assign dataBanks_0_perm_wdata_read_0_0_MPORT_addr = io_raddr_0[0];
  assign dataBanks_0_perm_wdata_read_0_0_MPORT_data = dataBanks_0_perm_w[dataBanks_0_perm_wdata_read_0_0_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_0_perm_wdata_read_1_0_MPORT_en = 1'h1;
  assign dataBanks_0_perm_wdata_read_1_0_MPORT_addr = io_raddr_0[0];
  assign dataBanks_0_perm_wdata_read_1_0_MPORT_data = dataBanks_0_perm_w[dataBanks_0_perm_wdata_read_1_0_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_0_perm_wdata_read_0_0_MPORT_1_en = 1'h1;
  assign dataBanks_0_perm_wdata_read_0_0_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_0_perm_wdata_read_0_0_MPORT_1_data =
    dataBanks_0_perm_w[dataBanks_0_perm_wdata_read_0_0_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_0_perm_wdata_read_1_0_MPORT_1_en = 1'h1;
  assign dataBanks_0_perm_wdata_read_1_0_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_0_perm_wdata_read_1_0_MPORT_1_data =
    dataBanks_0_perm_w[dataBanks_0_perm_wdata_read_1_0_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_0_perm_wMPORT_data = io_wdata_perm_w;
  assign dataBanks_0_perm_wMPORT_addr = io_waddr[0];
  assign dataBanks_0_perm_wMPORT_mask = 1'h1;
  assign dataBanks_0_perm_wMPORT_en = io_wen & _T_1;
  assign dataBanks_0_perm_rdata_read_0_0_MPORT_en = 1'h1;
  assign dataBanks_0_perm_rdata_read_0_0_MPORT_addr = io_raddr_0[0];
  assign dataBanks_0_perm_rdata_read_0_0_MPORT_data = dataBanks_0_perm_r[dataBanks_0_perm_rdata_read_0_0_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_0_perm_rdata_read_1_0_MPORT_en = 1'h1;
  assign dataBanks_0_perm_rdata_read_1_0_MPORT_addr = io_raddr_0[0];
  assign dataBanks_0_perm_rdata_read_1_0_MPORT_data = dataBanks_0_perm_r[dataBanks_0_perm_rdata_read_1_0_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_0_perm_rdata_read_0_0_MPORT_1_en = 1'h1;
  assign dataBanks_0_perm_rdata_read_0_0_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_0_perm_rdata_read_0_0_MPORT_1_data =
    dataBanks_0_perm_r[dataBanks_0_perm_rdata_read_0_0_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_0_perm_rdata_read_1_0_MPORT_1_en = 1'h1;
  assign dataBanks_0_perm_rdata_read_1_0_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_0_perm_rdata_read_1_0_MPORT_1_data =
    dataBanks_0_perm_r[dataBanks_0_perm_rdata_read_1_0_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_0_perm_rMPORT_data = io_wdata_perm_r;
  assign dataBanks_0_perm_rMPORT_addr = io_waddr[0];
  assign dataBanks_0_perm_rMPORT_mask = 1'h1;
  assign dataBanks_0_perm_rMPORT_en = io_wen & _T_1;
  assign dataBanks_0_perm_pm_rdata_read_0_0_MPORT_en = 1'h1;
  assign dataBanks_0_perm_pm_rdata_read_0_0_MPORT_addr = io_raddr_0[0];
  assign dataBanks_0_perm_pm_rdata_read_0_0_MPORT_data =
    dataBanks_0_perm_pm_r[dataBanks_0_perm_pm_rdata_read_0_0_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_0_perm_pm_rdata_read_1_0_MPORT_en = 1'h1;
  assign dataBanks_0_perm_pm_rdata_read_1_0_MPORT_addr = io_raddr_0[0];
  assign dataBanks_0_perm_pm_rdata_read_1_0_MPORT_data =
    dataBanks_0_perm_pm_r[dataBanks_0_perm_pm_rdata_read_1_0_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_0_perm_pm_rdata_read_0_0_MPORT_1_en = 1'h1;
  assign dataBanks_0_perm_pm_rdata_read_0_0_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_0_perm_pm_rdata_read_0_0_MPORT_1_data =
    dataBanks_0_perm_pm_r[dataBanks_0_perm_pm_rdata_read_0_0_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_0_perm_pm_rdata_read_1_0_MPORT_1_en = 1'h1;
  assign dataBanks_0_perm_pm_rdata_read_1_0_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_0_perm_pm_rdata_read_1_0_MPORT_1_data =
    dataBanks_0_perm_pm_r[dataBanks_0_perm_pm_rdata_read_1_0_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_0_perm_pm_rMPORT_data = io_wdata_perm_pm_r;
  assign dataBanks_0_perm_pm_rMPORT_addr = io_waddr[0];
  assign dataBanks_0_perm_pm_rMPORT_mask = 1'h1;
  assign dataBanks_0_perm_pm_rMPORT_en = io_wen & _T_1;
  assign dataBanks_0_perm_pm_wdata_read_0_0_MPORT_en = 1'h1;
  assign dataBanks_0_perm_pm_wdata_read_0_0_MPORT_addr = io_raddr_0[0];
  assign dataBanks_0_perm_pm_wdata_read_0_0_MPORT_data =
    dataBanks_0_perm_pm_w[dataBanks_0_perm_pm_wdata_read_0_0_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_0_perm_pm_wdata_read_1_0_MPORT_en = 1'h1;
  assign dataBanks_0_perm_pm_wdata_read_1_0_MPORT_addr = io_raddr_0[0];
  assign dataBanks_0_perm_pm_wdata_read_1_0_MPORT_data =
    dataBanks_0_perm_pm_w[dataBanks_0_perm_pm_wdata_read_1_0_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_0_perm_pm_wdata_read_0_0_MPORT_1_en = 1'h1;
  assign dataBanks_0_perm_pm_wdata_read_0_0_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_0_perm_pm_wdata_read_0_0_MPORT_1_data =
    dataBanks_0_perm_pm_w[dataBanks_0_perm_pm_wdata_read_0_0_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_0_perm_pm_wdata_read_1_0_MPORT_1_en = 1'h1;
  assign dataBanks_0_perm_pm_wdata_read_1_0_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_0_perm_pm_wdata_read_1_0_MPORT_1_data =
    dataBanks_0_perm_pm_w[dataBanks_0_perm_pm_wdata_read_1_0_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_0_perm_pm_wMPORT_data = io_wdata_perm_pm_w;
  assign dataBanks_0_perm_pm_wMPORT_addr = io_waddr[0];
  assign dataBanks_0_perm_pm_wMPORT_mask = 1'h1;
  assign dataBanks_0_perm_pm_wMPORT_en = io_wen & _T_1;
  assign dataBanks_0_perm_pm_c_data_read_0_0_MPORT_en = 1'h1;
  assign dataBanks_0_perm_pm_c_data_read_0_0_MPORT_addr = io_raddr_0[0];
  assign dataBanks_0_perm_pm_c_data_read_0_0_MPORT_data =
    dataBanks_0_perm_pm_c[dataBanks_0_perm_pm_c_data_read_0_0_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_0_perm_pm_c_data_read_1_0_MPORT_en = 1'h1;
  assign dataBanks_0_perm_pm_c_data_read_1_0_MPORT_addr = io_raddr_0[0];
  assign dataBanks_0_perm_pm_c_data_read_1_0_MPORT_data =
    dataBanks_0_perm_pm_c[dataBanks_0_perm_pm_c_data_read_1_0_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_0_perm_pm_c_data_read_0_0_MPORT_1_en = 1'h1;
  assign dataBanks_0_perm_pm_c_data_read_0_0_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_0_perm_pm_c_data_read_0_0_MPORT_1_data =
    dataBanks_0_perm_pm_c[dataBanks_0_perm_pm_c_data_read_0_0_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_0_perm_pm_c_data_read_1_0_MPORT_1_en = 1'h1;
  assign dataBanks_0_perm_pm_c_data_read_1_0_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_0_perm_pm_c_data_read_1_0_MPORT_1_data =
    dataBanks_0_perm_pm_c[dataBanks_0_perm_pm_c_data_read_1_0_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_0_perm_pm_c_MPORT_data = io_wdata_perm_pm_c;
  assign dataBanks_0_perm_pm_c_MPORT_addr = io_waddr[0];
  assign dataBanks_0_perm_pm_c_MPORT_mask = 1'h1;
  assign dataBanks_0_perm_pm_c_MPORT_en = io_wen & _T_1;
  assign dataBanks_1_tag_data_read_0_1_MPORT_en = 1'h1;
  assign dataBanks_1_tag_data_read_0_1_MPORT_addr = io_raddr_0[0];
  assign dataBanks_1_tag_data_read_0_1_MPORT_data = dataBanks_1_tag[dataBanks_1_tag_data_read_0_1_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_1_tag_data_read_1_1_MPORT_en = 1'h1;
  assign dataBanks_1_tag_data_read_1_1_MPORT_addr = io_raddr_0[0];
  assign dataBanks_1_tag_data_read_1_1_MPORT_data = dataBanks_1_tag[dataBanks_1_tag_data_read_1_1_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_1_tag_data_read_0_1_MPORT_1_en = 1'h1;
  assign dataBanks_1_tag_data_read_0_1_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_1_tag_data_read_0_1_MPORT_1_data = dataBanks_1_tag[dataBanks_1_tag_data_read_0_1_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_1_tag_data_read_1_1_MPORT_1_en = 1'h1;
  assign dataBanks_1_tag_data_read_1_1_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_1_tag_data_read_1_1_MPORT_1_data = dataBanks_1_tag[dataBanks_1_tag_data_read_1_1_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_1_tag_MPORT_1_data = io_wdata_tag;
  assign dataBanks_1_tag_MPORT_1_addr = io_waddr[0];
  assign dataBanks_1_tag_MPORT_1_mask = 1'h1;
  assign dataBanks_1_tag_MPORT_1_en = io_wen & _T_5;
  assign dataBanks_1_asid_data_read_0_1_MPORT_en = 1'h1;
  assign dataBanks_1_asid_data_read_0_1_MPORT_addr = io_raddr_0[0];
  assign dataBanks_1_asid_data_read_0_1_MPORT_data = dataBanks_1_asid[dataBanks_1_asid_data_read_0_1_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_1_asid_data_read_1_1_MPORT_en = 1'h1;
  assign dataBanks_1_asid_data_read_1_1_MPORT_addr = io_raddr_0[0];
  assign dataBanks_1_asid_data_read_1_1_MPORT_data = dataBanks_1_asid[dataBanks_1_asid_data_read_1_1_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_1_asid_data_read_0_1_MPORT_1_en = 1'h1;
  assign dataBanks_1_asid_data_read_0_1_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_1_asid_data_read_0_1_MPORT_1_data = dataBanks_1_asid[dataBanks_1_asid_data_read_0_1_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_1_asid_data_read_1_1_MPORT_1_en = 1'h1;
  assign dataBanks_1_asid_data_read_1_1_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_1_asid_data_read_1_1_MPORT_1_data = dataBanks_1_asid[dataBanks_1_asid_data_read_1_1_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_1_asid_MPORT_1_data = io_wdata_asid;
  assign dataBanks_1_asid_MPORT_1_addr = io_waddr[0];
  assign dataBanks_1_asid_MPORT_1_mask = 1'h1;
  assign dataBanks_1_asid_MPORT_1_en = io_wen & _T_5;
  assign dataBanks_1_ppn_data_read_0_1_MPORT_en = 1'h1;
  assign dataBanks_1_ppn_data_read_0_1_MPORT_addr = io_raddr_0[0];
  assign dataBanks_1_ppn_data_read_0_1_MPORT_data = dataBanks_1_ppn[dataBanks_1_ppn_data_read_0_1_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_1_ppn_data_read_1_1_MPORT_en = 1'h1;
  assign dataBanks_1_ppn_data_read_1_1_MPORT_addr = io_raddr_0[0];
  assign dataBanks_1_ppn_data_read_1_1_MPORT_data = dataBanks_1_ppn[dataBanks_1_ppn_data_read_1_1_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_1_ppn_data_read_0_1_MPORT_1_en = 1'h1;
  assign dataBanks_1_ppn_data_read_0_1_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_1_ppn_data_read_0_1_MPORT_1_data = dataBanks_1_ppn[dataBanks_1_ppn_data_read_0_1_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_1_ppn_data_read_1_1_MPORT_1_en = 1'h1;
  assign dataBanks_1_ppn_data_read_1_1_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_1_ppn_data_read_1_1_MPORT_1_data = dataBanks_1_ppn[dataBanks_1_ppn_data_read_1_1_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_1_ppn_MPORT_1_data = io_wdata_ppn;
  assign dataBanks_1_ppn_MPORT_1_addr = io_waddr[0];
  assign dataBanks_1_ppn_MPORT_1_mask = 1'h1;
  assign dataBanks_1_ppn_MPORT_1_en = io_wen & _T_5;
  assign dataBanks_1_perm_pf_data_read_0_1_MPORT_en = 1'h1;
  assign dataBanks_1_perm_pf_data_read_0_1_MPORT_addr = io_raddr_0[0];
  assign dataBanks_1_perm_pf_data_read_0_1_MPORT_data =
    dataBanks_1_perm_pf[dataBanks_1_perm_pf_data_read_0_1_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_1_perm_pf_data_read_1_1_MPORT_en = 1'h1;
  assign dataBanks_1_perm_pf_data_read_1_1_MPORT_addr = io_raddr_0[0];
  assign dataBanks_1_perm_pf_data_read_1_1_MPORT_data =
    dataBanks_1_perm_pf[dataBanks_1_perm_pf_data_read_1_1_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_1_perm_pf_data_read_0_1_MPORT_1_en = 1'h1;
  assign dataBanks_1_perm_pf_data_read_0_1_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_1_perm_pf_data_read_0_1_MPORT_1_data =
    dataBanks_1_perm_pf[dataBanks_1_perm_pf_data_read_0_1_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_1_perm_pf_data_read_1_1_MPORT_1_en = 1'h1;
  assign dataBanks_1_perm_pf_data_read_1_1_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_1_perm_pf_data_read_1_1_MPORT_1_data =
    dataBanks_1_perm_pf[dataBanks_1_perm_pf_data_read_1_1_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_1_perm_pf_MPORT_1_data = io_wdata_perm_pf;
  assign dataBanks_1_perm_pf_MPORT_1_addr = io_waddr[0];
  assign dataBanks_1_perm_pf_MPORT_1_mask = 1'h1;
  assign dataBanks_1_perm_pf_MPORT_1_en = io_wen & _T_5;
  assign dataBanks_1_perm_af_data_read_0_1_MPORT_en = 1'h1;
  assign dataBanks_1_perm_af_data_read_0_1_MPORT_addr = io_raddr_0[0];
  assign dataBanks_1_perm_af_data_read_0_1_MPORT_data =
    dataBanks_1_perm_af[dataBanks_1_perm_af_data_read_0_1_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_1_perm_af_data_read_1_1_MPORT_en = 1'h1;
  assign dataBanks_1_perm_af_data_read_1_1_MPORT_addr = io_raddr_0[0];
  assign dataBanks_1_perm_af_data_read_1_1_MPORT_data =
    dataBanks_1_perm_af[dataBanks_1_perm_af_data_read_1_1_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_1_perm_af_data_read_0_1_MPORT_1_en = 1'h1;
  assign dataBanks_1_perm_af_data_read_0_1_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_1_perm_af_data_read_0_1_MPORT_1_data =
    dataBanks_1_perm_af[dataBanks_1_perm_af_data_read_0_1_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_1_perm_af_data_read_1_1_MPORT_1_en = 1'h1;
  assign dataBanks_1_perm_af_data_read_1_1_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_1_perm_af_data_read_1_1_MPORT_1_data =
    dataBanks_1_perm_af[dataBanks_1_perm_af_data_read_1_1_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_1_perm_af_MPORT_1_data = io_wdata_perm_af;
  assign dataBanks_1_perm_af_MPORT_1_addr = io_waddr[0];
  assign dataBanks_1_perm_af_MPORT_1_mask = 1'h1;
  assign dataBanks_1_perm_af_MPORT_1_en = io_wen & _T_5;
  assign dataBanks_1_perm_d_data_read_0_1_MPORT_en = 1'h1;
  assign dataBanks_1_perm_d_data_read_0_1_MPORT_addr = io_raddr_0[0];
  assign dataBanks_1_perm_d_data_read_0_1_MPORT_data = dataBanks_1_perm_d[dataBanks_1_perm_d_data_read_0_1_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_1_perm_d_data_read_1_1_MPORT_en = 1'h1;
  assign dataBanks_1_perm_d_data_read_1_1_MPORT_addr = io_raddr_0[0];
  assign dataBanks_1_perm_d_data_read_1_1_MPORT_data = dataBanks_1_perm_d[dataBanks_1_perm_d_data_read_1_1_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_1_perm_d_data_read_0_1_MPORT_1_en = 1'h1;
  assign dataBanks_1_perm_d_data_read_0_1_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_1_perm_d_data_read_0_1_MPORT_1_data =
    dataBanks_1_perm_d[dataBanks_1_perm_d_data_read_0_1_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_1_perm_d_data_read_1_1_MPORT_1_en = 1'h1;
  assign dataBanks_1_perm_d_data_read_1_1_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_1_perm_d_data_read_1_1_MPORT_1_data =
    dataBanks_1_perm_d[dataBanks_1_perm_d_data_read_1_1_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_1_perm_d_MPORT_1_data = io_wdata_perm_d;
  assign dataBanks_1_perm_d_MPORT_1_addr = io_waddr[0];
  assign dataBanks_1_perm_d_MPORT_1_mask = 1'h1;
  assign dataBanks_1_perm_d_MPORT_1_en = io_wen & _T_5;
  assign dataBanks_1_perm_a_data_read_0_1_MPORT_en = 1'h1;
  assign dataBanks_1_perm_a_data_read_0_1_MPORT_addr = io_raddr_0[0];
  assign dataBanks_1_perm_a_data_read_0_1_MPORT_data = dataBanks_1_perm_a[dataBanks_1_perm_a_data_read_0_1_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_1_perm_a_data_read_1_1_MPORT_en = 1'h1;
  assign dataBanks_1_perm_a_data_read_1_1_MPORT_addr = io_raddr_0[0];
  assign dataBanks_1_perm_a_data_read_1_1_MPORT_data = dataBanks_1_perm_a[dataBanks_1_perm_a_data_read_1_1_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_1_perm_a_data_read_0_1_MPORT_1_en = 1'h1;
  assign dataBanks_1_perm_a_data_read_0_1_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_1_perm_a_data_read_0_1_MPORT_1_data =
    dataBanks_1_perm_a[dataBanks_1_perm_a_data_read_0_1_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_1_perm_a_data_read_1_1_MPORT_1_en = 1'h1;
  assign dataBanks_1_perm_a_data_read_1_1_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_1_perm_a_data_read_1_1_MPORT_1_data =
    dataBanks_1_perm_a[dataBanks_1_perm_a_data_read_1_1_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_1_perm_a_MPORT_1_data = io_wdata_perm_a;
  assign dataBanks_1_perm_a_MPORT_1_addr = io_waddr[0];
  assign dataBanks_1_perm_a_MPORT_1_mask = 1'h1;
  assign dataBanks_1_perm_a_MPORT_1_en = io_wen & _T_5;
  assign dataBanks_1_perm_u_data_read_0_1_MPORT_en = 1'h1;
  assign dataBanks_1_perm_u_data_read_0_1_MPORT_addr = io_raddr_0[0];
  assign dataBanks_1_perm_u_data_read_0_1_MPORT_data = dataBanks_1_perm_u[dataBanks_1_perm_u_data_read_0_1_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_1_perm_u_data_read_1_1_MPORT_en = 1'h1;
  assign dataBanks_1_perm_u_data_read_1_1_MPORT_addr = io_raddr_0[0];
  assign dataBanks_1_perm_u_data_read_1_1_MPORT_data = dataBanks_1_perm_u[dataBanks_1_perm_u_data_read_1_1_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_1_perm_u_data_read_0_1_MPORT_1_en = 1'h1;
  assign dataBanks_1_perm_u_data_read_0_1_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_1_perm_u_data_read_0_1_MPORT_1_data =
    dataBanks_1_perm_u[dataBanks_1_perm_u_data_read_0_1_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_1_perm_u_data_read_1_1_MPORT_1_en = 1'h1;
  assign dataBanks_1_perm_u_data_read_1_1_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_1_perm_u_data_read_1_1_MPORT_1_data =
    dataBanks_1_perm_u[dataBanks_1_perm_u_data_read_1_1_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_1_perm_u_MPORT_1_data = io_wdata_perm_u;
  assign dataBanks_1_perm_u_MPORT_1_addr = io_waddr[0];
  assign dataBanks_1_perm_u_MPORT_1_mask = 1'h1;
  assign dataBanks_1_perm_u_MPORT_1_en = io_wen & _T_5;
  assign dataBanks_1_perm_x_data_read_0_1_MPORT_en = 1'h1;
  assign dataBanks_1_perm_x_data_read_0_1_MPORT_addr = io_raddr_0[0];
  assign dataBanks_1_perm_x_data_read_0_1_MPORT_data = dataBanks_1_perm_x[dataBanks_1_perm_x_data_read_0_1_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_1_perm_x_data_read_1_1_MPORT_en = 1'h1;
  assign dataBanks_1_perm_x_data_read_1_1_MPORT_addr = io_raddr_0[0];
  assign dataBanks_1_perm_x_data_read_1_1_MPORT_data = dataBanks_1_perm_x[dataBanks_1_perm_x_data_read_1_1_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_1_perm_x_data_read_0_1_MPORT_1_en = 1'h1;
  assign dataBanks_1_perm_x_data_read_0_1_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_1_perm_x_data_read_0_1_MPORT_1_data =
    dataBanks_1_perm_x[dataBanks_1_perm_x_data_read_0_1_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_1_perm_x_data_read_1_1_MPORT_1_en = 1'h1;
  assign dataBanks_1_perm_x_data_read_1_1_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_1_perm_x_data_read_1_1_MPORT_1_data =
    dataBanks_1_perm_x[dataBanks_1_perm_x_data_read_1_1_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_1_perm_x_MPORT_1_data = io_wdata_perm_x;
  assign dataBanks_1_perm_x_MPORT_1_addr = io_waddr[0];
  assign dataBanks_1_perm_x_MPORT_1_mask = 1'h1;
  assign dataBanks_1_perm_x_MPORT_1_en = io_wen & _T_5;
  assign dataBanks_1_perm_wdata_read_0_1_MPORT_en = 1'h1;
  assign dataBanks_1_perm_wdata_read_0_1_MPORT_addr = io_raddr_0[0];
  assign dataBanks_1_perm_wdata_read_0_1_MPORT_data = dataBanks_1_perm_w[dataBanks_1_perm_wdata_read_0_1_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_1_perm_wdata_read_1_1_MPORT_en = 1'h1;
  assign dataBanks_1_perm_wdata_read_1_1_MPORT_addr = io_raddr_0[0];
  assign dataBanks_1_perm_wdata_read_1_1_MPORT_data = dataBanks_1_perm_w[dataBanks_1_perm_wdata_read_1_1_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_1_perm_wdata_read_0_1_MPORT_1_en = 1'h1;
  assign dataBanks_1_perm_wdata_read_0_1_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_1_perm_wdata_read_0_1_MPORT_1_data =
    dataBanks_1_perm_w[dataBanks_1_perm_wdata_read_0_1_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_1_perm_wdata_read_1_1_MPORT_1_en = 1'h1;
  assign dataBanks_1_perm_wdata_read_1_1_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_1_perm_wdata_read_1_1_MPORT_1_data =
    dataBanks_1_perm_w[dataBanks_1_perm_wdata_read_1_1_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_1_perm_wMPORT_1_data = io_wdata_perm_w;
  assign dataBanks_1_perm_wMPORT_1_addr = io_waddr[0];
  assign dataBanks_1_perm_wMPORT_1_mask = 1'h1;
  assign dataBanks_1_perm_wMPORT_1_en = io_wen & _T_5;
  assign dataBanks_1_perm_rdata_read_0_1_MPORT_en = 1'h1;
  assign dataBanks_1_perm_rdata_read_0_1_MPORT_addr = io_raddr_0[0];
  assign dataBanks_1_perm_rdata_read_0_1_MPORT_data = dataBanks_1_perm_r[dataBanks_1_perm_rdata_read_0_1_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_1_perm_rdata_read_1_1_MPORT_en = 1'h1;
  assign dataBanks_1_perm_rdata_read_1_1_MPORT_addr = io_raddr_0[0];
  assign dataBanks_1_perm_rdata_read_1_1_MPORT_data = dataBanks_1_perm_r[dataBanks_1_perm_rdata_read_1_1_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_1_perm_rdata_read_0_1_MPORT_1_en = 1'h1;
  assign dataBanks_1_perm_rdata_read_0_1_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_1_perm_rdata_read_0_1_MPORT_1_data =
    dataBanks_1_perm_r[dataBanks_1_perm_rdata_read_0_1_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_1_perm_rdata_read_1_1_MPORT_1_en = 1'h1;
  assign dataBanks_1_perm_rdata_read_1_1_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_1_perm_rdata_read_1_1_MPORT_1_data =
    dataBanks_1_perm_r[dataBanks_1_perm_rdata_read_1_1_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_1_perm_rMPORT_1_data = io_wdata_perm_r;
  assign dataBanks_1_perm_rMPORT_1_addr = io_waddr[0];
  assign dataBanks_1_perm_rMPORT_1_mask = 1'h1;
  assign dataBanks_1_perm_rMPORT_1_en = io_wen & _T_5;
  assign dataBanks_1_perm_pm_rdata_read_0_1_MPORT_en = 1'h1;
  assign dataBanks_1_perm_pm_rdata_read_0_1_MPORT_addr = io_raddr_0[0];
  assign dataBanks_1_perm_pm_rdata_read_0_1_MPORT_data =
    dataBanks_1_perm_pm_r[dataBanks_1_perm_pm_rdata_read_0_1_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_1_perm_pm_rdata_read_1_1_MPORT_en = 1'h1;
  assign dataBanks_1_perm_pm_rdata_read_1_1_MPORT_addr = io_raddr_0[0];
  assign dataBanks_1_perm_pm_rdata_read_1_1_MPORT_data =
    dataBanks_1_perm_pm_r[dataBanks_1_perm_pm_rdata_read_1_1_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_1_perm_pm_rdata_read_0_1_MPORT_1_en = 1'h1;
  assign dataBanks_1_perm_pm_rdata_read_0_1_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_1_perm_pm_rdata_read_0_1_MPORT_1_data =
    dataBanks_1_perm_pm_r[dataBanks_1_perm_pm_rdata_read_0_1_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_1_perm_pm_rdata_read_1_1_MPORT_1_en = 1'h1;
  assign dataBanks_1_perm_pm_rdata_read_1_1_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_1_perm_pm_rdata_read_1_1_MPORT_1_data =
    dataBanks_1_perm_pm_r[dataBanks_1_perm_pm_rdata_read_1_1_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_1_perm_pm_rMPORT_1_data = io_wdata_perm_pm_r;
  assign dataBanks_1_perm_pm_rMPORT_1_addr = io_waddr[0];
  assign dataBanks_1_perm_pm_rMPORT_1_mask = 1'h1;
  assign dataBanks_1_perm_pm_rMPORT_1_en = io_wen & _T_5;
  assign dataBanks_1_perm_pm_wdata_read_0_1_MPORT_en = 1'h1;
  assign dataBanks_1_perm_pm_wdata_read_0_1_MPORT_addr = io_raddr_0[0];
  assign dataBanks_1_perm_pm_wdata_read_0_1_MPORT_data =
    dataBanks_1_perm_pm_w[dataBanks_1_perm_pm_wdata_read_0_1_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_1_perm_pm_wdata_read_1_1_MPORT_en = 1'h1;
  assign dataBanks_1_perm_pm_wdata_read_1_1_MPORT_addr = io_raddr_0[0];
  assign dataBanks_1_perm_pm_wdata_read_1_1_MPORT_data =
    dataBanks_1_perm_pm_w[dataBanks_1_perm_pm_wdata_read_1_1_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_1_perm_pm_wdata_read_0_1_MPORT_1_en = 1'h1;
  assign dataBanks_1_perm_pm_wdata_read_0_1_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_1_perm_pm_wdata_read_0_1_MPORT_1_data =
    dataBanks_1_perm_pm_w[dataBanks_1_perm_pm_wdata_read_0_1_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_1_perm_pm_wdata_read_1_1_MPORT_1_en = 1'h1;
  assign dataBanks_1_perm_pm_wdata_read_1_1_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_1_perm_pm_wdata_read_1_1_MPORT_1_data =
    dataBanks_1_perm_pm_w[dataBanks_1_perm_pm_wdata_read_1_1_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_1_perm_pm_wMPORT_1_data = io_wdata_perm_pm_w;
  assign dataBanks_1_perm_pm_wMPORT_1_addr = io_waddr[0];
  assign dataBanks_1_perm_pm_wMPORT_1_mask = 1'h1;
  assign dataBanks_1_perm_pm_wMPORT_1_en = io_wen & _T_5;
  assign dataBanks_1_perm_pm_c_data_read_0_1_MPORT_en = 1'h1;
  assign dataBanks_1_perm_pm_c_data_read_0_1_MPORT_addr = io_raddr_0[0];
  assign dataBanks_1_perm_pm_c_data_read_0_1_MPORT_data =
    dataBanks_1_perm_pm_c[dataBanks_1_perm_pm_c_data_read_0_1_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_1_perm_pm_c_data_read_1_1_MPORT_en = 1'h1;
  assign dataBanks_1_perm_pm_c_data_read_1_1_MPORT_addr = io_raddr_0[0];
  assign dataBanks_1_perm_pm_c_data_read_1_1_MPORT_data =
    dataBanks_1_perm_pm_c[dataBanks_1_perm_pm_c_data_read_1_1_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_1_perm_pm_c_data_read_0_1_MPORT_1_en = 1'h1;
  assign dataBanks_1_perm_pm_c_data_read_0_1_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_1_perm_pm_c_data_read_0_1_MPORT_1_data =
    dataBanks_1_perm_pm_c[dataBanks_1_perm_pm_c_data_read_0_1_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_1_perm_pm_c_data_read_1_1_MPORT_1_en = 1'h1;
  assign dataBanks_1_perm_pm_c_data_read_1_1_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_1_perm_pm_c_data_read_1_1_MPORT_1_data =
    dataBanks_1_perm_pm_c[dataBanks_1_perm_pm_c_data_read_1_1_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_1_perm_pm_c_MPORT_1_data = io_wdata_perm_pm_c;
  assign dataBanks_1_perm_pm_c_MPORT_1_addr = io_waddr[0];
  assign dataBanks_1_perm_pm_c_MPORT_1_mask = 1'h1;
  assign dataBanks_1_perm_pm_c_MPORT_1_en = io_wen & _T_5;
  assign dataBanks_2_tag_data_read_0_2_MPORT_en = 1'h1;
  assign dataBanks_2_tag_data_read_0_2_MPORT_addr = io_raddr_0[0];
  assign dataBanks_2_tag_data_read_0_2_MPORT_data = dataBanks_2_tag[dataBanks_2_tag_data_read_0_2_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_2_tag_data_read_1_2_MPORT_en = 1'h1;
  assign dataBanks_2_tag_data_read_1_2_MPORT_addr = io_raddr_0[0];
  assign dataBanks_2_tag_data_read_1_2_MPORT_data = dataBanks_2_tag[dataBanks_2_tag_data_read_1_2_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_2_tag_data_read_0_2_MPORT_1_en = 1'h1;
  assign dataBanks_2_tag_data_read_0_2_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_2_tag_data_read_0_2_MPORT_1_data = dataBanks_2_tag[dataBanks_2_tag_data_read_0_2_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_2_tag_data_read_1_2_MPORT_1_en = 1'h1;
  assign dataBanks_2_tag_data_read_1_2_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_2_tag_data_read_1_2_MPORT_1_data = dataBanks_2_tag[dataBanks_2_tag_data_read_1_2_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_2_tag_MPORT_2_data = io_wdata_tag;
  assign dataBanks_2_tag_MPORT_2_addr = io_waddr[0];
  assign dataBanks_2_tag_MPORT_2_mask = 1'h1;
  assign dataBanks_2_tag_MPORT_2_en = io_wen & _T_9;
  assign dataBanks_2_asid_data_read_0_2_MPORT_en = 1'h1;
  assign dataBanks_2_asid_data_read_0_2_MPORT_addr = io_raddr_0[0];
  assign dataBanks_2_asid_data_read_0_2_MPORT_data = dataBanks_2_asid[dataBanks_2_asid_data_read_0_2_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_2_asid_data_read_1_2_MPORT_en = 1'h1;
  assign dataBanks_2_asid_data_read_1_2_MPORT_addr = io_raddr_0[0];
  assign dataBanks_2_asid_data_read_1_2_MPORT_data = dataBanks_2_asid[dataBanks_2_asid_data_read_1_2_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_2_asid_data_read_0_2_MPORT_1_en = 1'h1;
  assign dataBanks_2_asid_data_read_0_2_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_2_asid_data_read_0_2_MPORT_1_data = dataBanks_2_asid[dataBanks_2_asid_data_read_0_2_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_2_asid_data_read_1_2_MPORT_1_en = 1'h1;
  assign dataBanks_2_asid_data_read_1_2_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_2_asid_data_read_1_2_MPORT_1_data = dataBanks_2_asid[dataBanks_2_asid_data_read_1_2_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_2_asid_MPORT_2_data = io_wdata_asid;
  assign dataBanks_2_asid_MPORT_2_addr = io_waddr[0];
  assign dataBanks_2_asid_MPORT_2_mask = 1'h1;
  assign dataBanks_2_asid_MPORT_2_en = io_wen & _T_9;
  assign dataBanks_2_ppn_data_read_0_2_MPORT_en = 1'h1;
  assign dataBanks_2_ppn_data_read_0_2_MPORT_addr = io_raddr_0[0];
  assign dataBanks_2_ppn_data_read_0_2_MPORT_data = dataBanks_2_ppn[dataBanks_2_ppn_data_read_0_2_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_2_ppn_data_read_1_2_MPORT_en = 1'h1;
  assign dataBanks_2_ppn_data_read_1_2_MPORT_addr = io_raddr_0[0];
  assign dataBanks_2_ppn_data_read_1_2_MPORT_data = dataBanks_2_ppn[dataBanks_2_ppn_data_read_1_2_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_2_ppn_data_read_0_2_MPORT_1_en = 1'h1;
  assign dataBanks_2_ppn_data_read_0_2_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_2_ppn_data_read_0_2_MPORT_1_data = dataBanks_2_ppn[dataBanks_2_ppn_data_read_0_2_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_2_ppn_data_read_1_2_MPORT_1_en = 1'h1;
  assign dataBanks_2_ppn_data_read_1_2_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_2_ppn_data_read_1_2_MPORT_1_data = dataBanks_2_ppn[dataBanks_2_ppn_data_read_1_2_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_2_ppn_MPORT_2_data = io_wdata_ppn;
  assign dataBanks_2_ppn_MPORT_2_addr = io_waddr[0];
  assign dataBanks_2_ppn_MPORT_2_mask = 1'h1;
  assign dataBanks_2_ppn_MPORT_2_en = io_wen & _T_9;
  assign dataBanks_2_perm_pf_data_read_0_2_MPORT_en = 1'h1;
  assign dataBanks_2_perm_pf_data_read_0_2_MPORT_addr = io_raddr_0[0];
  assign dataBanks_2_perm_pf_data_read_0_2_MPORT_data =
    dataBanks_2_perm_pf[dataBanks_2_perm_pf_data_read_0_2_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_2_perm_pf_data_read_1_2_MPORT_en = 1'h1;
  assign dataBanks_2_perm_pf_data_read_1_2_MPORT_addr = io_raddr_0[0];
  assign dataBanks_2_perm_pf_data_read_1_2_MPORT_data =
    dataBanks_2_perm_pf[dataBanks_2_perm_pf_data_read_1_2_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_2_perm_pf_data_read_0_2_MPORT_1_en = 1'h1;
  assign dataBanks_2_perm_pf_data_read_0_2_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_2_perm_pf_data_read_0_2_MPORT_1_data =
    dataBanks_2_perm_pf[dataBanks_2_perm_pf_data_read_0_2_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_2_perm_pf_data_read_1_2_MPORT_1_en = 1'h1;
  assign dataBanks_2_perm_pf_data_read_1_2_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_2_perm_pf_data_read_1_2_MPORT_1_data =
    dataBanks_2_perm_pf[dataBanks_2_perm_pf_data_read_1_2_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_2_perm_pf_MPORT_2_data = io_wdata_perm_pf;
  assign dataBanks_2_perm_pf_MPORT_2_addr = io_waddr[0];
  assign dataBanks_2_perm_pf_MPORT_2_mask = 1'h1;
  assign dataBanks_2_perm_pf_MPORT_2_en = io_wen & _T_9;
  assign dataBanks_2_perm_af_data_read_0_2_MPORT_en = 1'h1;
  assign dataBanks_2_perm_af_data_read_0_2_MPORT_addr = io_raddr_0[0];
  assign dataBanks_2_perm_af_data_read_0_2_MPORT_data =
    dataBanks_2_perm_af[dataBanks_2_perm_af_data_read_0_2_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_2_perm_af_data_read_1_2_MPORT_en = 1'h1;
  assign dataBanks_2_perm_af_data_read_1_2_MPORT_addr = io_raddr_0[0];
  assign dataBanks_2_perm_af_data_read_1_2_MPORT_data =
    dataBanks_2_perm_af[dataBanks_2_perm_af_data_read_1_2_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_2_perm_af_data_read_0_2_MPORT_1_en = 1'h1;
  assign dataBanks_2_perm_af_data_read_0_2_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_2_perm_af_data_read_0_2_MPORT_1_data =
    dataBanks_2_perm_af[dataBanks_2_perm_af_data_read_0_2_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_2_perm_af_data_read_1_2_MPORT_1_en = 1'h1;
  assign dataBanks_2_perm_af_data_read_1_2_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_2_perm_af_data_read_1_2_MPORT_1_data =
    dataBanks_2_perm_af[dataBanks_2_perm_af_data_read_1_2_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_2_perm_af_MPORT_2_data = io_wdata_perm_af;
  assign dataBanks_2_perm_af_MPORT_2_addr = io_waddr[0];
  assign dataBanks_2_perm_af_MPORT_2_mask = 1'h1;
  assign dataBanks_2_perm_af_MPORT_2_en = io_wen & _T_9;
  assign dataBanks_2_perm_d_data_read_0_2_MPORT_en = 1'h1;
  assign dataBanks_2_perm_d_data_read_0_2_MPORT_addr = io_raddr_0[0];
  assign dataBanks_2_perm_d_data_read_0_2_MPORT_data = dataBanks_2_perm_d[dataBanks_2_perm_d_data_read_0_2_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_2_perm_d_data_read_1_2_MPORT_en = 1'h1;
  assign dataBanks_2_perm_d_data_read_1_2_MPORT_addr = io_raddr_0[0];
  assign dataBanks_2_perm_d_data_read_1_2_MPORT_data = dataBanks_2_perm_d[dataBanks_2_perm_d_data_read_1_2_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_2_perm_d_data_read_0_2_MPORT_1_en = 1'h1;
  assign dataBanks_2_perm_d_data_read_0_2_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_2_perm_d_data_read_0_2_MPORT_1_data =
    dataBanks_2_perm_d[dataBanks_2_perm_d_data_read_0_2_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_2_perm_d_data_read_1_2_MPORT_1_en = 1'h1;
  assign dataBanks_2_perm_d_data_read_1_2_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_2_perm_d_data_read_1_2_MPORT_1_data =
    dataBanks_2_perm_d[dataBanks_2_perm_d_data_read_1_2_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_2_perm_d_MPORT_2_data = io_wdata_perm_d;
  assign dataBanks_2_perm_d_MPORT_2_addr = io_waddr[0];
  assign dataBanks_2_perm_d_MPORT_2_mask = 1'h1;
  assign dataBanks_2_perm_d_MPORT_2_en = io_wen & _T_9;
  assign dataBanks_2_perm_a_data_read_0_2_MPORT_en = 1'h1;
  assign dataBanks_2_perm_a_data_read_0_2_MPORT_addr = io_raddr_0[0];
  assign dataBanks_2_perm_a_data_read_0_2_MPORT_data = dataBanks_2_perm_a[dataBanks_2_perm_a_data_read_0_2_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_2_perm_a_data_read_1_2_MPORT_en = 1'h1;
  assign dataBanks_2_perm_a_data_read_1_2_MPORT_addr = io_raddr_0[0];
  assign dataBanks_2_perm_a_data_read_1_2_MPORT_data = dataBanks_2_perm_a[dataBanks_2_perm_a_data_read_1_2_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_2_perm_a_data_read_0_2_MPORT_1_en = 1'h1;
  assign dataBanks_2_perm_a_data_read_0_2_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_2_perm_a_data_read_0_2_MPORT_1_data =
    dataBanks_2_perm_a[dataBanks_2_perm_a_data_read_0_2_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_2_perm_a_data_read_1_2_MPORT_1_en = 1'h1;
  assign dataBanks_2_perm_a_data_read_1_2_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_2_perm_a_data_read_1_2_MPORT_1_data =
    dataBanks_2_perm_a[dataBanks_2_perm_a_data_read_1_2_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_2_perm_a_MPORT_2_data = io_wdata_perm_a;
  assign dataBanks_2_perm_a_MPORT_2_addr = io_waddr[0];
  assign dataBanks_2_perm_a_MPORT_2_mask = 1'h1;
  assign dataBanks_2_perm_a_MPORT_2_en = io_wen & _T_9;
  assign dataBanks_2_perm_u_data_read_0_2_MPORT_en = 1'h1;
  assign dataBanks_2_perm_u_data_read_0_2_MPORT_addr = io_raddr_0[0];
  assign dataBanks_2_perm_u_data_read_0_2_MPORT_data = dataBanks_2_perm_u[dataBanks_2_perm_u_data_read_0_2_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_2_perm_u_data_read_1_2_MPORT_en = 1'h1;
  assign dataBanks_2_perm_u_data_read_1_2_MPORT_addr = io_raddr_0[0];
  assign dataBanks_2_perm_u_data_read_1_2_MPORT_data = dataBanks_2_perm_u[dataBanks_2_perm_u_data_read_1_2_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_2_perm_u_data_read_0_2_MPORT_1_en = 1'h1;
  assign dataBanks_2_perm_u_data_read_0_2_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_2_perm_u_data_read_0_2_MPORT_1_data =
    dataBanks_2_perm_u[dataBanks_2_perm_u_data_read_0_2_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_2_perm_u_data_read_1_2_MPORT_1_en = 1'h1;
  assign dataBanks_2_perm_u_data_read_1_2_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_2_perm_u_data_read_1_2_MPORT_1_data =
    dataBanks_2_perm_u[dataBanks_2_perm_u_data_read_1_2_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_2_perm_u_MPORT_2_data = io_wdata_perm_u;
  assign dataBanks_2_perm_u_MPORT_2_addr = io_waddr[0];
  assign dataBanks_2_perm_u_MPORT_2_mask = 1'h1;
  assign dataBanks_2_perm_u_MPORT_2_en = io_wen & _T_9;
  assign dataBanks_2_perm_x_data_read_0_2_MPORT_en = 1'h1;
  assign dataBanks_2_perm_x_data_read_0_2_MPORT_addr = io_raddr_0[0];
  assign dataBanks_2_perm_x_data_read_0_2_MPORT_data = dataBanks_2_perm_x[dataBanks_2_perm_x_data_read_0_2_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_2_perm_x_data_read_1_2_MPORT_en = 1'h1;
  assign dataBanks_2_perm_x_data_read_1_2_MPORT_addr = io_raddr_0[0];
  assign dataBanks_2_perm_x_data_read_1_2_MPORT_data = dataBanks_2_perm_x[dataBanks_2_perm_x_data_read_1_2_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_2_perm_x_data_read_0_2_MPORT_1_en = 1'h1;
  assign dataBanks_2_perm_x_data_read_0_2_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_2_perm_x_data_read_0_2_MPORT_1_data =
    dataBanks_2_perm_x[dataBanks_2_perm_x_data_read_0_2_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_2_perm_x_data_read_1_2_MPORT_1_en = 1'h1;
  assign dataBanks_2_perm_x_data_read_1_2_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_2_perm_x_data_read_1_2_MPORT_1_data =
    dataBanks_2_perm_x[dataBanks_2_perm_x_data_read_1_2_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_2_perm_x_MPORT_2_data = io_wdata_perm_x;
  assign dataBanks_2_perm_x_MPORT_2_addr = io_waddr[0];
  assign dataBanks_2_perm_x_MPORT_2_mask = 1'h1;
  assign dataBanks_2_perm_x_MPORT_2_en = io_wen & _T_9;
  assign dataBanks_2_perm_wdata_read_0_2_MPORT_en = 1'h1;
  assign dataBanks_2_perm_wdata_read_0_2_MPORT_addr = io_raddr_0[0];
  assign dataBanks_2_perm_wdata_read_0_2_MPORT_data = dataBanks_2_perm_w[dataBanks_2_perm_wdata_read_0_2_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_2_perm_wdata_read_1_2_MPORT_en = 1'h1;
  assign dataBanks_2_perm_wdata_read_1_2_MPORT_addr = io_raddr_0[0];
  assign dataBanks_2_perm_wdata_read_1_2_MPORT_data = dataBanks_2_perm_w[dataBanks_2_perm_wdata_read_1_2_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_2_perm_wdata_read_0_2_MPORT_1_en = 1'h1;
  assign dataBanks_2_perm_wdata_read_0_2_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_2_perm_wdata_read_0_2_MPORT_1_data =
    dataBanks_2_perm_w[dataBanks_2_perm_wdata_read_0_2_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_2_perm_wdata_read_1_2_MPORT_1_en = 1'h1;
  assign dataBanks_2_perm_wdata_read_1_2_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_2_perm_wdata_read_1_2_MPORT_1_data =
    dataBanks_2_perm_w[dataBanks_2_perm_wdata_read_1_2_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_2_perm_wMPORT_2_data = io_wdata_perm_w;
  assign dataBanks_2_perm_wMPORT_2_addr = io_waddr[0];
  assign dataBanks_2_perm_wMPORT_2_mask = 1'h1;
  assign dataBanks_2_perm_wMPORT_2_en = io_wen & _T_9;
  assign dataBanks_2_perm_rdata_read_0_2_MPORT_en = 1'h1;
  assign dataBanks_2_perm_rdata_read_0_2_MPORT_addr = io_raddr_0[0];
  assign dataBanks_2_perm_rdata_read_0_2_MPORT_data = dataBanks_2_perm_r[dataBanks_2_perm_rdata_read_0_2_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_2_perm_rdata_read_1_2_MPORT_en = 1'h1;
  assign dataBanks_2_perm_rdata_read_1_2_MPORT_addr = io_raddr_0[0];
  assign dataBanks_2_perm_rdata_read_1_2_MPORT_data = dataBanks_2_perm_r[dataBanks_2_perm_rdata_read_1_2_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_2_perm_rdata_read_0_2_MPORT_1_en = 1'h1;
  assign dataBanks_2_perm_rdata_read_0_2_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_2_perm_rdata_read_0_2_MPORT_1_data =
    dataBanks_2_perm_r[dataBanks_2_perm_rdata_read_0_2_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_2_perm_rdata_read_1_2_MPORT_1_en = 1'h1;
  assign dataBanks_2_perm_rdata_read_1_2_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_2_perm_rdata_read_1_2_MPORT_1_data =
    dataBanks_2_perm_r[dataBanks_2_perm_rdata_read_1_2_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_2_perm_rMPORT_2_data = io_wdata_perm_r;
  assign dataBanks_2_perm_rMPORT_2_addr = io_waddr[0];
  assign dataBanks_2_perm_rMPORT_2_mask = 1'h1;
  assign dataBanks_2_perm_rMPORT_2_en = io_wen & _T_9;
  assign dataBanks_2_perm_pm_rdata_read_0_2_MPORT_en = 1'h1;
  assign dataBanks_2_perm_pm_rdata_read_0_2_MPORT_addr = io_raddr_0[0];
  assign dataBanks_2_perm_pm_rdata_read_0_2_MPORT_data =
    dataBanks_2_perm_pm_r[dataBanks_2_perm_pm_rdata_read_0_2_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_2_perm_pm_rdata_read_1_2_MPORT_en = 1'h1;
  assign dataBanks_2_perm_pm_rdata_read_1_2_MPORT_addr = io_raddr_0[0];
  assign dataBanks_2_perm_pm_rdata_read_1_2_MPORT_data =
    dataBanks_2_perm_pm_r[dataBanks_2_perm_pm_rdata_read_1_2_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_2_perm_pm_rdata_read_0_2_MPORT_1_en = 1'h1;
  assign dataBanks_2_perm_pm_rdata_read_0_2_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_2_perm_pm_rdata_read_0_2_MPORT_1_data =
    dataBanks_2_perm_pm_r[dataBanks_2_perm_pm_rdata_read_0_2_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_2_perm_pm_rdata_read_1_2_MPORT_1_en = 1'h1;
  assign dataBanks_2_perm_pm_rdata_read_1_2_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_2_perm_pm_rdata_read_1_2_MPORT_1_data =
    dataBanks_2_perm_pm_r[dataBanks_2_perm_pm_rdata_read_1_2_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_2_perm_pm_rMPORT_2_data = io_wdata_perm_pm_r;
  assign dataBanks_2_perm_pm_rMPORT_2_addr = io_waddr[0];
  assign dataBanks_2_perm_pm_rMPORT_2_mask = 1'h1;
  assign dataBanks_2_perm_pm_rMPORT_2_en = io_wen & _T_9;
  assign dataBanks_2_perm_pm_wdata_read_0_2_MPORT_en = 1'h1;
  assign dataBanks_2_perm_pm_wdata_read_0_2_MPORT_addr = io_raddr_0[0];
  assign dataBanks_2_perm_pm_wdata_read_0_2_MPORT_data =
    dataBanks_2_perm_pm_w[dataBanks_2_perm_pm_wdata_read_0_2_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_2_perm_pm_wdata_read_1_2_MPORT_en = 1'h1;
  assign dataBanks_2_perm_pm_wdata_read_1_2_MPORT_addr = io_raddr_0[0];
  assign dataBanks_2_perm_pm_wdata_read_1_2_MPORT_data =
    dataBanks_2_perm_pm_w[dataBanks_2_perm_pm_wdata_read_1_2_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_2_perm_pm_wdata_read_0_2_MPORT_1_en = 1'h1;
  assign dataBanks_2_perm_pm_wdata_read_0_2_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_2_perm_pm_wdata_read_0_2_MPORT_1_data =
    dataBanks_2_perm_pm_w[dataBanks_2_perm_pm_wdata_read_0_2_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_2_perm_pm_wdata_read_1_2_MPORT_1_en = 1'h1;
  assign dataBanks_2_perm_pm_wdata_read_1_2_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_2_perm_pm_wdata_read_1_2_MPORT_1_data =
    dataBanks_2_perm_pm_w[dataBanks_2_perm_pm_wdata_read_1_2_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_2_perm_pm_wMPORT_2_data = io_wdata_perm_pm_w;
  assign dataBanks_2_perm_pm_wMPORT_2_addr = io_waddr[0];
  assign dataBanks_2_perm_pm_wMPORT_2_mask = 1'h1;
  assign dataBanks_2_perm_pm_wMPORT_2_en = io_wen & _T_9;
  assign dataBanks_2_perm_pm_c_data_read_0_2_MPORT_en = 1'h1;
  assign dataBanks_2_perm_pm_c_data_read_0_2_MPORT_addr = io_raddr_0[0];
  assign dataBanks_2_perm_pm_c_data_read_0_2_MPORT_data =
    dataBanks_2_perm_pm_c[dataBanks_2_perm_pm_c_data_read_0_2_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_2_perm_pm_c_data_read_1_2_MPORT_en = 1'h1;
  assign dataBanks_2_perm_pm_c_data_read_1_2_MPORT_addr = io_raddr_0[0];
  assign dataBanks_2_perm_pm_c_data_read_1_2_MPORT_data =
    dataBanks_2_perm_pm_c[dataBanks_2_perm_pm_c_data_read_1_2_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_2_perm_pm_c_data_read_0_2_MPORT_1_en = 1'h1;
  assign dataBanks_2_perm_pm_c_data_read_0_2_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_2_perm_pm_c_data_read_0_2_MPORT_1_data =
    dataBanks_2_perm_pm_c[dataBanks_2_perm_pm_c_data_read_0_2_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_2_perm_pm_c_data_read_1_2_MPORT_1_en = 1'h1;
  assign dataBanks_2_perm_pm_c_data_read_1_2_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_2_perm_pm_c_data_read_1_2_MPORT_1_data =
    dataBanks_2_perm_pm_c[dataBanks_2_perm_pm_c_data_read_1_2_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_2_perm_pm_c_MPORT_2_data = io_wdata_perm_pm_c;
  assign dataBanks_2_perm_pm_c_MPORT_2_addr = io_waddr[0];
  assign dataBanks_2_perm_pm_c_MPORT_2_mask = 1'h1;
  assign dataBanks_2_perm_pm_c_MPORT_2_en = io_wen & _T_9;
  assign dataBanks_3_tag_data_read_0_3_MPORT_en = 1'h1;
  assign dataBanks_3_tag_data_read_0_3_MPORT_addr = io_raddr_0[0];
  assign dataBanks_3_tag_data_read_0_3_MPORT_data = dataBanks_3_tag[dataBanks_3_tag_data_read_0_3_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_3_tag_data_read_1_3_MPORT_en = 1'h1;
  assign dataBanks_3_tag_data_read_1_3_MPORT_addr = io_raddr_0[0];
  assign dataBanks_3_tag_data_read_1_3_MPORT_data = dataBanks_3_tag[dataBanks_3_tag_data_read_1_3_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_3_tag_data_read_0_3_MPORT_1_en = 1'h1;
  assign dataBanks_3_tag_data_read_0_3_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_3_tag_data_read_0_3_MPORT_1_data = dataBanks_3_tag[dataBanks_3_tag_data_read_0_3_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_3_tag_data_read_1_3_MPORT_1_en = 1'h1;
  assign dataBanks_3_tag_data_read_1_3_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_3_tag_data_read_1_3_MPORT_1_data = dataBanks_3_tag[dataBanks_3_tag_data_read_1_3_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_3_tag_MPORT_3_data = io_wdata_tag;
  assign dataBanks_3_tag_MPORT_3_addr = io_waddr[0];
  assign dataBanks_3_tag_MPORT_3_mask = 1'h1;
  assign dataBanks_3_tag_MPORT_3_en = io_wen & _T_13;
  assign dataBanks_3_asid_data_read_0_3_MPORT_en = 1'h1;
  assign dataBanks_3_asid_data_read_0_3_MPORT_addr = io_raddr_0[0];
  assign dataBanks_3_asid_data_read_0_3_MPORT_data = dataBanks_3_asid[dataBanks_3_asid_data_read_0_3_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_3_asid_data_read_1_3_MPORT_en = 1'h1;
  assign dataBanks_3_asid_data_read_1_3_MPORT_addr = io_raddr_0[0];
  assign dataBanks_3_asid_data_read_1_3_MPORT_data = dataBanks_3_asid[dataBanks_3_asid_data_read_1_3_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_3_asid_data_read_0_3_MPORT_1_en = 1'h1;
  assign dataBanks_3_asid_data_read_0_3_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_3_asid_data_read_0_3_MPORT_1_data = dataBanks_3_asid[dataBanks_3_asid_data_read_0_3_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_3_asid_data_read_1_3_MPORT_1_en = 1'h1;
  assign dataBanks_3_asid_data_read_1_3_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_3_asid_data_read_1_3_MPORT_1_data = dataBanks_3_asid[dataBanks_3_asid_data_read_1_3_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_3_asid_MPORT_3_data = io_wdata_asid;
  assign dataBanks_3_asid_MPORT_3_addr = io_waddr[0];
  assign dataBanks_3_asid_MPORT_3_mask = 1'h1;
  assign dataBanks_3_asid_MPORT_3_en = io_wen & _T_13;
  assign dataBanks_3_ppn_data_read_0_3_MPORT_en = 1'h1;
  assign dataBanks_3_ppn_data_read_0_3_MPORT_addr = io_raddr_0[0];
  assign dataBanks_3_ppn_data_read_0_3_MPORT_data = dataBanks_3_ppn[dataBanks_3_ppn_data_read_0_3_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_3_ppn_data_read_1_3_MPORT_en = 1'h1;
  assign dataBanks_3_ppn_data_read_1_3_MPORT_addr = io_raddr_0[0];
  assign dataBanks_3_ppn_data_read_1_3_MPORT_data = dataBanks_3_ppn[dataBanks_3_ppn_data_read_1_3_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_3_ppn_data_read_0_3_MPORT_1_en = 1'h1;
  assign dataBanks_3_ppn_data_read_0_3_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_3_ppn_data_read_0_3_MPORT_1_data = dataBanks_3_ppn[dataBanks_3_ppn_data_read_0_3_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_3_ppn_data_read_1_3_MPORT_1_en = 1'h1;
  assign dataBanks_3_ppn_data_read_1_3_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_3_ppn_data_read_1_3_MPORT_1_data = dataBanks_3_ppn[dataBanks_3_ppn_data_read_1_3_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_3_ppn_MPORT_3_data = io_wdata_ppn;
  assign dataBanks_3_ppn_MPORT_3_addr = io_waddr[0];
  assign dataBanks_3_ppn_MPORT_3_mask = 1'h1;
  assign dataBanks_3_ppn_MPORT_3_en = io_wen & _T_13;
  assign dataBanks_3_perm_pf_data_read_0_3_MPORT_en = 1'h1;
  assign dataBanks_3_perm_pf_data_read_0_3_MPORT_addr = io_raddr_0[0];
  assign dataBanks_3_perm_pf_data_read_0_3_MPORT_data =
    dataBanks_3_perm_pf[dataBanks_3_perm_pf_data_read_0_3_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_3_perm_pf_data_read_1_3_MPORT_en = 1'h1;
  assign dataBanks_3_perm_pf_data_read_1_3_MPORT_addr = io_raddr_0[0];
  assign dataBanks_3_perm_pf_data_read_1_3_MPORT_data =
    dataBanks_3_perm_pf[dataBanks_3_perm_pf_data_read_1_3_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_3_perm_pf_data_read_0_3_MPORT_1_en = 1'h1;
  assign dataBanks_3_perm_pf_data_read_0_3_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_3_perm_pf_data_read_0_3_MPORT_1_data =
    dataBanks_3_perm_pf[dataBanks_3_perm_pf_data_read_0_3_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_3_perm_pf_data_read_1_3_MPORT_1_en = 1'h1;
  assign dataBanks_3_perm_pf_data_read_1_3_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_3_perm_pf_data_read_1_3_MPORT_1_data =
    dataBanks_3_perm_pf[dataBanks_3_perm_pf_data_read_1_3_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_3_perm_pf_MPORT_3_data = io_wdata_perm_pf;
  assign dataBanks_3_perm_pf_MPORT_3_addr = io_waddr[0];
  assign dataBanks_3_perm_pf_MPORT_3_mask = 1'h1;
  assign dataBanks_3_perm_pf_MPORT_3_en = io_wen & _T_13;
  assign dataBanks_3_perm_af_data_read_0_3_MPORT_en = 1'h1;
  assign dataBanks_3_perm_af_data_read_0_3_MPORT_addr = io_raddr_0[0];
  assign dataBanks_3_perm_af_data_read_0_3_MPORT_data =
    dataBanks_3_perm_af[dataBanks_3_perm_af_data_read_0_3_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_3_perm_af_data_read_1_3_MPORT_en = 1'h1;
  assign dataBanks_3_perm_af_data_read_1_3_MPORT_addr = io_raddr_0[0];
  assign dataBanks_3_perm_af_data_read_1_3_MPORT_data =
    dataBanks_3_perm_af[dataBanks_3_perm_af_data_read_1_3_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_3_perm_af_data_read_0_3_MPORT_1_en = 1'h1;
  assign dataBanks_3_perm_af_data_read_0_3_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_3_perm_af_data_read_0_3_MPORT_1_data =
    dataBanks_3_perm_af[dataBanks_3_perm_af_data_read_0_3_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_3_perm_af_data_read_1_3_MPORT_1_en = 1'h1;
  assign dataBanks_3_perm_af_data_read_1_3_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_3_perm_af_data_read_1_3_MPORT_1_data =
    dataBanks_3_perm_af[dataBanks_3_perm_af_data_read_1_3_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_3_perm_af_MPORT_3_data = io_wdata_perm_af;
  assign dataBanks_3_perm_af_MPORT_3_addr = io_waddr[0];
  assign dataBanks_3_perm_af_MPORT_3_mask = 1'h1;
  assign dataBanks_3_perm_af_MPORT_3_en = io_wen & _T_13;
  assign dataBanks_3_perm_d_data_read_0_3_MPORT_en = 1'h1;
  assign dataBanks_3_perm_d_data_read_0_3_MPORT_addr = io_raddr_0[0];
  assign dataBanks_3_perm_d_data_read_0_3_MPORT_data = dataBanks_3_perm_d[dataBanks_3_perm_d_data_read_0_3_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_3_perm_d_data_read_1_3_MPORT_en = 1'h1;
  assign dataBanks_3_perm_d_data_read_1_3_MPORT_addr = io_raddr_0[0];
  assign dataBanks_3_perm_d_data_read_1_3_MPORT_data = dataBanks_3_perm_d[dataBanks_3_perm_d_data_read_1_3_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_3_perm_d_data_read_0_3_MPORT_1_en = 1'h1;
  assign dataBanks_3_perm_d_data_read_0_3_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_3_perm_d_data_read_0_3_MPORT_1_data =
    dataBanks_3_perm_d[dataBanks_3_perm_d_data_read_0_3_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_3_perm_d_data_read_1_3_MPORT_1_en = 1'h1;
  assign dataBanks_3_perm_d_data_read_1_3_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_3_perm_d_data_read_1_3_MPORT_1_data =
    dataBanks_3_perm_d[dataBanks_3_perm_d_data_read_1_3_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_3_perm_d_MPORT_3_data = io_wdata_perm_d;
  assign dataBanks_3_perm_d_MPORT_3_addr = io_waddr[0];
  assign dataBanks_3_perm_d_MPORT_3_mask = 1'h1;
  assign dataBanks_3_perm_d_MPORT_3_en = io_wen & _T_13;
  assign dataBanks_3_perm_a_data_read_0_3_MPORT_en = 1'h1;
  assign dataBanks_3_perm_a_data_read_0_3_MPORT_addr = io_raddr_0[0];
  assign dataBanks_3_perm_a_data_read_0_3_MPORT_data = dataBanks_3_perm_a[dataBanks_3_perm_a_data_read_0_3_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_3_perm_a_data_read_1_3_MPORT_en = 1'h1;
  assign dataBanks_3_perm_a_data_read_1_3_MPORT_addr = io_raddr_0[0];
  assign dataBanks_3_perm_a_data_read_1_3_MPORT_data = dataBanks_3_perm_a[dataBanks_3_perm_a_data_read_1_3_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_3_perm_a_data_read_0_3_MPORT_1_en = 1'h1;
  assign dataBanks_3_perm_a_data_read_0_3_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_3_perm_a_data_read_0_3_MPORT_1_data =
    dataBanks_3_perm_a[dataBanks_3_perm_a_data_read_0_3_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_3_perm_a_data_read_1_3_MPORT_1_en = 1'h1;
  assign dataBanks_3_perm_a_data_read_1_3_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_3_perm_a_data_read_1_3_MPORT_1_data =
    dataBanks_3_perm_a[dataBanks_3_perm_a_data_read_1_3_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_3_perm_a_MPORT_3_data = io_wdata_perm_a;
  assign dataBanks_3_perm_a_MPORT_3_addr = io_waddr[0];
  assign dataBanks_3_perm_a_MPORT_3_mask = 1'h1;
  assign dataBanks_3_perm_a_MPORT_3_en = io_wen & _T_13;
  assign dataBanks_3_perm_u_data_read_0_3_MPORT_en = 1'h1;
  assign dataBanks_3_perm_u_data_read_0_3_MPORT_addr = io_raddr_0[0];
  assign dataBanks_3_perm_u_data_read_0_3_MPORT_data = dataBanks_3_perm_u[dataBanks_3_perm_u_data_read_0_3_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_3_perm_u_data_read_1_3_MPORT_en = 1'h1;
  assign dataBanks_3_perm_u_data_read_1_3_MPORT_addr = io_raddr_0[0];
  assign dataBanks_3_perm_u_data_read_1_3_MPORT_data = dataBanks_3_perm_u[dataBanks_3_perm_u_data_read_1_3_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_3_perm_u_data_read_0_3_MPORT_1_en = 1'h1;
  assign dataBanks_3_perm_u_data_read_0_3_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_3_perm_u_data_read_0_3_MPORT_1_data =
    dataBanks_3_perm_u[dataBanks_3_perm_u_data_read_0_3_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_3_perm_u_data_read_1_3_MPORT_1_en = 1'h1;
  assign dataBanks_3_perm_u_data_read_1_3_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_3_perm_u_data_read_1_3_MPORT_1_data =
    dataBanks_3_perm_u[dataBanks_3_perm_u_data_read_1_3_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_3_perm_u_MPORT_3_data = io_wdata_perm_u;
  assign dataBanks_3_perm_u_MPORT_3_addr = io_waddr[0];
  assign dataBanks_3_perm_u_MPORT_3_mask = 1'h1;
  assign dataBanks_3_perm_u_MPORT_3_en = io_wen & _T_13;
  assign dataBanks_3_perm_x_data_read_0_3_MPORT_en = 1'h1;
  assign dataBanks_3_perm_x_data_read_0_3_MPORT_addr = io_raddr_0[0];
  assign dataBanks_3_perm_x_data_read_0_3_MPORT_data = dataBanks_3_perm_x[dataBanks_3_perm_x_data_read_0_3_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_3_perm_x_data_read_1_3_MPORT_en = 1'h1;
  assign dataBanks_3_perm_x_data_read_1_3_MPORT_addr = io_raddr_0[0];
  assign dataBanks_3_perm_x_data_read_1_3_MPORT_data = dataBanks_3_perm_x[dataBanks_3_perm_x_data_read_1_3_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_3_perm_x_data_read_0_3_MPORT_1_en = 1'h1;
  assign dataBanks_3_perm_x_data_read_0_3_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_3_perm_x_data_read_0_3_MPORT_1_data =
    dataBanks_3_perm_x[dataBanks_3_perm_x_data_read_0_3_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_3_perm_x_data_read_1_3_MPORT_1_en = 1'h1;
  assign dataBanks_3_perm_x_data_read_1_3_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_3_perm_x_data_read_1_3_MPORT_1_data =
    dataBanks_3_perm_x[dataBanks_3_perm_x_data_read_1_3_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_3_perm_x_MPORT_3_data = io_wdata_perm_x;
  assign dataBanks_3_perm_x_MPORT_3_addr = io_waddr[0];
  assign dataBanks_3_perm_x_MPORT_3_mask = 1'h1;
  assign dataBanks_3_perm_x_MPORT_3_en = io_wen & _T_13;
  assign dataBanks_3_perm_wdata_read_0_3_MPORT_en = 1'h1;
  assign dataBanks_3_perm_wdata_read_0_3_MPORT_addr = io_raddr_0[0];
  assign dataBanks_3_perm_wdata_read_0_3_MPORT_data = dataBanks_3_perm_w[dataBanks_3_perm_wdata_read_0_3_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_3_perm_wdata_read_1_3_MPORT_en = 1'h1;
  assign dataBanks_3_perm_wdata_read_1_3_MPORT_addr = io_raddr_0[0];
  assign dataBanks_3_perm_wdata_read_1_3_MPORT_data = dataBanks_3_perm_w[dataBanks_3_perm_wdata_read_1_3_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_3_perm_wdata_read_0_3_MPORT_1_en = 1'h1;
  assign dataBanks_3_perm_wdata_read_0_3_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_3_perm_wdata_read_0_3_MPORT_1_data =
    dataBanks_3_perm_w[dataBanks_3_perm_wdata_read_0_3_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_3_perm_wdata_read_1_3_MPORT_1_en = 1'h1;
  assign dataBanks_3_perm_wdata_read_1_3_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_3_perm_wdata_read_1_3_MPORT_1_data =
    dataBanks_3_perm_w[dataBanks_3_perm_wdata_read_1_3_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_3_perm_wMPORT_3_data = io_wdata_perm_w;
  assign dataBanks_3_perm_wMPORT_3_addr = io_waddr[0];
  assign dataBanks_3_perm_wMPORT_3_mask = 1'h1;
  assign dataBanks_3_perm_wMPORT_3_en = io_wen & _T_13;
  assign dataBanks_3_perm_rdata_read_0_3_MPORT_en = 1'h1;
  assign dataBanks_3_perm_rdata_read_0_3_MPORT_addr = io_raddr_0[0];
  assign dataBanks_3_perm_rdata_read_0_3_MPORT_data = dataBanks_3_perm_r[dataBanks_3_perm_rdata_read_0_3_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_3_perm_rdata_read_1_3_MPORT_en = 1'h1;
  assign dataBanks_3_perm_rdata_read_1_3_MPORT_addr = io_raddr_0[0];
  assign dataBanks_3_perm_rdata_read_1_3_MPORT_data = dataBanks_3_perm_r[dataBanks_3_perm_rdata_read_1_3_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_3_perm_rdata_read_0_3_MPORT_1_en = 1'h1;
  assign dataBanks_3_perm_rdata_read_0_3_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_3_perm_rdata_read_0_3_MPORT_1_data =
    dataBanks_3_perm_r[dataBanks_3_perm_rdata_read_0_3_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_3_perm_rdata_read_1_3_MPORT_1_en = 1'h1;
  assign dataBanks_3_perm_rdata_read_1_3_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_3_perm_rdata_read_1_3_MPORT_1_data =
    dataBanks_3_perm_r[dataBanks_3_perm_rdata_read_1_3_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_3_perm_rMPORT_3_data = io_wdata_perm_r;
  assign dataBanks_3_perm_rMPORT_3_addr = io_waddr[0];
  assign dataBanks_3_perm_rMPORT_3_mask = 1'h1;
  assign dataBanks_3_perm_rMPORT_3_en = io_wen & _T_13;
  assign dataBanks_3_perm_pm_rdata_read_0_3_MPORT_en = 1'h1;
  assign dataBanks_3_perm_pm_rdata_read_0_3_MPORT_addr = io_raddr_0[0];
  assign dataBanks_3_perm_pm_rdata_read_0_3_MPORT_data =
    dataBanks_3_perm_pm_r[dataBanks_3_perm_pm_rdata_read_0_3_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_3_perm_pm_rdata_read_1_3_MPORT_en = 1'h1;
  assign dataBanks_3_perm_pm_rdata_read_1_3_MPORT_addr = io_raddr_0[0];
  assign dataBanks_3_perm_pm_rdata_read_1_3_MPORT_data =
    dataBanks_3_perm_pm_r[dataBanks_3_perm_pm_rdata_read_1_3_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_3_perm_pm_rdata_read_0_3_MPORT_1_en = 1'h1;
  assign dataBanks_3_perm_pm_rdata_read_0_3_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_3_perm_pm_rdata_read_0_3_MPORT_1_data =
    dataBanks_3_perm_pm_r[dataBanks_3_perm_pm_rdata_read_0_3_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_3_perm_pm_rdata_read_1_3_MPORT_1_en = 1'h1;
  assign dataBanks_3_perm_pm_rdata_read_1_3_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_3_perm_pm_rdata_read_1_3_MPORT_1_data =
    dataBanks_3_perm_pm_r[dataBanks_3_perm_pm_rdata_read_1_3_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_3_perm_pm_rMPORT_3_data = io_wdata_perm_pm_r;
  assign dataBanks_3_perm_pm_rMPORT_3_addr = io_waddr[0];
  assign dataBanks_3_perm_pm_rMPORT_3_mask = 1'h1;
  assign dataBanks_3_perm_pm_rMPORT_3_en = io_wen & _T_13;
  assign dataBanks_3_perm_pm_wdata_read_0_3_MPORT_en = 1'h1;
  assign dataBanks_3_perm_pm_wdata_read_0_3_MPORT_addr = io_raddr_0[0];
  assign dataBanks_3_perm_pm_wdata_read_0_3_MPORT_data =
    dataBanks_3_perm_pm_w[dataBanks_3_perm_pm_wdata_read_0_3_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_3_perm_pm_wdata_read_1_3_MPORT_en = 1'h1;
  assign dataBanks_3_perm_pm_wdata_read_1_3_MPORT_addr = io_raddr_0[0];
  assign dataBanks_3_perm_pm_wdata_read_1_3_MPORT_data =
    dataBanks_3_perm_pm_w[dataBanks_3_perm_pm_wdata_read_1_3_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_3_perm_pm_wdata_read_0_3_MPORT_1_en = 1'h1;
  assign dataBanks_3_perm_pm_wdata_read_0_3_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_3_perm_pm_wdata_read_0_3_MPORT_1_data =
    dataBanks_3_perm_pm_w[dataBanks_3_perm_pm_wdata_read_0_3_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_3_perm_pm_wdata_read_1_3_MPORT_1_en = 1'h1;
  assign dataBanks_3_perm_pm_wdata_read_1_3_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_3_perm_pm_wdata_read_1_3_MPORT_1_data =
    dataBanks_3_perm_pm_w[dataBanks_3_perm_pm_wdata_read_1_3_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_3_perm_pm_wMPORT_3_data = io_wdata_perm_pm_w;
  assign dataBanks_3_perm_pm_wMPORT_3_addr = io_waddr[0];
  assign dataBanks_3_perm_pm_wMPORT_3_mask = 1'h1;
  assign dataBanks_3_perm_pm_wMPORT_3_en = io_wen & _T_13;
  assign dataBanks_3_perm_pm_c_data_read_0_3_MPORT_en = 1'h1;
  assign dataBanks_3_perm_pm_c_data_read_0_3_MPORT_addr = io_raddr_0[0];
  assign dataBanks_3_perm_pm_c_data_read_0_3_MPORT_data =
    dataBanks_3_perm_pm_c[dataBanks_3_perm_pm_c_data_read_0_3_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_3_perm_pm_c_data_read_1_3_MPORT_en = 1'h1;
  assign dataBanks_3_perm_pm_c_data_read_1_3_MPORT_addr = io_raddr_0[0];
  assign dataBanks_3_perm_pm_c_data_read_1_3_MPORT_data =
    dataBanks_3_perm_pm_c[dataBanks_3_perm_pm_c_data_read_1_3_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_3_perm_pm_c_data_read_0_3_MPORT_1_en = 1'h1;
  assign dataBanks_3_perm_pm_c_data_read_0_3_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_3_perm_pm_c_data_read_0_3_MPORT_1_data =
    dataBanks_3_perm_pm_c[dataBanks_3_perm_pm_c_data_read_0_3_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_3_perm_pm_c_data_read_1_3_MPORT_1_en = 1'h1;
  assign dataBanks_3_perm_pm_c_data_read_1_3_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_3_perm_pm_c_data_read_1_3_MPORT_1_data =
    dataBanks_3_perm_pm_c[dataBanks_3_perm_pm_c_data_read_1_3_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_3_perm_pm_c_MPORT_3_data = io_wdata_perm_pm_c;
  assign dataBanks_3_perm_pm_c_MPORT_3_addr = io_waddr[0];
  assign dataBanks_3_perm_pm_c_MPORT_3_mask = 1'h1;
  assign dataBanks_3_perm_pm_c_MPORT_3_en = io_wen & _T_13;
  assign dataBanks_4_tag_data_read_0_4_MPORT_en = 1'h1;
  assign dataBanks_4_tag_data_read_0_4_MPORT_addr = io_raddr_0[0];
  assign dataBanks_4_tag_data_read_0_4_MPORT_data = dataBanks_4_tag[dataBanks_4_tag_data_read_0_4_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_4_tag_data_read_1_4_MPORT_en = 1'h1;
  assign dataBanks_4_tag_data_read_1_4_MPORT_addr = io_raddr_0[0];
  assign dataBanks_4_tag_data_read_1_4_MPORT_data = dataBanks_4_tag[dataBanks_4_tag_data_read_1_4_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_4_tag_data_read_0_4_MPORT_1_en = 1'h1;
  assign dataBanks_4_tag_data_read_0_4_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_4_tag_data_read_0_4_MPORT_1_data = dataBanks_4_tag[dataBanks_4_tag_data_read_0_4_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_4_tag_data_read_1_4_MPORT_1_en = 1'h1;
  assign dataBanks_4_tag_data_read_1_4_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_4_tag_data_read_1_4_MPORT_1_data = dataBanks_4_tag[dataBanks_4_tag_data_read_1_4_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_4_tag_MPORT_4_data = io_wdata_tag;
  assign dataBanks_4_tag_MPORT_4_addr = io_waddr[0];
  assign dataBanks_4_tag_MPORT_4_mask = 1'h1;
  assign dataBanks_4_tag_MPORT_4_en = io_wen & _T_17;
  assign dataBanks_4_asid_data_read_0_4_MPORT_en = 1'h1;
  assign dataBanks_4_asid_data_read_0_4_MPORT_addr = io_raddr_0[0];
  assign dataBanks_4_asid_data_read_0_4_MPORT_data = dataBanks_4_asid[dataBanks_4_asid_data_read_0_4_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_4_asid_data_read_1_4_MPORT_en = 1'h1;
  assign dataBanks_4_asid_data_read_1_4_MPORT_addr = io_raddr_0[0];
  assign dataBanks_4_asid_data_read_1_4_MPORT_data = dataBanks_4_asid[dataBanks_4_asid_data_read_1_4_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_4_asid_data_read_0_4_MPORT_1_en = 1'h1;
  assign dataBanks_4_asid_data_read_0_4_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_4_asid_data_read_0_4_MPORT_1_data = dataBanks_4_asid[dataBanks_4_asid_data_read_0_4_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_4_asid_data_read_1_4_MPORT_1_en = 1'h1;
  assign dataBanks_4_asid_data_read_1_4_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_4_asid_data_read_1_4_MPORT_1_data = dataBanks_4_asid[dataBanks_4_asid_data_read_1_4_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_4_asid_MPORT_4_data = io_wdata_asid;
  assign dataBanks_4_asid_MPORT_4_addr = io_waddr[0];
  assign dataBanks_4_asid_MPORT_4_mask = 1'h1;
  assign dataBanks_4_asid_MPORT_4_en = io_wen & _T_17;
  assign dataBanks_4_ppn_data_read_0_4_MPORT_en = 1'h1;
  assign dataBanks_4_ppn_data_read_0_4_MPORT_addr = io_raddr_0[0];
  assign dataBanks_4_ppn_data_read_0_4_MPORT_data = dataBanks_4_ppn[dataBanks_4_ppn_data_read_0_4_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_4_ppn_data_read_1_4_MPORT_en = 1'h1;
  assign dataBanks_4_ppn_data_read_1_4_MPORT_addr = io_raddr_0[0];
  assign dataBanks_4_ppn_data_read_1_4_MPORT_data = dataBanks_4_ppn[dataBanks_4_ppn_data_read_1_4_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_4_ppn_data_read_0_4_MPORT_1_en = 1'h1;
  assign dataBanks_4_ppn_data_read_0_4_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_4_ppn_data_read_0_4_MPORT_1_data = dataBanks_4_ppn[dataBanks_4_ppn_data_read_0_4_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_4_ppn_data_read_1_4_MPORT_1_en = 1'h1;
  assign dataBanks_4_ppn_data_read_1_4_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_4_ppn_data_read_1_4_MPORT_1_data = dataBanks_4_ppn[dataBanks_4_ppn_data_read_1_4_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_4_ppn_MPORT_4_data = io_wdata_ppn;
  assign dataBanks_4_ppn_MPORT_4_addr = io_waddr[0];
  assign dataBanks_4_ppn_MPORT_4_mask = 1'h1;
  assign dataBanks_4_ppn_MPORT_4_en = io_wen & _T_17;
  assign dataBanks_4_perm_pf_data_read_0_4_MPORT_en = 1'h1;
  assign dataBanks_4_perm_pf_data_read_0_4_MPORT_addr = io_raddr_0[0];
  assign dataBanks_4_perm_pf_data_read_0_4_MPORT_data =
    dataBanks_4_perm_pf[dataBanks_4_perm_pf_data_read_0_4_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_4_perm_pf_data_read_1_4_MPORT_en = 1'h1;
  assign dataBanks_4_perm_pf_data_read_1_4_MPORT_addr = io_raddr_0[0];
  assign dataBanks_4_perm_pf_data_read_1_4_MPORT_data =
    dataBanks_4_perm_pf[dataBanks_4_perm_pf_data_read_1_4_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_4_perm_pf_data_read_0_4_MPORT_1_en = 1'h1;
  assign dataBanks_4_perm_pf_data_read_0_4_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_4_perm_pf_data_read_0_4_MPORT_1_data =
    dataBanks_4_perm_pf[dataBanks_4_perm_pf_data_read_0_4_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_4_perm_pf_data_read_1_4_MPORT_1_en = 1'h1;
  assign dataBanks_4_perm_pf_data_read_1_4_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_4_perm_pf_data_read_1_4_MPORT_1_data =
    dataBanks_4_perm_pf[dataBanks_4_perm_pf_data_read_1_4_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_4_perm_pf_MPORT_4_data = io_wdata_perm_pf;
  assign dataBanks_4_perm_pf_MPORT_4_addr = io_waddr[0];
  assign dataBanks_4_perm_pf_MPORT_4_mask = 1'h1;
  assign dataBanks_4_perm_pf_MPORT_4_en = io_wen & _T_17;
  assign dataBanks_4_perm_af_data_read_0_4_MPORT_en = 1'h1;
  assign dataBanks_4_perm_af_data_read_0_4_MPORT_addr = io_raddr_0[0];
  assign dataBanks_4_perm_af_data_read_0_4_MPORT_data =
    dataBanks_4_perm_af[dataBanks_4_perm_af_data_read_0_4_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_4_perm_af_data_read_1_4_MPORT_en = 1'h1;
  assign dataBanks_4_perm_af_data_read_1_4_MPORT_addr = io_raddr_0[0];
  assign dataBanks_4_perm_af_data_read_1_4_MPORT_data =
    dataBanks_4_perm_af[dataBanks_4_perm_af_data_read_1_4_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_4_perm_af_data_read_0_4_MPORT_1_en = 1'h1;
  assign dataBanks_4_perm_af_data_read_0_4_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_4_perm_af_data_read_0_4_MPORT_1_data =
    dataBanks_4_perm_af[dataBanks_4_perm_af_data_read_0_4_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_4_perm_af_data_read_1_4_MPORT_1_en = 1'h1;
  assign dataBanks_4_perm_af_data_read_1_4_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_4_perm_af_data_read_1_4_MPORT_1_data =
    dataBanks_4_perm_af[dataBanks_4_perm_af_data_read_1_4_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_4_perm_af_MPORT_4_data = io_wdata_perm_af;
  assign dataBanks_4_perm_af_MPORT_4_addr = io_waddr[0];
  assign dataBanks_4_perm_af_MPORT_4_mask = 1'h1;
  assign dataBanks_4_perm_af_MPORT_4_en = io_wen & _T_17;
  assign dataBanks_4_perm_d_data_read_0_4_MPORT_en = 1'h1;
  assign dataBanks_4_perm_d_data_read_0_4_MPORT_addr = io_raddr_0[0];
  assign dataBanks_4_perm_d_data_read_0_4_MPORT_data = dataBanks_4_perm_d[dataBanks_4_perm_d_data_read_0_4_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_4_perm_d_data_read_1_4_MPORT_en = 1'h1;
  assign dataBanks_4_perm_d_data_read_1_4_MPORT_addr = io_raddr_0[0];
  assign dataBanks_4_perm_d_data_read_1_4_MPORT_data = dataBanks_4_perm_d[dataBanks_4_perm_d_data_read_1_4_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_4_perm_d_data_read_0_4_MPORT_1_en = 1'h1;
  assign dataBanks_4_perm_d_data_read_0_4_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_4_perm_d_data_read_0_4_MPORT_1_data =
    dataBanks_4_perm_d[dataBanks_4_perm_d_data_read_0_4_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_4_perm_d_data_read_1_4_MPORT_1_en = 1'h1;
  assign dataBanks_4_perm_d_data_read_1_4_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_4_perm_d_data_read_1_4_MPORT_1_data =
    dataBanks_4_perm_d[dataBanks_4_perm_d_data_read_1_4_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_4_perm_d_MPORT_4_data = io_wdata_perm_d;
  assign dataBanks_4_perm_d_MPORT_4_addr = io_waddr[0];
  assign dataBanks_4_perm_d_MPORT_4_mask = 1'h1;
  assign dataBanks_4_perm_d_MPORT_4_en = io_wen & _T_17;
  assign dataBanks_4_perm_a_data_read_0_4_MPORT_en = 1'h1;
  assign dataBanks_4_perm_a_data_read_0_4_MPORT_addr = io_raddr_0[0];
  assign dataBanks_4_perm_a_data_read_0_4_MPORT_data = dataBanks_4_perm_a[dataBanks_4_perm_a_data_read_0_4_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_4_perm_a_data_read_1_4_MPORT_en = 1'h1;
  assign dataBanks_4_perm_a_data_read_1_4_MPORT_addr = io_raddr_0[0];
  assign dataBanks_4_perm_a_data_read_1_4_MPORT_data = dataBanks_4_perm_a[dataBanks_4_perm_a_data_read_1_4_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_4_perm_a_data_read_0_4_MPORT_1_en = 1'h1;
  assign dataBanks_4_perm_a_data_read_0_4_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_4_perm_a_data_read_0_4_MPORT_1_data =
    dataBanks_4_perm_a[dataBanks_4_perm_a_data_read_0_4_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_4_perm_a_data_read_1_4_MPORT_1_en = 1'h1;
  assign dataBanks_4_perm_a_data_read_1_4_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_4_perm_a_data_read_1_4_MPORT_1_data =
    dataBanks_4_perm_a[dataBanks_4_perm_a_data_read_1_4_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_4_perm_a_MPORT_4_data = io_wdata_perm_a;
  assign dataBanks_4_perm_a_MPORT_4_addr = io_waddr[0];
  assign dataBanks_4_perm_a_MPORT_4_mask = 1'h1;
  assign dataBanks_4_perm_a_MPORT_4_en = io_wen & _T_17;
  assign dataBanks_4_perm_u_data_read_0_4_MPORT_en = 1'h1;
  assign dataBanks_4_perm_u_data_read_0_4_MPORT_addr = io_raddr_0[0];
  assign dataBanks_4_perm_u_data_read_0_4_MPORT_data = dataBanks_4_perm_u[dataBanks_4_perm_u_data_read_0_4_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_4_perm_u_data_read_1_4_MPORT_en = 1'h1;
  assign dataBanks_4_perm_u_data_read_1_4_MPORT_addr = io_raddr_0[0];
  assign dataBanks_4_perm_u_data_read_1_4_MPORT_data = dataBanks_4_perm_u[dataBanks_4_perm_u_data_read_1_4_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_4_perm_u_data_read_0_4_MPORT_1_en = 1'h1;
  assign dataBanks_4_perm_u_data_read_0_4_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_4_perm_u_data_read_0_4_MPORT_1_data =
    dataBanks_4_perm_u[dataBanks_4_perm_u_data_read_0_4_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_4_perm_u_data_read_1_4_MPORT_1_en = 1'h1;
  assign dataBanks_4_perm_u_data_read_1_4_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_4_perm_u_data_read_1_4_MPORT_1_data =
    dataBanks_4_perm_u[dataBanks_4_perm_u_data_read_1_4_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_4_perm_u_MPORT_4_data = io_wdata_perm_u;
  assign dataBanks_4_perm_u_MPORT_4_addr = io_waddr[0];
  assign dataBanks_4_perm_u_MPORT_4_mask = 1'h1;
  assign dataBanks_4_perm_u_MPORT_4_en = io_wen & _T_17;
  assign dataBanks_4_perm_x_data_read_0_4_MPORT_en = 1'h1;
  assign dataBanks_4_perm_x_data_read_0_4_MPORT_addr = io_raddr_0[0];
  assign dataBanks_4_perm_x_data_read_0_4_MPORT_data = dataBanks_4_perm_x[dataBanks_4_perm_x_data_read_0_4_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_4_perm_x_data_read_1_4_MPORT_en = 1'h1;
  assign dataBanks_4_perm_x_data_read_1_4_MPORT_addr = io_raddr_0[0];
  assign dataBanks_4_perm_x_data_read_1_4_MPORT_data = dataBanks_4_perm_x[dataBanks_4_perm_x_data_read_1_4_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_4_perm_x_data_read_0_4_MPORT_1_en = 1'h1;
  assign dataBanks_4_perm_x_data_read_0_4_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_4_perm_x_data_read_0_4_MPORT_1_data =
    dataBanks_4_perm_x[dataBanks_4_perm_x_data_read_0_4_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_4_perm_x_data_read_1_4_MPORT_1_en = 1'h1;
  assign dataBanks_4_perm_x_data_read_1_4_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_4_perm_x_data_read_1_4_MPORT_1_data =
    dataBanks_4_perm_x[dataBanks_4_perm_x_data_read_1_4_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_4_perm_x_MPORT_4_data = io_wdata_perm_x;
  assign dataBanks_4_perm_x_MPORT_4_addr = io_waddr[0];
  assign dataBanks_4_perm_x_MPORT_4_mask = 1'h1;
  assign dataBanks_4_perm_x_MPORT_4_en = io_wen & _T_17;
  assign dataBanks_4_perm_wdata_read_0_4_MPORT_en = 1'h1;
  assign dataBanks_4_perm_wdata_read_0_4_MPORT_addr = io_raddr_0[0];
  assign dataBanks_4_perm_wdata_read_0_4_MPORT_data = dataBanks_4_perm_w[dataBanks_4_perm_wdata_read_0_4_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_4_perm_wdata_read_1_4_MPORT_en = 1'h1;
  assign dataBanks_4_perm_wdata_read_1_4_MPORT_addr = io_raddr_0[0];
  assign dataBanks_4_perm_wdata_read_1_4_MPORT_data = dataBanks_4_perm_w[dataBanks_4_perm_wdata_read_1_4_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_4_perm_wdata_read_0_4_MPORT_1_en = 1'h1;
  assign dataBanks_4_perm_wdata_read_0_4_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_4_perm_wdata_read_0_4_MPORT_1_data =
    dataBanks_4_perm_w[dataBanks_4_perm_wdata_read_0_4_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_4_perm_wdata_read_1_4_MPORT_1_en = 1'h1;
  assign dataBanks_4_perm_wdata_read_1_4_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_4_perm_wdata_read_1_4_MPORT_1_data =
    dataBanks_4_perm_w[dataBanks_4_perm_wdata_read_1_4_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_4_perm_wMPORT_4_data = io_wdata_perm_w;
  assign dataBanks_4_perm_wMPORT_4_addr = io_waddr[0];
  assign dataBanks_4_perm_wMPORT_4_mask = 1'h1;
  assign dataBanks_4_perm_wMPORT_4_en = io_wen & _T_17;
  assign dataBanks_4_perm_rdata_read_0_4_MPORT_en = 1'h1;
  assign dataBanks_4_perm_rdata_read_0_4_MPORT_addr = io_raddr_0[0];
  assign dataBanks_4_perm_rdata_read_0_4_MPORT_data = dataBanks_4_perm_r[dataBanks_4_perm_rdata_read_0_4_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_4_perm_rdata_read_1_4_MPORT_en = 1'h1;
  assign dataBanks_4_perm_rdata_read_1_4_MPORT_addr = io_raddr_0[0];
  assign dataBanks_4_perm_rdata_read_1_4_MPORT_data = dataBanks_4_perm_r[dataBanks_4_perm_rdata_read_1_4_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_4_perm_rdata_read_0_4_MPORT_1_en = 1'h1;
  assign dataBanks_4_perm_rdata_read_0_4_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_4_perm_rdata_read_0_4_MPORT_1_data =
    dataBanks_4_perm_r[dataBanks_4_perm_rdata_read_0_4_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_4_perm_rdata_read_1_4_MPORT_1_en = 1'h1;
  assign dataBanks_4_perm_rdata_read_1_4_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_4_perm_rdata_read_1_4_MPORT_1_data =
    dataBanks_4_perm_r[dataBanks_4_perm_rdata_read_1_4_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_4_perm_rMPORT_4_data = io_wdata_perm_r;
  assign dataBanks_4_perm_rMPORT_4_addr = io_waddr[0];
  assign dataBanks_4_perm_rMPORT_4_mask = 1'h1;
  assign dataBanks_4_perm_rMPORT_4_en = io_wen & _T_17;
  assign dataBanks_4_perm_pm_rdata_read_0_4_MPORT_en = 1'h1;
  assign dataBanks_4_perm_pm_rdata_read_0_4_MPORT_addr = io_raddr_0[0];
  assign dataBanks_4_perm_pm_rdata_read_0_4_MPORT_data =
    dataBanks_4_perm_pm_r[dataBanks_4_perm_pm_rdata_read_0_4_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_4_perm_pm_rdata_read_1_4_MPORT_en = 1'h1;
  assign dataBanks_4_perm_pm_rdata_read_1_4_MPORT_addr = io_raddr_0[0];
  assign dataBanks_4_perm_pm_rdata_read_1_4_MPORT_data =
    dataBanks_4_perm_pm_r[dataBanks_4_perm_pm_rdata_read_1_4_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_4_perm_pm_rdata_read_0_4_MPORT_1_en = 1'h1;
  assign dataBanks_4_perm_pm_rdata_read_0_4_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_4_perm_pm_rdata_read_0_4_MPORT_1_data =
    dataBanks_4_perm_pm_r[dataBanks_4_perm_pm_rdata_read_0_4_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_4_perm_pm_rdata_read_1_4_MPORT_1_en = 1'h1;
  assign dataBanks_4_perm_pm_rdata_read_1_4_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_4_perm_pm_rdata_read_1_4_MPORT_1_data =
    dataBanks_4_perm_pm_r[dataBanks_4_perm_pm_rdata_read_1_4_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_4_perm_pm_rMPORT_4_data = io_wdata_perm_pm_r;
  assign dataBanks_4_perm_pm_rMPORT_4_addr = io_waddr[0];
  assign dataBanks_4_perm_pm_rMPORT_4_mask = 1'h1;
  assign dataBanks_4_perm_pm_rMPORT_4_en = io_wen & _T_17;
  assign dataBanks_4_perm_pm_wdata_read_0_4_MPORT_en = 1'h1;
  assign dataBanks_4_perm_pm_wdata_read_0_4_MPORT_addr = io_raddr_0[0];
  assign dataBanks_4_perm_pm_wdata_read_0_4_MPORT_data =
    dataBanks_4_perm_pm_w[dataBanks_4_perm_pm_wdata_read_0_4_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_4_perm_pm_wdata_read_1_4_MPORT_en = 1'h1;
  assign dataBanks_4_perm_pm_wdata_read_1_4_MPORT_addr = io_raddr_0[0];
  assign dataBanks_4_perm_pm_wdata_read_1_4_MPORT_data =
    dataBanks_4_perm_pm_w[dataBanks_4_perm_pm_wdata_read_1_4_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_4_perm_pm_wdata_read_0_4_MPORT_1_en = 1'h1;
  assign dataBanks_4_perm_pm_wdata_read_0_4_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_4_perm_pm_wdata_read_0_4_MPORT_1_data =
    dataBanks_4_perm_pm_w[dataBanks_4_perm_pm_wdata_read_0_4_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_4_perm_pm_wdata_read_1_4_MPORT_1_en = 1'h1;
  assign dataBanks_4_perm_pm_wdata_read_1_4_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_4_perm_pm_wdata_read_1_4_MPORT_1_data =
    dataBanks_4_perm_pm_w[dataBanks_4_perm_pm_wdata_read_1_4_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_4_perm_pm_wMPORT_4_data = io_wdata_perm_pm_w;
  assign dataBanks_4_perm_pm_wMPORT_4_addr = io_waddr[0];
  assign dataBanks_4_perm_pm_wMPORT_4_mask = 1'h1;
  assign dataBanks_4_perm_pm_wMPORT_4_en = io_wen & _T_17;
  assign dataBanks_4_perm_pm_c_data_read_0_4_MPORT_en = 1'h1;
  assign dataBanks_4_perm_pm_c_data_read_0_4_MPORT_addr = io_raddr_0[0];
  assign dataBanks_4_perm_pm_c_data_read_0_4_MPORT_data =
    dataBanks_4_perm_pm_c[dataBanks_4_perm_pm_c_data_read_0_4_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_4_perm_pm_c_data_read_1_4_MPORT_en = 1'h1;
  assign dataBanks_4_perm_pm_c_data_read_1_4_MPORT_addr = io_raddr_0[0];
  assign dataBanks_4_perm_pm_c_data_read_1_4_MPORT_data =
    dataBanks_4_perm_pm_c[dataBanks_4_perm_pm_c_data_read_1_4_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_4_perm_pm_c_data_read_0_4_MPORT_1_en = 1'h1;
  assign dataBanks_4_perm_pm_c_data_read_0_4_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_4_perm_pm_c_data_read_0_4_MPORT_1_data =
    dataBanks_4_perm_pm_c[dataBanks_4_perm_pm_c_data_read_0_4_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_4_perm_pm_c_data_read_1_4_MPORT_1_en = 1'h1;
  assign dataBanks_4_perm_pm_c_data_read_1_4_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_4_perm_pm_c_data_read_1_4_MPORT_1_data =
    dataBanks_4_perm_pm_c[dataBanks_4_perm_pm_c_data_read_1_4_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_4_perm_pm_c_MPORT_4_data = io_wdata_perm_pm_c;
  assign dataBanks_4_perm_pm_c_MPORT_4_addr = io_waddr[0];
  assign dataBanks_4_perm_pm_c_MPORT_4_mask = 1'h1;
  assign dataBanks_4_perm_pm_c_MPORT_4_en = io_wen & _T_17;
  assign dataBanks_5_tag_data_read_0_5_MPORT_en = 1'h1;
  assign dataBanks_5_tag_data_read_0_5_MPORT_addr = io_raddr_0[0];
  assign dataBanks_5_tag_data_read_0_5_MPORT_data = dataBanks_5_tag[dataBanks_5_tag_data_read_0_5_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_5_tag_data_read_1_5_MPORT_en = 1'h1;
  assign dataBanks_5_tag_data_read_1_5_MPORT_addr = io_raddr_0[0];
  assign dataBanks_5_tag_data_read_1_5_MPORT_data = dataBanks_5_tag[dataBanks_5_tag_data_read_1_5_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_5_tag_data_read_0_5_MPORT_1_en = 1'h1;
  assign dataBanks_5_tag_data_read_0_5_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_5_tag_data_read_0_5_MPORT_1_data = dataBanks_5_tag[dataBanks_5_tag_data_read_0_5_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_5_tag_data_read_1_5_MPORT_1_en = 1'h1;
  assign dataBanks_5_tag_data_read_1_5_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_5_tag_data_read_1_5_MPORT_1_data = dataBanks_5_tag[dataBanks_5_tag_data_read_1_5_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_5_tag_MPORT_5_data = io_wdata_tag;
  assign dataBanks_5_tag_MPORT_5_addr = io_waddr[0];
  assign dataBanks_5_tag_MPORT_5_mask = 1'h1;
  assign dataBanks_5_tag_MPORT_5_en = io_wen & _T_21;
  assign dataBanks_5_asid_data_read_0_5_MPORT_en = 1'h1;
  assign dataBanks_5_asid_data_read_0_5_MPORT_addr = io_raddr_0[0];
  assign dataBanks_5_asid_data_read_0_5_MPORT_data = dataBanks_5_asid[dataBanks_5_asid_data_read_0_5_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_5_asid_data_read_1_5_MPORT_en = 1'h1;
  assign dataBanks_5_asid_data_read_1_5_MPORT_addr = io_raddr_0[0];
  assign dataBanks_5_asid_data_read_1_5_MPORT_data = dataBanks_5_asid[dataBanks_5_asid_data_read_1_5_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_5_asid_data_read_0_5_MPORT_1_en = 1'h1;
  assign dataBanks_5_asid_data_read_0_5_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_5_asid_data_read_0_5_MPORT_1_data = dataBanks_5_asid[dataBanks_5_asid_data_read_0_5_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_5_asid_data_read_1_5_MPORT_1_en = 1'h1;
  assign dataBanks_5_asid_data_read_1_5_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_5_asid_data_read_1_5_MPORT_1_data = dataBanks_5_asid[dataBanks_5_asid_data_read_1_5_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_5_asid_MPORT_5_data = io_wdata_asid;
  assign dataBanks_5_asid_MPORT_5_addr = io_waddr[0];
  assign dataBanks_5_asid_MPORT_5_mask = 1'h1;
  assign dataBanks_5_asid_MPORT_5_en = io_wen & _T_21;
  assign dataBanks_5_ppn_data_read_0_5_MPORT_en = 1'h1;
  assign dataBanks_5_ppn_data_read_0_5_MPORT_addr = io_raddr_0[0];
  assign dataBanks_5_ppn_data_read_0_5_MPORT_data = dataBanks_5_ppn[dataBanks_5_ppn_data_read_0_5_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_5_ppn_data_read_1_5_MPORT_en = 1'h1;
  assign dataBanks_5_ppn_data_read_1_5_MPORT_addr = io_raddr_0[0];
  assign dataBanks_5_ppn_data_read_1_5_MPORT_data = dataBanks_5_ppn[dataBanks_5_ppn_data_read_1_5_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_5_ppn_data_read_0_5_MPORT_1_en = 1'h1;
  assign dataBanks_5_ppn_data_read_0_5_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_5_ppn_data_read_0_5_MPORT_1_data = dataBanks_5_ppn[dataBanks_5_ppn_data_read_0_5_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_5_ppn_data_read_1_5_MPORT_1_en = 1'h1;
  assign dataBanks_5_ppn_data_read_1_5_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_5_ppn_data_read_1_5_MPORT_1_data = dataBanks_5_ppn[dataBanks_5_ppn_data_read_1_5_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_5_ppn_MPORT_5_data = io_wdata_ppn;
  assign dataBanks_5_ppn_MPORT_5_addr = io_waddr[0];
  assign dataBanks_5_ppn_MPORT_5_mask = 1'h1;
  assign dataBanks_5_ppn_MPORT_5_en = io_wen & _T_21;
  assign dataBanks_5_perm_pf_data_read_0_5_MPORT_en = 1'h1;
  assign dataBanks_5_perm_pf_data_read_0_5_MPORT_addr = io_raddr_0[0];
  assign dataBanks_5_perm_pf_data_read_0_5_MPORT_data =
    dataBanks_5_perm_pf[dataBanks_5_perm_pf_data_read_0_5_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_5_perm_pf_data_read_1_5_MPORT_en = 1'h1;
  assign dataBanks_5_perm_pf_data_read_1_5_MPORT_addr = io_raddr_0[0];
  assign dataBanks_5_perm_pf_data_read_1_5_MPORT_data =
    dataBanks_5_perm_pf[dataBanks_5_perm_pf_data_read_1_5_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_5_perm_pf_data_read_0_5_MPORT_1_en = 1'h1;
  assign dataBanks_5_perm_pf_data_read_0_5_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_5_perm_pf_data_read_0_5_MPORT_1_data =
    dataBanks_5_perm_pf[dataBanks_5_perm_pf_data_read_0_5_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_5_perm_pf_data_read_1_5_MPORT_1_en = 1'h1;
  assign dataBanks_5_perm_pf_data_read_1_5_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_5_perm_pf_data_read_1_5_MPORT_1_data =
    dataBanks_5_perm_pf[dataBanks_5_perm_pf_data_read_1_5_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_5_perm_pf_MPORT_5_data = io_wdata_perm_pf;
  assign dataBanks_5_perm_pf_MPORT_5_addr = io_waddr[0];
  assign dataBanks_5_perm_pf_MPORT_5_mask = 1'h1;
  assign dataBanks_5_perm_pf_MPORT_5_en = io_wen & _T_21;
  assign dataBanks_5_perm_af_data_read_0_5_MPORT_en = 1'h1;
  assign dataBanks_5_perm_af_data_read_0_5_MPORT_addr = io_raddr_0[0];
  assign dataBanks_5_perm_af_data_read_0_5_MPORT_data =
    dataBanks_5_perm_af[dataBanks_5_perm_af_data_read_0_5_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_5_perm_af_data_read_1_5_MPORT_en = 1'h1;
  assign dataBanks_5_perm_af_data_read_1_5_MPORT_addr = io_raddr_0[0];
  assign dataBanks_5_perm_af_data_read_1_5_MPORT_data =
    dataBanks_5_perm_af[dataBanks_5_perm_af_data_read_1_5_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_5_perm_af_data_read_0_5_MPORT_1_en = 1'h1;
  assign dataBanks_5_perm_af_data_read_0_5_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_5_perm_af_data_read_0_5_MPORT_1_data =
    dataBanks_5_perm_af[dataBanks_5_perm_af_data_read_0_5_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_5_perm_af_data_read_1_5_MPORT_1_en = 1'h1;
  assign dataBanks_5_perm_af_data_read_1_5_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_5_perm_af_data_read_1_5_MPORT_1_data =
    dataBanks_5_perm_af[dataBanks_5_perm_af_data_read_1_5_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_5_perm_af_MPORT_5_data = io_wdata_perm_af;
  assign dataBanks_5_perm_af_MPORT_5_addr = io_waddr[0];
  assign dataBanks_5_perm_af_MPORT_5_mask = 1'h1;
  assign dataBanks_5_perm_af_MPORT_5_en = io_wen & _T_21;
  assign dataBanks_5_perm_d_data_read_0_5_MPORT_en = 1'h1;
  assign dataBanks_5_perm_d_data_read_0_5_MPORT_addr = io_raddr_0[0];
  assign dataBanks_5_perm_d_data_read_0_5_MPORT_data = dataBanks_5_perm_d[dataBanks_5_perm_d_data_read_0_5_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_5_perm_d_data_read_1_5_MPORT_en = 1'h1;
  assign dataBanks_5_perm_d_data_read_1_5_MPORT_addr = io_raddr_0[0];
  assign dataBanks_5_perm_d_data_read_1_5_MPORT_data = dataBanks_5_perm_d[dataBanks_5_perm_d_data_read_1_5_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_5_perm_d_data_read_0_5_MPORT_1_en = 1'h1;
  assign dataBanks_5_perm_d_data_read_0_5_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_5_perm_d_data_read_0_5_MPORT_1_data =
    dataBanks_5_perm_d[dataBanks_5_perm_d_data_read_0_5_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_5_perm_d_data_read_1_5_MPORT_1_en = 1'h1;
  assign dataBanks_5_perm_d_data_read_1_5_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_5_perm_d_data_read_1_5_MPORT_1_data =
    dataBanks_5_perm_d[dataBanks_5_perm_d_data_read_1_5_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_5_perm_d_MPORT_5_data = io_wdata_perm_d;
  assign dataBanks_5_perm_d_MPORT_5_addr = io_waddr[0];
  assign dataBanks_5_perm_d_MPORT_5_mask = 1'h1;
  assign dataBanks_5_perm_d_MPORT_5_en = io_wen & _T_21;
  assign dataBanks_5_perm_a_data_read_0_5_MPORT_en = 1'h1;
  assign dataBanks_5_perm_a_data_read_0_5_MPORT_addr = io_raddr_0[0];
  assign dataBanks_5_perm_a_data_read_0_5_MPORT_data = dataBanks_5_perm_a[dataBanks_5_perm_a_data_read_0_5_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_5_perm_a_data_read_1_5_MPORT_en = 1'h1;
  assign dataBanks_5_perm_a_data_read_1_5_MPORT_addr = io_raddr_0[0];
  assign dataBanks_5_perm_a_data_read_1_5_MPORT_data = dataBanks_5_perm_a[dataBanks_5_perm_a_data_read_1_5_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_5_perm_a_data_read_0_5_MPORT_1_en = 1'h1;
  assign dataBanks_5_perm_a_data_read_0_5_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_5_perm_a_data_read_0_5_MPORT_1_data =
    dataBanks_5_perm_a[dataBanks_5_perm_a_data_read_0_5_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_5_perm_a_data_read_1_5_MPORT_1_en = 1'h1;
  assign dataBanks_5_perm_a_data_read_1_5_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_5_perm_a_data_read_1_5_MPORT_1_data =
    dataBanks_5_perm_a[dataBanks_5_perm_a_data_read_1_5_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_5_perm_a_MPORT_5_data = io_wdata_perm_a;
  assign dataBanks_5_perm_a_MPORT_5_addr = io_waddr[0];
  assign dataBanks_5_perm_a_MPORT_5_mask = 1'h1;
  assign dataBanks_5_perm_a_MPORT_5_en = io_wen & _T_21;
  assign dataBanks_5_perm_u_data_read_0_5_MPORT_en = 1'h1;
  assign dataBanks_5_perm_u_data_read_0_5_MPORT_addr = io_raddr_0[0];
  assign dataBanks_5_perm_u_data_read_0_5_MPORT_data = dataBanks_5_perm_u[dataBanks_5_perm_u_data_read_0_5_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_5_perm_u_data_read_1_5_MPORT_en = 1'h1;
  assign dataBanks_5_perm_u_data_read_1_5_MPORT_addr = io_raddr_0[0];
  assign dataBanks_5_perm_u_data_read_1_5_MPORT_data = dataBanks_5_perm_u[dataBanks_5_perm_u_data_read_1_5_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_5_perm_u_data_read_0_5_MPORT_1_en = 1'h1;
  assign dataBanks_5_perm_u_data_read_0_5_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_5_perm_u_data_read_0_5_MPORT_1_data =
    dataBanks_5_perm_u[dataBanks_5_perm_u_data_read_0_5_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_5_perm_u_data_read_1_5_MPORT_1_en = 1'h1;
  assign dataBanks_5_perm_u_data_read_1_5_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_5_perm_u_data_read_1_5_MPORT_1_data =
    dataBanks_5_perm_u[dataBanks_5_perm_u_data_read_1_5_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_5_perm_u_MPORT_5_data = io_wdata_perm_u;
  assign dataBanks_5_perm_u_MPORT_5_addr = io_waddr[0];
  assign dataBanks_5_perm_u_MPORT_5_mask = 1'h1;
  assign dataBanks_5_perm_u_MPORT_5_en = io_wen & _T_21;
  assign dataBanks_5_perm_x_data_read_0_5_MPORT_en = 1'h1;
  assign dataBanks_5_perm_x_data_read_0_5_MPORT_addr = io_raddr_0[0];
  assign dataBanks_5_perm_x_data_read_0_5_MPORT_data = dataBanks_5_perm_x[dataBanks_5_perm_x_data_read_0_5_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_5_perm_x_data_read_1_5_MPORT_en = 1'h1;
  assign dataBanks_5_perm_x_data_read_1_5_MPORT_addr = io_raddr_0[0];
  assign dataBanks_5_perm_x_data_read_1_5_MPORT_data = dataBanks_5_perm_x[dataBanks_5_perm_x_data_read_1_5_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_5_perm_x_data_read_0_5_MPORT_1_en = 1'h1;
  assign dataBanks_5_perm_x_data_read_0_5_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_5_perm_x_data_read_0_5_MPORT_1_data =
    dataBanks_5_perm_x[dataBanks_5_perm_x_data_read_0_5_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_5_perm_x_data_read_1_5_MPORT_1_en = 1'h1;
  assign dataBanks_5_perm_x_data_read_1_5_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_5_perm_x_data_read_1_5_MPORT_1_data =
    dataBanks_5_perm_x[dataBanks_5_perm_x_data_read_1_5_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_5_perm_x_MPORT_5_data = io_wdata_perm_x;
  assign dataBanks_5_perm_x_MPORT_5_addr = io_waddr[0];
  assign dataBanks_5_perm_x_MPORT_5_mask = 1'h1;
  assign dataBanks_5_perm_x_MPORT_5_en = io_wen & _T_21;
  assign dataBanks_5_perm_wdata_read_0_5_MPORT_en = 1'h1;
  assign dataBanks_5_perm_wdata_read_0_5_MPORT_addr = io_raddr_0[0];
  assign dataBanks_5_perm_wdata_read_0_5_MPORT_data = dataBanks_5_perm_w[dataBanks_5_perm_wdata_read_0_5_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_5_perm_wdata_read_1_5_MPORT_en = 1'h1;
  assign dataBanks_5_perm_wdata_read_1_5_MPORT_addr = io_raddr_0[0];
  assign dataBanks_5_perm_wdata_read_1_5_MPORT_data = dataBanks_5_perm_w[dataBanks_5_perm_wdata_read_1_5_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_5_perm_wdata_read_0_5_MPORT_1_en = 1'h1;
  assign dataBanks_5_perm_wdata_read_0_5_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_5_perm_wdata_read_0_5_MPORT_1_data =
    dataBanks_5_perm_w[dataBanks_5_perm_wdata_read_0_5_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_5_perm_wdata_read_1_5_MPORT_1_en = 1'h1;
  assign dataBanks_5_perm_wdata_read_1_5_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_5_perm_wdata_read_1_5_MPORT_1_data =
    dataBanks_5_perm_w[dataBanks_5_perm_wdata_read_1_5_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_5_perm_wMPORT_5_data = io_wdata_perm_w;
  assign dataBanks_5_perm_wMPORT_5_addr = io_waddr[0];
  assign dataBanks_5_perm_wMPORT_5_mask = 1'h1;
  assign dataBanks_5_perm_wMPORT_5_en = io_wen & _T_21;
  assign dataBanks_5_perm_rdata_read_0_5_MPORT_en = 1'h1;
  assign dataBanks_5_perm_rdata_read_0_5_MPORT_addr = io_raddr_0[0];
  assign dataBanks_5_perm_rdata_read_0_5_MPORT_data = dataBanks_5_perm_r[dataBanks_5_perm_rdata_read_0_5_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_5_perm_rdata_read_1_5_MPORT_en = 1'h1;
  assign dataBanks_5_perm_rdata_read_1_5_MPORT_addr = io_raddr_0[0];
  assign dataBanks_5_perm_rdata_read_1_5_MPORT_data = dataBanks_5_perm_r[dataBanks_5_perm_rdata_read_1_5_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_5_perm_rdata_read_0_5_MPORT_1_en = 1'h1;
  assign dataBanks_5_perm_rdata_read_0_5_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_5_perm_rdata_read_0_5_MPORT_1_data =
    dataBanks_5_perm_r[dataBanks_5_perm_rdata_read_0_5_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_5_perm_rdata_read_1_5_MPORT_1_en = 1'h1;
  assign dataBanks_5_perm_rdata_read_1_5_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_5_perm_rdata_read_1_5_MPORT_1_data =
    dataBanks_5_perm_r[dataBanks_5_perm_rdata_read_1_5_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_5_perm_rMPORT_5_data = io_wdata_perm_r;
  assign dataBanks_5_perm_rMPORT_5_addr = io_waddr[0];
  assign dataBanks_5_perm_rMPORT_5_mask = 1'h1;
  assign dataBanks_5_perm_rMPORT_5_en = io_wen & _T_21;
  assign dataBanks_5_perm_pm_rdata_read_0_5_MPORT_en = 1'h1;
  assign dataBanks_5_perm_pm_rdata_read_0_5_MPORT_addr = io_raddr_0[0];
  assign dataBanks_5_perm_pm_rdata_read_0_5_MPORT_data =
    dataBanks_5_perm_pm_r[dataBanks_5_perm_pm_rdata_read_0_5_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_5_perm_pm_rdata_read_1_5_MPORT_en = 1'h1;
  assign dataBanks_5_perm_pm_rdata_read_1_5_MPORT_addr = io_raddr_0[0];
  assign dataBanks_5_perm_pm_rdata_read_1_5_MPORT_data =
    dataBanks_5_perm_pm_r[dataBanks_5_perm_pm_rdata_read_1_5_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_5_perm_pm_rdata_read_0_5_MPORT_1_en = 1'h1;
  assign dataBanks_5_perm_pm_rdata_read_0_5_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_5_perm_pm_rdata_read_0_5_MPORT_1_data =
    dataBanks_5_perm_pm_r[dataBanks_5_perm_pm_rdata_read_0_5_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_5_perm_pm_rdata_read_1_5_MPORT_1_en = 1'h1;
  assign dataBanks_5_perm_pm_rdata_read_1_5_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_5_perm_pm_rdata_read_1_5_MPORT_1_data =
    dataBanks_5_perm_pm_r[dataBanks_5_perm_pm_rdata_read_1_5_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_5_perm_pm_rMPORT_5_data = io_wdata_perm_pm_r;
  assign dataBanks_5_perm_pm_rMPORT_5_addr = io_waddr[0];
  assign dataBanks_5_perm_pm_rMPORT_5_mask = 1'h1;
  assign dataBanks_5_perm_pm_rMPORT_5_en = io_wen & _T_21;
  assign dataBanks_5_perm_pm_wdata_read_0_5_MPORT_en = 1'h1;
  assign dataBanks_5_perm_pm_wdata_read_0_5_MPORT_addr = io_raddr_0[0];
  assign dataBanks_5_perm_pm_wdata_read_0_5_MPORT_data =
    dataBanks_5_perm_pm_w[dataBanks_5_perm_pm_wdata_read_0_5_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_5_perm_pm_wdata_read_1_5_MPORT_en = 1'h1;
  assign dataBanks_5_perm_pm_wdata_read_1_5_MPORT_addr = io_raddr_0[0];
  assign dataBanks_5_perm_pm_wdata_read_1_5_MPORT_data =
    dataBanks_5_perm_pm_w[dataBanks_5_perm_pm_wdata_read_1_5_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_5_perm_pm_wdata_read_0_5_MPORT_1_en = 1'h1;
  assign dataBanks_5_perm_pm_wdata_read_0_5_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_5_perm_pm_wdata_read_0_5_MPORT_1_data =
    dataBanks_5_perm_pm_w[dataBanks_5_perm_pm_wdata_read_0_5_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_5_perm_pm_wdata_read_1_5_MPORT_1_en = 1'h1;
  assign dataBanks_5_perm_pm_wdata_read_1_5_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_5_perm_pm_wdata_read_1_5_MPORT_1_data =
    dataBanks_5_perm_pm_w[dataBanks_5_perm_pm_wdata_read_1_5_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_5_perm_pm_wMPORT_5_data = io_wdata_perm_pm_w;
  assign dataBanks_5_perm_pm_wMPORT_5_addr = io_waddr[0];
  assign dataBanks_5_perm_pm_wMPORT_5_mask = 1'h1;
  assign dataBanks_5_perm_pm_wMPORT_5_en = io_wen & _T_21;
  assign dataBanks_5_perm_pm_c_data_read_0_5_MPORT_en = 1'h1;
  assign dataBanks_5_perm_pm_c_data_read_0_5_MPORT_addr = io_raddr_0[0];
  assign dataBanks_5_perm_pm_c_data_read_0_5_MPORT_data =
    dataBanks_5_perm_pm_c[dataBanks_5_perm_pm_c_data_read_0_5_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_5_perm_pm_c_data_read_1_5_MPORT_en = 1'h1;
  assign dataBanks_5_perm_pm_c_data_read_1_5_MPORT_addr = io_raddr_0[0];
  assign dataBanks_5_perm_pm_c_data_read_1_5_MPORT_data =
    dataBanks_5_perm_pm_c[dataBanks_5_perm_pm_c_data_read_1_5_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_5_perm_pm_c_data_read_0_5_MPORT_1_en = 1'h1;
  assign dataBanks_5_perm_pm_c_data_read_0_5_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_5_perm_pm_c_data_read_0_5_MPORT_1_data =
    dataBanks_5_perm_pm_c[dataBanks_5_perm_pm_c_data_read_0_5_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_5_perm_pm_c_data_read_1_5_MPORT_1_en = 1'h1;
  assign dataBanks_5_perm_pm_c_data_read_1_5_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_5_perm_pm_c_data_read_1_5_MPORT_1_data =
    dataBanks_5_perm_pm_c[dataBanks_5_perm_pm_c_data_read_1_5_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_5_perm_pm_c_MPORT_5_data = io_wdata_perm_pm_c;
  assign dataBanks_5_perm_pm_c_MPORT_5_addr = io_waddr[0];
  assign dataBanks_5_perm_pm_c_MPORT_5_mask = 1'h1;
  assign dataBanks_5_perm_pm_c_MPORT_5_en = io_wen & _T_21;
  assign dataBanks_6_tag_data_read_0_6_MPORT_en = 1'h1;
  assign dataBanks_6_tag_data_read_0_6_MPORT_addr = io_raddr_0[0];
  assign dataBanks_6_tag_data_read_0_6_MPORT_data = dataBanks_6_tag[dataBanks_6_tag_data_read_0_6_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_6_tag_data_read_1_6_MPORT_en = 1'h1;
  assign dataBanks_6_tag_data_read_1_6_MPORT_addr = io_raddr_0[0];
  assign dataBanks_6_tag_data_read_1_6_MPORT_data = dataBanks_6_tag[dataBanks_6_tag_data_read_1_6_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_6_tag_data_read_0_6_MPORT_1_en = 1'h1;
  assign dataBanks_6_tag_data_read_0_6_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_6_tag_data_read_0_6_MPORT_1_data = dataBanks_6_tag[dataBanks_6_tag_data_read_0_6_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_6_tag_data_read_1_6_MPORT_1_en = 1'h1;
  assign dataBanks_6_tag_data_read_1_6_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_6_tag_data_read_1_6_MPORT_1_data = dataBanks_6_tag[dataBanks_6_tag_data_read_1_6_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_6_tag_MPORT_6_data = io_wdata_tag;
  assign dataBanks_6_tag_MPORT_6_addr = io_waddr[0];
  assign dataBanks_6_tag_MPORT_6_mask = 1'h1;
  assign dataBanks_6_tag_MPORT_6_en = io_wen & _T_25;
  assign dataBanks_6_asid_data_read_0_6_MPORT_en = 1'h1;
  assign dataBanks_6_asid_data_read_0_6_MPORT_addr = io_raddr_0[0];
  assign dataBanks_6_asid_data_read_0_6_MPORT_data = dataBanks_6_asid[dataBanks_6_asid_data_read_0_6_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_6_asid_data_read_1_6_MPORT_en = 1'h1;
  assign dataBanks_6_asid_data_read_1_6_MPORT_addr = io_raddr_0[0];
  assign dataBanks_6_asid_data_read_1_6_MPORT_data = dataBanks_6_asid[dataBanks_6_asid_data_read_1_6_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_6_asid_data_read_0_6_MPORT_1_en = 1'h1;
  assign dataBanks_6_asid_data_read_0_6_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_6_asid_data_read_0_6_MPORT_1_data = dataBanks_6_asid[dataBanks_6_asid_data_read_0_6_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_6_asid_data_read_1_6_MPORT_1_en = 1'h1;
  assign dataBanks_6_asid_data_read_1_6_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_6_asid_data_read_1_6_MPORT_1_data = dataBanks_6_asid[dataBanks_6_asid_data_read_1_6_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_6_asid_MPORT_6_data = io_wdata_asid;
  assign dataBanks_6_asid_MPORT_6_addr = io_waddr[0];
  assign dataBanks_6_asid_MPORT_6_mask = 1'h1;
  assign dataBanks_6_asid_MPORT_6_en = io_wen & _T_25;
  assign dataBanks_6_ppn_data_read_0_6_MPORT_en = 1'h1;
  assign dataBanks_6_ppn_data_read_0_6_MPORT_addr = io_raddr_0[0];
  assign dataBanks_6_ppn_data_read_0_6_MPORT_data = dataBanks_6_ppn[dataBanks_6_ppn_data_read_0_6_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_6_ppn_data_read_1_6_MPORT_en = 1'h1;
  assign dataBanks_6_ppn_data_read_1_6_MPORT_addr = io_raddr_0[0];
  assign dataBanks_6_ppn_data_read_1_6_MPORT_data = dataBanks_6_ppn[dataBanks_6_ppn_data_read_1_6_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_6_ppn_data_read_0_6_MPORT_1_en = 1'h1;
  assign dataBanks_6_ppn_data_read_0_6_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_6_ppn_data_read_0_6_MPORT_1_data = dataBanks_6_ppn[dataBanks_6_ppn_data_read_0_6_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_6_ppn_data_read_1_6_MPORT_1_en = 1'h1;
  assign dataBanks_6_ppn_data_read_1_6_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_6_ppn_data_read_1_6_MPORT_1_data = dataBanks_6_ppn[dataBanks_6_ppn_data_read_1_6_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_6_ppn_MPORT_6_data = io_wdata_ppn;
  assign dataBanks_6_ppn_MPORT_6_addr = io_waddr[0];
  assign dataBanks_6_ppn_MPORT_6_mask = 1'h1;
  assign dataBanks_6_ppn_MPORT_6_en = io_wen & _T_25;
  assign dataBanks_6_perm_pf_data_read_0_6_MPORT_en = 1'h1;
  assign dataBanks_6_perm_pf_data_read_0_6_MPORT_addr = io_raddr_0[0];
  assign dataBanks_6_perm_pf_data_read_0_6_MPORT_data =
    dataBanks_6_perm_pf[dataBanks_6_perm_pf_data_read_0_6_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_6_perm_pf_data_read_1_6_MPORT_en = 1'h1;
  assign dataBanks_6_perm_pf_data_read_1_6_MPORT_addr = io_raddr_0[0];
  assign dataBanks_6_perm_pf_data_read_1_6_MPORT_data =
    dataBanks_6_perm_pf[dataBanks_6_perm_pf_data_read_1_6_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_6_perm_pf_data_read_0_6_MPORT_1_en = 1'h1;
  assign dataBanks_6_perm_pf_data_read_0_6_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_6_perm_pf_data_read_0_6_MPORT_1_data =
    dataBanks_6_perm_pf[dataBanks_6_perm_pf_data_read_0_6_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_6_perm_pf_data_read_1_6_MPORT_1_en = 1'h1;
  assign dataBanks_6_perm_pf_data_read_1_6_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_6_perm_pf_data_read_1_6_MPORT_1_data =
    dataBanks_6_perm_pf[dataBanks_6_perm_pf_data_read_1_6_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_6_perm_pf_MPORT_6_data = io_wdata_perm_pf;
  assign dataBanks_6_perm_pf_MPORT_6_addr = io_waddr[0];
  assign dataBanks_6_perm_pf_MPORT_6_mask = 1'h1;
  assign dataBanks_6_perm_pf_MPORT_6_en = io_wen & _T_25;
  assign dataBanks_6_perm_af_data_read_0_6_MPORT_en = 1'h1;
  assign dataBanks_6_perm_af_data_read_0_6_MPORT_addr = io_raddr_0[0];
  assign dataBanks_6_perm_af_data_read_0_6_MPORT_data =
    dataBanks_6_perm_af[dataBanks_6_perm_af_data_read_0_6_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_6_perm_af_data_read_1_6_MPORT_en = 1'h1;
  assign dataBanks_6_perm_af_data_read_1_6_MPORT_addr = io_raddr_0[0];
  assign dataBanks_6_perm_af_data_read_1_6_MPORT_data =
    dataBanks_6_perm_af[dataBanks_6_perm_af_data_read_1_6_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_6_perm_af_data_read_0_6_MPORT_1_en = 1'h1;
  assign dataBanks_6_perm_af_data_read_0_6_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_6_perm_af_data_read_0_6_MPORT_1_data =
    dataBanks_6_perm_af[dataBanks_6_perm_af_data_read_0_6_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_6_perm_af_data_read_1_6_MPORT_1_en = 1'h1;
  assign dataBanks_6_perm_af_data_read_1_6_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_6_perm_af_data_read_1_6_MPORT_1_data =
    dataBanks_6_perm_af[dataBanks_6_perm_af_data_read_1_6_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_6_perm_af_MPORT_6_data = io_wdata_perm_af;
  assign dataBanks_6_perm_af_MPORT_6_addr = io_waddr[0];
  assign dataBanks_6_perm_af_MPORT_6_mask = 1'h1;
  assign dataBanks_6_perm_af_MPORT_6_en = io_wen & _T_25;
  assign dataBanks_6_perm_d_data_read_0_6_MPORT_en = 1'h1;
  assign dataBanks_6_perm_d_data_read_0_6_MPORT_addr = io_raddr_0[0];
  assign dataBanks_6_perm_d_data_read_0_6_MPORT_data = dataBanks_6_perm_d[dataBanks_6_perm_d_data_read_0_6_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_6_perm_d_data_read_1_6_MPORT_en = 1'h1;
  assign dataBanks_6_perm_d_data_read_1_6_MPORT_addr = io_raddr_0[0];
  assign dataBanks_6_perm_d_data_read_1_6_MPORT_data = dataBanks_6_perm_d[dataBanks_6_perm_d_data_read_1_6_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_6_perm_d_data_read_0_6_MPORT_1_en = 1'h1;
  assign dataBanks_6_perm_d_data_read_0_6_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_6_perm_d_data_read_0_6_MPORT_1_data =
    dataBanks_6_perm_d[dataBanks_6_perm_d_data_read_0_6_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_6_perm_d_data_read_1_6_MPORT_1_en = 1'h1;
  assign dataBanks_6_perm_d_data_read_1_6_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_6_perm_d_data_read_1_6_MPORT_1_data =
    dataBanks_6_perm_d[dataBanks_6_perm_d_data_read_1_6_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_6_perm_d_MPORT_6_data = io_wdata_perm_d;
  assign dataBanks_6_perm_d_MPORT_6_addr = io_waddr[0];
  assign dataBanks_6_perm_d_MPORT_6_mask = 1'h1;
  assign dataBanks_6_perm_d_MPORT_6_en = io_wen & _T_25;
  assign dataBanks_6_perm_a_data_read_0_6_MPORT_en = 1'h1;
  assign dataBanks_6_perm_a_data_read_0_6_MPORT_addr = io_raddr_0[0];
  assign dataBanks_6_perm_a_data_read_0_6_MPORT_data = dataBanks_6_perm_a[dataBanks_6_perm_a_data_read_0_6_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_6_perm_a_data_read_1_6_MPORT_en = 1'h1;
  assign dataBanks_6_perm_a_data_read_1_6_MPORT_addr = io_raddr_0[0];
  assign dataBanks_6_perm_a_data_read_1_6_MPORT_data = dataBanks_6_perm_a[dataBanks_6_perm_a_data_read_1_6_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_6_perm_a_data_read_0_6_MPORT_1_en = 1'h1;
  assign dataBanks_6_perm_a_data_read_0_6_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_6_perm_a_data_read_0_6_MPORT_1_data =
    dataBanks_6_perm_a[dataBanks_6_perm_a_data_read_0_6_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_6_perm_a_data_read_1_6_MPORT_1_en = 1'h1;
  assign dataBanks_6_perm_a_data_read_1_6_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_6_perm_a_data_read_1_6_MPORT_1_data =
    dataBanks_6_perm_a[dataBanks_6_perm_a_data_read_1_6_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_6_perm_a_MPORT_6_data = io_wdata_perm_a;
  assign dataBanks_6_perm_a_MPORT_6_addr = io_waddr[0];
  assign dataBanks_6_perm_a_MPORT_6_mask = 1'h1;
  assign dataBanks_6_perm_a_MPORT_6_en = io_wen & _T_25;
  assign dataBanks_6_perm_u_data_read_0_6_MPORT_en = 1'h1;
  assign dataBanks_6_perm_u_data_read_0_6_MPORT_addr = io_raddr_0[0];
  assign dataBanks_6_perm_u_data_read_0_6_MPORT_data = dataBanks_6_perm_u[dataBanks_6_perm_u_data_read_0_6_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_6_perm_u_data_read_1_6_MPORT_en = 1'h1;
  assign dataBanks_6_perm_u_data_read_1_6_MPORT_addr = io_raddr_0[0];
  assign dataBanks_6_perm_u_data_read_1_6_MPORT_data = dataBanks_6_perm_u[dataBanks_6_perm_u_data_read_1_6_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_6_perm_u_data_read_0_6_MPORT_1_en = 1'h1;
  assign dataBanks_6_perm_u_data_read_0_6_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_6_perm_u_data_read_0_6_MPORT_1_data =
    dataBanks_6_perm_u[dataBanks_6_perm_u_data_read_0_6_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_6_perm_u_data_read_1_6_MPORT_1_en = 1'h1;
  assign dataBanks_6_perm_u_data_read_1_6_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_6_perm_u_data_read_1_6_MPORT_1_data =
    dataBanks_6_perm_u[dataBanks_6_perm_u_data_read_1_6_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_6_perm_u_MPORT_6_data = io_wdata_perm_u;
  assign dataBanks_6_perm_u_MPORT_6_addr = io_waddr[0];
  assign dataBanks_6_perm_u_MPORT_6_mask = 1'h1;
  assign dataBanks_6_perm_u_MPORT_6_en = io_wen & _T_25;
  assign dataBanks_6_perm_x_data_read_0_6_MPORT_en = 1'h1;
  assign dataBanks_6_perm_x_data_read_0_6_MPORT_addr = io_raddr_0[0];
  assign dataBanks_6_perm_x_data_read_0_6_MPORT_data = dataBanks_6_perm_x[dataBanks_6_perm_x_data_read_0_6_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_6_perm_x_data_read_1_6_MPORT_en = 1'h1;
  assign dataBanks_6_perm_x_data_read_1_6_MPORT_addr = io_raddr_0[0];
  assign dataBanks_6_perm_x_data_read_1_6_MPORT_data = dataBanks_6_perm_x[dataBanks_6_perm_x_data_read_1_6_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_6_perm_x_data_read_0_6_MPORT_1_en = 1'h1;
  assign dataBanks_6_perm_x_data_read_0_6_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_6_perm_x_data_read_0_6_MPORT_1_data =
    dataBanks_6_perm_x[dataBanks_6_perm_x_data_read_0_6_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_6_perm_x_data_read_1_6_MPORT_1_en = 1'h1;
  assign dataBanks_6_perm_x_data_read_1_6_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_6_perm_x_data_read_1_6_MPORT_1_data =
    dataBanks_6_perm_x[dataBanks_6_perm_x_data_read_1_6_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_6_perm_x_MPORT_6_data = io_wdata_perm_x;
  assign dataBanks_6_perm_x_MPORT_6_addr = io_waddr[0];
  assign dataBanks_6_perm_x_MPORT_6_mask = 1'h1;
  assign dataBanks_6_perm_x_MPORT_6_en = io_wen & _T_25;
  assign dataBanks_6_perm_wdata_read_0_6_MPORT_en = 1'h1;
  assign dataBanks_6_perm_wdata_read_0_6_MPORT_addr = io_raddr_0[0];
  assign dataBanks_6_perm_wdata_read_0_6_MPORT_data = dataBanks_6_perm_w[dataBanks_6_perm_wdata_read_0_6_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_6_perm_wdata_read_1_6_MPORT_en = 1'h1;
  assign dataBanks_6_perm_wdata_read_1_6_MPORT_addr = io_raddr_0[0];
  assign dataBanks_6_perm_wdata_read_1_6_MPORT_data = dataBanks_6_perm_w[dataBanks_6_perm_wdata_read_1_6_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_6_perm_wdata_read_0_6_MPORT_1_en = 1'h1;
  assign dataBanks_6_perm_wdata_read_0_6_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_6_perm_wdata_read_0_6_MPORT_1_data =
    dataBanks_6_perm_w[dataBanks_6_perm_wdata_read_0_6_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_6_perm_wdata_read_1_6_MPORT_1_en = 1'h1;
  assign dataBanks_6_perm_wdata_read_1_6_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_6_perm_wdata_read_1_6_MPORT_1_data =
    dataBanks_6_perm_w[dataBanks_6_perm_wdata_read_1_6_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_6_perm_wMPORT_6_data = io_wdata_perm_w;
  assign dataBanks_6_perm_wMPORT_6_addr = io_waddr[0];
  assign dataBanks_6_perm_wMPORT_6_mask = 1'h1;
  assign dataBanks_6_perm_wMPORT_6_en = io_wen & _T_25;
  assign dataBanks_6_perm_rdata_read_0_6_MPORT_en = 1'h1;
  assign dataBanks_6_perm_rdata_read_0_6_MPORT_addr = io_raddr_0[0];
  assign dataBanks_6_perm_rdata_read_0_6_MPORT_data = dataBanks_6_perm_r[dataBanks_6_perm_rdata_read_0_6_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_6_perm_rdata_read_1_6_MPORT_en = 1'h1;
  assign dataBanks_6_perm_rdata_read_1_6_MPORT_addr = io_raddr_0[0];
  assign dataBanks_6_perm_rdata_read_1_6_MPORT_data = dataBanks_6_perm_r[dataBanks_6_perm_rdata_read_1_6_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_6_perm_rdata_read_0_6_MPORT_1_en = 1'h1;
  assign dataBanks_6_perm_rdata_read_0_6_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_6_perm_rdata_read_0_6_MPORT_1_data =
    dataBanks_6_perm_r[dataBanks_6_perm_rdata_read_0_6_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_6_perm_rdata_read_1_6_MPORT_1_en = 1'h1;
  assign dataBanks_6_perm_rdata_read_1_6_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_6_perm_rdata_read_1_6_MPORT_1_data =
    dataBanks_6_perm_r[dataBanks_6_perm_rdata_read_1_6_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_6_perm_rMPORT_6_data = io_wdata_perm_r;
  assign dataBanks_6_perm_rMPORT_6_addr = io_waddr[0];
  assign dataBanks_6_perm_rMPORT_6_mask = 1'h1;
  assign dataBanks_6_perm_rMPORT_6_en = io_wen & _T_25;
  assign dataBanks_6_perm_pm_rdata_read_0_6_MPORT_en = 1'h1;
  assign dataBanks_6_perm_pm_rdata_read_0_6_MPORT_addr = io_raddr_0[0];
  assign dataBanks_6_perm_pm_rdata_read_0_6_MPORT_data =
    dataBanks_6_perm_pm_r[dataBanks_6_perm_pm_rdata_read_0_6_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_6_perm_pm_rdata_read_1_6_MPORT_en = 1'h1;
  assign dataBanks_6_perm_pm_rdata_read_1_6_MPORT_addr = io_raddr_0[0];
  assign dataBanks_6_perm_pm_rdata_read_1_6_MPORT_data =
    dataBanks_6_perm_pm_r[dataBanks_6_perm_pm_rdata_read_1_6_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_6_perm_pm_rdata_read_0_6_MPORT_1_en = 1'h1;
  assign dataBanks_6_perm_pm_rdata_read_0_6_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_6_perm_pm_rdata_read_0_6_MPORT_1_data =
    dataBanks_6_perm_pm_r[dataBanks_6_perm_pm_rdata_read_0_6_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_6_perm_pm_rdata_read_1_6_MPORT_1_en = 1'h1;
  assign dataBanks_6_perm_pm_rdata_read_1_6_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_6_perm_pm_rdata_read_1_6_MPORT_1_data =
    dataBanks_6_perm_pm_r[dataBanks_6_perm_pm_rdata_read_1_6_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_6_perm_pm_rMPORT_6_data = io_wdata_perm_pm_r;
  assign dataBanks_6_perm_pm_rMPORT_6_addr = io_waddr[0];
  assign dataBanks_6_perm_pm_rMPORT_6_mask = 1'h1;
  assign dataBanks_6_perm_pm_rMPORT_6_en = io_wen & _T_25;
  assign dataBanks_6_perm_pm_wdata_read_0_6_MPORT_en = 1'h1;
  assign dataBanks_6_perm_pm_wdata_read_0_6_MPORT_addr = io_raddr_0[0];
  assign dataBanks_6_perm_pm_wdata_read_0_6_MPORT_data =
    dataBanks_6_perm_pm_w[dataBanks_6_perm_pm_wdata_read_0_6_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_6_perm_pm_wdata_read_1_6_MPORT_en = 1'h1;
  assign dataBanks_6_perm_pm_wdata_read_1_6_MPORT_addr = io_raddr_0[0];
  assign dataBanks_6_perm_pm_wdata_read_1_6_MPORT_data =
    dataBanks_6_perm_pm_w[dataBanks_6_perm_pm_wdata_read_1_6_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_6_perm_pm_wdata_read_0_6_MPORT_1_en = 1'h1;
  assign dataBanks_6_perm_pm_wdata_read_0_6_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_6_perm_pm_wdata_read_0_6_MPORT_1_data =
    dataBanks_6_perm_pm_w[dataBanks_6_perm_pm_wdata_read_0_6_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_6_perm_pm_wdata_read_1_6_MPORT_1_en = 1'h1;
  assign dataBanks_6_perm_pm_wdata_read_1_6_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_6_perm_pm_wdata_read_1_6_MPORT_1_data =
    dataBanks_6_perm_pm_w[dataBanks_6_perm_pm_wdata_read_1_6_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_6_perm_pm_wMPORT_6_data = io_wdata_perm_pm_w;
  assign dataBanks_6_perm_pm_wMPORT_6_addr = io_waddr[0];
  assign dataBanks_6_perm_pm_wMPORT_6_mask = 1'h1;
  assign dataBanks_6_perm_pm_wMPORT_6_en = io_wen & _T_25;
  assign dataBanks_6_perm_pm_c_data_read_0_6_MPORT_en = 1'h1;
  assign dataBanks_6_perm_pm_c_data_read_0_6_MPORT_addr = io_raddr_0[0];
  assign dataBanks_6_perm_pm_c_data_read_0_6_MPORT_data =
    dataBanks_6_perm_pm_c[dataBanks_6_perm_pm_c_data_read_0_6_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_6_perm_pm_c_data_read_1_6_MPORT_en = 1'h1;
  assign dataBanks_6_perm_pm_c_data_read_1_6_MPORT_addr = io_raddr_0[0];
  assign dataBanks_6_perm_pm_c_data_read_1_6_MPORT_data =
    dataBanks_6_perm_pm_c[dataBanks_6_perm_pm_c_data_read_1_6_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_6_perm_pm_c_data_read_0_6_MPORT_1_en = 1'h1;
  assign dataBanks_6_perm_pm_c_data_read_0_6_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_6_perm_pm_c_data_read_0_6_MPORT_1_data =
    dataBanks_6_perm_pm_c[dataBanks_6_perm_pm_c_data_read_0_6_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_6_perm_pm_c_data_read_1_6_MPORT_1_en = 1'h1;
  assign dataBanks_6_perm_pm_c_data_read_1_6_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_6_perm_pm_c_data_read_1_6_MPORT_1_data =
    dataBanks_6_perm_pm_c[dataBanks_6_perm_pm_c_data_read_1_6_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_6_perm_pm_c_MPORT_6_data = io_wdata_perm_pm_c;
  assign dataBanks_6_perm_pm_c_MPORT_6_addr = io_waddr[0];
  assign dataBanks_6_perm_pm_c_MPORT_6_mask = 1'h1;
  assign dataBanks_6_perm_pm_c_MPORT_6_en = io_wen & _T_25;
  assign dataBanks_7_tag_data_read_0_7_MPORT_en = 1'h1;
  assign dataBanks_7_tag_data_read_0_7_MPORT_addr = io_raddr_0[0];
  assign dataBanks_7_tag_data_read_0_7_MPORT_data = dataBanks_7_tag[dataBanks_7_tag_data_read_0_7_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_7_tag_data_read_1_7_MPORT_en = 1'h1;
  assign dataBanks_7_tag_data_read_1_7_MPORT_addr = io_raddr_0[0];
  assign dataBanks_7_tag_data_read_1_7_MPORT_data = dataBanks_7_tag[dataBanks_7_tag_data_read_1_7_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_7_tag_data_read_0_7_MPORT_1_en = 1'h1;
  assign dataBanks_7_tag_data_read_0_7_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_7_tag_data_read_0_7_MPORT_1_data = dataBanks_7_tag[dataBanks_7_tag_data_read_0_7_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_7_tag_data_read_1_7_MPORT_1_en = 1'h1;
  assign dataBanks_7_tag_data_read_1_7_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_7_tag_data_read_1_7_MPORT_1_data = dataBanks_7_tag[dataBanks_7_tag_data_read_1_7_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_7_tag_MPORT_7_data = io_wdata_tag;
  assign dataBanks_7_tag_MPORT_7_addr = io_waddr[0];
  assign dataBanks_7_tag_MPORT_7_mask = 1'h1;
  assign dataBanks_7_tag_MPORT_7_en = io_wen & _T_29;
  assign dataBanks_7_asid_data_read_0_7_MPORT_en = 1'h1;
  assign dataBanks_7_asid_data_read_0_7_MPORT_addr = io_raddr_0[0];
  assign dataBanks_7_asid_data_read_0_7_MPORT_data = dataBanks_7_asid[dataBanks_7_asid_data_read_0_7_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_7_asid_data_read_1_7_MPORT_en = 1'h1;
  assign dataBanks_7_asid_data_read_1_7_MPORT_addr = io_raddr_0[0];
  assign dataBanks_7_asid_data_read_1_7_MPORT_data = dataBanks_7_asid[dataBanks_7_asid_data_read_1_7_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_7_asid_data_read_0_7_MPORT_1_en = 1'h1;
  assign dataBanks_7_asid_data_read_0_7_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_7_asid_data_read_0_7_MPORT_1_data = dataBanks_7_asid[dataBanks_7_asid_data_read_0_7_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_7_asid_data_read_1_7_MPORT_1_en = 1'h1;
  assign dataBanks_7_asid_data_read_1_7_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_7_asid_data_read_1_7_MPORT_1_data = dataBanks_7_asid[dataBanks_7_asid_data_read_1_7_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_7_asid_MPORT_7_data = io_wdata_asid;
  assign dataBanks_7_asid_MPORT_7_addr = io_waddr[0];
  assign dataBanks_7_asid_MPORT_7_mask = 1'h1;
  assign dataBanks_7_asid_MPORT_7_en = io_wen & _T_29;
  assign dataBanks_7_ppn_data_read_0_7_MPORT_en = 1'h1;
  assign dataBanks_7_ppn_data_read_0_7_MPORT_addr = io_raddr_0[0];
  assign dataBanks_7_ppn_data_read_0_7_MPORT_data = dataBanks_7_ppn[dataBanks_7_ppn_data_read_0_7_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_7_ppn_data_read_1_7_MPORT_en = 1'h1;
  assign dataBanks_7_ppn_data_read_1_7_MPORT_addr = io_raddr_0[0];
  assign dataBanks_7_ppn_data_read_1_7_MPORT_data = dataBanks_7_ppn[dataBanks_7_ppn_data_read_1_7_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_7_ppn_data_read_0_7_MPORT_1_en = 1'h1;
  assign dataBanks_7_ppn_data_read_0_7_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_7_ppn_data_read_0_7_MPORT_1_data = dataBanks_7_ppn[dataBanks_7_ppn_data_read_0_7_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_7_ppn_data_read_1_7_MPORT_1_en = 1'h1;
  assign dataBanks_7_ppn_data_read_1_7_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_7_ppn_data_read_1_7_MPORT_1_data = dataBanks_7_ppn[dataBanks_7_ppn_data_read_1_7_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_7_ppn_MPORT_7_data = io_wdata_ppn;
  assign dataBanks_7_ppn_MPORT_7_addr = io_waddr[0];
  assign dataBanks_7_ppn_MPORT_7_mask = 1'h1;
  assign dataBanks_7_ppn_MPORT_7_en = io_wen & _T_29;
  assign dataBanks_7_perm_pf_data_read_0_7_MPORT_en = 1'h1;
  assign dataBanks_7_perm_pf_data_read_0_7_MPORT_addr = io_raddr_0[0];
  assign dataBanks_7_perm_pf_data_read_0_7_MPORT_data =
    dataBanks_7_perm_pf[dataBanks_7_perm_pf_data_read_0_7_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_7_perm_pf_data_read_1_7_MPORT_en = 1'h1;
  assign dataBanks_7_perm_pf_data_read_1_7_MPORT_addr = io_raddr_0[0];
  assign dataBanks_7_perm_pf_data_read_1_7_MPORT_data =
    dataBanks_7_perm_pf[dataBanks_7_perm_pf_data_read_1_7_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_7_perm_pf_data_read_0_7_MPORT_1_en = 1'h1;
  assign dataBanks_7_perm_pf_data_read_0_7_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_7_perm_pf_data_read_0_7_MPORT_1_data =
    dataBanks_7_perm_pf[dataBanks_7_perm_pf_data_read_0_7_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_7_perm_pf_data_read_1_7_MPORT_1_en = 1'h1;
  assign dataBanks_7_perm_pf_data_read_1_7_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_7_perm_pf_data_read_1_7_MPORT_1_data =
    dataBanks_7_perm_pf[dataBanks_7_perm_pf_data_read_1_7_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_7_perm_pf_MPORT_7_data = io_wdata_perm_pf;
  assign dataBanks_7_perm_pf_MPORT_7_addr = io_waddr[0];
  assign dataBanks_7_perm_pf_MPORT_7_mask = 1'h1;
  assign dataBanks_7_perm_pf_MPORT_7_en = io_wen & _T_29;
  assign dataBanks_7_perm_af_data_read_0_7_MPORT_en = 1'h1;
  assign dataBanks_7_perm_af_data_read_0_7_MPORT_addr = io_raddr_0[0];
  assign dataBanks_7_perm_af_data_read_0_7_MPORT_data =
    dataBanks_7_perm_af[dataBanks_7_perm_af_data_read_0_7_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_7_perm_af_data_read_1_7_MPORT_en = 1'h1;
  assign dataBanks_7_perm_af_data_read_1_7_MPORT_addr = io_raddr_0[0];
  assign dataBanks_7_perm_af_data_read_1_7_MPORT_data =
    dataBanks_7_perm_af[dataBanks_7_perm_af_data_read_1_7_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_7_perm_af_data_read_0_7_MPORT_1_en = 1'h1;
  assign dataBanks_7_perm_af_data_read_0_7_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_7_perm_af_data_read_0_7_MPORT_1_data =
    dataBanks_7_perm_af[dataBanks_7_perm_af_data_read_0_7_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_7_perm_af_data_read_1_7_MPORT_1_en = 1'h1;
  assign dataBanks_7_perm_af_data_read_1_7_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_7_perm_af_data_read_1_7_MPORT_1_data =
    dataBanks_7_perm_af[dataBanks_7_perm_af_data_read_1_7_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_7_perm_af_MPORT_7_data = io_wdata_perm_af;
  assign dataBanks_7_perm_af_MPORT_7_addr = io_waddr[0];
  assign dataBanks_7_perm_af_MPORT_7_mask = 1'h1;
  assign dataBanks_7_perm_af_MPORT_7_en = io_wen & _T_29;
  assign dataBanks_7_perm_d_data_read_0_7_MPORT_en = 1'h1;
  assign dataBanks_7_perm_d_data_read_0_7_MPORT_addr = io_raddr_0[0];
  assign dataBanks_7_perm_d_data_read_0_7_MPORT_data = dataBanks_7_perm_d[dataBanks_7_perm_d_data_read_0_7_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_7_perm_d_data_read_1_7_MPORT_en = 1'h1;
  assign dataBanks_7_perm_d_data_read_1_7_MPORT_addr = io_raddr_0[0];
  assign dataBanks_7_perm_d_data_read_1_7_MPORT_data = dataBanks_7_perm_d[dataBanks_7_perm_d_data_read_1_7_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_7_perm_d_data_read_0_7_MPORT_1_en = 1'h1;
  assign dataBanks_7_perm_d_data_read_0_7_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_7_perm_d_data_read_0_7_MPORT_1_data =
    dataBanks_7_perm_d[dataBanks_7_perm_d_data_read_0_7_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_7_perm_d_data_read_1_7_MPORT_1_en = 1'h1;
  assign dataBanks_7_perm_d_data_read_1_7_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_7_perm_d_data_read_1_7_MPORT_1_data =
    dataBanks_7_perm_d[dataBanks_7_perm_d_data_read_1_7_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_7_perm_d_MPORT_7_data = io_wdata_perm_d;
  assign dataBanks_7_perm_d_MPORT_7_addr = io_waddr[0];
  assign dataBanks_7_perm_d_MPORT_7_mask = 1'h1;
  assign dataBanks_7_perm_d_MPORT_7_en = io_wen & _T_29;
  assign dataBanks_7_perm_a_data_read_0_7_MPORT_en = 1'h1;
  assign dataBanks_7_perm_a_data_read_0_7_MPORT_addr = io_raddr_0[0];
  assign dataBanks_7_perm_a_data_read_0_7_MPORT_data = dataBanks_7_perm_a[dataBanks_7_perm_a_data_read_0_7_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_7_perm_a_data_read_1_7_MPORT_en = 1'h1;
  assign dataBanks_7_perm_a_data_read_1_7_MPORT_addr = io_raddr_0[0];
  assign dataBanks_7_perm_a_data_read_1_7_MPORT_data = dataBanks_7_perm_a[dataBanks_7_perm_a_data_read_1_7_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_7_perm_a_data_read_0_7_MPORT_1_en = 1'h1;
  assign dataBanks_7_perm_a_data_read_0_7_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_7_perm_a_data_read_0_7_MPORT_1_data =
    dataBanks_7_perm_a[dataBanks_7_perm_a_data_read_0_7_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_7_perm_a_data_read_1_7_MPORT_1_en = 1'h1;
  assign dataBanks_7_perm_a_data_read_1_7_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_7_perm_a_data_read_1_7_MPORT_1_data =
    dataBanks_7_perm_a[dataBanks_7_perm_a_data_read_1_7_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_7_perm_a_MPORT_7_data = io_wdata_perm_a;
  assign dataBanks_7_perm_a_MPORT_7_addr = io_waddr[0];
  assign dataBanks_7_perm_a_MPORT_7_mask = 1'h1;
  assign dataBanks_7_perm_a_MPORT_7_en = io_wen & _T_29;
  assign dataBanks_7_perm_u_data_read_0_7_MPORT_en = 1'h1;
  assign dataBanks_7_perm_u_data_read_0_7_MPORT_addr = io_raddr_0[0];
  assign dataBanks_7_perm_u_data_read_0_7_MPORT_data = dataBanks_7_perm_u[dataBanks_7_perm_u_data_read_0_7_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_7_perm_u_data_read_1_7_MPORT_en = 1'h1;
  assign dataBanks_7_perm_u_data_read_1_7_MPORT_addr = io_raddr_0[0];
  assign dataBanks_7_perm_u_data_read_1_7_MPORT_data = dataBanks_7_perm_u[dataBanks_7_perm_u_data_read_1_7_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_7_perm_u_data_read_0_7_MPORT_1_en = 1'h1;
  assign dataBanks_7_perm_u_data_read_0_7_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_7_perm_u_data_read_0_7_MPORT_1_data =
    dataBanks_7_perm_u[dataBanks_7_perm_u_data_read_0_7_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_7_perm_u_data_read_1_7_MPORT_1_en = 1'h1;
  assign dataBanks_7_perm_u_data_read_1_7_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_7_perm_u_data_read_1_7_MPORT_1_data =
    dataBanks_7_perm_u[dataBanks_7_perm_u_data_read_1_7_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_7_perm_u_MPORT_7_data = io_wdata_perm_u;
  assign dataBanks_7_perm_u_MPORT_7_addr = io_waddr[0];
  assign dataBanks_7_perm_u_MPORT_7_mask = 1'h1;
  assign dataBanks_7_perm_u_MPORT_7_en = io_wen & _T_29;
  assign dataBanks_7_perm_x_data_read_0_7_MPORT_en = 1'h1;
  assign dataBanks_7_perm_x_data_read_0_7_MPORT_addr = io_raddr_0[0];
  assign dataBanks_7_perm_x_data_read_0_7_MPORT_data = dataBanks_7_perm_x[dataBanks_7_perm_x_data_read_0_7_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_7_perm_x_data_read_1_7_MPORT_en = 1'h1;
  assign dataBanks_7_perm_x_data_read_1_7_MPORT_addr = io_raddr_0[0];
  assign dataBanks_7_perm_x_data_read_1_7_MPORT_data = dataBanks_7_perm_x[dataBanks_7_perm_x_data_read_1_7_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_7_perm_x_data_read_0_7_MPORT_1_en = 1'h1;
  assign dataBanks_7_perm_x_data_read_0_7_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_7_perm_x_data_read_0_7_MPORT_1_data =
    dataBanks_7_perm_x[dataBanks_7_perm_x_data_read_0_7_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_7_perm_x_data_read_1_7_MPORT_1_en = 1'h1;
  assign dataBanks_7_perm_x_data_read_1_7_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_7_perm_x_data_read_1_7_MPORT_1_data =
    dataBanks_7_perm_x[dataBanks_7_perm_x_data_read_1_7_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_7_perm_x_MPORT_7_data = io_wdata_perm_x;
  assign dataBanks_7_perm_x_MPORT_7_addr = io_waddr[0];
  assign dataBanks_7_perm_x_MPORT_7_mask = 1'h1;
  assign dataBanks_7_perm_x_MPORT_7_en = io_wen & _T_29;
  assign dataBanks_7_perm_wdata_read_0_7_MPORT_en = 1'h1;
  assign dataBanks_7_perm_wdata_read_0_7_MPORT_addr = io_raddr_0[0];
  assign dataBanks_7_perm_wdata_read_0_7_MPORT_data = dataBanks_7_perm_w[dataBanks_7_perm_wdata_read_0_7_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_7_perm_wdata_read_1_7_MPORT_en = 1'h1;
  assign dataBanks_7_perm_wdata_read_1_7_MPORT_addr = io_raddr_0[0];
  assign dataBanks_7_perm_wdata_read_1_7_MPORT_data = dataBanks_7_perm_w[dataBanks_7_perm_wdata_read_1_7_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_7_perm_wdata_read_0_7_MPORT_1_en = 1'h1;
  assign dataBanks_7_perm_wdata_read_0_7_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_7_perm_wdata_read_0_7_MPORT_1_data =
    dataBanks_7_perm_w[dataBanks_7_perm_wdata_read_0_7_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_7_perm_wdata_read_1_7_MPORT_1_en = 1'h1;
  assign dataBanks_7_perm_wdata_read_1_7_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_7_perm_wdata_read_1_7_MPORT_1_data =
    dataBanks_7_perm_w[dataBanks_7_perm_wdata_read_1_7_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_7_perm_wMPORT_7_data = io_wdata_perm_w;
  assign dataBanks_7_perm_wMPORT_7_addr = io_waddr[0];
  assign dataBanks_7_perm_wMPORT_7_mask = 1'h1;
  assign dataBanks_7_perm_wMPORT_7_en = io_wen & _T_29;
  assign dataBanks_7_perm_rdata_read_0_7_MPORT_en = 1'h1;
  assign dataBanks_7_perm_rdata_read_0_7_MPORT_addr = io_raddr_0[0];
  assign dataBanks_7_perm_rdata_read_0_7_MPORT_data = dataBanks_7_perm_r[dataBanks_7_perm_rdata_read_0_7_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_7_perm_rdata_read_1_7_MPORT_en = 1'h1;
  assign dataBanks_7_perm_rdata_read_1_7_MPORT_addr = io_raddr_0[0];
  assign dataBanks_7_perm_rdata_read_1_7_MPORT_data = dataBanks_7_perm_r[dataBanks_7_perm_rdata_read_1_7_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_7_perm_rdata_read_0_7_MPORT_1_en = 1'h1;
  assign dataBanks_7_perm_rdata_read_0_7_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_7_perm_rdata_read_0_7_MPORT_1_data =
    dataBanks_7_perm_r[dataBanks_7_perm_rdata_read_0_7_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_7_perm_rdata_read_1_7_MPORT_1_en = 1'h1;
  assign dataBanks_7_perm_rdata_read_1_7_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_7_perm_rdata_read_1_7_MPORT_1_data =
    dataBanks_7_perm_r[dataBanks_7_perm_rdata_read_1_7_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_7_perm_rMPORT_7_data = io_wdata_perm_r;
  assign dataBanks_7_perm_rMPORT_7_addr = io_waddr[0];
  assign dataBanks_7_perm_rMPORT_7_mask = 1'h1;
  assign dataBanks_7_perm_rMPORT_7_en = io_wen & _T_29;
  assign dataBanks_7_perm_pm_rdata_read_0_7_MPORT_en = 1'h1;
  assign dataBanks_7_perm_pm_rdata_read_0_7_MPORT_addr = io_raddr_0[0];
  assign dataBanks_7_perm_pm_rdata_read_0_7_MPORT_data =
    dataBanks_7_perm_pm_r[dataBanks_7_perm_pm_rdata_read_0_7_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_7_perm_pm_rdata_read_1_7_MPORT_en = 1'h1;
  assign dataBanks_7_perm_pm_rdata_read_1_7_MPORT_addr = io_raddr_0[0];
  assign dataBanks_7_perm_pm_rdata_read_1_7_MPORT_data =
    dataBanks_7_perm_pm_r[dataBanks_7_perm_pm_rdata_read_1_7_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_7_perm_pm_rdata_read_0_7_MPORT_1_en = 1'h1;
  assign dataBanks_7_perm_pm_rdata_read_0_7_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_7_perm_pm_rdata_read_0_7_MPORT_1_data =
    dataBanks_7_perm_pm_r[dataBanks_7_perm_pm_rdata_read_0_7_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_7_perm_pm_rdata_read_1_7_MPORT_1_en = 1'h1;
  assign dataBanks_7_perm_pm_rdata_read_1_7_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_7_perm_pm_rdata_read_1_7_MPORT_1_data =
    dataBanks_7_perm_pm_r[dataBanks_7_perm_pm_rdata_read_1_7_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_7_perm_pm_rMPORT_7_data = io_wdata_perm_pm_r;
  assign dataBanks_7_perm_pm_rMPORT_7_addr = io_waddr[0];
  assign dataBanks_7_perm_pm_rMPORT_7_mask = 1'h1;
  assign dataBanks_7_perm_pm_rMPORT_7_en = io_wen & _T_29;
  assign dataBanks_7_perm_pm_wdata_read_0_7_MPORT_en = 1'h1;
  assign dataBanks_7_perm_pm_wdata_read_0_7_MPORT_addr = io_raddr_0[0];
  assign dataBanks_7_perm_pm_wdata_read_0_7_MPORT_data =
    dataBanks_7_perm_pm_w[dataBanks_7_perm_pm_wdata_read_0_7_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_7_perm_pm_wdata_read_1_7_MPORT_en = 1'h1;
  assign dataBanks_7_perm_pm_wdata_read_1_7_MPORT_addr = io_raddr_0[0];
  assign dataBanks_7_perm_pm_wdata_read_1_7_MPORT_data =
    dataBanks_7_perm_pm_w[dataBanks_7_perm_pm_wdata_read_1_7_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_7_perm_pm_wdata_read_0_7_MPORT_1_en = 1'h1;
  assign dataBanks_7_perm_pm_wdata_read_0_7_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_7_perm_pm_wdata_read_0_7_MPORT_1_data =
    dataBanks_7_perm_pm_w[dataBanks_7_perm_pm_wdata_read_0_7_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_7_perm_pm_wdata_read_1_7_MPORT_1_en = 1'h1;
  assign dataBanks_7_perm_pm_wdata_read_1_7_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_7_perm_pm_wdata_read_1_7_MPORT_1_data =
    dataBanks_7_perm_pm_w[dataBanks_7_perm_pm_wdata_read_1_7_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_7_perm_pm_wMPORT_7_data = io_wdata_perm_pm_w;
  assign dataBanks_7_perm_pm_wMPORT_7_addr = io_waddr[0];
  assign dataBanks_7_perm_pm_wMPORT_7_mask = 1'h1;
  assign dataBanks_7_perm_pm_wMPORT_7_en = io_wen & _T_29;
  assign dataBanks_7_perm_pm_c_data_read_0_7_MPORT_en = 1'h1;
  assign dataBanks_7_perm_pm_c_data_read_0_7_MPORT_addr = io_raddr_0[0];
  assign dataBanks_7_perm_pm_c_data_read_0_7_MPORT_data =
    dataBanks_7_perm_pm_c[dataBanks_7_perm_pm_c_data_read_0_7_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_7_perm_pm_c_data_read_1_7_MPORT_en = 1'h1;
  assign dataBanks_7_perm_pm_c_data_read_1_7_MPORT_addr = io_raddr_0[0];
  assign dataBanks_7_perm_pm_c_data_read_1_7_MPORT_data =
    dataBanks_7_perm_pm_c[dataBanks_7_perm_pm_c_data_read_1_7_MPORT_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_7_perm_pm_c_data_read_0_7_MPORT_1_en = 1'h1;
  assign dataBanks_7_perm_pm_c_data_read_0_7_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_7_perm_pm_c_data_read_0_7_MPORT_1_data =
    dataBanks_7_perm_pm_c[dataBanks_7_perm_pm_c_data_read_0_7_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_7_perm_pm_c_data_read_1_7_MPORT_1_en = 1'h1;
  assign dataBanks_7_perm_pm_c_data_read_1_7_MPORT_1_addr = io_raddr_1[0];
  assign dataBanks_7_perm_pm_c_data_read_1_7_MPORT_1_data =
    dataBanks_7_perm_pm_c[dataBanks_7_perm_pm_c_data_read_1_7_MPORT_1_addr]; // @[TLBStorage.scala 58:8]
  assign dataBanks_7_perm_pm_c_MPORT_7_data = io_wdata_perm_pm_c;
  assign dataBanks_7_perm_pm_c_MPORT_7_addr = io_waddr[0];
  assign dataBanks_7_perm_pm_c_MPORT_7_mask = 1'h1;
  assign dataBanks_7_perm_pm_c_MPORT_7_en = io_wen & _T_29;
  assign io_rdata_0_0_tag = _io_rdata_0_0_T_261 | _io_rdata_0_0_T_255; // @[Mux.scala 27:73]
  assign io_rdata_0_0_asid = _io_rdata_0_0_T_246 | _io_rdata_0_0_T_240; // @[Mux.scala 27:73]
  assign io_rdata_0_0_ppn = _io_rdata_0_0_T_231 | _io_rdata_0_0_T_225; // @[Mux.scala 27:73]
  assign io_rdata_0_0_perm_pf = bank_index__0[0] & data_read__0_0_perm_pf | bank_index__0[1] & data_read__0_1_perm_pf |
    bank_index__0[2] & data_read__0_2_perm_pf | bank_index__0[3] & data_read__0_3_perm_pf | bank_index__0[4] &
    data_read__0_4_perm_pf | bank_index__0[5] & data_read__0_5_perm_pf | bank_index__0[6] & data_read__0_6_perm_pf |
    bank_index__0[7] & data_read__0_7_perm_pf; // @[Mux.scala 27:73]
  assign io_rdata_0_0_perm_af = bank_index__0[0] & data_read__0_0_perm_af | bank_index__0[1] & data_read__0_1_perm_af |
    bank_index__0[2] & data_read__0_2_perm_af | bank_index__0[3] & data_read__0_3_perm_af | bank_index__0[4] &
    data_read__0_4_perm_af | bank_index__0[5] & data_read__0_5_perm_af | bank_index__0[6] & data_read__0_6_perm_af |
    bank_index__0[7] & data_read__0_7_perm_af; // @[Mux.scala 27:73]
  assign io_rdata_0_0_perm_d = bank_index__0[0] & data_read__0_0_perm_d | bank_index__0[1] & data_read__0_1_perm_d |
    bank_index__0[2] & data_read__0_2_perm_d | bank_index__0[3] & data_read__0_3_perm_d | bank_index__0[4] &
    data_read__0_4_perm_d | bank_index__0[5] & data_read__0_5_perm_d | bank_index__0[6] & data_read__0_6_perm_d |
    bank_index__0[7] & data_read__0_7_perm_d; // @[Mux.scala 27:73]
  assign io_rdata_0_0_perm_a = bank_index__0[0] & data_read__0_0_perm_a | bank_index__0[1] & data_read__0_1_perm_a |
    bank_index__0[2] & data_read__0_2_perm_a | bank_index__0[3] & data_read__0_3_perm_a | bank_index__0[4] &
    data_read__0_4_perm_a | bank_index__0[5] & data_read__0_5_perm_a | bank_index__0[6] & data_read__0_6_perm_a |
    bank_index__0[7] & data_read__0_7_perm_a; // @[Mux.scala 27:73]
  assign io_rdata_0_0_perm_u = bank_index__0[0] & data_read__0_0_perm_u | bank_index__0[1] & data_read__0_1_perm_u |
    bank_index__0[2] & data_read__0_2_perm_u | bank_index__0[3] & data_read__0_3_perm_u | bank_index__0[4] &
    data_read__0_4_perm_u | bank_index__0[5] & data_read__0_5_perm_u | bank_index__0[6] & data_read__0_6_perm_u |
    bank_index__0[7] & data_read__0_7_perm_u; // @[Mux.scala 27:73]
  assign io_rdata_0_0_perm_x = bank_index__0[0] & data_read__0_0_perm_x | bank_index__0[1] & data_read__0_1_perm_x |
    bank_index__0[2] & data_read__0_2_perm_x | bank_index__0[3] & data_read__0_3_perm_x | bank_index__0[4] &
    data_read__0_4_perm_x | bank_index__0[5] & data_read__0_5_perm_x | bank_index__0[6] & data_read__0_6_perm_x |
    bank_index__0[7] & data_read__0_7_perm_x; // @[Mux.scala 27:73]
  assign io_rdata_0_0_perm_w = bank_index__0[0] & data_read__0_0_perm_w | bank_index__0[1] & data_read__0_1_perm_w |
    bank_index__0[2] & data_read__0_2_perm_w | bank_index__0[3] & data_read__0_3_perm_w | bank_index__0[4] &
    data_read__0_4_perm_w | bank_index__0[5] & data_read__0_5_perm_w | bank_index__0[6] & data_read__0_6_perm_w |
    bank_index__0[7] & data_read__0_7_perm_w; // @[Mux.scala 27:73]
  assign io_rdata_0_0_perm_r = bank_index__0[0] & data_read__0_0_perm_r | bank_index__0[1] & data_read__0_1_perm_r |
    bank_index__0[2] & data_read__0_2_perm_r | bank_index__0[3] & data_read__0_3_perm_r | bank_index__0[4] &
    data_read__0_4_perm_r | bank_index__0[5] & data_read__0_5_perm_r | bank_index__0[6] & data_read__0_6_perm_r |
    bank_index__0[7] & data_read__0_7_perm_r; // @[Mux.scala 27:73]
  assign io_rdata_0_0_perm_pm_r = bank_index__0[0] & data_read__0_0_perm_pm_r | bank_index__0[1] &
    data_read__0_1_perm_pm_r | bank_index__0[2] & data_read__0_2_perm_pm_r | bank_index__0[3] & data_read__0_3_perm_pm_r
     | bank_index__0[4] & data_read__0_4_perm_pm_r | bank_index__0[5] & data_read__0_5_perm_pm_r | bank_index__0[6] &
    data_read__0_6_perm_pm_r | bank_index__0[7] & data_read__0_7_perm_pm_r; // @[Mux.scala 27:73]
  assign io_rdata_0_0_perm_pm_w = bank_index__0[0] & data_read__0_0_perm_pm_w | bank_index__0[1] &
    data_read__0_1_perm_pm_w | bank_index__0[2] & data_read__0_2_perm_pm_w | bank_index__0[3] & data_read__0_3_perm_pm_w
     | bank_index__0[4] & data_read__0_4_perm_pm_w | bank_index__0[5] & data_read__0_5_perm_pm_w | bank_index__0[6] &
    data_read__0_6_perm_pm_w | bank_index__0[7] & data_read__0_7_perm_pm_w; // @[Mux.scala 27:73]
  assign io_rdata_0_0_perm_pm_c = bank_index__0[0] & data_read__0_0_perm_pm_c | bank_index__0[1] &
    data_read__0_1_perm_pm_c | bank_index__0[2] & data_read__0_2_perm_pm_c | bank_index__0[3] & data_read__0_3_perm_pm_c
     | bank_index__0[4] & data_read__0_4_perm_pm_c | bank_index__0[5] & data_read__0_5_perm_pm_c | bank_index__0[6] &
    data_read__0_6_perm_pm_c | bank_index__0[7] & data_read__0_7_perm_pm_c; // @[Mux.scala 27:73]
  assign io_rdata_0_1_ppn = _io_rdata_0_1_T_231 | _io_rdata_0_1_T_225; // @[Mux.scala 27:73]
  assign io_rdata_1_0_tag = _io_rdata_1_0_T_261 | _io_rdata_1_0_T_255; // @[Mux.scala 27:73]
  assign io_rdata_1_0_asid = _io_rdata_1_0_T_246 | _io_rdata_1_0_T_240; // @[Mux.scala 27:73]
  assign io_rdata_1_0_ppn = _io_rdata_1_0_T_231 | _io_rdata_1_0_T_225; // @[Mux.scala 27:73]
  assign io_rdata_1_0_perm_pf = bank_index_1_0[0] & data_read_1_0_0_perm_pf | bank_index_1_0[1] &
    data_read_1_0_1_perm_pf | bank_index_1_0[2] & data_read_1_0_2_perm_pf | bank_index_1_0[3] & data_read_1_0_3_perm_pf
     | bank_index_1_0[4] & data_read_1_0_4_perm_pf | bank_index_1_0[5] & data_read_1_0_5_perm_pf | bank_index_1_0[6] &
    data_read_1_0_6_perm_pf | bank_index_1_0[7] & data_read_1_0_7_perm_pf; // @[Mux.scala 27:73]
  assign io_rdata_1_0_perm_af = bank_index_1_0[0] & data_read_1_0_0_perm_af | bank_index_1_0[1] &
    data_read_1_0_1_perm_af | bank_index_1_0[2] & data_read_1_0_2_perm_af | bank_index_1_0[3] & data_read_1_0_3_perm_af
     | bank_index_1_0[4] & data_read_1_0_4_perm_af | bank_index_1_0[5] & data_read_1_0_5_perm_af | bank_index_1_0[6] &
    data_read_1_0_6_perm_af | bank_index_1_0[7] & data_read_1_0_7_perm_af; // @[Mux.scala 27:73]
  assign io_rdata_1_0_perm_a = bank_index_1_0[0] & data_read_1_0_0_perm_a | bank_index_1_0[1] & data_read_1_0_1_perm_a
     | bank_index_1_0[2] & data_read_1_0_2_perm_a | bank_index_1_0[3] & data_read_1_0_3_perm_a | bank_index_1_0[4] &
    data_read_1_0_4_perm_a | bank_index_1_0[5] & data_read_1_0_5_perm_a | bank_index_1_0[6] & data_read_1_0_6_perm_a |
    bank_index_1_0[7] & data_read_1_0_7_perm_a; // @[Mux.scala 27:73]
  assign io_rdata_1_0_perm_u = bank_index_1_0[0] & data_read_1_0_0_perm_u | bank_index_1_0[1] & data_read_1_0_1_perm_u
     | bank_index_1_0[2] & data_read_1_0_2_perm_u | bank_index_1_0[3] & data_read_1_0_3_perm_u | bank_index_1_0[4] &
    data_read_1_0_4_perm_u | bank_index_1_0[5] & data_read_1_0_5_perm_u | bank_index_1_0[6] & data_read_1_0_6_perm_u |
    bank_index_1_0[7] & data_read_1_0_7_perm_u; // @[Mux.scala 27:73]
  assign io_rdata_1_0_perm_x = bank_index_1_0[0] & data_read_1_0_0_perm_x | bank_index_1_0[1] & data_read_1_0_1_perm_x
     | bank_index_1_0[2] & data_read_1_0_2_perm_x | bank_index_1_0[3] & data_read_1_0_3_perm_x | bank_index_1_0[4] &
    data_read_1_0_4_perm_x | bank_index_1_0[5] & data_read_1_0_5_perm_x | bank_index_1_0[6] & data_read_1_0_6_perm_x |
    bank_index_1_0[7] & data_read_1_0_7_perm_x; // @[Mux.scala 27:73]
  assign io_rdata_1_0_perm_r = bank_index_1_0[0] & data_read_1_0_0_perm_r | bank_index_1_0[1] & data_read_1_0_1_perm_r
     | bank_index_1_0[2] & data_read_1_0_2_perm_r | bank_index_1_0[3] & data_read_1_0_3_perm_r | bank_index_1_0[4] &
    data_read_1_0_4_perm_r | bank_index_1_0[5] & data_read_1_0_5_perm_r | bank_index_1_0[6] & data_read_1_0_6_perm_r |
    bank_index_1_0[7] & data_read_1_0_7_perm_r; // @[Mux.scala 27:73]
  assign io_rdata_1_0_perm_pm_r = bank_index_1_0[0] & data_read_1_0_0_perm_pm_r | bank_index_1_0[1] &
    data_read_1_0_1_perm_pm_r | bank_index_1_0[2] & data_read_1_0_2_perm_pm_r | bank_index_1_0[3] &
    data_read_1_0_3_perm_pm_r | bank_index_1_0[4] & data_read_1_0_4_perm_pm_r | bank_index_1_0[5] &
    data_read_1_0_5_perm_pm_r | bank_index_1_0[6] & data_read_1_0_6_perm_pm_r | bank_index_1_0[7] &
    data_read_1_0_7_perm_pm_r; // @[Mux.scala 27:73]
  assign io_rdata_1_0_perm_pm_c = bank_index_1_0[0] & data_read_1_0_0_perm_pm_c | bank_index_1_0[1] &
    data_read_1_0_1_perm_pm_c | bank_index_1_0[2] & data_read_1_0_2_perm_pm_c | bank_index_1_0[3] &
    data_read_1_0_3_perm_pm_c | bank_index_1_0[4] & data_read_1_0_4_perm_pm_c | bank_index_1_0[5] &
    data_read_1_0_5_perm_pm_c | bank_index_1_0[6] & data_read_1_0_6_perm_pm_c | bank_index_1_0[7] &
    data_read_1_0_7_perm_pm_c; // @[Mux.scala 27:73]
  assign io_rdata_1_1_ppn = _io_rdata_1_1_T_231 | _io_rdata_1_1_T_225; // @[Mux.scala 27:73]
  always @(posedge clock) begin
    if (dataBanks_0_tag_MPORT_en & dataBanks_0_tag_MPORT_mask) begin
      dataBanks_0_tag[dataBanks_0_tag_MPORT_addr] <= dataBanks_0_tag_MPORT_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_0_asid_MPORT_en & dataBanks_0_asid_MPORT_mask) begin
      dataBanks_0_asid[dataBanks_0_asid_MPORT_addr] <= dataBanks_0_asid_MPORT_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_0_ppn_MPORT_en & dataBanks_0_ppn_MPORT_mask) begin
      dataBanks_0_ppn[dataBanks_0_ppn_MPORT_addr] <= dataBanks_0_ppn_MPORT_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_0_perm_pf_MPORT_en & dataBanks_0_perm_pf_MPORT_mask) begin
      dataBanks_0_perm_pf[dataBanks_0_perm_pf_MPORT_addr] <= dataBanks_0_perm_pf_MPORT_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_0_perm_af_MPORT_en & dataBanks_0_perm_af_MPORT_mask) begin
      dataBanks_0_perm_af[dataBanks_0_perm_af_MPORT_addr] <= dataBanks_0_perm_af_MPORT_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_0_perm_d_MPORT_en & dataBanks_0_perm_d_MPORT_mask) begin
      dataBanks_0_perm_d[dataBanks_0_perm_d_MPORT_addr] <= dataBanks_0_perm_d_MPORT_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_0_perm_a_MPORT_en & dataBanks_0_perm_a_MPORT_mask) begin
      dataBanks_0_perm_a[dataBanks_0_perm_a_MPORT_addr] <= dataBanks_0_perm_a_MPORT_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_0_perm_u_MPORT_en & dataBanks_0_perm_u_MPORT_mask) begin
      dataBanks_0_perm_u[dataBanks_0_perm_u_MPORT_addr] <= dataBanks_0_perm_u_MPORT_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_0_perm_x_MPORT_en & dataBanks_0_perm_x_MPORT_mask) begin
      dataBanks_0_perm_x[dataBanks_0_perm_x_MPORT_addr] <= dataBanks_0_perm_x_MPORT_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_0_perm_wMPORT_en & dataBanks_0_perm_wMPORT_mask) begin
      dataBanks_0_perm_w[dataBanks_0_perm_wMPORT_addr] <= dataBanks_0_perm_wMPORT_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_0_perm_rMPORT_en & dataBanks_0_perm_rMPORT_mask) begin
      dataBanks_0_perm_r[dataBanks_0_perm_rMPORT_addr] <= dataBanks_0_perm_rMPORT_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_0_perm_pm_rMPORT_en & dataBanks_0_perm_pm_rMPORT_mask) begin
      dataBanks_0_perm_pm_r[dataBanks_0_perm_pm_rMPORT_addr] <= dataBanks_0_perm_pm_rMPORT_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_0_perm_pm_wMPORT_en & dataBanks_0_perm_pm_wMPORT_mask) begin
      dataBanks_0_perm_pm_w[dataBanks_0_perm_pm_wMPORT_addr] <= dataBanks_0_perm_pm_wMPORT_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_0_perm_pm_c_MPORT_en & dataBanks_0_perm_pm_c_MPORT_mask) begin
      dataBanks_0_perm_pm_c[dataBanks_0_perm_pm_c_MPORT_addr] <= dataBanks_0_perm_pm_c_MPORT_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_1_tag_MPORT_1_en & dataBanks_1_tag_MPORT_1_mask) begin
      dataBanks_1_tag[dataBanks_1_tag_MPORT_1_addr] <= dataBanks_1_tag_MPORT_1_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_1_asid_MPORT_1_en & dataBanks_1_asid_MPORT_1_mask) begin
      dataBanks_1_asid[dataBanks_1_asid_MPORT_1_addr] <= dataBanks_1_asid_MPORT_1_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_1_ppn_MPORT_1_en & dataBanks_1_ppn_MPORT_1_mask) begin
      dataBanks_1_ppn[dataBanks_1_ppn_MPORT_1_addr] <= dataBanks_1_ppn_MPORT_1_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_1_perm_pf_MPORT_1_en & dataBanks_1_perm_pf_MPORT_1_mask) begin
      dataBanks_1_perm_pf[dataBanks_1_perm_pf_MPORT_1_addr] <= dataBanks_1_perm_pf_MPORT_1_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_1_perm_af_MPORT_1_en & dataBanks_1_perm_af_MPORT_1_mask) begin
      dataBanks_1_perm_af[dataBanks_1_perm_af_MPORT_1_addr] <= dataBanks_1_perm_af_MPORT_1_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_1_perm_d_MPORT_1_en & dataBanks_1_perm_d_MPORT_1_mask) begin
      dataBanks_1_perm_d[dataBanks_1_perm_d_MPORT_1_addr] <= dataBanks_1_perm_d_MPORT_1_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_1_perm_a_MPORT_1_en & dataBanks_1_perm_a_MPORT_1_mask) begin
      dataBanks_1_perm_a[dataBanks_1_perm_a_MPORT_1_addr] <= dataBanks_1_perm_a_MPORT_1_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_1_perm_u_MPORT_1_en & dataBanks_1_perm_u_MPORT_1_mask) begin
      dataBanks_1_perm_u[dataBanks_1_perm_u_MPORT_1_addr] <= dataBanks_1_perm_u_MPORT_1_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_1_perm_x_MPORT_1_en & dataBanks_1_perm_x_MPORT_1_mask) begin
      dataBanks_1_perm_x[dataBanks_1_perm_x_MPORT_1_addr] <= dataBanks_1_perm_x_MPORT_1_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_1_perm_wMPORT_1_en & dataBanks_1_perm_wMPORT_1_mask) begin
      dataBanks_1_perm_w[dataBanks_1_perm_wMPORT_1_addr] <= dataBanks_1_perm_wMPORT_1_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_1_perm_rMPORT_1_en & dataBanks_1_perm_rMPORT_1_mask) begin
      dataBanks_1_perm_r[dataBanks_1_perm_rMPORT_1_addr] <= dataBanks_1_perm_rMPORT_1_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_1_perm_pm_rMPORT_1_en & dataBanks_1_perm_pm_rMPORT_1_mask) begin
      dataBanks_1_perm_pm_r[dataBanks_1_perm_pm_rMPORT_1_addr] <= dataBanks_1_perm_pm_rMPORT_1_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_1_perm_pm_wMPORT_1_en & dataBanks_1_perm_pm_wMPORT_1_mask) begin
      dataBanks_1_perm_pm_w[dataBanks_1_perm_pm_wMPORT_1_addr] <= dataBanks_1_perm_pm_wMPORT_1_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_1_perm_pm_c_MPORT_1_en & dataBanks_1_perm_pm_c_MPORT_1_mask) begin
      dataBanks_1_perm_pm_c[dataBanks_1_perm_pm_c_MPORT_1_addr] <= dataBanks_1_perm_pm_c_MPORT_1_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_2_tag_MPORT_2_en & dataBanks_2_tag_MPORT_2_mask) begin
      dataBanks_2_tag[dataBanks_2_tag_MPORT_2_addr] <= dataBanks_2_tag_MPORT_2_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_2_asid_MPORT_2_en & dataBanks_2_asid_MPORT_2_mask) begin
      dataBanks_2_asid[dataBanks_2_asid_MPORT_2_addr] <= dataBanks_2_asid_MPORT_2_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_2_ppn_MPORT_2_en & dataBanks_2_ppn_MPORT_2_mask) begin
      dataBanks_2_ppn[dataBanks_2_ppn_MPORT_2_addr] <= dataBanks_2_ppn_MPORT_2_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_2_perm_pf_MPORT_2_en & dataBanks_2_perm_pf_MPORT_2_mask) begin
      dataBanks_2_perm_pf[dataBanks_2_perm_pf_MPORT_2_addr] <= dataBanks_2_perm_pf_MPORT_2_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_2_perm_af_MPORT_2_en & dataBanks_2_perm_af_MPORT_2_mask) begin
      dataBanks_2_perm_af[dataBanks_2_perm_af_MPORT_2_addr] <= dataBanks_2_perm_af_MPORT_2_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_2_perm_d_MPORT_2_en & dataBanks_2_perm_d_MPORT_2_mask) begin
      dataBanks_2_perm_d[dataBanks_2_perm_d_MPORT_2_addr] <= dataBanks_2_perm_d_MPORT_2_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_2_perm_a_MPORT_2_en & dataBanks_2_perm_a_MPORT_2_mask) begin
      dataBanks_2_perm_a[dataBanks_2_perm_a_MPORT_2_addr] <= dataBanks_2_perm_a_MPORT_2_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_2_perm_u_MPORT_2_en & dataBanks_2_perm_u_MPORT_2_mask) begin
      dataBanks_2_perm_u[dataBanks_2_perm_u_MPORT_2_addr] <= dataBanks_2_perm_u_MPORT_2_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_2_perm_x_MPORT_2_en & dataBanks_2_perm_x_MPORT_2_mask) begin
      dataBanks_2_perm_x[dataBanks_2_perm_x_MPORT_2_addr] <= dataBanks_2_perm_x_MPORT_2_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_2_perm_wMPORT_2_en & dataBanks_2_perm_wMPORT_2_mask) begin
      dataBanks_2_perm_w[dataBanks_2_perm_wMPORT_2_addr] <= dataBanks_2_perm_wMPORT_2_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_2_perm_rMPORT_2_en & dataBanks_2_perm_rMPORT_2_mask) begin
      dataBanks_2_perm_r[dataBanks_2_perm_rMPORT_2_addr] <= dataBanks_2_perm_rMPORT_2_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_2_perm_pm_rMPORT_2_en & dataBanks_2_perm_pm_rMPORT_2_mask) begin
      dataBanks_2_perm_pm_r[dataBanks_2_perm_pm_rMPORT_2_addr] <= dataBanks_2_perm_pm_rMPORT_2_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_2_perm_pm_wMPORT_2_en & dataBanks_2_perm_pm_wMPORT_2_mask) begin
      dataBanks_2_perm_pm_w[dataBanks_2_perm_pm_wMPORT_2_addr] <= dataBanks_2_perm_pm_wMPORT_2_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_2_perm_pm_c_MPORT_2_en & dataBanks_2_perm_pm_c_MPORT_2_mask) begin
      dataBanks_2_perm_pm_c[dataBanks_2_perm_pm_c_MPORT_2_addr] <= dataBanks_2_perm_pm_c_MPORT_2_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_3_tag_MPORT_3_en & dataBanks_3_tag_MPORT_3_mask) begin
      dataBanks_3_tag[dataBanks_3_tag_MPORT_3_addr] <= dataBanks_3_tag_MPORT_3_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_3_asid_MPORT_3_en & dataBanks_3_asid_MPORT_3_mask) begin
      dataBanks_3_asid[dataBanks_3_asid_MPORT_3_addr] <= dataBanks_3_asid_MPORT_3_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_3_ppn_MPORT_3_en & dataBanks_3_ppn_MPORT_3_mask) begin
      dataBanks_3_ppn[dataBanks_3_ppn_MPORT_3_addr] <= dataBanks_3_ppn_MPORT_3_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_3_perm_pf_MPORT_3_en & dataBanks_3_perm_pf_MPORT_3_mask) begin
      dataBanks_3_perm_pf[dataBanks_3_perm_pf_MPORT_3_addr] <= dataBanks_3_perm_pf_MPORT_3_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_3_perm_af_MPORT_3_en & dataBanks_3_perm_af_MPORT_3_mask) begin
      dataBanks_3_perm_af[dataBanks_3_perm_af_MPORT_3_addr] <= dataBanks_3_perm_af_MPORT_3_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_3_perm_d_MPORT_3_en & dataBanks_3_perm_d_MPORT_3_mask) begin
      dataBanks_3_perm_d[dataBanks_3_perm_d_MPORT_3_addr] <= dataBanks_3_perm_d_MPORT_3_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_3_perm_a_MPORT_3_en & dataBanks_3_perm_a_MPORT_3_mask) begin
      dataBanks_3_perm_a[dataBanks_3_perm_a_MPORT_3_addr] <= dataBanks_3_perm_a_MPORT_3_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_3_perm_u_MPORT_3_en & dataBanks_3_perm_u_MPORT_3_mask) begin
      dataBanks_3_perm_u[dataBanks_3_perm_u_MPORT_3_addr] <= dataBanks_3_perm_u_MPORT_3_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_3_perm_x_MPORT_3_en & dataBanks_3_perm_x_MPORT_3_mask) begin
      dataBanks_3_perm_x[dataBanks_3_perm_x_MPORT_3_addr] <= dataBanks_3_perm_x_MPORT_3_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_3_perm_wMPORT_3_en & dataBanks_3_perm_wMPORT_3_mask) begin
      dataBanks_3_perm_w[dataBanks_3_perm_wMPORT_3_addr] <= dataBanks_3_perm_wMPORT_3_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_3_perm_rMPORT_3_en & dataBanks_3_perm_rMPORT_3_mask) begin
      dataBanks_3_perm_r[dataBanks_3_perm_rMPORT_3_addr] <= dataBanks_3_perm_rMPORT_3_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_3_perm_pm_rMPORT_3_en & dataBanks_3_perm_pm_rMPORT_3_mask) begin
      dataBanks_3_perm_pm_r[dataBanks_3_perm_pm_rMPORT_3_addr] <= dataBanks_3_perm_pm_rMPORT_3_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_3_perm_pm_wMPORT_3_en & dataBanks_3_perm_pm_wMPORT_3_mask) begin
      dataBanks_3_perm_pm_w[dataBanks_3_perm_pm_wMPORT_3_addr] <= dataBanks_3_perm_pm_wMPORT_3_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_3_perm_pm_c_MPORT_3_en & dataBanks_3_perm_pm_c_MPORT_3_mask) begin
      dataBanks_3_perm_pm_c[dataBanks_3_perm_pm_c_MPORT_3_addr] <= dataBanks_3_perm_pm_c_MPORT_3_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_4_tag_MPORT_4_en & dataBanks_4_tag_MPORT_4_mask) begin
      dataBanks_4_tag[dataBanks_4_tag_MPORT_4_addr] <= dataBanks_4_tag_MPORT_4_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_4_asid_MPORT_4_en & dataBanks_4_asid_MPORT_4_mask) begin
      dataBanks_4_asid[dataBanks_4_asid_MPORT_4_addr] <= dataBanks_4_asid_MPORT_4_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_4_ppn_MPORT_4_en & dataBanks_4_ppn_MPORT_4_mask) begin
      dataBanks_4_ppn[dataBanks_4_ppn_MPORT_4_addr] <= dataBanks_4_ppn_MPORT_4_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_4_perm_pf_MPORT_4_en & dataBanks_4_perm_pf_MPORT_4_mask) begin
      dataBanks_4_perm_pf[dataBanks_4_perm_pf_MPORT_4_addr] <= dataBanks_4_perm_pf_MPORT_4_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_4_perm_af_MPORT_4_en & dataBanks_4_perm_af_MPORT_4_mask) begin
      dataBanks_4_perm_af[dataBanks_4_perm_af_MPORT_4_addr] <= dataBanks_4_perm_af_MPORT_4_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_4_perm_d_MPORT_4_en & dataBanks_4_perm_d_MPORT_4_mask) begin
      dataBanks_4_perm_d[dataBanks_4_perm_d_MPORT_4_addr] <= dataBanks_4_perm_d_MPORT_4_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_4_perm_a_MPORT_4_en & dataBanks_4_perm_a_MPORT_4_mask) begin
      dataBanks_4_perm_a[dataBanks_4_perm_a_MPORT_4_addr] <= dataBanks_4_perm_a_MPORT_4_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_4_perm_u_MPORT_4_en & dataBanks_4_perm_u_MPORT_4_mask) begin
      dataBanks_4_perm_u[dataBanks_4_perm_u_MPORT_4_addr] <= dataBanks_4_perm_u_MPORT_4_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_4_perm_x_MPORT_4_en & dataBanks_4_perm_x_MPORT_4_mask) begin
      dataBanks_4_perm_x[dataBanks_4_perm_x_MPORT_4_addr] <= dataBanks_4_perm_x_MPORT_4_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_4_perm_wMPORT_4_en & dataBanks_4_perm_wMPORT_4_mask) begin
      dataBanks_4_perm_w[dataBanks_4_perm_wMPORT_4_addr] <= dataBanks_4_perm_wMPORT_4_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_4_perm_rMPORT_4_en & dataBanks_4_perm_rMPORT_4_mask) begin
      dataBanks_4_perm_r[dataBanks_4_perm_rMPORT_4_addr] <= dataBanks_4_perm_rMPORT_4_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_4_perm_pm_rMPORT_4_en & dataBanks_4_perm_pm_rMPORT_4_mask) begin
      dataBanks_4_perm_pm_r[dataBanks_4_perm_pm_rMPORT_4_addr] <= dataBanks_4_perm_pm_rMPORT_4_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_4_perm_pm_wMPORT_4_en & dataBanks_4_perm_pm_wMPORT_4_mask) begin
      dataBanks_4_perm_pm_w[dataBanks_4_perm_pm_wMPORT_4_addr] <= dataBanks_4_perm_pm_wMPORT_4_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_4_perm_pm_c_MPORT_4_en & dataBanks_4_perm_pm_c_MPORT_4_mask) begin
      dataBanks_4_perm_pm_c[dataBanks_4_perm_pm_c_MPORT_4_addr] <= dataBanks_4_perm_pm_c_MPORT_4_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_5_tag_MPORT_5_en & dataBanks_5_tag_MPORT_5_mask) begin
      dataBanks_5_tag[dataBanks_5_tag_MPORT_5_addr] <= dataBanks_5_tag_MPORT_5_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_5_asid_MPORT_5_en & dataBanks_5_asid_MPORT_5_mask) begin
      dataBanks_5_asid[dataBanks_5_asid_MPORT_5_addr] <= dataBanks_5_asid_MPORT_5_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_5_ppn_MPORT_5_en & dataBanks_5_ppn_MPORT_5_mask) begin
      dataBanks_5_ppn[dataBanks_5_ppn_MPORT_5_addr] <= dataBanks_5_ppn_MPORT_5_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_5_perm_pf_MPORT_5_en & dataBanks_5_perm_pf_MPORT_5_mask) begin
      dataBanks_5_perm_pf[dataBanks_5_perm_pf_MPORT_5_addr] <= dataBanks_5_perm_pf_MPORT_5_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_5_perm_af_MPORT_5_en & dataBanks_5_perm_af_MPORT_5_mask) begin
      dataBanks_5_perm_af[dataBanks_5_perm_af_MPORT_5_addr] <= dataBanks_5_perm_af_MPORT_5_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_5_perm_d_MPORT_5_en & dataBanks_5_perm_d_MPORT_5_mask) begin
      dataBanks_5_perm_d[dataBanks_5_perm_d_MPORT_5_addr] <= dataBanks_5_perm_d_MPORT_5_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_5_perm_a_MPORT_5_en & dataBanks_5_perm_a_MPORT_5_mask) begin
      dataBanks_5_perm_a[dataBanks_5_perm_a_MPORT_5_addr] <= dataBanks_5_perm_a_MPORT_5_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_5_perm_u_MPORT_5_en & dataBanks_5_perm_u_MPORT_5_mask) begin
      dataBanks_5_perm_u[dataBanks_5_perm_u_MPORT_5_addr] <= dataBanks_5_perm_u_MPORT_5_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_5_perm_x_MPORT_5_en & dataBanks_5_perm_x_MPORT_5_mask) begin
      dataBanks_5_perm_x[dataBanks_5_perm_x_MPORT_5_addr] <= dataBanks_5_perm_x_MPORT_5_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_5_perm_wMPORT_5_en & dataBanks_5_perm_wMPORT_5_mask) begin
      dataBanks_5_perm_w[dataBanks_5_perm_wMPORT_5_addr] <= dataBanks_5_perm_wMPORT_5_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_5_perm_rMPORT_5_en & dataBanks_5_perm_rMPORT_5_mask) begin
      dataBanks_5_perm_r[dataBanks_5_perm_rMPORT_5_addr] <= dataBanks_5_perm_rMPORT_5_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_5_perm_pm_rMPORT_5_en & dataBanks_5_perm_pm_rMPORT_5_mask) begin
      dataBanks_5_perm_pm_r[dataBanks_5_perm_pm_rMPORT_5_addr] <= dataBanks_5_perm_pm_rMPORT_5_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_5_perm_pm_wMPORT_5_en & dataBanks_5_perm_pm_wMPORT_5_mask) begin
      dataBanks_5_perm_pm_w[dataBanks_5_perm_pm_wMPORT_5_addr] <= dataBanks_5_perm_pm_wMPORT_5_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_5_perm_pm_c_MPORT_5_en & dataBanks_5_perm_pm_c_MPORT_5_mask) begin
      dataBanks_5_perm_pm_c[dataBanks_5_perm_pm_c_MPORT_5_addr] <= dataBanks_5_perm_pm_c_MPORT_5_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_6_tag_MPORT_6_en & dataBanks_6_tag_MPORT_6_mask) begin
      dataBanks_6_tag[dataBanks_6_tag_MPORT_6_addr] <= dataBanks_6_tag_MPORT_6_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_6_asid_MPORT_6_en & dataBanks_6_asid_MPORT_6_mask) begin
      dataBanks_6_asid[dataBanks_6_asid_MPORT_6_addr] <= dataBanks_6_asid_MPORT_6_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_6_ppn_MPORT_6_en & dataBanks_6_ppn_MPORT_6_mask) begin
      dataBanks_6_ppn[dataBanks_6_ppn_MPORT_6_addr] <= dataBanks_6_ppn_MPORT_6_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_6_perm_pf_MPORT_6_en & dataBanks_6_perm_pf_MPORT_6_mask) begin
      dataBanks_6_perm_pf[dataBanks_6_perm_pf_MPORT_6_addr] <= dataBanks_6_perm_pf_MPORT_6_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_6_perm_af_MPORT_6_en & dataBanks_6_perm_af_MPORT_6_mask) begin
      dataBanks_6_perm_af[dataBanks_6_perm_af_MPORT_6_addr] <= dataBanks_6_perm_af_MPORT_6_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_6_perm_d_MPORT_6_en & dataBanks_6_perm_d_MPORT_6_mask) begin
      dataBanks_6_perm_d[dataBanks_6_perm_d_MPORT_6_addr] <= dataBanks_6_perm_d_MPORT_6_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_6_perm_a_MPORT_6_en & dataBanks_6_perm_a_MPORT_6_mask) begin
      dataBanks_6_perm_a[dataBanks_6_perm_a_MPORT_6_addr] <= dataBanks_6_perm_a_MPORT_6_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_6_perm_u_MPORT_6_en & dataBanks_6_perm_u_MPORT_6_mask) begin
      dataBanks_6_perm_u[dataBanks_6_perm_u_MPORT_6_addr] <= dataBanks_6_perm_u_MPORT_6_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_6_perm_x_MPORT_6_en & dataBanks_6_perm_x_MPORT_6_mask) begin
      dataBanks_6_perm_x[dataBanks_6_perm_x_MPORT_6_addr] <= dataBanks_6_perm_x_MPORT_6_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_6_perm_wMPORT_6_en & dataBanks_6_perm_wMPORT_6_mask) begin
      dataBanks_6_perm_w[dataBanks_6_perm_wMPORT_6_addr] <= dataBanks_6_perm_wMPORT_6_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_6_perm_rMPORT_6_en & dataBanks_6_perm_rMPORT_6_mask) begin
      dataBanks_6_perm_r[dataBanks_6_perm_rMPORT_6_addr] <= dataBanks_6_perm_rMPORT_6_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_6_perm_pm_rMPORT_6_en & dataBanks_6_perm_pm_rMPORT_6_mask) begin
      dataBanks_6_perm_pm_r[dataBanks_6_perm_pm_rMPORT_6_addr] <= dataBanks_6_perm_pm_rMPORT_6_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_6_perm_pm_wMPORT_6_en & dataBanks_6_perm_pm_wMPORT_6_mask) begin
      dataBanks_6_perm_pm_w[dataBanks_6_perm_pm_wMPORT_6_addr] <= dataBanks_6_perm_pm_wMPORT_6_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_6_perm_pm_c_MPORT_6_en & dataBanks_6_perm_pm_c_MPORT_6_mask) begin
      dataBanks_6_perm_pm_c[dataBanks_6_perm_pm_c_MPORT_6_addr] <= dataBanks_6_perm_pm_c_MPORT_6_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_7_tag_MPORT_7_en & dataBanks_7_tag_MPORT_7_mask) begin
      dataBanks_7_tag[dataBanks_7_tag_MPORT_7_addr] <= dataBanks_7_tag_MPORT_7_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_7_asid_MPORT_7_en & dataBanks_7_asid_MPORT_7_mask) begin
      dataBanks_7_asid[dataBanks_7_asid_MPORT_7_addr] <= dataBanks_7_asid_MPORT_7_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_7_ppn_MPORT_7_en & dataBanks_7_ppn_MPORT_7_mask) begin
      dataBanks_7_ppn[dataBanks_7_ppn_MPORT_7_addr] <= dataBanks_7_ppn_MPORT_7_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_7_perm_pf_MPORT_7_en & dataBanks_7_perm_pf_MPORT_7_mask) begin
      dataBanks_7_perm_pf[dataBanks_7_perm_pf_MPORT_7_addr] <= dataBanks_7_perm_pf_MPORT_7_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_7_perm_af_MPORT_7_en & dataBanks_7_perm_af_MPORT_7_mask) begin
      dataBanks_7_perm_af[dataBanks_7_perm_af_MPORT_7_addr] <= dataBanks_7_perm_af_MPORT_7_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_7_perm_d_MPORT_7_en & dataBanks_7_perm_d_MPORT_7_mask) begin
      dataBanks_7_perm_d[dataBanks_7_perm_d_MPORT_7_addr] <= dataBanks_7_perm_d_MPORT_7_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_7_perm_a_MPORT_7_en & dataBanks_7_perm_a_MPORT_7_mask) begin
      dataBanks_7_perm_a[dataBanks_7_perm_a_MPORT_7_addr] <= dataBanks_7_perm_a_MPORT_7_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_7_perm_u_MPORT_7_en & dataBanks_7_perm_u_MPORT_7_mask) begin
      dataBanks_7_perm_u[dataBanks_7_perm_u_MPORT_7_addr] <= dataBanks_7_perm_u_MPORT_7_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_7_perm_x_MPORT_7_en & dataBanks_7_perm_x_MPORT_7_mask) begin
      dataBanks_7_perm_x[dataBanks_7_perm_x_MPORT_7_addr] <= dataBanks_7_perm_x_MPORT_7_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_7_perm_wMPORT_7_en & dataBanks_7_perm_wMPORT_7_mask) begin
      dataBanks_7_perm_w[dataBanks_7_perm_wMPORT_7_addr] <= dataBanks_7_perm_wMPORT_7_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_7_perm_rMPORT_7_en & dataBanks_7_perm_rMPORT_7_mask) begin
      dataBanks_7_perm_r[dataBanks_7_perm_rMPORT_7_addr] <= dataBanks_7_perm_rMPORT_7_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_7_perm_pm_rMPORT_7_en & dataBanks_7_perm_pm_rMPORT_7_mask) begin
      dataBanks_7_perm_pm_r[dataBanks_7_perm_pm_rMPORT_7_addr] <= dataBanks_7_perm_pm_rMPORT_7_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_7_perm_pm_wMPORT_7_en & dataBanks_7_perm_pm_wMPORT_7_mask) begin
      dataBanks_7_perm_pm_w[dataBanks_7_perm_pm_wMPORT_7_addr] <= dataBanks_7_perm_pm_wMPORT_7_data; // @[TLBStorage.scala 58:8]
    end
    if (dataBanks_7_perm_pm_c_MPORT_7_en & dataBanks_7_perm_pm_c_MPORT_7_mask) begin
      dataBanks_7_perm_pm_c[dataBanks_7_perm_pm_c_MPORT_7_addr] <= dataBanks_7_perm_pm_c_MPORT_7_data; // @[TLBStorage.scala 58:8]
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_0_tag <= io_wdata_tag;
    end else begin
      data_read__0_0_tag <= dataBanks_0_tag_data_read_0_0_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_0_asid <= io_wdata_asid;
    end else begin
      data_read__0_0_asid <= dataBanks_0_asid_data_read_0_0_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_0_ppn <= io_wdata_ppn;
    end else begin
      data_read__0_0_ppn <= dataBanks_0_ppn_data_read_0_0_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_0_perm_pf <= io_wdata_perm_pf;
    end else begin
      data_read__0_0_perm_pf <= dataBanks_0_perm_pf_data_read_0_0_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_0_perm_af <= io_wdata_perm_af;
    end else begin
      data_read__0_0_perm_af <= dataBanks_0_perm_af_data_read_0_0_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_0_perm_d <= io_wdata_perm_d;
    end else begin
      data_read__0_0_perm_d <= dataBanks_0_perm_d_data_read_0_0_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_0_perm_a <= io_wdata_perm_a;
    end else begin
      data_read__0_0_perm_a <= dataBanks_0_perm_a_data_read_0_0_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_0_perm_u <= io_wdata_perm_u;
    end else begin
      data_read__0_0_perm_u <= dataBanks_0_perm_u_data_read_0_0_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_0_perm_x <= io_wdata_perm_x;
    end else begin
      data_read__0_0_perm_x <= dataBanks_0_perm_x_data_read_0_0_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_0_perm_w <= io_wdata_perm_w;
    end else begin
      data_read__0_0_perm_w <= dataBanks_0_perm_wdata_read_0_0_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_0_perm_r <= io_wdata_perm_r;
    end else begin
      data_read__0_0_perm_r <= dataBanks_0_perm_rdata_read_0_0_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_0_perm_pm_r <= io_wdata_perm_pm_r;
    end else begin
      data_read__0_0_perm_pm_r <= dataBanks_0_perm_pm_rdata_read_0_0_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_0_perm_pm_w <= io_wdata_perm_pm_w;
    end else begin
      data_read__0_0_perm_pm_w <= dataBanks_0_perm_pm_wdata_read_0_0_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_0_perm_pm_c <= io_wdata_perm_pm_c;
    end else begin
      data_read__0_0_perm_pm_c <= dataBanks_0_perm_pm_c_data_read_0_0_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_1_tag <= io_wdata_tag;
    end else begin
      data_read__0_1_tag <= dataBanks_1_tag_data_read_0_1_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_1_asid <= io_wdata_asid;
    end else begin
      data_read__0_1_asid <= dataBanks_1_asid_data_read_0_1_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_1_ppn <= io_wdata_ppn;
    end else begin
      data_read__0_1_ppn <= dataBanks_1_ppn_data_read_0_1_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_1_perm_pf <= io_wdata_perm_pf;
    end else begin
      data_read__0_1_perm_pf <= dataBanks_1_perm_pf_data_read_0_1_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_1_perm_af <= io_wdata_perm_af;
    end else begin
      data_read__0_1_perm_af <= dataBanks_1_perm_af_data_read_0_1_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_1_perm_d <= io_wdata_perm_d;
    end else begin
      data_read__0_1_perm_d <= dataBanks_1_perm_d_data_read_0_1_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_1_perm_a <= io_wdata_perm_a;
    end else begin
      data_read__0_1_perm_a <= dataBanks_1_perm_a_data_read_0_1_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_1_perm_u <= io_wdata_perm_u;
    end else begin
      data_read__0_1_perm_u <= dataBanks_1_perm_u_data_read_0_1_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_1_perm_x <= io_wdata_perm_x;
    end else begin
      data_read__0_1_perm_x <= dataBanks_1_perm_x_data_read_0_1_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_1_perm_w <= io_wdata_perm_w;
    end else begin
      data_read__0_1_perm_w <= dataBanks_1_perm_wdata_read_0_1_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_1_perm_r <= io_wdata_perm_r;
    end else begin
      data_read__0_1_perm_r <= dataBanks_1_perm_rdata_read_0_1_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_1_perm_pm_r <= io_wdata_perm_pm_r;
    end else begin
      data_read__0_1_perm_pm_r <= dataBanks_1_perm_pm_rdata_read_0_1_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_1_perm_pm_w <= io_wdata_perm_pm_w;
    end else begin
      data_read__0_1_perm_pm_w <= dataBanks_1_perm_pm_wdata_read_0_1_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_1_perm_pm_c <= io_wdata_perm_pm_c;
    end else begin
      data_read__0_1_perm_pm_c <= dataBanks_1_perm_pm_c_data_read_0_1_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_2_tag <= io_wdata_tag;
    end else begin
      data_read__0_2_tag <= dataBanks_2_tag_data_read_0_2_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_2_asid <= io_wdata_asid;
    end else begin
      data_read__0_2_asid <= dataBanks_2_asid_data_read_0_2_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_2_ppn <= io_wdata_ppn;
    end else begin
      data_read__0_2_ppn <= dataBanks_2_ppn_data_read_0_2_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_2_perm_pf <= io_wdata_perm_pf;
    end else begin
      data_read__0_2_perm_pf <= dataBanks_2_perm_pf_data_read_0_2_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_2_perm_af <= io_wdata_perm_af;
    end else begin
      data_read__0_2_perm_af <= dataBanks_2_perm_af_data_read_0_2_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_2_perm_d <= io_wdata_perm_d;
    end else begin
      data_read__0_2_perm_d <= dataBanks_2_perm_d_data_read_0_2_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_2_perm_a <= io_wdata_perm_a;
    end else begin
      data_read__0_2_perm_a <= dataBanks_2_perm_a_data_read_0_2_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_2_perm_u <= io_wdata_perm_u;
    end else begin
      data_read__0_2_perm_u <= dataBanks_2_perm_u_data_read_0_2_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_2_perm_x <= io_wdata_perm_x;
    end else begin
      data_read__0_2_perm_x <= dataBanks_2_perm_x_data_read_0_2_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_2_perm_w <= io_wdata_perm_w;
    end else begin
      data_read__0_2_perm_w <= dataBanks_2_perm_wdata_read_0_2_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_2_perm_r <= io_wdata_perm_r;
    end else begin
      data_read__0_2_perm_r <= dataBanks_2_perm_rdata_read_0_2_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_2_perm_pm_r <= io_wdata_perm_pm_r;
    end else begin
      data_read__0_2_perm_pm_r <= dataBanks_2_perm_pm_rdata_read_0_2_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_2_perm_pm_w <= io_wdata_perm_pm_w;
    end else begin
      data_read__0_2_perm_pm_w <= dataBanks_2_perm_pm_wdata_read_0_2_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_2_perm_pm_c <= io_wdata_perm_pm_c;
    end else begin
      data_read__0_2_perm_pm_c <= dataBanks_2_perm_pm_c_data_read_0_2_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_3_tag <= io_wdata_tag;
    end else begin
      data_read__0_3_tag <= dataBanks_3_tag_data_read_0_3_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_3_asid <= io_wdata_asid;
    end else begin
      data_read__0_3_asid <= dataBanks_3_asid_data_read_0_3_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_3_ppn <= io_wdata_ppn;
    end else begin
      data_read__0_3_ppn <= dataBanks_3_ppn_data_read_0_3_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_3_perm_pf <= io_wdata_perm_pf;
    end else begin
      data_read__0_3_perm_pf <= dataBanks_3_perm_pf_data_read_0_3_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_3_perm_af <= io_wdata_perm_af;
    end else begin
      data_read__0_3_perm_af <= dataBanks_3_perm_af_data_read_0_3_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_3_perm_d <= io_wdata_perm_d;
    end else begin
      data_read__0_3_perm_d <= dataBanks_3_perm_d_data_read_0_3_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_3_perm_a <= io_wdata_perm_a;
    end else begin
      data_read__0_3_perm_a <= dataBanks_3_perm_a_data_read_0_3_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_3_perm_u <= io_wdata_perm_u;
    end else begin
      data_read__0_3_perm_u <= dataBanks_3_perm_u_data_read_0_3_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_3_perm_x <= io_wdata_perm_x;
    end else begin
      data_read__0_3_perm_x <= dataBanks_3_perm_x_data_read_0_3_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_3_perm_w <= io_wdata_perm_w;
    end else begin
      data_read__0_3_perm_w <= dataBanks_3_perm_wdata_read_0_3_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_3_perm_r <= io_wdata_perm_r;
    end else begin
      data_read__0_3_perm_r <= dataBanks_3_perm_rdata_read_0_3_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_3_perm_pm_r <= io_wdata_perm_pm_r;
    end else begin
      data_read__0_3_perm_pm_r <= dataBanks_3_perm_pm_rdata_read_0_3_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_3_perm_pm_w <= io_wdata_perm_pm_w;
    end else begin
      data_read__0_3_perm_pm_w <= dataBanks_3_perm_pm_wdata_read_0_3_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_3_perm_pm_c <= io_wdata_perm_pm_c;
    end else begin
      data_read__0_3_perm_pm_c <= dataBanks_3_perm_pm_c_data_read_0_3_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_4_tag <= io_wdata_tag;
    end else begin
      data_read__0_4_tag <= dataBanks_4_tag_data_read_0_4_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_4_asid <= io_wdata_asid;
    end else begin
      data_read__0_4_asid <= dataBanks_4_asid_data_read_0_4_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_4_ppn <= io_wdata_ppn;
    end else begin
      data_read__0_4_ppn <= dataBanks_4_ppn_data_read_0_4_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_4_perm_pf <= io_wdata_perm_pf;
    end else begin
      data_read__0_4_perm_pf <= dataBanks_4_perm_pf_data_read_0_4_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_4_perm_af <= io_wdata_perm_af;
    end else begin
      data_read__0_4_perm_af <= dataBanks_4_perm_af_data_read_0_4_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_4_perm_d <= io_wdata_perm_d;
    end else begin
      data_read__0_4_perm_d <= dataBanks_4_perm_d_data_read_0_4_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_4_perm_a <= io_wdata_perm_a;
    end else begin
      data_read__0_4_perm_a <= dataBanks_4_perm_a_data_read_0_4_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_4_perm_u <= io_wdata_perm_u;
    end else begin
      data_read__0_4_perm_u <= dataBanks_4_perm_u_data_read_0_4_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_4_perm_x <= io_wdata_perm_x;
    end else begin
      data_read__0_4_perm_x <= dataBanks_4_perm_x_data_read_0_4_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_4_perm_w <= io_wdata_perm_w;
    end else begin
      data_read__0_4_perm_w <= dataBanks_4_perm_wdata_read_0_4_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_4_perm_r <= io_wdata_perm_r;
    end else begin
      data_read__0_4_perm_r <= dataBanks_4_perm_rdata_read_0_4_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_4_perm_pm_r <= io_wdata_perm_pm_r;
    end else begin
      data_read__0_4_perm_pm_r <= dataBanks_4_perm_pm_rdata_read_0_4_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_4_perm_pm_w <= io_wdata_perm_pm_w;
    end else begin
      data_read__0_4_perm_pm_w <= dataBanks_4_perm_pm_wdata_read_0_4_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_4_perm_pm_c <= io_wdata_perm_pm_c;
    end else begin
      data_read__0_4_perm_pm_c <= dataBanks_4_perm_pm_c_data_read_0_4_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_5_tag <= io_wdata_tag;
    end else begin
      data_read__0_5_tag <= dataBanks_5_tag_data_read_0_5_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_5_asid <= io_wdata_asid;
    end else begin
      data_read__0_5_asid <= dataBanks_5_asid_data_read_0_5_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_5_ppn <= io_wdata_ppn;
    end else begin
      data_read__0_5_ppn <= dataBanks_5_ppn_data_read_0_5_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_5_perm_pf <= io_wdata_perm_pf;
    end else begin
      data_read__0_5_perm_pf <= dataBanks_5_perm_pf_data_read_0_5_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_5_perm_af <= io_wdata_perm_af;
    end else begin
      data_read__0_5_perm_af <= dataBanks_5_perm_af_data_read_0_5_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_5_perm_d <= io_wdata_perm_d;
    end else begin
      data_read__0_5_perm_d <= dataBanks_5_perm_d_data_read_0_5_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_5_perm_a <= io_wdata_perm_a;
    end else begin
      data_read__0_5_perm_a <= dataBanks_5_perm_a_data_read_0_5_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_5_perm_u <= io_wdata_perm_u;
    end else begin
      data_read__0_5_perm_u <= dataBanks_5_perm_u_data_read_0_5_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_5_perm_x <= io_wdata_perm_x;
    end else begin
      data_read__0_5_perm_x <= dataBanks_5_perm_x_data_read_0_5_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_5_perm_w <= io_wdata_perm_w;
    end else begin
      data_read__0_5_perm_w <= dataBanks_5_perm_wdata_read_0_5_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_5_perm_r <= io_wdata_perm_r;
    end else begin
      data_read__0_5_perm_r <= dataBanks_5_perm_rdata_read_0_5_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_5_perm_pm_r <= io_wdata_perm_pm_r;
    end else begin
      data_read__0_5_perm_pm_r <= dataBanks_5_perm_pm_rdata_read_0_5_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_5_perm_pm_w <= io_wdata_perm_pm_w;
    end else begin
      data_read__0_5_perm_pm_w <= dataBanks_5_perm_pm_wdata_read_0_5_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_5_perm_pm_c <= io_wdata_perm_pm_c;
    end else begin
      data_read__0_5_perm_pm_c <= dataBanks_5_perm_pm_c_data_read_0_5_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_6_tag <= io_wdata_tag;
    end else begin
      data_read__0_6_tag <= dataBanks_6_tag_data_read_0_6_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_6_asid <= io_wdata_asid;
    end else begin
      data_read__0_6_asid <= dataBanks_6_asid_data_read_0_6_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_6_ppn <= io_wdata_ppn;
    end else begin
      data_read__0_6_ppn <= dataBanks_6_ppn_data_read_0_6_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_6_perm_pf <= io_wdata_perm_pf;
    end else begin
      data_read__0_6_perm_pf <= dataBanks_6_perm_pf_data_read_0_6_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_6_perm_af <= io_wdata_perm_af;
    end else begin
      data_read__0_6_perm_af <= dataBanks_6_perm_af_data_read_0_6_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_6_perm_d <= io_wdata_perm_d;
    end else begin
      data_read__0_6_perm_d <= dataBanks_6_perm_d_data_read_0_6_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_6_perm_a <= io_wdata_perm_a;
    end else begin
      data_read__0_6_perm_a <= dataBanks_6_perm_a_data_read_0_6_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_6_perm_u <= io_wdata_perm_u;
    end else begin
      data_read__0_6_perm_u <= dataBanks_6_perm_u_data_read_0_6_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_6_perm_x <= io_wdata_perm_x;
    end else begin
      data_read__0_6_perm_x <= dataBanks_6_perm_x_data_read_0_6_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_6_perm_w <= io_wdata_perm_w;
    end else begin
      data_read__0_6_perm_w <= dataBanks_6_perm_wdata_read_0_6_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_6_perm_r <= io_wdata_perm_r;
    end else begin
      data_read__0_6_perm_r <= dataBanks_6_perm_rdata_read_0_6_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_6_perm_pm_r <= io_wdata_perm_pm_r;
    end else begin
      data_read__0_6_perm_pm_r <= dataBanks_6_perm_pm_rdata_read_0_6_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_6_perm_pm_w <= io_wdata_perm_pm_w;
    end else begin
      data_read__0_6_perm_pm_w <= dataBanks_6_perm_pm_wdata_read_0_6_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_6_perm_pm_c <= io_wdata_perm_pm_c;
    end else begin
      data_read__0_6_perm_pm_c <= dataBanks_6_perm_pm_c_data_read_0_6_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_7_tag <= io_wdata_tag;
    end else begin
      data_read__0_7_tag <= dataBanks_7_tag_data_read_0_7_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_7_asid <= io_wdata_asid;
    end else begin
      data_read__0_7_asid <= dataBanks_7_asid_data_read_0_7_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_7_ppn <= io_wdata_ppn;
    end else begin
      data_read__0_7_ppn <= dataBanks_7_ppn_data_read_0_7_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_7_perm_pf <= io_wdata_perm_pf;
    end else begin
      data_read__0_7_perm_pf <= dataBanks_7_perm_pf_data_read_0_7_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_7_perm_af <= io_wdata_perm_af;
    end else begin
      data_read__0_7_perm_af <= dataBanks_7_perm_af_data_read_0_7_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_7_perm_d <= io_wdata_perm_d;
    end else begin
      data_read__0_7_perm_d <= dataBanks_7_perm_d_data_read_0_7_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_7_perm_a <= io_wdata_perm_a;
    end else begin
      data_read__0_7_perm_a <= dataBanks_7_perm_a_data_read_0_7_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_7_perm_u <= io_wdata_perm_u;
    end else begin
      data_read__0_7_perm_u <= dataBanks_7_perm_u_data_read_0_7_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_7_perm_x <= io_wdata_perm_x;
    end else begin
      data_read__0_7_perm_x <= dataBanks_7_perm_x_data_read_0_7_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_7_perm_w <= io_wdata_perm_w;
    end else begin
      data_read__0_7_perm_w <= dataBanks_7_perm_wdata_read_0_7_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_7_perm_r <= io_wdata_perm_r;
    end else begin
      data_read__0_7_perm_r <= dataBanks_7_perm_rdata_read_0_7_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_7_perm_pm_r <= io_wdata_perm_pm_r;
    end else begin
      data_read__0_7_perm_pm_r <= dataBanks_7_perm_pm_rdata_read_0_7_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_7_perm_pm_w <= io_wdata_perm_pm_w;
    end else begin
      data_read__0_7_perm_pm_w <= dataBanks_7_perm_pm_wdata_read_0_7_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__0_7_perm_pm_c <= io_wdata_perm_pm_c;
    end else begin
      data_read__0_7_perm_pm_c <= dataBanks_7_perm_pm_c_data_read_0_7_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__1_0_ppn <= io_wdata_ppn;
    end else begin
      data_read__1_0_ppn <= dataBanks_0_ppn_data_read_1_0_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__1_1_ppn <= io_wdata_ppn;
    end else begin
      data_read__1_1_ppn <= dataBanks_1_ppn_data_read_1_1_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__1_2_ppn <= io_wdata_ppn;
    end else begin
      data_read__1_2_ppn <= dataBanks_2_ppn_data_read_1_2_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__1_3_ppn <= io_wdata_ppn;
    end else begin
      data_read__1_3_ppn <= dataBanks_3_ppn_data_read_1_3_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__1_4_ppn <= io_wdata_ppn;
    end else begin
      data_read__1_4_ppn <= dataBanks_4_ppn_data_read_1_4_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__1_5_ppn <= io_wdata_ppn;
    end else begin
      data_read__1_5_ppn <= dataBanks_5_ppn_data_read_1_5_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__1_6_ppn <= io_wdata_ppn;
    end else begin
      data_read__1_6_ppn <= dataBanks_6_ppn_data_read_1_6_MPORT_data;
    end
    if (io_wen & io_waddr == io_raddr_0) begin // @[TLBStorage.scala 68:31]
      data_read__1_7_ppn <= io_wdata_ppn;
    end else begin
      data_read__1_7_ppn <= dataBanks_7_ppn_data_read_1_7_MPORT_data;
    end
    bank_index__0 <= 8'h1 << io_raddr_0[3:1]; // @[OneHot.scala 57:35]
    bank_index__1 <= 8'h1 << io_raddr_0[3:1]; // @[OneHot.scala 57:35]
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_0_0_tag <= io_wdata_tag;
    end else begin
      data_read_1_0_0_tag <= dataBanks_0_tag_data_read_0_0_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_0_0_asid <= io_wdata_asid;
    end else begin
      data_read_1_0_0_asid <= dataBanks_0_asid_data_read_0_0_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_0_0_ppn <= io_wdata_ppn;
    end else begin
      data_read_1_0_0_ppn <= dataBanks_0_ppn_data_read_0_0_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_0_0_perm_pf <= io_wdata_perm_pf;
    end else begin
      data_read_1_0_0_perm_pf <= dataBanks_0_perm_pf_data_read_0_0_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_0_0_perm_af <= io_wdata_perm_af;
    end else begin
      data_read_1_0_0_perm_af <= dataBanks_0_perm_af_data_read_0_0_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_0_0_perm_a <= io_wdata_perm_a;
    end else begin
      data_read_1_0_0_perm_a <= dataBanks_0_perm_a_data_read_0_0_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_0_0_perm_u <= io_wdata_perm_u;
    end else begin
      data_read_1_0_0_perm_u <= dataBanks_0_perm_u_data_read_0_0_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_0_0_perm_x <= io_wdata_perm_x;
    end else begin
      data_read_1_0_0_perm_x <= dataBanks_0_perm_x_data_read_0_0_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_0_0_perm_r <= io_wdata_perm_r;
    end else begin
      data_read_1_0_0_perm_r <= dataBanks_0_perm_rdata_read_0_0_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_0_0_perm_pm_r <= io_wdata_perm_pm_r;
    end else begin
      data_read_1_0_0_perm_pm_r <= dataBanks_0_perm_pm_rdata_read_0_0_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_0_0_perm_pm_c <= io_wdata_perm_pm_c;
    end else begin
      data_read_1_0_0_perm_pm_c <= dataBanks_0_perm_pm_c_data_read_0_0_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_0_1_tag <= io_wdata_tag;
    end else begin
      data_read_1_0_1_tag <= dataBanks_1_tag_data_read_0_1_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_0_1_asid <= io_wdata_asid;
    end else begin
      data_read_1_0_1_asid <= dataBanks_1_asid_data_read_0_1_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_0_1_ppn <= io_wdata_ppn;
    end else begin
      data_read_1_0_1_ppn <= dataBanks_1_ppn_data_read_0_1_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_0_1_perm_pf <= io_wdata_perm_pf;
    end else begin
      data_read_1_0_1_perm_pf <= dataBanks_1_perm_pf_data_read_0_1_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_0_1_perm_af <= io_wdata_perm_af;
    end else begin
      data_read_1_0_1_perm_af <= dataBanks_1_perm_af_data_read_0_1_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_0_1_perm_a <= io_wdata_perm_a;
    end else begin
      data_read_1_0_1_perm_a <= dataBanks_1_perm_a_data_read_0_1_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_0_1_perm_u <= io_wdata_perm_u;
    end else begin
      data_read_1_0_1_perm_u <= dataBanks_1_perm_u_data_read_0_1_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_0_1_perm_x <= io_wdata_perm_x;
    end else begin
      data_read_1_0_1_perm_x <= dataBanks_1_perm_x_data_read_0_1_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_0_1_perm_r <= io_wdata_perm_r;
    end else begin
      data_read_1_0_1_perm_r <= dataBanks_1_perm_rdata_read_0_1_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_0_1_perm_pm_r <= io_wdata_perm_pm_r;
    end else begin
      data_read_1_0_1_perm_pm_r <= dataBanks_1_perm_pm_rdata_read_0_1_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_0_1_perm_pm_c <= io_wdata_perm_pm_c;
    end else begin
      data_read_1_0_1_perm_pm_c <= dataBanks_1_perm_pm_c_data_read_0_1_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_0_2_tag <= io_wdata_tag;
    end else begin
      data_read_1_0_2_tag <= dataBanks_2_tag_data_read_0_2_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_0_2_asid <= io_wdata_asid;
    end else begin
      data_read_1_0_2_asid <= dataBanks_2_asid_data_read_0_2_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_0_2_ppn <= io_wdata_ppn;
    end else begin
      data_read_1_0_2_ppn <= dataBanks_2_ppn_data_read_0_2_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_0_2_perm_pf <= io_wdata_perm_pf;
    end else begin
      data_read_1_0_2_perm_pf <= dataBanks_2_perm_pf_data_read_0_2_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_0_2_perm_af <= io_wdata_perm_af;
    end else begin
      data_read_1_0_2_perm_af <= dataBanks_2_perm_af_data_read_0_2_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_0_2_perm_a <= io_wdata_perm_a;
    end else begin
      data_read_1_0_2_perm_a <= dataBanks_2_perm_a_data_read_0_2_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_0_2_perm_u <= io_wdata_perm_u;
    end else begin
      data_read_1_0_2_perm_u <= dataBanks_2_perm_u_data_read_0_2_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_0_2_perm_x <= io_wdata_perm_x;
    end else begin
      data_read_1_0_2_perm_x <= dataBanks_2_perm_x_data_read_0_2_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_0_2_perm_r <= io_wdata_perm_r;
    end else begin
      data_read_1_0_2_perm_r <= dataBanks_2_perm_rdata_read_0_2_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_0_2_perm_pm_r <= io_wdata_perm_pm_r;
    end else begin
      data_read_1_0_2_perm_pm_r <= dataBanks_2_perm_pm_rdata_read_0_2_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_0_2_perm_pm_c <= io_wdata_perm_pm_c;
    end else begin
      data_read_1_0_2_perm_pm_c <= dataBanks_2_perm_pm_c_data_read_0_2_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_0_3_tag <= io_wdata_tag;
    end else begin
      data_read_1_0_3_tag <= dataBanks_3_tag_data_read_0_3_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_0_3_asid <= io_wdata_asid;
    end else begin
      data_read_1_0_3_asid <= dataBanks_3_asid_data_read_0_3_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_0_3_ppn <= io_wdata_ppn;
    end else begin
      data_read_1_0_3_ppn <= dataBanks_3_ppn_data_read_0_3_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_0_3_perm_pf <= io_wdata_perm_pf;
    end else begin
      data_read_1_0_3_perm_pf <= dataBanks_3_perm_pf_data_read_0_3_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_0_3_perm_af <= io_wdata_perm_af;
    end else begin
      data_read_1_0_3_perm_af <= dataBanks_3_perm_af_data_read_0_3_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_0_3_perm_a <= io_wdata_perm_a;
    end else begin
      data_read_1_0_3_perm_a <= dataBanks_3_perm_a_data_read_0_3_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_0_3_perm_u <= io_wdata_perm_u;
    end else begin
      data_read_1_0_3_perm_u <= dataBanks_3_perm_u_data_read_0_3_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_0_3_perm_x <= io_wdata_perm_x;
    end else begin
      data_read_1_0_3_perm_x <= dataBanks_3_perm_x_data_read_0_3_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_0_3_perm_r <= io_wdata_perm_r;
    end else begin
      data_read_1_0_3_perm_r <= dataBanks_3_perm_rdata_read_0_3_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_0_3_perm_pm_r <= io_wdata_perm_pm_r;
    end else begin
      data_read_1_0_3_perm_pm_r <= dataBanks_3_perm_pm_rdata_read_0_3_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_0_3_perm_pm_c <= io_wdata_perm_pm_c;
    end else begin
      data_read_1_0_3_perm_pm_c <= dataBanks_3_perm_pm_c_data_read_0_3_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_0_4_tag <= io_wdata_tag;
    end else begin
      data_read_1_0_4_tag <= dataBanks_4_tag_data_read_0_4_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_0_4_asid <= io_wdata_asid;
    end else begin
      data_read_1_0_4_asid <= dataBanks_4_asid_data_read_0_4_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_0_4_ppn <= io_wdata_ppn;
    end else begin
      data_read_1_0_4_ppn <= dataBanks_4_ppn_data_read_0_4_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_0_4_perm_pf <= io_wdata_perm_pf;
    end else begin
      data_read_1_0_4_perm_pf <= dataBanks_4_perm_pf_data_read_0_4_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_0_4_perm_af <= io_wdata_perm_af;
    end else begin
      data_read_1_0_4_perm_af <= dataBanks_4_perm_af_data_read_0_4_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_0_4_perm_a <= io_wdata_perm_a;
    end else begin
      data_read_1_0_4_perm_a <= dataBanks_4_perm_a_data_read_0_4_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_0_4_perm_u <= io_wdata_perm_u;
    end else begin
      data_read_1_0_4_perm_u <= dataBanks_4_perm_u_data_read_0_4_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_0_4_perm_x <= io_wdata_perm_x;
    end else begin
      data_read_1_0_4_perm_x <= dataBanks_4_perm_x_data_read_0_4_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_0_4_perm_r <= io_wdata_perm_r;
    end else begin
      data_read_1_0_4_perm_r <= dataBanks_4_perm_rdata_read_0_4_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_0_4_perm_pm_r <= io_wdata_perm_pm_r;
    end else begin
      data_read_1_0_4_perm_pm_r <= dataBanks_4_perm_pm_rdata_read_0_4_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_0_4_perm_pm_c <= io_wdata_perm_pm_c;
    end else begin
      data_read_1_0_4_perm_pm_c <= dataBanks_4_perm_pm_c_data_read_0_4_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_0_5_tag <= io_wdata_tag;
    end else begin
      data_read_1_0_5_tag <= dataBanks_5_tag_data_read_0_5_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_0_5_asid <= io_wdata_asid;
    end else begin
      data_read_1_0_5_asid <= dataBanks_5_asid_data_read_0_5_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_0_5_ppn <= io_wdata_ppn;
    end else begin
      data_read_1_0_5_ppn <= dataBanks_5_ppn_data_read_0_5_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_0_5_perm_pf <= io_wdata_perm_pf;
    end else begin
      data_read_1_0_5_perm_pf <= dataBanks_5_perm_pf_data_read_0_5_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_0_5_perm_af <= io_wdata_perm_af;
    end else begin
      data_read_1_0_5_perm_af <= dataBanks_5_perm_af_data_read_0_5_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_0_5_perm_a <= io_wdata_perm_a;
    end else begin
      data_read_1_0_5_perm_a <= dataBanks_5_perm_a_data_read_0_5_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_0_5_perm_u <= io_wdata_perm_u;
    end else begin
      data_read_1_0_5_perm_u <= dataBanks_5_perm_u_data_read_0_5_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_0_5_perm_x <= io_wdata_perm_x;
    end else begin
      data_read_1_0_5_perm_x <= dataBanks_5_perm_x_data_read_0_5_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_0_5_perm_r <= io_wdata_perm_r;
    end else begin
      data_read_1_0_5_perm_r <= dataBanks_5_perm_rdata_read_0_5_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_0_5_perm_pm_r <= io_wdata_perm_pm_r;
    end else begin
      data_read_1_0_5_perm_pm_r <= dataBanks_5_perm_pm_rdata_read_0_5_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_0_5_perm_pm_c <= io_wdata_perm_pm_c;
    end else begin
      data_read_1_0_5_perm_pm_c <= dataBanks_5_perm_pm_c_data_read_0_5_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_0_6_tag <= io_wdata_tag;
    end else begin
      data_read_1_0_6_tag <= dataBanks_6_tag_data_read_0_6_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_0_6_asid <= io_wdata_asid;
    end else begin
      data_read_1_0_6_asid <= dataBanks_6_asid_data_read_0_6_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_0_6_ppn <= io_wdata_ppn;
    end else begin
      data_read_1_0_6_ppn <= dataBanks_6_ppn_data_read_0_6_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_0_6_perm_pf <= io_wdata_perm_pf;
    end else begin
      data_read_1_0_6_perm_pf <= dataBanks_6_perm_pf_data_read_0_6_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_0_6_perm_af <= io_wdata_perm_af;
    end else begin
      data_read_1_0_6_perm_af <= dataBanks_6_perm_af_data_read_0_6_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_0_6_perm_a <= io_wdata_perm_a;
    end else begin
      data_read_1_0_6_perm_a <= dataBanks_6_perm_a_data_read_0_6_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_0_6_perm_u <= io_wdata_perm_u;
    end else begin
      data_read_1_0_6_perm_u <= dataBanks_6_perm_u_data_read_0_6_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_0_6_perm_x <= io_wdata_perm_x;
    end else begin
      data_read_1_0_6_perm_x <= dataBanks_6_perm_x_data_read_0_6_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_0_6_perm_r <= io_wdata_perm_r;
    end else begin
      data_read_1_0_6_perm_r <= dataBanks_6_perm_rdata_read_0_6_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_0_6_perm_pm_r <= io_wdata_perm_pm_r;
    end else begin
      data_read_1_0_6_perm_pm_r <= dataBanks_6_perm_pm_rdata_read_0_6_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_0_6_perm_pm_c <= io_wdata_perm_pm_c;
    end else begin
      data_read_1_0_6_perm_pm_c <= dataBanks_6_perm_pm_c_data_read_0_6_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_0_7_tag <= io_wdata_tag;
    end else begin
      data_read_1_0_7_tag <= dataBanks_7_tag_data_read_0_7_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_0_7_asid <= io_wdata_asid;
    end else begin
      data_read_1_0_7_asid <= dataBanks_7_asid_data_read_0_7_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_0_7_ppn <= io_wdata_ppn;
    end else begin
      data_read_1_0_7_ppn <= dataBanks_7_ppn_data_read_0_7_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_0_7_perm_pf <= io_wdata_perm_pf;
    end else begin
      data_read_1_0_7_perm_pf <= dataBanks_7_perm_pf_data_read_0_7_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_0_7_perm_af <= io_wdata_perm_af;
    end else begin
      data_read_1_0_7_perm_af <= dataBanks_7_perm_af_data_read_0_7_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_0_7_perm_a <= io_wdata_perm_a;
    end else begin
      data_read_1_0_7_perm_a <= dataBanks_7_perm_a_data_read_0_7_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_0_7_perm_u <= io_wdata_perm_u;
    end else begin
      data_read_1_0_7_perm_u <= dataBanks_7_perm_u_data_read_0_7_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_0_7_perm_x <= io_wdata_perm_x;
    end else begin
      data_read_1_0_7_perm_x <= dataBanks_7_perm_x_data_read_0_7_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_0_7_perm_r <= io_wdata_perm_r;
    end else begin
      data_read_1_0_7_perm_r <= dataBanks_7_perm_rdata_read_0_7_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_0_7_perm_pm_r <= io_wdata_perm_pm_r;
    end else begin
      data_read_1_0_7_perm_pm_r <= dataBanks_7_perm_pm_rdata_read_0_7_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_0_7_perm_pm_c <= io_wdata_perm_pm_c;
    end else begin
      data_read_1_0_7_perm_pm_c <= dataBanks_7_perm_pm_c_data_read_0_7_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_1_0_ppn <= io_wdata_ppn;
    end else begin
      data_read_1_1_0_ppn <= dataBanks_0_ppn_data_read_1_0_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_1_1_ppn <= io_wdata_ppn;
    end else begin
      data_read_1_1_1_ppn <= dataBanks_1_ppn_data_read_1_1_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_1_2_ppn <= io_wdata_ppn;
    end else begin
      data_read_1_1_2_ppn <= dataBanks_2_ppn_data_read_1_2_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_1_3_ppn <= io_wdata_ppn;
    end else begin
      data_read_1_1_3_ppn <= dataBanks_3_ppn_data_read_1_3_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_1_4_ppn <= io_wdata_ppn;
    end else begin
      data_read_1_1_4_ppn <= dataBanks_4_ppn_data_read_1_4_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_1_5_ppn <= io_wdata_ppn;
    end else begin
      data_read_1_1_5_ppn <= dataBanks_5_ppn_data_read_1_5_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_1_6_ppn <= io_wdata_ppn;
    end else begin
      data_read_1_1_6_ppn <= dataBanks_6_ppn_data_read_1_6_MPORT_1_data;
    end
    if (io_wen & io_waddr == io_raddr_1) begin // @[TLBStorage.scala 68:31]
      data_read_1_1_7_ppn <= io_wdata_ppn;
    end else begin
      data_read_1_1_7_ppn <= dataBanks_7_ppn_data_read_1_7_MPORT_1_data;
    end
    bank_index_1_0 <= 8'h1 << io_raddr_1[3:1]; // @[OneHot.scala 57:35]
    bank_index_1_1 <= 8'h1 << io_raddr_1[3:1]; // @[OneHot.scala 57:35]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_0_tag[initvar] = _RAND_0[26:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_0_asid[initvar] = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_0_ppn[initvar] = _RAND_2[23:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_0_perm_pf[initvar] = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_0_perm_af[initvar] = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_0_perm_d[initvar] = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_0_perm_a[initvar] = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_0_perm_u[initvar] = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_0_perm_x[initvar] = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_0_perm_w[initvar] = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_0_perm_r[initvar] = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_0_perm_pm_r[initvar] = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_0_perm_pm_w[initvar] = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_0_perm_pm_c[initvar] = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_1_tag[initvar] = _RAND_14[26:0];
  _RAND_15 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_1_asid[initvar] = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_1_ppn[initvar] = _RAND_16[23:0];
  _RAND_17 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_1_perm_pf[initvar] = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_1_perm_af[initvar] = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_1_perm_d[initvar] = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_1_perm_a[initvar] = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_1_perm_u[initvar] = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_1_perm_x[initvar] = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_1_perm_w[initvar] = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_1_perm_r[initvar] = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_1_perm_pm_r[initvar] = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_1_perm_pm_w[initvar] = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_1_perm_pm_c[initvar] = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_2_tag[initvar] = _RAND_28[26:0];
  _RAND_29 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_2_asid[initvar] = _RAND_29[15:0];
  _RAND_30 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_2_ppn[initvar] = _RAND_30[23:0];
  _RAND_31 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_2_perm_pf[initvar] = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_2_perm_af[initvar] = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_2_perm_d[initvar] = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_2_perm_a[initvar] = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_2_perm_u[initvar] = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_2_perm_x[initvar] = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_2_perm_w[initvar] = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_2_perm_r[initvar] = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_2_perm_pm_r[initvar] = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_2_perm_pm_w[initvar] = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_2_perm_pm_c[initvar] = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_3_tag[initvar] = _RAND_42[26:0];
  _RAND_43 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_3_asid[initvar] = _RAND_43[15:0];
  _RAND_44 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_3_ppn[initvar] = _RAND_44[23:0];
  _RAND_45 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_3_perm_pf[initvar] = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_3_perm_af[initvar] = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_3_perm_d[initvar] = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_3_perm_a[initvar] = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_3_perm_u[initvar] = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_3_perm_x[initvar] = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_3_perm_w[initvar] = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_3_perm_r[initvar] = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_3_perm_pm_r[initvar] = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_3_perm_pm_w[initvar] = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_3_perm_pm_c[initvar] = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_4_tag[initvar] = _RAND_56[26:0];
  _RAND_57 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_4_asid[initvar] = _RAND_57[15:0];
  _RAND_58 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_4_ppn[initvar] = _RAND_58[23:0];
  _RAND_59 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_4_perm_pf[initvar] = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_4_perm_af[initvar] = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_4_perm_d[initvar] = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_4_perm_a[initvar] = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_4_perm_u[initvar] = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_4_perm_x[initvar] = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_4_perm_w[initvar] = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_4_perm_r[initvar] = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_4_perm_pm_r[initvar] = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_4_perm_pm_w[initvar] = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_4_perm_pm_c[initvar] = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_5_tag[initvar] = _RAND_70[26:0];
  _RAND_71 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_5_asid[initvar] = _RAND_71[15:0];
  _RAND_72 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_5_ppn[initvar] = _RAND_72[23:0];
  _RAND_73 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_5_perm_pf[initvar] = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_5_perm_af[initvar] = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_5_perm_d[initvar] = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_5_perm_a[initvar] = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_5_perm_u[initvar] = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_5_perm_x[initvar] = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_5_perm_w[initvar] = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_5_perm_r[initvar] = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_5_perm_pm_r[initvar] = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_5_perm_pm_w[initvar] = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_5_perm_pm_c[initvar] = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_6_tag[initvar] = _RAND_84[26:0];
  _RAND_85 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_6_asid[initvar] = _RAND_85[15:0];
  _RAND_86 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_6_ppn[initvar] = _RAND_86[23:0];
  _RAND_87 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_6_perm_pf[initvar] = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_6_perm_af[initvar] = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_6_perm_d[initvar] = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_6_perm_a[initvar] = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_6_perm_u[initvar] = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_6_perm_x[initvar] = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_6_perm_w[initvar] = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_6_perm_r[initvar] = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_6_perm_pm_r[initvar] = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_6_perm_pm_w[initvar] = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_6_perm_pm_c[initvar] = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_7_tag[initvar] = _RAND_98[26:0];
  _RAND_99 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_7_asid[initvar] = _RAND_99[15:0];
  _RAND_100 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_7_ppn[initvar] = _RAND_100[23:0];
  _RAND_101 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_7_perm_pf[initvar] = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_7_perm_af[initvar] = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_7_perm_d[initvar] = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_7_perm_a[initvar] = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_7_perm_u[initvar] = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_7_perm_x[initvar] = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_7_perm_w[initvar] = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_7_perm_r[initvar] = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_7_perm_pm_r[initvar] = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_7_perm_pm_w[initvar] = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    dataBanks_7_perm_pm_c[initvar] = _RAND_111[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  data_read__0_0_tag = _RAND_112[26:0];
  _RAND_113 = {1{`RANDOM}};
  data_read__0_0_asid = _RAND_113[15:0];
  _RAND_114 = {1{`RANDOM}};
  data_read__0_0_ppn = _RAND_114[23:0];
  _RAND_115 = {1{`RANDOM}};
  data_read__0_0_perm_pf = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  data_read__0_0_perm_af = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  data_read__0_0_perm_d = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  data_read__0_0_perm_a = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  data_read__0_0_perm_u = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  data_read__0_0_perm_x = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  data_read__0_0_perm_w = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  data_read__0_0_perm_r = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  data_read__0_0_perm_pm_r = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  data_read__0_0_perm_pm_w = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  data_read__0_0_perm_pm_c = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  data_read__0_1_tag = _RAND_126[26:0];
  _RAND_127 = {1{`RANDOM}};
  data_read__0_1_asid = _RAND_127[15:0];
  _RAND_128 = {1{`RANDOM}};
  data_read__0_1_ppn = _RAND_128[23:0];
  _RAND_129 = {1{`RANDOM}};
  data_read__0_1_perm_pf = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  data_read__0_1_perm_af = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  data_read__0_1_perm_d = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  data_read__0_1_perm_a = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  data_read__0_1_perm_u = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  data_read__0_1_perm_x = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  data_read__0_1_perm_w = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  data_read__0_1_perm_r = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  data_read__0_1_perm_pm_r = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  data_read__0_1_perm_pm_w = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  data_read__0_1_perm_pm_c = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  data_read__0_2_tag = _RAND_140[26:0];
  _RAND_141 = {1{`RANDOM}};
  data_read__0_2_asid = _RAND_141[15:0];
  _RAND_142 = {1{`RANDOM}};
  data_read__0_2_ppn = _RAND_142[23:0];
  _RAND_143 = {1{`RANDOM}};
  data_read__0_2_perm_pf = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  data_read__0_2_perm_af = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  data_read__0_2_perm_d = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  data_read__0_2_perm_a = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  data_read__0_2_perm_u = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  data_read__0_2_perm_x = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  data_read__0_2_perm_w = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  data_read__0_2_perm_r = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  data_read__0_2_perm_pm_r = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  data_read__0_2_perm_pm_w = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  data_read__0_2_perm_pm_c = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  data_read__0_3_tag = _RAND_154[26:0];
  _RAND_155 = {1{`RANDOM}};
  data_read__0_3_asid = _RAND_155[15:0];
  _RAND_156 = {1{`RANDOM}};
  data_read__0_3_ppn = _RAND_156[23:0];
  _RAND_157 = {1{`RANDOM}};
  data_read__0_3_perm_pf = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  data_read__0_3_perm_af = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  data_read__0_3_perm_d = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  data_read__0_3_perm_a = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  data_read__0_3_perm_u = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  data_read__0_3_perm_x = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  data_read__0_3_perm_w = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  data_read__0_3_perm_r = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  data_read__0_3_perm_pm_r = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  data_read__0_3_perm_pm_w = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  data_read__0_3_perm_pm_c = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  data_read__0_4_tag = _RAND_168[26:0];
  _RAND_169 = {1{`RANDOM}};
  data_read__0_4_asid = _RAND_169[15:0];
  _RAND_170 = {1{`RANDOM}};
  data_read__0_4_ppn = _RAND_170[23:0];
  _RAND_171 = {1{`RANDOM}};
  data_read__0_4_perm_pf = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  data_read__0_4_perm_af = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  data_read__0_4_perm_d = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  data_read__0_4_perm_a = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  data_read__0_4_perm_u = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  data_read__0_4_perm_x = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  data_read__0_4_perm_w = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  data_read__0_4_perm_r = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  data_read__0_4_perm_pm_r = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  data_read__0_4_perm_pm_w = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  data_read__0_4_perm_pm_c = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  data_read__0_5_tag = _RAND_182[26:0];
  _RAND_183 = {1{`RANDOM}};
  data_read__0_5_asid = _RAND_183[15:0];
  _RAND_184 = {1{`RANDOM}};
  data_read__0_5_ppn = _RAND_184[23:0];
  _RAND_185 = {1{`RANDOM}};
  data_read__0_5_perm_pf = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  data_read__0_5_perm_af = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  data_read__0_5_perm_d = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  data_read__0_5_perm_a = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  data_read__0_5_perm_u = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  data_read__0_5_perm_x = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  data_read__0_5_perm_w = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  data_read__0_5_perm_r = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  data_read__0_5_perm_pm_r = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  data_read__0_5_perm_pm_w = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  data_read__0_5_perm_pm_c = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  data_read__0_6_tag = _RAND_196[26:0];
  _RAND_197 = {1{`RANDOM}};
  data_read__0_6_asid = _RAND_197[15:0];
  _RAND_198 = {1{`RANDOM}};
  data_read__0_6_ppn = _RAND_198[23:0];
  _RAND_199 = {1{`RANDOM}};
  data_read__0_6_perm_pf = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  data_read__0_6_perm_af = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  data_read__0_6_perm_d = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  data_read__0_6_perm_a = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  data_read__0_6_perm_u = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  data_read__0_6_perm_x = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  data_read__0_6_perm_w = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  data_read__0_6_perm_r = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  data_read__0_6_perm_pm_r = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  data_read__0_6_perm_pm_w = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  data_read__0_6_perm_pm_c = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  data_read__0_7_tag = _RAND_210[26:0];
  _RAND_211 = {1{`RANDOM}};
  data_read__0_7_asid = _RAND_211[15:0];
  _RAND_212 = {1{`RANDOM}};
  data_read__0_7_ppn = _RAND_212[23:0];
  _RAND_213 = {1{`RANDOM}};
  data_read__0_7_perm_pf = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  data_read__0_7_perm_af = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  data_read__0_7_perm_d = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  data_read__0_7_perm_a = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  data_read__0_7_perm_u = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  data_read__0_7_perm_x = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  data_read__0_7_perm_w = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  data_read__0_7_perm_r = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  data_read__0_7_perm_pm_r = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  data_read__0_7_perm_pm_w = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  data_read__0_7_perm_pm_c = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  data_read__1_0_ppn = _RAND_224[23:0];
  _RAND_225 = {1{`RANDOM}};
  data_read__1_1_ppn = _RAND_225[23:0];
  _RAND_226 = {1{`RANDOM}};
  data_read__1_2_ppn = _RAND_226[23:0];
  _RAND_227 = {1{`RANDOM}};
  data_read__1_3_ppn = _RAND_227[23:0];
  _RAND_228 = {1{`RANDOM}};
  data_read__1_4_ppn = _RAND_228[23:0];
  _RAND_229 = {1{`RANDOM}};
  data_read__1_5_ppn = _RAND_229[23:0];
  _RAND_230 = {1{`RANDOM}};
  data_read__1_6_ppn = _RAND_230[23:0];
  _RAND_231 = {1{`RANDOM}};
  data_read__1_7_ppn = _RAND_231[23:0];
  _RAND_232 = {1{`RANDOM}};
  bank_index__0 = _RAND_232[7:0];
  _RAND_233 = {1{`RANDOM}};
  bank_index__1 = _RAND_233[7:0];
  _RAND_234 = {1{`RANDOM}};
  data_read_1_0_0_tag = _RAND_234[26:0];
  _RAND_235 = {1{`RANDOM}};
  data_read_1_0_0_asid = _RAND_235[15:0];
  _RAND_236 = {1{`RANDOM}};
  data_read_1_0_0_ppn = _RAND_236[23:0];
  _RAND_237 = {1{`RANDOM}};
  data_read_1_0_0_perm_pf = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  data_read_1_0_0_perm_af = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  data_read_1_0_0_perm_a = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  data_read_1_0_0_perm_u = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  data_read_1_0_0_perm_x = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  data_read_1_0_0_perm_r = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  data_read_1_0_0_perm_pm_r = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  data_read_1_0_0_perm_pm_c = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  data_read_1_0_1_tag = _RAND_245[26:0];
  _RAND_246 = {1{`RANDOM}};
  data_read_1_0_1_asid = _RAND_246[15:0];
  _RAND_247 = {1{`RANDOM}};
  data_read_1_0_1_ppn = _RAND_247[23:0];
  _RAND_248 = {1{`RANDOM}};
  data_read_1_0_1_perm_pf = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  data_read_1_0_1_perm_af = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  data_read_1_0_1_perm_a = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  data_read_1_0_1_perm_u = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  data_read_1_0_1_perm_x = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  data_read_1_0_1_perm_r = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  data_read_1_0_1_perm_pm_r = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  data_read_1_0_1_perm_pm_c = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  data_read_1_0_2_tag = _RAND_256[26:0];
  _RAND_257 = {1{`RANDOM}};
  data_read_1_0_2_asid = _RAND_257[15:0];
  _RAND_258 = {1{`RANDOM}};
  data_read_1_0_2_ppn = _RAND_258[23:0];
  _RAND_259 = {1{`RANDOM}};
  data_read_1_0_2_perm_pf = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  data_read_1_0_2_perm_af = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  data_read_1_0_2_perm_a = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  data_read_1_0_2_perm_u = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  data_read_1_0_2_perm_x = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  data_read_1_0_2_perm_r = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  data_read_1_0_2_perm_pm_r = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  data_read_1_0_2_perm_pm_c = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  data_read_1_0_3_tag = _RAND_267[26:0];
  _RAND_268 = {1{`RANDOM}};
  data_read_1_0_3_asid = _RAND_268[15:0];
  _RAND_269 = {1{`RANDOM}};
  data_read_1_0_3_ppn = _RAND_269[23:0];
  _RAND_270 = {1{`RANDOM}};
  data_read_1_0_3_perm_pf = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  data_read_1_0_3_perm_af = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  data_read_1_0_3_perm_a = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  data_read_1_0_3_perm_u = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  data_read_1_0_3_perm_x = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  data_read_1_0_3_perm_r = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  data_read_1_0_3_perm_pm_r = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  data_read_1_0_3_perm_pm_c = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  data_read_1_0_4_tag = _RAND_278[26:0];
  _RAND_279 = {1{`RANDOM}};
  data_read_1_0_4_asid = _RAND_279[15:0];
  _RAND_280 = {1{`RANDOM}};
  data_read_1_0_4_ppn = _RAND_280[23:0];
  _RAND_281 = {1{`RANDOM}};
  data_read_1_0_4_perm_pf = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  data_read_1_0_4_perm_af = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  data_read_1_0_4_perm_a = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  data_read_1_0_4_perm_u = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  data_read_1_0_4_perm_x = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  data_read_1_0_4_perm_r = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  data_read_1_0_4_perm_pm_r = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  data_read_1_0_4_perm_pm_c = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  data_read_1_0_5_tag = _RAND_289[26:0];
  _RAND_290 = {1{`RANDOM}};
  data_read_1_0_5_asid = _RAND_290[15:0];
  _RAND_291 = {1{`RANDOM}};
  data_read_1_0_5_ppn = _RAND_291[23:0];
  _RAND_292 = {1{`RANDOM}};
  data_read_1_0_5_perm_pf = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  data_read_1_0_5_perm_af = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  data_read_1_0_5_perm_a = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  data_read_1_0_5_perm_u = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  data_read_1_0_5_perm_x = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  data_read_1_0_5_perm_r = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  data_read_1_0_5_perm_pm_r = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  data_read_1_0_5_perm_pm_c = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  data_read_1_0_6_tag = _RAND_300[26:0];
  _RAND_301 = {1{`RANDOM}};
  data_read_1_0_6_asid = _RAND_301[15:0];
  _RAND_302 = {1{`RANDOM}};
  data_read_1_0_6_ppn = _RAND_302[23:0];
  _RAND_303 = {1{`RANDOM}};
  data_read_1_0_6_perm_pf = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  data_read_1_0_6_perm_af = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  data_read_1_0_6_perm_a = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  data_read_1_0_6_perm_u = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  data_read_1_0_6_perm_x = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  data_read_1_0_6_perm_r = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  data_read_1_0_6_perm_pm_r = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  data_read_1_0_6_perm_pm_c = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  data_read_1_0_7_tag = _RAND_311[26:0];
  _RAND_312 = {1{`RANDOM}};
  data_read_1_0_7_asid = _RAND_312[15:0];
  _RAND_313 = {1{`RANDOM}};
  data_read_1_0_7_ppn = _RAND_313[23:0];
  _RAND_314 = {1{`RANDOM}};
  data_read_1_0_7_perm_pf = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  data_read_1_0_7_perm_af = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  data_read_1_0_7_perm_a = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  data_read_1_0_7_perm_u = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  data_read_1_0_7_perm_x = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  data_read_1_0_7_perm_r = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  data_read_1_0_7_perm_pm_r = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  data_read_1_0_7_perm_pm_c = _RAND_321[0:0];
  _RAND_322 = {1{`RANDOM}};
  data_read_1_1_0_ppn = _RAND_322[23:0];
  _RAND_323 = {1{`RANDOM}};
  data_read_1_1_1_ppn = _RAND_323[23:0];
  _RAND_324 = {1{`RANDOM}};
  data_read_1_1_2_ppn = _RAND_324[23:0];
  _RAND_325 = {1{`RANDOM}};
  data_read_1_1_3_ppn = _RAND_325[23:0];
  _RAND_326 = {1{`RANDOM}};
  data_read_1_1_4_ppn = _RAND_326[23:0];
  _RAND_327 = {1{`RANDOM}};
  data_read_1_1_5_ppn = _RAND_327[23:0];
  _RAND_328 = {1{`RANDOM}};
  data_read_1_1_6_ppn = _RAND_328[23:0];
  _RAND_329 = {1{`RANDOM}};
  data_read_1_1_7_ppn = _RAND_329[23:0];
  _RAND_330 = {1{`RANDOM}};
  bank_index_1_0 = _RAND_330[7:0];
  _RAND_331 = {1{`RANDOM}};
  bank_index_1_1 = _RAND_331[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule

