module Slice(
  input          clock,
  input          reset,
  output         io_in_a_ready,
  input          io_in_a_valid,
  input  [2:0]   io_in_a_bits_opcode,
  input  [2:0]   io_in_a_bits_param,
  input  [2:0]   io_in_a_bits_size,
  input  [5:0]   io_in_a_bits_source,
  input  [35:0]  io_in_a_bits_address,
  input          io_in_a_bits_user_preferCache,
  input  [31:0]  io_in_a_bits_mask,
  input  [255:0] io_in_a_bits_data,
  input          io_in_bready,
  output         io_in_bvalid,
  output [1:0]   io_in_bparam,
  output [5:0]   io_in_bsource,
  output [35:0]  io_in_baddress,
  output [255:0] io_in_bdata,
  output         io_in_c_ready,
  input          io_in_c_valid,
  input  [2:0]   io_in_c_bits_opcode,
  input  [2:0]   io_in_c_bits_param,
  input  [2:0]   io_in_c_bits_size,
  input  [5:0]   io_in_c_bits_source,
  input  [35:0]  io_in_c_bits_address,
  input          io_in_c_bits_echo_blockisdirty,
  input  [255:0] io_in_c_bits_data,
  input          io_in_d_ready,
  output         io_in_d_valid,
  output [2:0]   io_in_d_bits_opcode,
  output [1:0]   io_in_d_bits_param,
  output [2:0]   io_in_d_bits_size,
  output [5:0]   io_in_d_bits_source,
  output [3:0]   io_in_d_bits_sink,
  output         io_in_d_bits_denied,
  output         io_in_d_bits_echo_blockisdirty,
  output [255:0] io_in_d_bits_data,
  output         io_in_d_bits_corrupt,
  input          io_in_e_valid,
  input  [3:0]   io_in_e_bits_sink,
  input          io_out_a_ready,
  output         io_out_a_valid,
  output [2:0]   io_out_a_bits_opcode,
  output [2:0]   io_out_a_bits_param,
  output [2:0]   io_out_a_bits_size,
  output [3:0]   io_out_a_bits_source,
  output [35:0]  io_out_a_bits_address,
  output [31:0]  io_out_a_bits_mask,
  output [255:0] io_out_a_bits_data,
  input          io_out_c_ready,
  output         io_out_c_valid,
  output [2:0]   io_out_c_bits_opcode,
  output [2:0]   io_out_c_bits_size,
  output [3:0]   io_out_c_bits_source,
  output [35:0]  io_out_c_bits_address,
  output [255:0] io_out_c_bits_data,
  output         io_out_d_ready,
  input          io_out_d_valid,
  input  [2:0]   io_out_d_bits_opcode,
  input  [1:0]   io_out_d_bits_param,
  input  [2:0]   io_out_d_bits_size,
  input  [3:0]   io_out_d_bits_source,
  input  [2:0]   io_out_d_bits_sink,
  input          io_out_d_bits_denied,
  input  [255:0] io_out_d_bits_data,
  output         io_out_e_valid,
  output [2:0]   io_out_e_bits_sink
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
`endif // RANDOMIZE_REG_INIT
  wire  sinkA_clock; // @[Slice.scala 56:21]
  wire  sinkA_reset; // @[Slice.scala 56:21]
  wire  sinkA_io_a_ready; // @[Slice.scala 56:21]
  wire  sinkA_io_a_valid; // @[Slice.scala 56:21]
  wire [2:0] sinkA_io_a_bits_opcode; // @[Slice.scala 56:21]
  wire [2:0] sinkA_io_a_bits_param; // @[Slice.scala 56:21]
  wire [2:0] sinkA_io_a_bits_size; // @[Slice.scala 56:21]
  wire [5:0] sinkA_io_a_bits_source; // @[Slice.scala 56:21]
  wire [35:0] sinkA_io_a_bits_address; // @[Slice.scala 56:21]
  wire  sinkA_io_a_bits_user_preferCache; // @[Slice.scala 56:21]
  wire [31:0] sinkA_io_a_bits_mask; // @[Slice.scala 56:21]
  wire [255:0] sinkA_io_a_bits_data; // @[Slice.scala 56:21]
  wire  sinkA_io_alloc_ready; // @[Slice.scala 56:21]
  wire  sinkA_io_alloc_valid; // @[Slice.scala 56:21]
  wire [2:0] sinkA_io_alloc_bits_opcode; // @[Slice.scala 56:21]
  wire [2:0] sinkA_io_alloc_bits_param; // @[Slice.scala 56:21]
  wire [2:0] sinkA_io_alloc_bits_size; // @[Slice.scala 56:21]
  wire [5:0] sinkA_io_alloc_bits_source; // @[Slice.scala 56:21]
  wire [9:0] sinkA_io_alloc_bits_set; // @[Slice.scala 56:21]
  wire [19:0] sinkA_io_alloc_bits_tag; // @[Slice.scala 56:21]
  wire [5:0] sinkA_io_alloc_bits_off; // @[Slice.scala 56:21]
  wire [31:0] sinkA_io_alloc_bits_mask; // @[Slice.scala 56:21]
  wire [2:0] sinkA_io_alloc_bits_bufIdx; // @[Slice.scala 56:21]
  wire  sinkA_io_alloc_bits_preferCache; // @[Slice.scala 56:21]
  wire  sinkA_io_d_pb_pop_ready; // @[Slice.scala 56:21]
  wire  sinkA_io_d_pb_pop_valid; // @[Slice.scala 56:21]
  wire [2:0] sinkA_io_d_pb_pop_bits_bufIdx; // @[Slice.scala 56:21]
  wire  sinkA_io_d_pb_pop_bits_count; // @[Slice.scala 56:21]
  wire  sinkA_io_d_pb_pop_bits_last; // @[Slice.scala 56:21]
  wire [255:0] sinkA_io_d_pb_beat_data; // @[Slice.scala 56:21]
  wire [31:0] sinkA_io_d_pb_beat_mask; // @[Slice.scala 56:21]
  wire  sinkA_io_a_pb_pop_ready; // @[Slice.scala 56:21]
  wire  sinkA_io_a_pb_pop_valid; // @[Slice.scala 56:21]
  wire [2:0] sinkA_io_a_pb_pop_bits_bufIdx; // @[Slice.scala 56:21]
  wire  sinkA_io_a_pb_pop_bits_count; // @[Slice.scala 56:21]
  wire  sinkA_io_a_pb_pop_bits_last; // @[Slice.scala 56:21]
  wire [255:0] sinkA_io_a_pb_beat_data; // @[Slice.scala 56:21]
  wire [31:0] sinkA_io_a_pb_beat_mask; // @[Slice.scala 56:21]
  wire  sourceB_clock; // @[Slice.scala 57:23]
  wire  sourceB_reset; // @[Slice.scala 57:23]
  wire  sourceB_io_bready; // @[Slice.scala 57:23]
  wire  sourceB_io_bvalid; // @[Slice.scala 57:23]
  wire [1:0] sourceB_io_bparam; // @[Slice.scala 57:23]
  wire [5:0] sourceB_io_bsource; // @[Slice.scala 57:23]
  wire [35:0] sourceB_io_baddress; // @[Slice.scala 57:23]
  wire [255:0] sourceB_io_bdata; // @[Slice.scala 57:23]
  wire  sourceB_io_task_ready; // @[Slice.scala 57:23]
  wire  sourceB_io_task_valid; // @[Slice.scala 57:23]
  wire [9:0] sourceB_io_task_bits_set; // @[Slice.scala 57:23]
  wire [19:0] sourceB_io_task_bits_tag; // @[Slice.scala 57:23]
  wire [2:0] sourceB_io_task_bits_param; // @[Slice.scala 57:23]
  wire [1:0] sourceB_io_task_bits_clients; // @[Slice.scala 57:23]
  wire  sourceB_io_task_bits_needData; // @[Slice.scala 57:23]
  wire  sinkC_clock; // @[Slice.scala 58:21]
  wire  sinkC_reset; // @[Slice.scala 58:21]
  wire  sinkC_io_c_ready; // @[Slice.scala 58:21]
  wire  sinkC_io_c_valid; // @[Slice.scala 58:21]
  wire [2:0] sinkC_io_c_bits_opcode; // @[Slice.scala 58:21]
  wire [2:0] sinkC_io_c_bits_param; // @[Slice.scala 58:21]
  wire [2:0] sinkC_io_c_bits_size; // @[Slice.scala 58:21]
  wire [5:0] sinkC_io_c_bits_source; // @[Slice.scala 58:21]
  wire [35:0] sinkC_io_c_bits_address; // @[Slice.scala 58:21]
  wire  sinkC_io_c_bits_echo_blockisdirty; // @[Slice.scala 58:21]
  wire [255:0] sinkC_io_c_bits_data; // @[Slice.scala 58:21]
  wire  sinkC_io_alloc_ready; // @[Slice.scala 58:21]
  wire  sinkC_io_alloc_valid; // @[Slice.scala 58:21]
  wire [2:0] sinkC_io_alloc_bits_opcode; // @[Slice.scala 58:21]
  wire [2:0] sinkC_io_alloc_bits_param; // @[Slice.scala 58:21]
  wire [2:0] sinkC_io_alloc_bits_size; // @[Slice.scala 58:21]
  wire [5:0] sinkC_io_alloc_bits_source; // @[Slice.scala 58:21]
  wire [9:0] sinkC_io_alloc_bits_set; // @[Slice.scala 58:21]
  wire [19:0] sinkC_io_alloc_bits_tag; // @[Slice.scala 58:21]
  wire [5:0] sinkC_io_alloc_bits_off; // @[Slice.scala 58:21]
  wire [2:0] sinkC_io_alloc_bits_bufIdx; // @[Slice.scala 58:21]
  wire  sinkC_io_alloc_bits_dirty; // @[Slice.scala 58:21]
  wire  sinkC_io_resp_valid; // @[Slice.scala 58:21]
  wire  sinkC_io_resp_bits_hasData; // @[Slice.scala 58:21]
  wire [2:0] sinkC_io_resp_bits_param; // @[Slice.scala 58:21]
  wire [5:0] sinkC_io_resp_bits_source; // @[Slice.scala 58:21]
  wire  sinkC_io_resp_bits_last; // @[Slice.scala 58:21]
  wire [9:0] sinkC_io_resp_bits_set; // @[Slice.scala 58:21]
  wire [2:0] sinkC_io_resp_bits_bufIdx; // @[Slice.scala 58:21]
  wire  sinkC_io_task_ready; // @[Slice.scala 58:21]
  wire  sinkC_io_task_valid; // @[Slice.scala 58:21]
  wire [9:0] sinkC_io_task_bits_set; // @[Slice.scala 58:21]
  wire [19:0] sinkC_io_task_bits_tag; // @[Slice.scala 58:21]
  wire [2:0] sinkC_io_task_bits_way; // @[Slice.scala 58:21]
  wire [2:0] sinkC_io_task_bits_bufIdx; // @[Slice.scala 58:21]
  wire [2:0] sinkC_io_task_bits_opcode; // @[Slice.scala 58:21]
  wire [3:0] sinkC_io_task_bits_source; // @[Slice.scala 58:21]
  wire  sinkC_io_task_bits_save; // @[Slice.scala 58:21]
  wire  sinkC_io_task_bits_drop; // @[Slice.scala 58:21]
  wire  sinkC_io_task_bits_release; // @[Slice.scala 58:21]
  wire  sinkC_io_bs_waddr_ready; // @[Slice.scala 58:21]
  wire  sinkC_io_bs_waddr_valid; // @[Slice.scala 58:21]
  wire [2:0] sinkC_io_bs_waddr_bits_way; // @[Slice.scala 58:21]
  wire [9:0] sinkC_io_bs_waddr_bits_set; // @[Slice.scala 58:21]
  wire  sinkC_io_bs_waddr_bits_beat; // @[Slice.scala 58:21]
  wire  sinkC_io_bs_waddr_bits_noop; // @[Slice.scala 58:21]
  wire [255:0] sinkC_io_bs_wdata_data; // @[Slice.scala 58:21]
  wire  sinkC_io_sourceD_rhazard_valid; // @[Slice.scala 58:21]
  wire [2:0] sinkC_io_sourceD_rhazard_bits_way; // @[Slice.scala 58:21]
  wire [9:0] sinkC_io_sourceD_rhazard_bits_set; // @[Slice.scala 58:21]
  wire  sinkC_io_release_ready; // @[Slice.scala 58:21]
  wire  sinkC_io_release_valid; // @[Slice.scala 58:21]
  wire [2:0] sinkC_io_release_bits_opcode; // @[Slice.scala 58:21]
  wire [3:0] sinkC_io_release_bits_source; // @[Slice.scala 58:21]
  wire [35:0] sinkC_io_release_bits_address; // @[Slice.scala 58:21]
  wire [255:0] sinkC_io_release_bits_data; // @[Slice.scala 58:21]
  wire  sourceD_clock; // @[Slice.scala 59:23]
  wire  sourceD_reset; // @[Slice.scala 59:23]
  wire  sourceD_io_d_ready; // @[Slice.scala 59:23]
  wire  sourceD_io_d_valid; // @[Slice.scala 59:23]
  wire [2:0] sourceD_io_d_bits_opcode; // @[Slice.scala 59:23]
  wire [1:0] sourceD_io_d_bits_param; // @[Slice.scala 59:23]
  wire [2:0] sourceD_io_d_bits_size; // @[Slice.scala 59:23]
  wire [5:0] sourceD_io_d_bits_source; // @[Slice.scala 59:23]
  wire [3:0] sourceD_io_d_bits_sink; // @[Slice.scala 59:23]
  wire  sourceD_io_d_bits_denied; // @[Slice.scala 59:23]
  wire  sourceD_io_d_bits_echo_blockisdirty; // @[Slice.scala 59:23]
  wire [255:0] sourceD_io_d_bits_data; // @[Slice.scala 59:23]
  wire  sourceD_io_d_bits_corrupt; // @[Slice.scala 59:23]
  wire  sourceD_io_task_ready; // @[Slice.scala 59:23]
  wire  sourceD_io_task_valid; // @[Slice.scala 59:23]
  wire [5:0] sourceD_io_task_bits_sourceId; // @[Slice.scala 59:23]
  wire [9:0] sourceD_io_task_bits_set; // @[Slice.scala 59:23]
  wire [2:0] sourceD_io_task_bits_channel; // @[Slice.scala 59:23]
  wire [2:0] sourceD_io_task_bits_opcode; // @[Slice.scala 59:23]
  wire [2:0] sourceD_io_task_bits_param; // @[Slice.scala 59:23]
  wire [2:0] sourceD_io_task_bits_size; // @[Slice.scala 59:23]
  wire [2:0] sourceD_io_task_bits_way; // @[Slice.scala 59:23]
  wire [5:0] sourceD_io_task_bits_off; // @[Slice.scala 59:23]
  wire  sourceD_io_task_bits_useBypass; // @[Slice.scala 59:23]
  wire [2:0] sourceD_io_task_bits_bufIdx; // @[Slice.scala 59:23]
  wire  sourceD_io_task_bits_denied; // @[Slice.scala 59:23]
  wire [3:0] sourceD_io_task_bits_sinkId; // @[Slice.scala 59:23]
  wire  sourceD_io_task_bits_bypassPut; // @[Slice.scala 59:23]
  wire  sourceD_io_task_bits_dirty; // @[Slice.scala 59:23]
  wire  sourceD_io_bs_raddr_ready; // @[Slice.scala 59:23]
  wire  sourceD_io_bs_raddr_valid; // @[Slice.scala 59:23]
  wire [2:0] sourceD_io_bs_raddr_bits_way; // @[Slice.scala 59:23]
  wire [9:0] sourceD_io_bs_raddr_bits_set; // @[Slice.scala 59:23]
  wire  sourceD_io_bs_raddr_bits_beat; // @[Slice.scala 59:23]
  wire [255:0] sourceD_io_bs_rdata_data; // @[Slice.scala 59:23]
  wire  sourceD_io_bypass_read_valid; // @[Slice.scala 59:23]
  wire  sourceD_io_bypass_read_beat; // @[Slice.scala 59:23]
  wire [2:0] sourceD_io_bypass_read_id; // @[Slice.scala 59:23]
  wire  sourceD_io_bypass_read_ready; // @[Slice.scala 59:23]
  wire [255:0] sourceD_io_bypass_read_buffer_data_data; // @[Slice.scala 59:23]
  wire  sourceD_io_bypass_read_last; // @[Slice.scala 59:23]
  wire  sourceD_io_bs_waddr_ready; // @[Slice.scala 59:23]
  wire  sourceD_io_bs_waddr_valid; // @[Slice.scala 59:23]
  wire [2:0] sourceD_io_bs_waddr_bits_way; // @[Slice.scala 59:23]
  wire [9:0] sourceD_io_bs_waddr_bits_set; // @[Slice.scala 59:23]
  wire  sourceD_io_bs_waddr_bits_beat; // @[Slice.scala 59:23]
  wire [255:0] sourceD_io_bs_wdata_data; // @[Slice.scala 59:23]
  wire  sourceD_io_sourceD_rhazard_valid; // @[Slice.scala 59:23]
  wire [2:0] sourceD_io_sourceD_rhazard_bits_way; // @[Slice.scala 59:23]
  wire [9:0] sourceD_io_sourceD_rhazard_bits_set; // @[Slice.scala 59:23]
  wire  sourceD_io_pb_pop_ready; // @[Slice.scala 59:23]
  wire  sourceD_io_pb_pop_valid; // @[Slice.scala 59:23]
  wire [2:0] sourceD_io_pb_pop_bits_bufIdx; // @[Slice.scala 59:23]
  wire  sourceD_io_pb_pop_bits_count; // @[Slice.scala 59:23]
  wire  sourceD_io_pb_pop_bits_last; // @[Slice.scala 59:23]
  wire [255:0] sourceD_io_pb_beat_data; // @[Slice.scala 59:23]
  wire [31:0] sourceD_io_pb_beat_mask; // @[Slice.scala 59:23]
  wire  sourceD_io_resp_valid; // @[Slice.scala 59:23]
  wire [3:0] sourceD_io_resp_bits_sink; // @[Slice.scala 59:23]
  wire  sinkE_io_e_ready; // @[Slice.scala 60:21]
  wire  sinkE_io_e_valid; // @[Slice.scala 60:21]
  wire [3:0] sinkE_io_e_bits_sink; // @[Slice.scala 60:21]
  wire  sinkE_io_resp_valid; // @[Slice.scala 60:21]
  wire [3:0] sinkE_io_resp_bits_sink; // @[Slice.scala 60:21]
  wire  sourceA_clock; // @[Slice.scala 70:23]
  wire  sourceA_reset; // @[Slice.scala 70:23]
  wire  sourceA_io_a_ready; // @[Slice.scala 70:23]
  wire  sourceA_io_a_valid; // @[Slice.scala 70:23]
  wire [2:0] sourceA_io_a_bits_opcode; // @[Slice.scala 70:23]
  wire [2:0] sourceA_io_a_bits_param; // @[Slice.scala 70:23]
  wire [2:0] sourceA_io_a_bits_size; // @[Slice.scala 70:23]
  wire [3:0] sourceA_io_a_bits_source; // @[Slice.scala 70:23]
  wire [35:0] sourceA_io_a_bits_address; // @[Slice.scala 70:23]
  wire [31:0] sourceA_io_a_bits_mask; // @[Slice.scala 70:23]
  wire [255:0] sourceA_io_a_bits_data; // @[Slice.scala 70:23]
  wire  sourceA_io_task_ready; // @[Slice.scala 70:23]
  wire  sourceA_io_task_valid; // @[Slice.scala 70:23]
  wire [19:0] sourceA_io_task_bits_tag; // @[Slice.scala 70:23]
  wire [9:0] sourceA_io_task_bits_set; // @[Slice.scala 70:23]
  wire [5:0] sourceA_io_task_bits_off; // @[Slice.scala 70:23]
  wire [2:0] sourceA_io_task_bits_opcode; // @[Slice.scala 70:23]
  wire [2:0] sourceA_io_task_bits_param; // @[Slice.scala 70:23]
  wire [3:0] sourceA_io_task_bits_source; // @[Slice.scala 70:23]
  wire [2:0] sourceA_io_task_bits_bufIdx; // @[Slice.scala 70:23]
  wire [2:0] sourceA_io_task_bits_size; // @[Slice.scala 70:23]
  wire  sourceA_io_task_bits_putData; // @[Slice.scala 70:23]
  wire  sourceA_io_pb_pop_ready; // @[Slice.scala 70:23]
  wire  sourceA_io_pb_pop_valid; // @[Slice.scala 70:23]
  wire [2:0] sourceA_io_pb_pop_bits_bufIdx; // @[Slice.scala 70:23]
  wire  sourceA_io_pb_pop_bits_count; // @[Slice.scala 70:23]
  wire  sourceA_io_pb_pop_bits_last; // @[Slice.scala 70:23]
  wire [255:0] sourceA_io_pb_beat_data; // @[Slice.scala 70:23]
  wire [31:0] sourceA_io_pb_beat_mask; // @[Slice.scala 70:23]
  wire  sinkB_io_bready; // @[Slice.scala 71:21]
  wire  sinkB_io_bvalid; // @[Slice.scala 71:21]
  wire [2:0] sinkB_io_bopcode; // @[Slice.scala 71:21]
  wire [1:0] sinkB_io_bparam; // @[Slice.scala 71:21]
  wire [2:0] sinkB_io_bsize; // @[Slice.scala 71:21]
  wire [3:0] sinkB_io_bsource; // @[Slice.scala 71:21]
  wire [35:0] sinkB_io_baddress; // @[Slice.scala 71:21]
  wire [31:0] sinkB_io_bmask; // @[Slice.scala 71:21]
  wire [255:0] sinkB_io_bdata; // @[Slice.scala 71:21]
  wire  sinkB_io_alloc_ready; // @[Slice.scala 71:21]
  wire  sinkB_io_alloc_valid; // @[Slice.scala 71:21]
  wire [2:0] sinkB_io_alloc_bits_opcode; // @[Slice.scala 71:21]
  wire [2:0] sinkB_io_alloc_bits_param; // @[Slice.scala 71:21]
  wire [2:0] sinkB_io_alloc_bits_size; // @[Slice.scala 71:21]
  wire [5:0] sinkB_io_alloc_bits_source; // @[Slice.scala 71:21]
  wire [9:0] sinkB_io_alloc_bits_set; // @[Slice.scala 71:21]
  wire [19:0] sinkB_io_alloc_bits_tag; // @[Slice.scala 71:21]
  wire [5:0] sinkB_io_alloc_bits_off; // @[Slice.scala 71:21]
  wire [31:0] sinkB_io_alloc_bits_mask; // @[Slice.scala 71:21]
  wire  sinkB_io_alloc_bits_needProbeAckData; // @[Slice.scala 71:21]
  wire  sourceC_clock; // @[Slice.scala 72:23]
  wire  sourceC_reset; // @[Slice.scala 72:23]
  wire  sourceC_io_c_ready; // @[Slice.scala 72:23]
  wire  sourceC_io_c_valid; // @[Slice.scala 72:23]
  wire [2:0] sourceC_io_c_bits_opcode; // @[Slice.scala 72:23]
  wire [2:0] sourceC_io_c_bits_size; // @[Slice.scala 72:23]
  wire [3:0] sourceC_io_c_bits_source; // @[Slice.scala 72:23]
  wire [35:0] sourceC_io_c_bits_address; // @[Slice.scala 72:23]
  wire [255:0] sourceC_io_c_bits_data; // @[Slice.scala 72:23]
  wire  sourceC_io_bs_raddr_ready; // @[Slice.scala 72:23]
  wire  sourceC_io_bs_raddr_valid; // @[Slice.scala 72:23]
  wire [2:0] sourceC_io_bs_raddr_bits_way; // @[Slice.scala 72:23]
  wire [9:0] sourceC_io_bs_raddr_bits_set; // @[Slice.scala 72:23]
  wire  sourceC_io_bs_raddr_bits_beat; // @[Slice.scala 72:23]
  wire [255:0] sourceC_io_bs_rdata_data; // @[Slice.scala 72:23]
  wire  sourceC_io_task_ready; // @[Slice.scala 72:23]
  wire  sourceC_io_task_valid; // @[Slice.scala 72:23]
  wire [2:0] sourceC_io_task_bits_opcode; // @[Slice.scala 72:23]
  wire [19:0] sourceC_io_task_bits_tag; // @[Slice.scala 72:23]
  wire [9:0] sourceC_io_task_bits_set; // @[Slice.scala 72:23]
  wire [3:0] sourceC_io_task_bits_source; // @[Slice.scala 72:23]
  wire [2:0] sourceC_io_task_bits_way; // @[Slice.scala 72:23]
  wire  sinkD_clock; // @[Slice.scala 73:21]
  wire  sinkD_reset; // @[Slice.scala 73:21]
  wire  sinkD_io_d_ready; // @[Slice.scala 73:21]
  wire  sinkD_io_d_valid; // @[Slice.scala 73:21]
  wire [2:0] sinkD_io_d_bits_opcode; // @[Slice.scala 73:21]
  wire [1:0] sinkD_io_d_bits_param; // @[Slice.scala 73:21]
  wire [2:0] sinkD_io_d_bits_size; // @[Slice.scala 73:21]
  wire [3:0] sinkD_io_d_bits_source; // @[Slice.scala 73:21]
  wire [2:0] sinkD_io_d_bits_sink; // @[Slice.scala 73:21]
  wire  sinkD_io_d_bits_denied; // @[Slice.scala 73:21]
  wire [255:0] sinkD_io_d_bits_data; // @[Slice.scala 73:21]
  wire  sinkD_io_bs_waddr_ready; // @[Slice.scala 73:21]
  wire  sinkD_io_bs_waddr_valid; // @[Slice.scala 73:21]
  wire [2:0] sinkD_io_bs_waddr_bits_way; // @[Slice.scala 73:21]
  wire [9:0] sinkD_io_bs_waddr_bits_set; // @[Slice.scala 73:21]
  wire  sinkD_io_bs_waddr_bits_beat; // @[Slice.scala 73:21]
  wire  sinkD_io_bs_waddr_bits_noop; // @[Slice.scala 73:21]
  wire [255:0] sinkD_io_bs_wdata_data; // @[Slice.scala 73:21]
  wire  sinkD_io_bypass_write_valid; // @[Slice.scala 73:21]
  wire  sinkD_io_bypass_write_beat; // @[Slice.scala 73:21]
  wire [255:0] sinkD_io_bypass_write_data_data; // @[Slice.scala 73:21]
  wire  sinkD_io_bypass_write_ready; // @[Slice.scala 73:21]
  wire [2:0] sinkD_io_bypass_write_id; // @[Slice.scala 73:21]
  wire [2:0] sinkD_io_way; // @[Slice.scala 73:21]
  wire [9:0] sinkD_io_set; // @[Slice.scala 73:21]
  wire  sinkD_io_inner_grant; // @[Slice.scala 73:21]
  wire  sinkD_io_save_data_in_bs; // @[Slice.scala 73:21]
  wire  sinkD_io_resp_valid; // @[Slice.scala 73:21]
  wire [2:0] sinkD_io_resp_bits_opcode; // @[Slice.scala 73:21]
  wire [2:0] sinkD_io_resp_bits_param; // @[Slice.scala 73:21]
  wire [3:0] sinkD_io_resp_bits_source; // @[Slice.scala 73:21]
  wire [2:0] sinkD_io_resp_bits_sink; // @[Slice.scala 73:21]
  wire  sinkD_io_resp_bits_last; // @[Slice.scala 73:21]
  wire  sinkD_io_resp_bits_denied; // @[Slice.scala 73:21]
  wire [2:0] sinkD_io_resp_bits_bufIdx; // @[Slice.scala 73:21]
  wire  sinkD_io_sourceD_rhazard_valid; // @[Slice.scala 73:21]
  wire [2:0] sinkD_io_sourceD_rhazard_bits_way; // @[Slice.scala 73:21]
  wire [9:0] sinkD_io_sourceD_rhazard_bits_set; // @[Slice.scala 73:21]
  wire  sourceE_io_e_ready; // @[Slice.scala 74:23]
  wire  sourceE_io_e_valid; // @[Slice.scala 74:23]
  wire [2:0] sourceE_io_e_bits_sink; // @[Slice.scala 74:23]
  wire  sourceE_io_task_ready; // @[Slice.scala 74:23]
  wire  sourceE_io_task_valid; // @[Slice.scala 74:23]
  wire [2:0] sourceE_io_task_bits_sink; // @[Slice.scala 74:23]
  wire  refillBuffer_clock; // @[Slice.scala 76:28]
  wire  refillBuffer_reset; // @[Slice.scala 76:28]
  wire  refillBuffer_io_rvalid; // @[Slice.scala 76:28]
  wire  refillBuffer_io_rbeat; // @[Slice.scala 76:28]
  wire [2:0] refillBuffer_io_rid; // @[Slice.scala 76:28]
  wire  refillBuffer_io_rready; // @[Slice.scala 76:28]
  wire [255:0] refillBuffer_io_rbuffer_data_data; // @[Slice.scala 76:28]
  wire  refillBuffer_io_rlast; // @[Slice.scala 76:28]
  wire  refillBuffer_io_wvalid; // @[Slice.scala 76:28]
  wire  refillBuffer_io_wbeat; // @[Slice.scala 76:28]
  wire [255:0] refillBuffer_io_wdata_data; // @[Slice.scala 76:28]
  wire  refillBuffer_io_wready; // @[Slice.scala 76:28]
  wire [2:0] refillBuffer_io_wid; // @[Slice.scala 76:28]
  wire  io_out_a_q_clock; // @[Decoupled.scala 361:21]
  wire  io_out_a_q_reset; // @[Decoupled.scala 361:21]
  wire  io_out_a_q_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  io_out_a_q_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [2:0] io_out_a_q_io_enq_bits_opcode; // @[Decoupled.scala 361:21]
  wire [2:0] io_out_a_q_io_enq_bits_param; // @[Decoupled.scala 361:21]
  wire [2:0] io_out_a_q_io_enq_bits_size; // @[Decoupled.scala 361:21]
  wire [3:0] io_out_a_q_io_enq_bits_source; // @[Decoupled.scala 361:21]
  wire [35:0] io_out_a_q_io_enq_bits_address; // @[Decoupled.scala 361:21]
  wire [31:0] io_out_a_q_io_enq_bits_mask; // @[Decoupled.scala 361:21]
  wire [255:0] io_out_a_q_io_enq_bits_data; // @[Decoupled.scala 361:21]
  wire  io_out_a_q_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  io_out_a_q_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [2:0] io_out_a_q_io_deq_bits_opcode; // @[Decoupled.scala 361:21]
  wire [2:0] io_out_a_q_io_deq_bits_param; // @[Decoupled.scala 361:21]
  wire [2:0] io_out_a_q_io_deq_bits_size; // @[Decoupled.scala 361:21]
  wire [3:0] io_out_a_q_io_deq_bits_source; // @[Decoupled.scala 361:21]
  wire [35:0] io_out_a_q_io_deq_bits_address; // @[Decoupled.scala 361:21]
  wire [31:0] io_out_a_q_io_deq_bits_mask; // @[Decoupled.scala 361:21]
  wire [255:0] io_out_a_q_io_deq_bits_data; // @[Decoupled.scala 361:21]
  wire  sinkB_io_bq_clock; // @[Decoupled.scala 361:21]
  wire  sinkB_io_bq_reset; // @[Decoupled.scala 361:21]
  wire  sinkB_io_bq_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  sinkB_io_bq_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [2:0] sinkB_io_bq_io_enq_bits_opcode; // @[Decoupled.scala 361:21]
  wire [1:0] sinkB_io_bq_io_enq_bits_param; // @[Decoupled.scala 361:21]
  wire [2:0] sinkB_io_bq_io_enq_bits_size; // @[Decoupled.scala 361:21]
  wire [3:0] sinkB_io_bq_io_enq_bits_source; // @[Decoupled.scala 361:21]
  wire [35:0] sinkB_io_bq_io_enq_bits_address; // @[Decoupled.scala 361:21]
  wire [31:0] sinkB_io_bq_io_enq_bits_mask; // @[Decoupled.scala 361:21]
  wire [255:0] sinkB_io_bq_io_enq_bits_data; // @[Decoupled.scala 361:21]
  wire  sinkB_io_bq_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  sinkB_io_bq_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [2:0] sinkB_io_bq_io_deq_bits_opcode; // @[Decoupled.scala 361:21]
  wire [1:0] sinkB_io_bq_io_deq_bits_param; // @[Decoupled.scala 361:21]
  wire [2:0] sinkB_io_bq_io_deq_bits_size; // @[Decoupled.scala 361:21]
  wire [3:0] sinkB_io_bq_io_deq_bits_source; // @[Decoupled.scala 361:21]
  wire [35:0] sinkB_io_bq_io_deq_bits_address; // @[Decoupled.scala 361:21]
  wire [31:0] sinkB_io_bq_io_deq_bits_mask; // @[Decoupled.scala 361:21]
  wire [255:0] sinkB_io_bq_io_deq_bits_data; // @[Decoupled.scala 361:21]
  wire  io_out_c_q_clock; // @[Decoupled.scala 361:21]
  wire  io_out_c_q_reset; // @[Decoupled.scala 361:21]
  wire  io_out_c_q_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  io_out_c_q_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [2:0] io_out_c_q_io_enq_bits_opcode; // @[Decoupled.scala 361:21]
  wire [2:0] io_out_c_q_io_enq_bits_size; // @[Decoupled.scala 361:21]
  wire [3:0] io_out_c_q_io_enq_bits_source; // @[Decoupled.scala 361:21]
  wire [35:0] io_out_c_q_io_enq_bits_address; // @[Decoupled.scala 361:21]
  wire [255:0] io_out_c_q_io_enq_bits_data; // @[Decoupled.scala 361:21]
  wire  io_out_c_q_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  io_out_c_q_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [2:0] io_out_c_q_io_deq_bits_opcode; // @[Decoupled.scala 361:21]
  wire [2:0] io_out_c_q_io_deq_bits_size; // @[Decoupled.scala 361:21]
  wire [3:0] io_out_c_q_io_deq_bits_source; // @[Decoupled.scala 361:21]
  wire [35:0] io_out_c_q_io_deq_bits_address; // @[Decoupled.scala 361:21]
  wire [255:0] io_out_c_q_io_deq_bits_data; // @[Decoupled.scala 361:21]
  wire  sinkD_io_d_q_clock; // @[Decoupled.scala 361:21]
  wire  sinkD_io_d_q_reset; // @[Decoupled.scala 361:21]
  wire  sinkD_io_d_q_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  sinkD_io_d_q_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [2:0] sinkD_io_d_q_io_enq_bits_opcode; // @[Decoupled.scala 361:21]
  wire [1:0] sinkD_io_d_q_io_enq_bits_param; // @[Decoupled.scala 361:21]
  wire [2:0] sinkD_io_d_q_io_enq_bits_size; // @[Decoupled.scala 361:21]
  wire [3:0] sinkD_io_d_q_io_enq_bits_source; // @[Decoupled.scala 361:21]
  wire [2:0] sinkD_io_d_q_io_enq_bits_sink; // @[Decoupled.scala 361:21]
  wire  sinkD_io_d_q_io_enq_bits_denied; // @[Decoupled.scala 361:21]
  wire [255:0] sinkD_io_d_q_io_enq_bits_data; // @[Decoupled.scala 361:21]
  wire  sinkD_io_d_q_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  sinkD_io_d_q_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [2:0] sinkD_io_d_q_io_deq_bits_opcode; // @[Decoupled.scala 361:21]
  wire [1:0] sinkD_io_d_q_io_deq_bits_param; // @[Decoupled.scala 361:21]
  wire [2:0] sinkD_io_d_q_io_deq_bits_size; // @[Decoupled.scala 361:21]
  wire [3:0] sinkD_io_d_q_io_deq_bits_source; // @[Decoupled.scala 361:21]
  wire [2:0] sinkD_io_d_q_io_deq_bits_sink; // @[Decoupled.scala 361:21]
  wire  sinkD_io_d_q_io_deq_bits_denied; // @[Decoupled.scala 361:21]
  wire [255:0] sinkD_io_d_q_io_deq_bits_data; // @[Decoupled.scala 361:21]
  wire  io_out_e_q_clock; // @[Decoupled.scala 361:21]
  wire  io_out_e_q_reset; // @[Decoupled.scala 361:21]
  wire  io_out_e_q_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  io_out_e_q_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [2:0] io_out_e_q_io_enq_bits_sink; // @[Decoupled.scala 361:21]
  wire  io_out_e_q_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [2:0] io_out_e_q_io_deq_bits_sink; // @[Decoupled.scala 361:21]
  wire  abc_mshr_0_clock; // @[Slice.scala 94:16]
  wire  abc_mshr_0_reset; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_0_io_id; // @[Slice.scala 94:16]
  wire  abc_mshr_0_io_enable; // @[Slice.scala 94:16]
  wire  abc_mshr_0_io_alloc_valid; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_0_io_alloc_bits_channel; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_0_io_alloc_bits_opcode; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_0_io_alloc_bits_param; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_0_io_alloc_bits_size; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_0_io_alloc_bits_source; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_0_io_alloc_bits_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_0_io_alloc_bits_tag; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_0_io_alloc_bits_off; // @[Slice.scala 94:16]
  wire [31:0] abc_mshr_0_io_alloc_bits_mask; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_0_io_alloc_bits_bufIdx; // @[Slice.scala 94:16]
  wire  abc_mshr_0_io_alloc_bits_preferCache; // @[Slice.scala 94:16]
  wire  abc_mshr_0_io_alloc_bits_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_0_io_alloc_bits_fromProbeHelper; // @[Slice.scala 94:16]
  wire  abc_mshr_0_io_alloc_bits_fromCmoHelper; // @[Slice.scala 94:16]
  wire  abc_mshr_0_io_alloc_bits_needProbeAckData; // @[Slice.scala 94:16]
  wire  abc_mshr_0_io_status_valid; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_0_io_status_bits_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_0_io_status_bits_tag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_0_io_status_bits_way; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_0_io_status_bits_way_reg; // @[Slice.scala 94:16]
  wire  abc_mshr_0_io_status_bits_nestB; // @[Slice.scala 94:16]
  wire  abc_mshr_0_io_status_bits_nestC; // @[Slice.scala 94:16]
  wire  abc_mshr_0_io_status_bits_will_grant_data; // @[Slice.scala 94:16]
  wire  abc_mshr_0_io_status_bits_will_save_data; // @[Slice.scala 94:16]
  wire  abc_mshr_0_io_status_bits_will_free; // @[Slice.scala 94:16]
  wire  abc_mshr_0_io_resps_sink_c_valid; // @[Slice.scala 94:16]
  wire  abc_mshr_0_io_resps_sink_c_bits_hasData; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_0_io_resps_sink_c_bits_param; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_0_io_resps_sink_c_bits_source; // @[Slice.scala 94:16]
  wire  abc_mshr_0_io_resps_sink_c_bits_last; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_0_io_resps_sink_c_bits_bufIdx; // @[Slice.scala 94:16]
  wire  abc_mshr_0_io_resps_sink_d_valid; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_0_io_resps_sink_d_bits_opcode; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_0_io_resps_sink_d_bits_param; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_0_io_resps_sink_d_bits_sink; // @[Slice.scala 94:16]
  wire  abc_mshr_0_io_resps_sink_d_bits_last; // @[Slice.scala 94:16]
  wire  abc_mshr_0_io_resps_sink_d_bits_denied; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_0_io_resps_sink_d_bits_bufIdx; // @[Slice.scala 94:16]
  wire  abc_mshr_0_io_resps_sink_e_valid; // @[Slice.scala 94:16]
  wire  abc_mshr_0_io_resps_source_d_valid; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_0_io_nestedwb_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_0_io_nestedwb_tag; // @[Slice.scala 94:16]
  wire  abc_mshr_0_io_nestedwb_btoN; // @[Slice.scala 94:16]
  wire  abc_mshr_0_io_nestedwb_btoB; // @[Slice.scala 94:16]
  wire  abc_mshr_0_io_nestedwb_bclr_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_0_io_nestedwb_bset_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_0_io_nestedwb_c_set_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_0_io_nestedwb_c_set_hit; // @[Slice.scala 94:16]
  wire  abc_mshr_0_io_nestedwb_clients_0_isToN; // @[Slice.scala 94:16]
  wire  abc_mshr_0_io_nestedwb_clients_1_isToN; // @[Slice.scala 94:16]
  wire  abc_mshr_0_io_tasks_sink_a_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_0_io_tasks_sink_a_valid; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_0_io_tasks_sink_a_bits_sourceId; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_0_io_tasks_sink_a_bits_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_0_io_tasks_sink_a_bits_tag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_0_io_tasks_sink_a_bits_size; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_0_io_tasks_sink_a_bits_off; // @[Slice.scala 94:16]
  wire  abc_mshr_0_io_tasks_source_bready; // @[Slice.scala 94:16]
  wire  abc_mshr_0_io_tasks_source_bvalid; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_0_io_tasks_source_bset; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_0_io_tasks_source_btag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_0_io_tasks_source_bparam; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_0_io_tasks_source_bclients; // @[Slice.scala 94:16]
  wire  abc_mshr_0_io_tasks_source_bneedData; // @[Slice.scala 94:16]
  wire  abc_mshr_0_io_tasks_sink_c_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_0_io_tasks_sink_c_valid; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_0_io_tasks_sink_c_bits_sourceId; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_0_io_tasks_sink_c_bits_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_0_io_tasks_sink_c_bits_tag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_0_io_tasks_sink_c_bits_size; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_0_io_tasks_sink_c_bits_way; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_0_io_tasks_sink_c_bits_off; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_0_io_tasks_sink_c_bits_bufIdx; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_0_io_tasks_sink_c_bits_opcode; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_0_io_tasks_sink_c_bits_param; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_0_io_tasks_sink_c_bits_source; // @[Slice.scala 94:16]
  wire  abc_mshr_0_io_tasks_sink_c_bits_save; // @[Slice.scala 94:16]
  wire  abc_mshr_0_io_tasks_sink_c_bits_drop; // @[Slice.scala 94:16]
  wire  abc_mshr_0_io_tasks_sink_c_bits_release; // @[Slice.scala 94:16]
  wire  abc_mshr_0_io_tasks_sink_c_bits_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_0_io_tasks_source_d_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_0_io_tasks_source_d_valid; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_0_io_tasks_source_d_bits_sourceId; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_0_io_tasks_source_d_bits_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_0_io_tasks_source_d_bits_tag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_0_io_tasks_source_d_bits_channel; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_0_io_tasks_source_d_bits_opcode; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_0_io_tasks_source_d_bits_param; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_0_io_tasks_source_d_bits_size; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_0_io_tasks_source_d_bits_way; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_0_io_tasks_source_d_bits_off; // @[Slice.scala 94:16]
  wire  abc_mshr_0_io_tasks_source_d_bits_useBypass; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_0_io_tasks_source_d_bits_bufIdx; // @[Slice.scala 94:16]
  wire  abc_mshr_0_io_tasks_source_d_bits_denied; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_0_io_tasks_source_d_bits_sinkId; // @[Slice.scala 94:16]
  wire  abc_mshr_0_io_tasks_source_d_bits_bypassPut; // @[Slice.scala 94:16]
  wire  abc_mshr_0_io_tasks_source_d_bits_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_0_io_tasks_source_a_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_0_io_tasks_source_a_valid; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_0_io_tasks_source_a_bits_tag; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_0_io_tasks_source_a_bits_set; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_0_io_tasks_source_a_bits_off; // @[Slice.scala 94:16]
  wire [31:0] abc_mshr_0_io_tasks_source_a_bits_mask; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_0_io_tasks_source_a_bits_opcode; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_0_io_tasks_source_a_bits_param; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_0_io_tasks_source_a_bits_source; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_0_io_tasks_source_a_bits_bufIdx; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_0_io_tasks_source_a_bits_size; // @[Slice.scala 94:16]
  wire  abc_mshr_0_io_tasks_source_a_bits_needData; // @[Slice.scala 94:16]
  wire  abc_mshr_0_io_tasks_source_a_bits_putData; // @[Slice.scala 94:16]
  wire  abc_mshr_0_io_tasks_source_c_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_0_io_tasks_source_c_valid; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_0_io_tasks_source_c_bits_opcode; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_0_io_tasks_source_c_bits_tag; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_0_io_tasks_source_c_bits_set; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_0_io_tasks_source_c_bits_param; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_0_io_tasks_source_c_bits_source; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_0_io_tasks_source_c_bits_way; // @[Slice.scala 94:16]
  wire  abc_mshr_0_io_tasks_source_c_bits_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_0_io_tasks_source_e_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_0_io_tasks_source_e_valid; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_0_io_tasks_source_e_bits_sink; // @[Slice.scala 94:16]
  wire  abc_mshr_0_io_tasks_dir_write_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_0_io_tasks_dir_write_valid; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_0_io_tasks_dir_write_bits_set; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_0_io_tasks_dir_write_bits_way; // @[Slice.scala 94:16]
  wire  abc_mshr_0_io_tasks_dir_write_bits_data_dirty; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_0_io_tasks_dir_write_bits_data_state; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_0_io_tasks_dir_write_bits_data_clientStates_0; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_0_io_tasks_dir_write_bits_data_clientStates_1; // @[Slice.scala 94:16]
  wire  abc_mshr_0_io_tasks_tag_write_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_0_io_tasks_tag_write_valid; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_0_io_tasks_tag_write_bits_set; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_0_io_tasks_tag_write_bits_way; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_0_io_tasks_tag_write_bits_tag; // @[Slice.scala 94:16]
  wire  abc_mshr_0_io_tasks_client_dir_write_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_0_io_tasks_client_dir_write_valid; // @[Slice.scala 94:16]
  wire [6:0] abc_mshr_0_io_tasks_client_dir_write_bits_set; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_0_io_tasks_client_dir_write_bits_way; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_0_io_tasks_client_dir_write_bits_data_0_state; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_0_io_tasks_client_dir_write_bits_data_1_state; // @[Slice.scala 94:16]
  wire  abc_mshr_0_io_tasks_client_tag_write_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_0_io_tasks_client_tag_write_valid; // @[Slice.scala 94:16]
  wire [6:0] abc_mshr_0_io_tasks_client_tag_write_bits_set; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_0_io_tasks_client_tag_write_bits_way; // @[Slice.scala 94:16]
  wire [22:0] abc_mshr_0_io_tasks_client_tag_write_bits_tag; // @[Slice.scala 94:16]
  wire  abc_mshr_0_io_dirResult_valid; // @[Slice.scala 94:16]
  wire  abc_mshr_0_io_dirResult_bits_self_dirty; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_0_io_dirResult_bits_self_state; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_0_io_dirResult_bits_self_clientStates_0; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_0_io_dirResult_bits_self_clientStates_1; // @[Slice.scala 94:16]
  wire  abc_mshr_0_io_dirResult_bits_self_hit; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_0_io_dirResult_bits_self_way; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_0_io_dirResult_bits_self_tag; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_0_io_dirResult_bits_clients_states_0_state; // @[Slice.scala 94:16]
  wire  abc_mshr_0_io_dirResult_bits_clients_states_0_hit; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_0_io_dirResult_bits_clients_states_1_state; // @[Slice.scala 94:16]
  wire  abc_mshr_0_io_dirResult_bits_clients_states_1_hit; // @[Slice.scala 94:16]
  wire [22:0] abc_mshr_0_io_dirResult_bits_clients_tag; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_0_io_dirResult_bits_clients_way; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_0_io_c_status_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_0_io_c_status_tag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_0_io_c_status_way; // @[Slice.scala 94:16]
  wire  abc_mshr_0_io_c_status_nestedReleaseData; // @[Slice.scala 94:16]
  wire  abc_mshr_0_io_c_status_releaseThrough; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_0_io_bstatus_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_0_io_bstatus_tag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_0_io_bstatus_way; // @[Slice.scala 94:16]
  wire  abc_mshr_0_io_bstatus_nestedProbeAckData; // @[Slice.scala 94:16]
  wire  abc_mshr_0_io_bstatus_probeHelperFinish; // @[Slice.scala 94:16]
  wire  abc_mshr_0_io_bstatus_probeAckDataThrough; // @[Slice.scala 94:16]
  wire  abc_mshr_0_io_releaseThrough; // @[Slice.scala 94:16]
  wire  abc_mshr_0_io_probeAckDataThrough; // @[Slice.scala 94:16]
  wire  abc_mshr_0_io_is_nestedReleaseData; // @[Slice.scala 94:16]
  wire  abc_mshr_0_io_is_nestedProbeAckData; // @[Slice.scala 94:16]
  wire  abc_mshr_0_io_probeHelperFinish; // @[Slice.scala 94:16]
  wire  abc_mshr_1_clock; // @[Slice.scala 94:16]
  wire  abc_mshr_1_reset; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_1_io_id; // @[Slice.scala 94:16]
  wire  abc_mshr_1_io_enable; // @[Slice.scala 94:16]
  wire  abc_mshr_1_io_alloc_valid; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_1_io_alloc_bits_channel; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_1_io_alloc_bits_opcode; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_1_io_alloc_bits_param; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_1_io_alloc_bits_size; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_1_io_alloc_bits_source; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_1_io_alloc_bits_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_1_io_alloc_bits_tag; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_1_io_alloc_bits_off; // @[Slice.scala 94:16]
  wire [31:0] abc_mshr_1_io_alloc_bits_mask; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_1_io_alloc_bits_bufIdx; // @[Slice.scala 94:16]
  wire  abc_mshr_1_io_alloc_bits_preferCache; // @[Slice.scala 94:16]
  wire  abc_mshr_1_io_alloc_bits_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_1_io_alloc_bits_fromProbeHelper; // @[Slice.scala 94:16]
  wire  abc_mshr_1_io_alloc_bits_fromCmoHelper; // @[Slice.scala 94:16]
  wire  abc_mshr_1_io_alloc_bits_needProbeAckData; // @[Slice.scala 94:16]
  wire  abc_mshr_1_io_status_valid; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_1_io_status_bits_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_1_io_status_bits_tag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_1_io_status_bits_way; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_1_io_status_bits_way_reg; // @[Slice.scala 94:16]
  wire  abc_mshr_1_io_status_bits_nestB; // @[Slice.scala 94:16]
  wire  abc_mshr_1_io_status_bits_nestC; // @[Slice.scala 94:16]
  wire  abc_mshr_1_io_status_bits_will_grant_data; // @[Slice.scala 94:16]
  wire  abc_mshr_1_io_status_bits_will_save_data; // @[Slice.scala 94:16]
  wire  abc_mshr_1_io_status_bits_will_free; // @[Slice.scala 94:16]
  wire  abc_mshr_1_io_resps_sink_c_valid; // @[Slice.scala 94:16]
  wire  abc_mshr_1_io_resps_sink_c_bits_hasData; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_1_io_resps_sink_c_bits_param; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_1_io_resps_sink_c_bits_source; // @[Slice.scala 94:16]
  wire  abc_mshr_1_io_resps_sink_c_bits_last; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_1_io_resps_sink_c_bits_bufIdx; // @[Slice.scala 94:16]
  wire  abc_mshr_1_io_resps_sink_d_valid; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_1_io_resps_sink_d_bits_opcode; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_1_io_resps_sink_d_bits_param; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_1_io_resps_sink_d_bits_sink; // @[Slice.scala 94:16]
  wire  abc_mshr_1_io_resps_sink_d_bits_last; // @[Slice.scala 94:16]
  wire  abc_mshr_1_io_resps_sink_d_bits_denied; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_1_io_resps_sink_d_bits_bufIdx; // @[Slice.scala 94:16]
  wire  abc_mshr_1_io_resps_sink_e_valid; // @[Slice.scala 94:16]
  wire  abc_mshr_1_io_resps_source_d_valid; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_1_io_nestedwb_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_1_io_nestedwb_tag; // @[Slice.scala 94:16]
  wire  abc_mshr_1_io_nestedwb_btoN; // @[Slice.scala 94:16]
  wire  abc_mshr_1_io_nestedwb_btoB; // @[Slice.scala 94:16]
  wire  abc_mshr_1_io_nestedwb_bclr_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_1_io_nestedwb_bset_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_1_io_nestedwb_c_set_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_1_io_nestedwb_c_set_hit; // @[Slice.scala 94:16]
  wire  abc_mshr_1_io_nestedwb_clients_0_isToN; // @[Slice.scala 94:16]
  wire  abc_mshr_1_io_nestedwb_clients_1_isToN; // @[Slice.scala 94:16]
  wire  abc_mshr_1_io_tasks_sink_a_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_1_io_tasks_sink_a_valid; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_1_io_tasks_sink_a_bits_sourceId; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_1_io_tasks_sink_a_bits_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_1_io_tasks_sink_a_bits_tag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_1_io_tasks_sink_a_bits_size; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_1_io_tasks_sink_a_bits_off; // @[Slice.scala 94:16]
  wire  abc_mshr_1_io_tasks_source_bready; // @[Slice.scala 94:16]
  wire  abc_mshr_1_io_tasks_source_bvalid; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_1_io_tasks_source_bset; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_1_io_tasks_source_btag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_1_io_tasks_source_bparam; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_1_io_tasks_source_bclients; // @[Slice.scala 94:16]
  wire  abc_mshr_1_io_tasks_source_bneedData; // @[Slice.scala 94:16]
  wire  abc_mshr_1_io_tasks_sink_c_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_1_io_tasks_sink_c_valid; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_1_io_tasks_sink_c_bits_sourceId; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_1_io_tasks_sink_c_bits_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_1_io_tasks_sink_c_bits_tag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_1_io_tasks_sink_c_bits_size; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_1_io_tasks_sink_c_bits_way; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_1_io_tasks_sink_c_bits_off; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_1_io_tasks_sink_c_bits_bufIdx; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_1_io_tasks_sink_c_bits_opcode; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_1_io_tasks_sink_c_bits_param; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_1_io_tasks_sink_c_bits_source; // @[Slice.scala 94:16]
  wire  abc_mshr_1_io_tasks_sink_c_bits_save; // @[Slice.scala 94:16]
  wire  abc_mshr_1_io_tasks_sink_c_bits_drop; // @[Slice.scala 94:16]
  wire  abc_mshr_1_io_tasks_sink_c_bits_release; // @[Slice.scala 94:16]
  wire  abc_mshr_1_io_tasks_sink_c_bits_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_1_io_tasks_source_d_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_1_io_tasks_source_d_valid; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_1_io_tasks_source_d_bits_sourceId; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_1_io_tasks_source_d_bits_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_1_io_tasks_source_d_bits_tag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_1_io_tasks_source_d_bits_channel; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_1_io_tasks_source_d_bits_opcode; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_1_io_tasks_source_d_bits_param; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_1_io_tasks_source_d_bits_size; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_1_io_tasks_source_d_bits_way; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_1_io_tasks_source_d_bits_off; // @[Slice.scala 94:16]
  wire  abc_mshr_1_io_tasks_source_d_bits_useBypass; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_1_io_tasks_source_d_bits_bufIdx; // @[Slice.scala 94:16]
  wire  abc_mshr_1_io_tasks_source_d_bits_denied; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_1_io_tasks_source_d_bits_sinkId; // @[Slice.scala 94:16]
  wire  abc_mshr_1_io_tasks_source_d_bits_bypassPut; // @[Slice.scala 94:16]
  wire  abc_mshr_1_io_tasks_source_d_bits_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_1_io_tasks_source_a_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_1_io_tasks_source_a_valid; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_1_io_tasks_source_a_bits_tag; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_1_io_tasks_source_a_bits_set; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_1_io_tasks_source_a_bits_off; // @[Slice.scala 94:16]
  wire [31:0] abc_mshr_1_io_tasks_source_a_bits_mask; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_1_io_tasks_source_a_bits_opcode; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_1_io_tasks_source_a_bits_param; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_1_io_tasks_source_a_bits_source; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_1_io_tasks_source_a_bits_bufIdx; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_1_io_tasks_source_a_bits_size; // @[Slice.scala 94:16]
  wire  abc_mshr_1_io_tasks_source_a_bits_needData; // @[Slice.scala 94:16]
  wire  abc_mshr_1_io_tasks_source_a_bits_putData; // @[Slice.scala 94:16]
  wire  abc_mshr_1_io_tasks_source_c_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_1_io_tasks_source_c_valid; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_1_io_tasks_source_c_bits_opcode; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_1_io_tasks_source_c_bits_tag; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_1_io_tasks_source_c_bits_set; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_1_io_tasks_source_c_bits_param; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_1_io_tasks_source_c_bits_source; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_1_io_tasks_source_c_bits_way; // @[Slice.scala 94:16]
  wire  abc_mshr_1_io_tasks_source_c_bits_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_1_io_tasks_source_e_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_1_io_tasks_source_e_valid; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_1_io_tasks_source_e_bits_sink; // @[Slice.scala 94:16]
  wire  abc_mshr_1_io_tasks_dir_write_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_1_io_tasks_dir_write_valid; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_1_io_tasks_dir_write_bits_set; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_1_io_tasks_dir_write_bits_way; // @[Slice.scala 94:16]
  wire  abc_mshr_1_io_tasks_dir_write_bits_data_dirty; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_1_io_tasks_dir_write_bits_data_state; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_1_io_tasks_dir_write_bits_data_clientStates_0; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_1_io_tasks_dir_write_bits_data_clientStates_1; // @[Slice.scala 94:16]
  wire  abc_mshr_1_io_tasks_tag_write_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_1_io_tasks_tag_write_valid; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_1_io_tasks_tag_write_bits_set; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_1_io_tasks_tag_write_bits_way; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_1_io_tasks_tag_write_bits_tag; // @[Slice.scala 94:16]
  wire  abc_mshr_1_io_tasks_client_dir_write_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_1_io_tasks_client_dir_write_valid; // @[Slice.scala 94:16]
  wire [6:0] abc_mshr_1_io_tasks_client_dir_write_bits_set; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_1_io_tasks_client_dir_write_bits_way; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_1_io_tasks_client_dir_write_bits_data_0_state; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_1_io_tasks_client_dir_write_bits_data_1_state; // @[Slice.scala 94:16]
  wire  abc_mshr_1_io_tasks_client_tag_write_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_1_io_tasks_client_tag_write_valid; // @[Slice.scala 94:16]
  wire [6:0] abc_mshr_1_io_tasks_client_tag_write_bits_set; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_1_io_tasks_client_tag_write_bits_way; // @[Slice.scala 94:16]
  wire [22:0] abc_mshr_1_io_tasks_client_tag_write_bits_tag; // @[Slice.scala 94:16]
  wire  abc_mshr_1_io_dirResult_valid; // @[Slice.scala 94:16]
  wire  abc_mshr_1_io_dirResult_bits_self_dirty; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_1_io_dirResult_bits_self_state; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_1_io_dirResult_bits_self_clientStates_0; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_1_io_dirResult_bits_self_clientStates_1; // @[Slice.scala 94:16]
  wire  abc_mshr_1_io_dirResult_bits_self_hit; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_1_io_dirResult_bits_self_way; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_1_io_dirResult_bits_self_tag; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_1_io_dirResult_bits_clients_states_0_state; // @[Slice.scala 94:16]
  wire  abc_mshr_1_io_dirResult_bits_clients_states_0_hit; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_1_io_dirResult_bits_clients_states_1_state; // @[Slice.scala 94:16]
  wire  abc_mshr_1_io_dirResult_bits_clients_states_1_hit; // @[Slice.scala 94:16]
  wire [22:0] abc_mshr_1_io_dirResult_bits_clients_tag; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_1_io_dirResult_bits_clients_way; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_1_io_c_status_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_1_io_c_status_tag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_1_io_c_status_way; // @[Slice.scala 94:16]
  wire  abc_mshr_1_io_c_status_nestedReleaseData; // @[Slice.scala 94:16]
  wire  abc_mshr_1_io_c_status_releaseThrough; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_1_io_bstatus_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_1_io_bstatus_tag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_1_io_bstatus_way; // @[Slice.scala 94:16]
  wire  abc_mshr_1_io_bstatus_nestedProbeAckData; // @[Slice.scala 94:16]
  wire  abc_mshr_1_io_bstatus_probeHelperFinish; // @[Slice.scala 94:16]
  wire  abc_mshr_1_io_bstatus_probeAckDataThrough; // @[Slice.scala 94:16]
  wire  abc_mshr_1_io_releaseThrough; // @[Slice.scala 94:16]
  wire  abc_mshr_1_io_probeAckDataThrough; // @[Slice.scala 94:16]
  wire  abc_mshr_1_io_is_nestedReleaseData; // @[Slice.scala 94:16]
  wire  abc_mshr_1_io_is_nestedProbeAckData; // @[Slice.scala 94:16]
  wire  abc_mshr_1_io_probeHelperFinish; // @[Slice.scala 94:16]
  wire  abc_mshr_2_clock; // @[Slice.scala 94:16]
  wire  abc_mshr_2_reset; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_2_io_id; // @[Slice.scala 94:16]
  wire  abc_mshr_2_io_enable; // @[Slice.scala 94:16]
  wire  abc_mshr_2_io_alloc_valid; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_2_io_alloc_bits_channel; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_2_io_alloc_bits_opcode; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_2_io_alloc_bits_param; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_2_io_alloc_bits_size; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_2_io_alloc_bits_source; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_2_io_alloc_bits_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_2_io_alloc_bits_tag; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_2_io_alloc_bits_off; // @[Slice.scala 94:16]
  wire [31:0] abc_mshr_2_io_alloc_bits_mask; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_2_io_alloc_bits_bufIdx; // @[Slice.scala 94:16]
  wire  abc_mshr_2_io_alloc_bits_preferCache; // @[Slice.scala 94:16]
  wire  abc_mshr_2_io_alloc_bits_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_2_io_alloc_bits_fromProbeHelper; // @[Slice.scala 94:16]
  wire  abc_mshr_2_io_alloc_bits_fromCmoHelper; // @[Slice.scala 94:16]
  wire  abc_mshr_2_io_alloc_bits_needProbeAckData; // @[Slice.scala 94:16]
  wire  abc_mshr_2_io_status_valid; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_2_io_status_bits_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_2_io_status_bits_tag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_2_io_status_bits_way; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_2_io_status_bits_way_reg; // @[Slice.scala 94:16]
  wire  abc_mshr_2_io_status_bits_nestB; // @[Slice.scala 94:16]
  wire  abc_mshr_2_io_status_bits_nestC; // @[Slice.scala 94:16]
  wire  abc_mshr_2_io_status_bits_will_grant_data; // @[Slice.scala 94:16]
  wire  abc_mshr_2_io_status_bits_will_save_data; // @[Slice.scala 94:16]
  wire  abc_mshr_2_io_status_bits_will_free; // @[Slice.scala 94:16]
  wire  abc_mshr_2_io_resps_sink_c_valid; // @[Slice.scala 94:16]
  wire  abc_mshr_2_io_resps_sink_c_bits_hasData; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_2_io_resps_sink_c_bits_param; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_2_io_resps_sink_c_bits_source; // @[Slice.scala 94:16]
  wire  abc_mshr_2_io_resps_sink_c_bits_last; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_2_io_resps_sink_c_bits_bufIdx; // @[Slice.scala 94:16]
  wire  abc_mshr_2_io_resps_sink_d_valid; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_2_io_resps_sink_d_bits_opcode; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_2_io_resps_sink_d_bits_param; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_2_io_resps_sink_d_bits_sink; // @[Slice.scala 94:16]
  wire  abc_mshr_2_io_resps_sink_d_bits_last; // @[Slice.scala 94:16]
  wire  abc_mshr_2_io_resps_sink_d_bits_denied; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_2_io_resps_sink_d_bits_bufIdx; // @[Slice.scala 94:16]
  wire  abc_mshr_2_io_resps_sink_e_valid; // @[Slice.scala 94:16]
  wire  abc_mshr_2_io_resps_source_d_valid; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_2_io_nestedwb_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_2_io_nestedwb_tag; // @[Slice.scala 94:16]
  wire  abc_mshr_2_io_nestedwb_btoN; // @[Slice.scala 94:16]
  wire  abc_mshr_2_io_nestedwb_btoB; // @[Slice.scala 94:16]
  wire  abc_mshr_2_io_nestedwb_bclr_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_2_io_nestedwb_bset_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_2_io_nestedwb_c_set_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_2_io_nestedwb_c_set_hit; // @[Slice.scala 94:16]
  wire  abc_mshr_2_io_nestedwb_clients_0_isToN; // @[Slice.scala 94:16]
  wire  abc_mshr_2_io_nestedwb_clients_1_isToN; // @[Slice.scala 94:16]
  wire  abc_mshr_2_io_tasks_sink_a_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_2_io_tasks_sink_a_valid; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_2_io_tasks_sink_a_bits_sourceId; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_2_io_tasks_sink_a_bits_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_2_io_tasks_sink_a_bits_tag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_2_io_tasks_sink_a_bits_size; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_2_io_tasks_sink_a_bits_off; // @[Slice.scala 94:16]
  wire  abc_mshr_2_io_tasks_source_bready; // @[Slice.scala 94:16]
  wire  abc_mshr_2_io_tasks_source_bvalid; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_2_io_tasks_source_bset; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_2_io_tasks_source_btag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_2_io_tasks_source_bparam; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_2_io_tasks_source_bclients; // @[Slice.scala 94:16]
  wire  abc_mshr_2_io_tasks_source_bneedData; // @[Slice.scala 94:16]
  wire  abc_mshr_2_io_tasks_sink_c_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_2_io_tasks_sink_c_valid; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_2_io_tasks_sink_c_bits_sourceId; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_2_io_tasks_sink_c_bits_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_2_io_tasks_sink_c_bits_tag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_2_io_tasks_sink_c_bits_size; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_2_io_tasks_sink_c_bits_way; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_2_io_tasks_sink_c_bits_off; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_2_io_tasks_sink_c_bits_bufIdx; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_2_io_tasks_sink_c_bits_opcode; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_2_io_tasks_sink_c_bits_param; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_2_io_tasks_sink_c_bits_source; // @[Slice.scala 94:16]
  wire  abc_mshr_2_io_tasks_sink_c_bits_save; // @[Slice.scala 94:16]
  wire  abc_mshr_2_io_tasks_sink_c_bits_drop; // @[Slice.scala 94:16]
  wire  abc_mshr_2_io_tasks_sink_c_bits_release; // @[Slice.scala 94:16]
  wire  abc_mshr_2_io_tasks_sink_c_bits_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_2_io_tasks_source_d_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_2_io_tasks_source_d_valid; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_2_io_tasks_source_d_bits_sourceId; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_2_io_tasks_source_d_bits_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_2_io_tasks_source_d_bits_tag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_2_io_tasks_source_d_bits_channel; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_2_io_tasks_source_d_bits_opcode; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_2_io_tasks_source_d_bits_param; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_2_io_tasks_source_d_bits_size; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_2_io_tasks_source_d_bits_way; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_2_io_tasks_source_d_bits_off; // @[Slice.scala 94:16]
  wire  abc_mshr_2_io_tasks_source_d_bits_useBypass; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_2_io_tasks_source_d_bits_bufIdx; // @[Slice.scala 94:16]
  wire  abc_mshr_2_io_tasks_source_d_bits_denied; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_2_io_tasks_source_d_bits_sinkId; // @[Slice.scala 94:16]
  wire  abc_mshr_2_io_tasks_source_d_bits_bypassPut; // @[Slice.scala 94:16]
  wire  abc_mshr_2_io_tasks_source_d_bits_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_2_io_tasks_source_a_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_2_io_tasks_source_a_valid; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_2_io_tasks_source_a_bits_tag; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_2_io_tasks_source_a_bits_set; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_2_io_tasks_source_a_bits_off; // @[Slice.scala 94:16]
  wire [31:0] abc_mshr_2_io_tasks_source_a_bits_mask; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_2_io_tasks_source_a_bits_opcode; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_2_io_tasks_source_a_bits_param; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_2_io_tasks_source_a_bits_source; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_2_io_tasks_source_a_bits_bufIdx; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_2_io_tasks_source_a_bits_size; // @[Slice.scala 94:16]
  wire  abc_mshr_2_io_tasks_source_a_bits_needData; // @[Slice.scala 94:16]
  wire  abc_mshr_2_io_tasks_source_a_bits_putData; // @[Slice.scala 94:16]
  wire  abc_mshr_2_io_tasks_source_c_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_2_io_tasks_source_c_valid; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_2_io_tasks_source_c_bits_opcode; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_2_io_tasks_source_c_bits_tag; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_2_io_tasks_source_c_bits_set; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_2_io_tasks_source_c_bits_param; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_2_io_tasks_source_c_bits_source; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_2_io_tasks_source_c_bits_way; // @[Slice.scala 94:16]
  wire  abc_mshr_2_io_tasks_source_c_bits_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_2_io_tasks_source_e_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_2_io_tasks_source_e_valid; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_2_io_tasks_source_e_bits_sink; // @[Slice.scala 94:16]
  wire  abc_mshr_2_io_tasks_dir_write_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_2_io_tasks_dir_write_valid; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_2_io_tasks_dir_write_bits_set; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_2_io_tasks_dir_write_bits_way; // @[Slice.scala 94:16]
  wire  abc_mshr_2_io_tasks_dir_write_bits_data_dirty; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_2_io_tasks_dir_write_bits_data_state; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_2_io_tasks_dir_write_bits_data_clientStates_0; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_2_io_tasks_dir_write_bits_data_clientStates_1; // @[Slice.scala 94:16]
  wire  abc_mshr_2_io_tasks_tag_write_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_2_io_tasks_tag_write_valid; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_2_io_tasks_tag_write_bits_set; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_2_io_tasks_tag_write_bits_way; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_2_io_tasks_tag_write_bits_tag; // @[Slice.scala 94:16]
  wire  abc_mshr_2_io_tasks_client_dir_write_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_2_io_tasks_client_dir_write_valid; // @[Slice.scala 94:16]
  wire [6:0] abc_mshr_2_io_tasks_client_dir_write_bits_set; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_2_io_tasks_client_dir_write_bits_way; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_2_io_tasks_client_dir_write_bits_data_0_state; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_2_io_tasks_client_dir_write_bits_data_1_state; // @[Slice.scala 94:16]
  wire  abc_mshr_2_io_tasks_client_tag_write_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_2_io_tasks_client_tag_write_valid; // @[Slice.scala 94:16]
  wire [6:0] abc_mshr_2_io_tasks_client_tag_write_bits_set; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_2_io_tasks_client_tag_write_bits_way; // @[Slice.scala 94:16]
  wire [22:0] abc_mshr_2_io_tasks_client_tag_write_bits_tag; // @[Slice.scala 94:16]
  wire  abc_mshr_2_io_dirResult_valid; // @[Slice.scala 94:16]
  wire  abc_mshr_2_io_dirResult_bits_self_dirty; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_2_io_dirResult_bits_self_state; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_2_io_dirResult_bits_self_clientStates_0; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_2_io_dirResult_bits_self_clientStates_1; // @[Slice.scala 94:16]
  wire  abc_mshr_2_io_dirResult_bits_self_hit; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_2_io_dirResult_bits_self_way; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_2_io_dirResult_bits_self_tag; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_2_io_dirResult_bits_clients_states_0_state; // @[Slice.scala 94:16]
  wire  abc_mshr_2_io_dirResult_bits_clients_states_0_hit; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_2_io_dirResult_bits_clients_states_1_state; // @[Slice.scala 94:16]
  wire  abc_mshr_2_io_dirResult_bits_clients_states_1_hit; // @[Slice.scala 94:16]
  wire [22:0] abc_mshr_2_io_dirResult_bits_clients_tag; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_2_io_dirResult_bits_clients_way; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_2_io_c_status_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_2_io_c_status_tag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_2_io_c_status_way; // @[Slice.scala 94:16]
  wire  abc_mshr_2_io_c_status_nestedReleaseData; // @[Slice.scala 94:16]
  wire  abc_mshr_2_io_c_status_releaseThrough; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_2_io_bstatus_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_2_io_bstatus_tag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_2_io_bstatus_way; // @[Slice.scala 94:16]
  wire  abc_mshr_2_io_bstatus_nestedProbeAckData; // @[Slice.scala 94:16]
  wire  abc_mshr_2_io_bstatus_probeHelperFinish; // @[Slice.scala 94:16]
  wire  abc_mshr_2_io_bstatus_probeAckDataThrough; // @[Slice.scala 94:16]
  wire  abc_mshr_2_io_releaseThrough; // @[Slice.scala 94:16]
  wire  abc_mshr_2_io_probeAckDataThrough; // @[Slice.scala 94:16]
  wire  abc_mshr_2_io_is_nestedReleaseData; // @[Slice.scala 94:16]
  wire  abc_mshr_2_io_is_nestedProbeAckData; // @[Slice.scala 94:16]
  wire  abc_mshr_2_io_probeHelperFinish; // @[Slice.scala 94:16]
  wire  abc_mshr_3_clock; // @[Slice.scala 94:16]
  wire  abc_mshr_3_reset; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_3_io_id; // @[Slice.scala 94:16]
  wire  abc_mshr_3_io_enable; // @[Slice.scala 94:16]
  wire  abc_mshr_3_io_alloc_valid; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_3_io_alloc_bits_channel; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_3_io_alloc_bits_opcode; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_3_io_alloc_bits_param; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_3_io_alloc_bits_size; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_3_io_alloc_bits_source; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_3_io_alloc_bits_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_3_io_alloc_bits_tag; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_3_io_alloc_bits_off; // @[Slice.scala 94:16]
  wire [31:0] abc_mshr_3_io_alloc_bits_mask; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_3_io_alloc_bits_bufIdx; // @[Slice.scala 94:16]
  wire  abc_mshr_3_io_alloc_bits_preferCache; // @[Slice.scala 94:16]
  wire  abc_mshr_3_io_alloc_bits_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_3_io_alloc_bits_fromProbeHelper; // @[Slice.scala 94:16]
  wire  abc_mshr_3_io_alloc_bits_fromCmoHelper; // @[Slice.scala 94:16]
  wire  abc_mshr_3_io_alloc_bits_needProbeAckData; // @[Slice.scala 94:16]
  wire  abc_mshr_3_io_status_valid; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_3_io_status_bits_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_3_io_status_bits_tag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_3_io_status_bits_way; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_3_io_status_bits_way_reg; // @[Slice.scala 94:16]
  wire  abc_mshr_3_io_status_bits_nestB; // @[Slice.scala 94:16]
  wire  abc_mshr_3_io_status_bits_nestC; // @[Slice.scala 94:16]
  wire  abc_mshr_3_io_status_bits_will_grant_data; // @[Slice.scala 94:16]
  wire  abc_mshr_3_io_status_bits_will_save_data; // @[Slice.scala 94:16]
  wire  abc_mshr_3_io_status_bits_will_free; // @[Slice.scala 94:16]
  wire  abc_mshr_3_io_resps_sink_c_valid; // @[Slice.scala 94:16]
  wire  abc_mshr_3_io_resps_sink_c_bits_hasData; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_3_io_resps_sink_c_bits_param; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_3_io_resps_sink_c_bits_source; // @[Slice.scala 94:16]
  wire  abc_mshr_3_io_resps_sink_c_bits_last; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_3_io_resps_sink_c_bits_bufIdx; // @[Slice.scala 94:16]
  wire  abc_mshr_3_io_resps_sink_d_valid; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_3_io_resps_sink_d_bits_opcode; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_3_io_resps_sink_d_bits_param; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_3_io_resps_sink_d_bits_sink; // @[Slice.scala 94:16]
  wire  abc_mshr_3_io_resps_sink_d_bits_last; // @[Slice.scala 94:16]
  wire  abc_mshr_3_io_resps_sink_d_bits_denied; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_3_io_resps_sink_d_bits_bufIdx; // @[Slice.scala 94:16]
  wire  abc_mshr_3_io_resps_sink_e_valid; // @[Slice.scala 94:16]
  wire  abc_mshr_3_io_resps_source_d_valid; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_3_io_nestedwb_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_3_io_nestedwb_tag; // @[Slice.scala 94:16]
  wire  abc_mshr_3_io_nestedwb_btoN; // @[Slice.scala 94:16]
  wire  abc_mshr_3_io_nestedwb_btoB; // @[Slice.scala 94:16]
  wire  abc_mshr_3_io_nestedwb_bclr_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_3_io_nestedwb_bset_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_3_io_nestedwb_c_set_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_3_io_nestedwb_c_set_hit; // @[Slice.scala 94:16]
  wire  abc_mshr_3_io_nestedwb_clients_0_isToN; // @[Slice.scala 94:16]
  wire  abc_mshr_3_io_nestedwb_clients_1_isToN; // @[Slice.scala 94:16]
  wire  abc_mshr_3_io_tasks_sink_a_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_3_io_tasks_sink_a_valid; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_3_io_tasks_sink_a_bits_sourceId; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_3_io_tasks_sink_a_bits_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_3_io_tasks_sink_a_bits_tag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_3_io_tasks_sink_a_bits_size; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_3_io_tasks_sink_a_bits_off; // @[Slice.scala 94:16]
  wire  abc_mshr_3_io_tasks_source_bready; // @[Slice.scala 94:16]
  wire  abc_mshr_3_io_tasks_source_bvalid; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_3_io_tasks_source_bset; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_3_io_tasks_source_btag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_3_io_tasks_source_bparam; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_3_io_tasks_source_bclients; // @[Slice.scala 94:16]
  wire  abc_mshr_3_io_tasks_source_bneedData; // @[Slice.scala 94:16]
  wire  abc_mshr_3_io_tasks_sink_c_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_3_io_tasks_sink_c_valid; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_3_io_tasks_sink_c_bits_sourceId; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_3_io_tasks_sink_c_bits_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_3_io_tasks_sink_c_bits_tag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_3_io_tasks_sink_c_bits_size; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_3_io_tasks_sink_c_bits_way; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_3_io_tasks_sink_c_bits_off; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_3_io_tasks_sink_c_bits_bufIdx; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_3_io_tasks_sink_c_bits_opcode; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_3_io_tasks_sink_c_bits_param; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_3_io_tasks_sink_c_bits_source; // @[Slice.scala 94:16]
  wire  abc_mshr_3_io_tasks_sink_c_bits_save; // @[Slice.scala 94:16]
  wire  abc_mshr_3_io_tasks_sink_c_bits_drop; // @[Slice.scala 94:16]
  wire  abc_mshr_3_io_tasks_sink_c_bits_release; // @[Slice.scala 94:16]
  wire  abc_mshr_3_io_tasks_sink_c_bits_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_3_io_tasks_source_d_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_3_io_tasks_source_d_valid; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_3_io_tasks_source_d_bits_sourceId; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_3_io_tasks_source_d_bits_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_3_io_tasks_source_d_bits_tag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_3_io_tasks_source_d_bits_channel; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_3_io_tasks_source_d_bits_opcode; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_3_io_tasks_source_d_bits_param; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_3_io_tasks_source_d_bits_size; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_3_io_tasks_source_d_bits_way; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_3_io_tasks_source_d_bits_off; // @[Slice.scala 94:16]
  wire  abc_mshr_3_io_tasks_source_d_bits_useBypass; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_3_io_tasks_source_d_bits_bufIdx; // @[Slice.scala 94:16]
  wire  abc_mshr_3_io_tasks_source_d_bits_denied; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_3_io_tasks_source_d_bits_sinkId; // @[Slice.scala 94:16]
  wire  abc_mshr_3_io_tasks_source_d_bits_bypassPut; // @[Slice.scala 94:16]
  wire  abc_mshr_3_io_tasks_source_d_bits_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_3_io_tasks_source_a_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_3_io_tasks_source_a_valid; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_3_io_tasks_source_a_bits_tag; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_3_io_tasks_source_a_bits_set; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_3_io_tasks_source_a_bits_off; // @[Slice.scala 94:16]
  wire [31:0] abc_mshr_3_io_tasks_source_a_bits_mask; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_3_io_tasks_source_a_bits_opcode; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_3_io_tasks_source_a_bits_param; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_3_io_tasks_source_a_bits_source; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_3_io_tasks_source_a_bits_bufIdx; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_3_io_tasks_source_a_bits_size; // @[Slice.scala 94:16]
  wire  abc_mshr_3_io_tasks_source_a_bits_needData; // @[Slice.scala 94:16]
  wire  abc_mshr_3_io_tasks_source_a_bits_putData; // @[Slice.scala 94:16]
  wire  abc_mshr_3_io_tasks_source_c_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_3_io_tasks_source_c_valid; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_3_io_tasks_source_c_bits_opcode; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_3_io_tasks_source_c_bits_tag; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_3_io_tasks_source_c_bits_set; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_3_io_tasks_source_c_bits_param; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_3_io_tasks_source_c_bits_source; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_3_io_tasks_source_c_bits_way; // @[Slice.scala 94:16]
  wire  abc_mshr_3_io_tasks_source_c_bits_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_3_io_tasks_source_e_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_3_io_tasks_source_e_valid; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_3_io_tasks_source_e_bits_sink; // @[Slice.scala 94:16]
  wire  abc_mshr_3_io_tasks_dir_write_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_3_io_tasks_dir_write_valid; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_3_io_tasks_dir_write_bits_set; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_3_io_tasks_dir_write_bits_way; // @[Slice.scala 94:16]
  wire  abc_mshr_3_io_tasks_dir_write_bits_data_dirty; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_3_io_tasks_dir_write_bits_data_state; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_3_io_tasks_dir_write_bits_data_clientStates_0; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_3_io_tasks_dir_write_bits_data_clientStates_1; // @[Slice.scala 94:16]
  wire  abc_mshr_3_io_tasks_tag_write_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_3_io_tasks_tag_write_valid; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_3_io_tasks_tag_write_bits_set; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_3_io_tasks_tag_write_bits_way; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_3_io_tasks_tag_write_bits_tag; // @[Slice.scala 94:16]
  wire  abc_mshr_3_io_tasks_client_dir_write_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_3_io_tasks_client_dir_write_valid; // @[Slice.scala 94:16]
  wire [6:0] abc_mshr_3_io_tasks_client_dir_write_bits_set; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_3_io_tasks_client_dir_write_bits_way; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_3_io_tasks_client_dir_write_bits_data_0_state; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_3_io_tasks_client_dir_write_bits_data_1_state; // @[Slice.scala 94:16]
  wire  abc_mshr_3_io_tasks_client_tag_write_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_3_io_tasks_client_tag_write_valid; // @[Slice.scala 94:16]
  wire [6:0] abc_mshr_3_io_tasks_client_tag_write_bits_set; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_3_io_tasks_client_tag_write_bits_way; // @[Slice.scala 94:16]
  wire [22:0] abc_mshr_3_io_tasks_client_tag_write_bits_tag; // @[Slice.scala 94:16]
  wire  abc_mshr_3_io_dirResult_valid; // @[Slice.scala 94:16]
  wire  abc_mshr_3_io_dirResult_bits_self_dirty; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_3_io_dirResult_bits_self_state; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_3_io_dirResult_bits_self_clientStates_0; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_3_io_dirResult_bits_self_clientStates_1; // @[Slice.scala 94:16]
  wire  abc_mshr_3_io_dirResult_bits_self_hit; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_3_io_dirResult_bits_self_way; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_3_io_dirResult_bits_self_tag; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_3_io_dirResult_bits_clients_states_0_state; // @[Slice.scala 94:16]
  wire  abc_mshr_3_io_dirResult_bits_clients_states_0_hit; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_3_io_dirResult_bits_clients_states_1_state; // @[Slice.scala 94:16]
  wire  abc_mshr_3_io_dirResult_bits_clients_states_1_hit; // @[Slice.scala 94:16]
  wire [22:0] abc_mshr_3_io_dirResult_bits_clients_tag; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_3_io_dirResult_bits_clients_way; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_3_io_c_status_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_3_io_c_status_tag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_3_io_c_status_way; // @[Slice.scala 94:16]
  wire  abc_mshr_3_io_c_status_nestedReleaseData; // @[Slice.scala 94:16]
  wire  abc_mshr_3_io_c_status_releaseThrough; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_3_io_bstatus_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_3_io_bstatus_tag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_3_io_bstatus_way; // @[Slice.scala 94:16]
  wire  abc_mshr_3_io_bstatus_nestedProbeAckData; // @[Slice.scala 94:16]
  wire  abc_mshr_3_io_bstatus_probeHelperFinish; // @[Slice.scala 94:16]
  wire  abc_mshr_3_io_bstatus_probeAckDataThrough; // @[Slice.scala 94:16]
  wire  abc_mshr_3_io_releaseThrough; // @[Slice.scala 94:16]
  wire  abc_mshr_3_io_probeAckDataThrough; // @[Slice.scala 94:16]
  wire  abc_mshr_3_io_is_nestedReleaseData; // @[Slice.scala 94:16]
  wire  abc_mshr_3_io_is_nestedProbeAckData; // @[Slice.scala 94:16]
  wire  abc_mshr_3_io_probeHelperFinish; // @[Slice.scala 94:16]
  wire  abc_mshr_4_clock; // @[Slice.scala 94:16]
  wire  abc_mshr_4_reset; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_4_io_id; // @[Slice.scala 94:16]
  wire  abc_mshr_4_io_enable; // @[Slice.scala 94:16]
  wire  abc_mshr_4_io_alloc_valid; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_4_io_alloc_bits_channel; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_4_io_alloc_bits_opcode; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_4_io_alloc_bits_param; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_4_io_alloc_bits_size; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_4_io_alloc_bits_source; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_4_io_alloc_bits_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_4_io_alloc_bits_tag; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_4_io_alloc_bits_off; // @[Slice.scala 94:16]
  wire [31:0] abc_mshr_4_io_alloc_bits_mask; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_4_io_alloc_bits_bufIdx; // @[Slice.scala 94:16]
  wire  abc_mshr_4_io_alloc_bits_preferCache; // @[Slice.scala 94:16]
  wire  abc_mshr_4_io_alloc_bits_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_4_io_alloc_bits_fromProbeHelper; // @[Slice.scala 94:16]
  wire  abc_mshr_4_io_alloc_bits_fromCmoHelper; // @[Slice.scala 94:16]
  wire  abc_mshr_4_io_alloc_bits_needProbeAckData; // @[Slice.scala 94:16]
  wire  abc_mshr_4_io_status_valid; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_4_io_status_bits_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_4_io_status_bits_tag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_4_io_status_bits_way; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_4_io_status_bits_way_reg; // @[Slice.scala 94:16]
  wire  abc_mshr_4_io_status_bits_nestB; // @[Slice.scala 94:16]
  wire  abc_mshr_4_io_status_bits_nestC; // @[Slice.scala 94:16]
  wire  abc_mshr_4_io_status_bits_will_grant_data; // @[Slice.scala 94:16]
  wire  abc_mshr_4_io_status_bits_will_save_data; // @[Slice.scala 94:16]
  wire  abc_mshr_4_io_status_bits_will_free; // @[Slice.scala 94:16]
  wire  abc_mshr_4_io_resps_sink_c_valid; // @[Slice.scala 94:16]
  wire  abc_mshr_4_io_resps_sink_c_bits_hasData; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_4_io_resps_sink_c_bits_param; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_4_io_resps_sink_c_bits_source; // @[Slice.scala 94:16]
  wire  abc_mshr_4_io_resps_sink_c_bits_last; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_4_io_resps_sink_c_bits_bufIdx; // @[Slice.scala 94:16]
  wire  abc_mshr_4_io_resps_sink_d_valid; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_4_io_resps_sink_d_bits_opcode; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_4_io_resps_sink_d_bits_param; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_4_io_resps_sink_d_bits_sink; // @[Slice.scala 94:16]
  wire  abc_mshr_4_io_resps_sink_d_bits_last; // @[Slice.scala 94:16]
  wire  abc_mshr_4_io_resps_sink_d_bits_denied; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_4_io_resps_sink_d_bits_bufIdx; // @[Slice.scala 94:16]
  wire  abc_mshr_4_io_resps_sink_e_valid; // @[Slice.scala 94:16]
  wire  abc_mshr_4_io_resps_source_d_valid; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_4_io_nestedwb_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_4_io_nestedwb_tag; // @[Slice.scala 94:16]
  wire  abc_mshr_4_io_nestedwb_btoN; // @[Slice.scala 94:16]
  wire  abc_mshr_4_io_nestedwb_btoB; // @[Slice.scala 94:16]
  wire  abc_mshr_4_io_nestedwb_bclr_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_4_io_nestedwb_bset_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_4_io_nestedwb_c_set_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_4_io_nestedwb_c_set_hit; // @[Slice.scala 94:16]
  wire  abc_mshr_4_io_nestedwb_clients_0_isToN; // @[Slice.scala 94:16]
  wire  abc_mshr_4_io_nestedwb_clients_1_isToN; // @[Slice.scala 94:16]
  wire  abc_mshr_4_io_tasks_sink_a_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_4_io_tasks_sink_a_valid; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_4_io_tasks_sink_a_bits_sourceId; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_4_io_tasks_sink_a_bits_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_4_io_tasks_sink_a_bits_tag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_4_io_tasks_sink_a_bits_size; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_4_io_tasks_sink_a_bits_off; // @[Slice.scala 94:16]
  wire  abc_mshr_4_io_tasks_source_bready; // @[Slice.scala 94:16]
  wire  abc_mshr_4_io_tasks_source_bvalid; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_4_io_tasks_source_bset; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_4_io_tasks_source_btag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_4_io_tasks_source_bparam; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_4_io_tasks_source_bclients; // @[Slice.scala 94:16]
  wire  abc_mshr_4_io_tasks_source_bneedData; // @[Slice.scala 94:16]
  wire  abc_mshr_4_io_tasks_sink_c_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_4_io_tasks_sink_c_valid; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_4_io_tasks_sink_c_bits_sourceId; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_4_io_tasks_sink_c_bits_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_4_io_tasks_sink_c_bits_tag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_4_io_tasks_sink_c_bits_size; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_4_io_tasks_sink_c_bits_way; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_4_io_tasks_sink_c_bits_off; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_4_io_tasks_sink_c_bits_bufIdx; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_4_io_tasks_sink_c_bits_opcode; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_4_io_tasks_sink_c_bits_param; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_4_io_tasks_sink_c_bits_source; // @[Slice.scala 94:16]
  wire  abc_mshr_4_io_tasks_sink_c_bits_save; // @[Slice.scala 94:16]
  wire  abc_mshr_4_io_tasks_sink_c_bits_drop; // @[Slice.scala 94:16]
  wire  abc_mshr_4_io_tasks_sink_c_bits_release; // @[Slice.scala 94:16]
  wire  abc_mshr_4_io_tasks_sink_c_bits_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_4_io_tasks_source_d_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_4_io_tasks_source_d_valid; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_4_io_tasks_source_d_bits_sourceId; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_4_io_tasks_source_d_bits_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_4_io_tasks_source_d_bits_tag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_4_io_tasks_source_d_bits_channel; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_4_io_tasks_source_d_bits_opcode; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_4_io_tasks_source_d_bits_param; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_4_io_tasks_source_d_bits_size; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_4_io_tasks_source_d_bits_way; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_4_io_tasks_source_d_bits_off; // @[Slice.scala 94:16]
  wire  abc_mshr_4_io_tasks_source_d_bits_useBypass; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_4_io_tasks_source_d_bits_bufIdx; // @[Slice.scala 94:16]
  wire  abc_mshr_4_io_tasks_source_d_bits_denied; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_4_io_tasks_source_d_bits_sinkId; // @[Slice.scala 94:16]
  wire  abc_mshr_4_io_tasks_source_d_bits_bypassPut; // @[Slice.scala 94:16]
  wire  abc_mshr_4_io_tasks_source_d_bits_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_4_io_tasks_source_a_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_4_io_tasks_source_a_valid; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_4_io_tasks_source_a_bits_tag; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_4_io_tasks_source_a_bits_set; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_4_io_tasks_source_a_bits_off; // @[Slice.scala 94:16]
  wire [31:0] abc_mshr_4_io_tasks_source_a_bits_mask; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_4_io_tasks_source_a_bits_opcode; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_4_io_tasks_source_a_bits_param; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_4_io_tasks_source_a_bits_source; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_4_io_tasks_source_a_bits_bufIdx; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_4_io_tasks_source_a_bits_size; // @[Slice.scala 94:16]
  wire  abc_mshr_4_io_tasks_source_a_bits_needData; // @[Slice.scala 94:16]
  wire  abc_mshr_4_io_tasks_source_a_bits_putData; // @[Slice.scala 94:16]
  wire  abc_mshr_4_io_tasks_source_c_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_4_io_tasks_source_c_valid; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_4_io_tasks_source_c_bits_opcode; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_4_io_tasks_source_c_bits_tag; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_4_io_tasks_source_c_bits_set; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_4_io_tasks_source_c_bits_param; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_4_io_tasks_source_c_bits_source; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_4_io_tasks_source_c_bits_way; // @[Slice.scala 94:16]
  wire  abc_mshr_4_io_tasks_source_c_bits_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_4_io_tasks_source_e_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_4_io_tasks_source_e_valid; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_4_io_tasks_source_e_bits_sink; // @[Slice.scala 94:16]
  wire  abc_mshr_4_io_tasks_dir_write_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_4_io_tasks_dir_write_valid; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_4_io_tasks_dir_write_bits_set; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_4_io_tasks_dir_write_bits_way; // @[Slice.scala 94:16]
  wire  abc_mshr_4_io_tasks_dir_write_bits_data_dirty; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_4_io_tasks_dir_write_bits_data_state; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_4_io_tasks_dir_write_bits_data_clientStates_0; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_4_io_tasks_dir_write_bits_data_clientStates_1; // @[Slice.scala 94:16]
  wire  abc_mshr_4_io_tasks_tag_write_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_4_io_tasks_tag_write_valid; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_4_io_tasks_tag_write_bits_set; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_4_io_tasks_tag_write_bits_way; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_4_io_tasks_tag_write_bits_tag; // @[Slice.scala 94:16]
  wire  abc_mshr_4_io_tasks_client_dir_write_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_4_io_tasks_client_dir_write_valid; // @[Slice.scala 94:16]
  wire [6:0] abc_mshr_4_io_tasks_client_dir_write_bits_set; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_4_io_tasks_client_dir_write_bits_way; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_4_io_tasks_client_dir_write_bits_data_0_state; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_4_io_tasks_client_dir_write_bits_data_1_state; // @[Slice.scala 94:16]
  wire  abc_mshr_4_io_tasks_client_tag_write_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_4_io_tasks_client_tag_write_valid; // @[Slice.scala 94:16]
  wire [6:0] abc_mshr_4_io_tasks_client_tag_write_bits_set; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_4_io_tasks_client_tag_write_bits_way; // @[Slice.scala 94:16]
  wire [22:0] abc_mshr_4_io_tasks_client_tag_write_bits_tag; // @[Slice.scala 94:16]
  wire  abc_mshr_4_io_dirResult_valid; // @[Slice.scala 94:16]
  wire  abc_mshr_4_io_dirResult_bits_self_dirty; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_4_io_dirResult_bits_self_state; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_4_io_dirResult_bits_self_clientStates_0; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_4_io_dirResult_bits_self_clientStates_1; // @[Slice.scala 94:16]
  wire  abc_mshr_4_io_dirResult_bits_self_hit; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_4_io_dirResult_bits_self_way; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_4_io_dirResult_bits_self_tag; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_4_io_dirResult_bits_clients_states_0_state; // @[Slice.scala 94:16]
  wire  abc_mshr_4_io_dirResult_bits_clients_states_0_hit; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_4_io_dirResult_bits_clients_states_1_state; // @[Slice.scala 94:16]
  wire  abc_mshr_4_io_dirResult_bits_clients_states_1_hit; // @[Slice.scala 94:16]
  wire [22:0] abc_mshr_4_io_dirResult_bits_clients_tag; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_4_io_dirResult_bits_clients_way; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_4_io_c_status_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_4_io_c_status_tag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_4_io_c_status_way; // @[Slice.scala 94:16]
  wire  abc_mshr_4_io_c_status_nestedReleaseData; // @[Slice.scala 94:16]
  wire  abc_mshr_4_io_c_status_releaseThrough; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_4_io_bstatus_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_4_io_bstatus_tag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_4_io_bstatus_way; // @[Slice.scala 94:16]
  wire  abc_mshr_4_io_bstatus_nestedProbeAckData; // @[Slice.scala 94:16]
  wire  abc_mshr_4_io_bstatus_probeHelperFinish; // @[Slice.scala 94:16]
  wire  abc_mshr_4_io_bstatus_probeAckDataThrough; // @[Slice.scala 94:16]
  wire  abc_mshr_4_io_releaseThrough; // @[Slice.scala 94:16]
  wire  abc_mshr_4_io_probeAckDataThrough; // @[Slice.scala 94:16]
  wire  abc_mshr_4_io_is_nestedReleaseData; // @[Slice.scala 94:16]
  wire  abc_mshr_4_io_is_nestedProbeAckData; // @[Slice.scala 94:16]
  wire  abc_mshr_4_io_probeHelperFinish; // @[Slice.scala 94:16]
  wire  abc_mshr_5_clock; // @[Slice.scala 94:16]
  wire  abc_mshr_5_reset; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_5_io_id; // @[Slice.scala 94:16]
  wire  abc_mshr_5_io_enable; // @[Slice.scala 94:16]
  wire  abc_mshr_5_io_alloc_valid; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_5_io_alloc_bits_channel; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_5_io_alloc_bits_opcode; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_5_io_alloc_bits_param; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_5_io_alloc_bits_size; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_5_io_alloc_bits_source; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_5_io_alloc_bits_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_5_io_alloc_bits_tag; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_5_io_alloc_bits_off; // @[Slice.scala 94:16]
  wire [31:0] abc_mshr_5_io_alloc_bits_mask; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_5_io_alloc_bits_bufIdx; // @[Slice.scala 94:16]
  wire  abc_mshr_5_io_alloc_bits_preferCache; // @[Slice.scala 94:16]
  wire  abc_mshr_5_io_alloc_bits_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_5_io_alloc_bits_fromProbeHelper; // @[Slice.scala 94:16]
  wire  abc_mshr_5_io_alloc_bits_fromCmoHelper; // @[Slice.scala 94:16]
  wire  abc_mshr_5_io_alloc_bits_needProbeAckData; // @[Slice.scala 94:16]
  wire  abc_mshr_5_io_status_valid; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_5_io_status_bits_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_5_io_status_bits_tag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_5_io_status_bits_way; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_5_io_status_bits_way_reg; // @[Slice.scala 94:16]
  wire  abc_mshr_5_io_status_bits_nestB; // @[Slice.scala 94:16]
  wire  abc_mshr_5_io_status_bits_nestC; // @[Slice.scala 94:16]
  wire  abc_mshr_5_io_status_bits_will_grant_data; // @[Slice.scala 94:16]
  wire  abc_mshr_5_io_status_bits_will_save_data; // @[Slice.scala 94:16]
  wire  abc_mshr_5_io_status_bits_will_free; // @[Slice.scala 94:16]
  wire  abc_mshr_5_io_resps_sink_c_valid; // @[Slice.scala 94:16]
  wire  abc_mshr_5_io_resps_sink_c_bits_hasData; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_5_io_resps_sink_c_bits_param; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_5_io_resps_sink_c_bits_source; // @[Slice.scala 94:16]
  wire  abc_mshr_5_io_resps_sink_c_bits_last; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_5_io_resps_sink_c_bits_bufIdx; // @[Slice.scala 94:16]
  wire  abc_mshr_5_io_resps_sink_d_valid; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_5_io_resps_sink_d_bits_opcode; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_5_io_resps_sink_d_bits_param; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_5_io_resps_sink_d_bits_sink; // @[Slice.scala 94:16]
  wire  abc_mshr_5_io_resps_sink_d_bits_last; // @[Slice.scala 94:16]
  wire  abc_mshr_5_io_resps_sink_d_bits_denied; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_5_io_resps_sink_d_bits_bufIdx; // @[Slice.scala 94:16]
  wire  abc_mshr_5_io_resps_sink_e_valid; // @[Slice.scala 94:16]
  wire  abc_mshr_5_io_resps_source_d_valid; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_5_io_nestedwb_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_5_io_nestedwb_tag; // @[Slice.scala 94:16]
  wire  abc_mshr_5_io_nestedwb_btoN; // @[Slice.scala 94:16]
  wire  abc_mshr_5_io_nestedwb_btoB; // @[Slice.scala 94:16]
  wire  abc_mshr_5_io_nestedwb_bclr_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_5_io_nestedwb_bset_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_5_io_nestedwb_c_set_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_5_io_nestedwb_c_set_hit; // @[Slice.scala 94:16]
  wire  abc_mshr_5_io_nestedwb_clients_0_isToN; // @[Slice.scala 94:16]
  wire  abc_mshr_5_io_nestedwb_clients_1_isToN; // @[Slice.scala 94:16]
  wire  abc_mshr_5_io_tasks_sink_a_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_5_io_tasks_sink_a_valid; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_5_io_tasks_sink_a_bits_sourceId; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_5_io_tasks_sink_a_bits_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_5_io_tasks_sink_a_bits_tag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_5_io_tasks_sink_a_bits_size; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_5_io_tasks_sink_a_bits_off; // @[Slice.scala 94:16]
  wire  abc_mshr_5_io_tasks_source_bready; // @[Slice.scala 94:16]
  wire  abc_mshr_5_io_tasks_source_bvalid; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_5_io_tasks_source_bset; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_5_io_tasks_source_btag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_5_io_tasks_source_bparam; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_5_io_tasks_source_bclients; // @[Slice.scala 94:16]
  wire  abc_mshr_5_io_tasks_source_bneedData; // @[Slice.scala 94:16]
  wire  abc_mshr_5_io_tasks_sink_c_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_5_io_tasks_sink_c_valid; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_5_io_tasks_sink_c_bits_sourceId; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_5_io_tasks_sink_c_bits_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_5_io_tasks_sink_c_bits_tag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_5_io_tasks_sink_c_bits_size; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_5_io_tasks_sink_c_bits_way; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_5_io_tasks_sink_c_bits_off; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_5_io_tasks_sink_c_bits_bufIdx; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_5_io_tasks_sink_c_bits_opcode; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_5_io_tasks_sink_c_bits_param; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_5_io_tasks_sink_c_bits_source; // @[Slice.scala 94:16]
  wire  abc_mshr_5_io_tasks_sink_c_bits_save; // @[Slice.scala 94:16]
  wire  abc_mshr_5_io_tasks_sink_c_bits_drop; // @[Slice.scala 94:16]
  wire  abc_mshr_5_io_tasks_sink_c_bits_release; // @[Slice.scala 94:16]
  wire  abc_mshr_5_io_tasks_sink_c_bits_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_5_io_tasks_source_d_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_5_io_tasks_source_d_valid; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_5_io_tasks_source_d_bits_sourceId; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_5_io_tasks_source_d_bits_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_5_io_tasks_source_d_bits_tag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_5_io_tasks_source_d_bits_channel; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_5_io_tasks_source_d_bits_opcode; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_5_io_tasks_source_d_bits_param; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_5_io_tasks_source_d_bits_size; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_5_io_tasks_source_d_bits_way; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_5_io_tasks_source_d_bits_off; // @[Slice.scala 94:16]
  wire  abc_mshr_5_io_tasks_source_d_bits_useBypass; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_5_io_tasks_source_d_bits_bufIdx; // @[Slice.scala 94:16]
  wire  abc_mshr_5_io_tasks_source_d_bits_denied; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_5_io_tasks_source_d_bits_sinkId; // @[Slice.scala 94:16]
  wire  abc_mshr_5_io_tasks_source_d_bits_bypassPut; // @[Slice.scala 94:16]
  wire  abc_mshr_5_io_tasks_source_d_bits_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_5_io_tasks_source_a_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_5_io_tasks_source_a_valid; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_5_io_tasks_source_a_bits_tag; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_5_io_tasks_source_a_bits_set; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_5_io_tasks_source_a_bits_off; // @[Slice.scala 94:16]
  wire [31:0] abc_mshr_5_io_tasks_source_a_bits_mask; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_5_io_tasks_source_a_bits_opcode; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_5_io_tasks_source_a_bits_param; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_5_io_tasks_source_a_bits_source; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_5_io_tasks_source_a_bits_bufIdx; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_5_io_tasks_source_a_bits_size; // @[Slice.scala 94:16]
  wire  abc_mshr_5_io_tasks_source_a_bits_needData; // @[Slice.scala 94:16]
  wire  abc_mshr_5_io_tasks_source_a_bits_putData; // @[Slice.scala 94:16]
  wire  abc_mshr_5_io_tasks_source_c_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_5_io_tasks_source_c_valid; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_5_io_tasks_source_c_bits_opcode; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_5_io_tasks_source_c_bits_tag; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_5_io_tasks_source_c_bits_set; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_5_io_tasks_source_c_bits_param; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_5_io_tasks_source_c_bits_source; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_5_io_tasks_source_c_bits_way; // @[Slice.scala 94:16]
  wire  abc_mshr_5_io_tasks_source_c_bits_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_5_io_tasks_source_e_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_5_io_tasks_source_e_valid; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_5_io_tasks_source_e_bits_sink; // @[Slice.scala 94:16]
  wire  abc_mshr_5_io_tasks_dir_write_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_5_io_tasks_dir_write_valid; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_5_io_tasks_dir_write_bits_set; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_5_io_tasks_dir_write_bits_way; // @[Slice.scala 94:16]
  wire  abc_mshr_5_io_tasks_dir_write_bits_data_dirty; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_5_io_tasks_dir_write_bits_data_state; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_5_io_tasks_dir_write_bits_data_clientStates_0; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_5_io_tasks_dir_write_bits_data_clientStates_1; // @[Slice.scala 94:16]
  wire  abc_mshr_5_io_tasks_tag_write_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_5_io_tasks_tag_write_valid; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_5_io_tasks_tag_write_bits_set; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_5_io_tasks_tag_write_bits_way; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_5_io_tasks_tag_write_bits_tag; // @[Slice.scala 94:16]
  wire  abc_mshr_5_io_tasks_client_dir_write_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_5_io_tasks_client_dir_write_valid; // @[Slice.scala 94:16]
  wire [6:0] abc_mshr_5_io_tasks_client_dir_write_bits_set; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_5_io_tasks_client_dir_write_bits_way; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_5_io_tasks_client_dir_write_bits_data_0_state; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_5_io_tasks_client_dir_write_bits_data_1_state; // @[Slice.scala 94:16]
  wire  abc_mshr_5_io_tasks_client_tag_write_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_5_io_tasks_client_tag_write_valid; // @[Slice.scala 94:16]
  wire [6:0] abc_mshr_5_io_tasks_client_tag_write_bits_set; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_5_io_tasks_client_tag_write_bits_way; // @[Slice.scala 94:16]
  wire [22:0] abc_mshr_5_io_tasks_client_tag_write_bits_tag; // @[Slice.scala 94:16]
  wire  abc_mshr_5_io_dirResult_valid; // @[Slice.scala 94:16]
  wire  abc_mshr_5_io_dirResult_bits_self_dirty; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_5_io_dirResult_bits_self_state; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_5_io_dirResult_bits_self_clientStates_0; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_5_io_dirResult_bits_self_clientStates_1; // @[Slice.scala 94:16]
  wire  abc_mshr_5_io_dirResult_bits_self_hit; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_5_io_dirResult_bits_self_way; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_5_io_dirResult_bits_self_tag; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_5_io_dirResult_bits_clients_states_0_state; // @[Slice.scala 94:16]
  wire  abc_mshr_5_io_dirResult_bits_clients_states_0_hit; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_5_io_dirResult_bits_clients_states_1_state; // @[Slice.scala 94:16]
  wire  abc_mshr_5_io_dirResult_bits_clients_states_1_hit; // @[Slice.scala 94:16]
  wire [22:0] abc_mshr_5_io_dirResult_bits_clients_tag; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_5_io_dirResult_bits_clients_way; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_5_io_c_status_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_5_io_c_status_tag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_5_io_c_status_way; // @[Slice.scala 94:16]
  wire  abc_mshr_5_io_c_status_nestedReleaseData; // @[Slice.scala 94:16]
  wire  abc_mshr_5_io_c_status_releaseThrough; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_5_io_bstatus_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_5_io_bstatus_tag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_5_io_bstatus_way; // @[Slice.scala 94:16]
  wire  abc_mshr_5_io_bstatus_nestedProbeAckData; // @[Slice.scala 94:16]
  wire  abc_mshr_5_io_bstatus_probeHelperFinish; // @[Slice.scala 94:16]
  wire  abc_mshr_5_io_bstatus_probeAckDataThrough; // @[Slice.scala 94:16]
  wire  abc_mshr_5_io_releaseThrough; // @[Slice.scala 94:16]
  wire  abc_mshr_5_io_probeAckDataThrough; // @[Slice.scala 94:16]
  wire  abc_mshr_5_io_is_nestedReleaseData; // @[Slice.scala 94:16]
  wire  abc_mshr_5_io_is_nestedProbeAckData; // @[Slice.scala 94:16]
  wire  abc_mshr_5_io_probeHelperFinish; // @[Slice.scala 94:16]
  wire  abc_mshr_6_clock; // @[Slice.scala 94:16]
  wire  abc_mshr_6_reset; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_6_io_id; // @[Slice.scala 94:16]
  wire  abc_mshr_6_io_enable; // @[Slice.scala 94:16]
  wire  abc_mshr_6_io_alloc_valid; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_6_io_alloc_bits_channel; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_6_io_alloc_bits_opcode; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_6_io_alloc_bits_param; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_6_io_alloc_bits_size; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_6_io_alloc_bits_source; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_6_io_alloc_bits_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_6_io_alloc_bits_tag; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_6_io_alloc_bits_off; // @[Slice.scala 94:16]
  wire [31:0] abc_mshr_6_io_alloc_bits_mask; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_6_io_alloc_bits_bufIdx; // @[Slice.scala 94:16]
  wire  abc_mshr_6_io_alloc_bits_preferCache; // @[Slice.scala 94:16]
  wire  abc_mshr_6_io_alloc_bits_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_6_io_alloc_bits_fromProbeHelper; // @[Slice.scala 94:16]
  wire  abc_mshr_6_io_alloc_bits_fromCmoHelper; // @[Slice.scala 94:16]
  wire  abc_mshr_6_io_alloc_bits_needProbeAckData; // @[Slice.scala 94:16]
  wire  abc_mshr_6_io_status_valid; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_6_io_status_bits_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_6_io_status_bits_tag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_6_io_status_bits_way; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_6_io_status_bits_way_reg; // @[Slice.scala 94:16]
  wire  abc_mshr_6_io_status_bits_nestB; // @[Slice.scala 94:16]
  wire  abc_mshr_6_io_status_bits_nestC; // @[Slice.scala 94:16]
  wire  abc_mshr_6_io_status_bits_will_grant_data; // @[Slice.scala 94:16]
  wire  abc_mshr_6_io_status_bits_will_save_data; // @[Slice.scala 94:16]
  wire  abc_mshr_6_io_status_bits_will_free; // @[Slice.scala 94:16]
  wire  abc_mshr_6_io_resps_sink_c_valid; // @[Slice.scala 94:16]
  wire  abc_mshr_6_io_resps_sink_c_bits_hasData; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_6_io_resps_sink_c_bits_param; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_6_io_resps_sink_c_bits_source; // @[Slice.scala 94:16]
  wire  abc_mshr_6_io_resps_sink_c_bits_last; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_6_io_resps_sink_c_bits_bufIdx; // @[Slice.scala 94:16]
  wire  abc_mshr_6_io_resps_sink_d_valid; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_6_io_resps_sink_d_bits_opcode; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_6_io_resps_sink_d_bits_param; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_6_io_resps_sink_d_bits_sink; // @[Slice.scala 94:16]
  wire  abc_mshr_6_io_resps_sink_d_bits_last; // @[Slice.scala 94:16]
  wire  abc_mshr_6_io_resps_sink_d_bits_denied; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_6_io_resps_sink_d_bits_bufIdx; // @[Slice.scala 94:16]
  wire  abc_mshr_6_io_resps_sink_e_valid; // @[Slice.scala 94:16]
  wire  abc_mshr_6_io_resps_source_d_valid; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_6_io_nestedwb_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_6_io_nestedwb_tag; // @[Slice.scala 94:16]
  wire  abc_mshr_6_io_nestedwb_btoN; // @[Slice.scala 94:16]
  wire  abc_mshr_6_io_nestedwb_btoB; // @[Slice.scala 94:16]
  wire  abc_mshr_6_io_nestedwb_bclr_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_6_io_nestedwb_bset_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_6_io_nestedwb_c_set_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_6_io_nestedwb_c_set_hit; // @[Slice.scala 94:16]
  wire  abc_mshr_6_io_nestedwb_clients_0_isToN; // @[Slice.scala 94:16]
  wire  abc_mshr_6_io_nestedwb_clients_1_isToN; // @[Slice.scala 94:16]
  wire  abc_mshr_6_io_tasks_sink_a_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_6_io_tasks_sink_a_valid; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_6_io_tasks_sink_a_bits_sourceId; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_6_io_tasks_sink_a_bits_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_6_io_tasks_sink_a_bits_tag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_6_io_tasks_sink_a_bits_size; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_6_io_tasks_sink_a_bits_off; // @[Slice.scala 94:16]
  wire  abc_mshr_6_io_tasks_source_bready; // @[Slice.scala 94:16]
  wire  abc_mshr_6_io_tasks_source_bvalid; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_6_io_tasks_source_bset; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_6_io_tasks_source_btag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_6_io_tasks_source_bparam; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_6_io_tasks_source_bclients; // @[Slice.scala 94:16]
  wire  abc_mshr_6_io_tasks_source_bneedData; // @[Slice.scala 94:16]
  wire  abc_mshr_6_io_tasks_sink_c_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_6_io_tasks_sink_c_valid; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_6_io_tasks_sink_c_bits_sourceId; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_6_io_tasks_sink_c_bits_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_6_io_tasks_sink_c_bits_tag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_6_io_tasks_sink_c_bits_size; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_6_io_tasks_sink_c_bits_way; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_6_io_tasks_sink_c_bits_off; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_6_io_tasks_sink_c_bits_bufIdx; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_6_io_tasks_sink_c_bits_opcode; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_6_io_tasks_sink_c_bits_param; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_6_io_tasks_sink_c_bits_source; // @[Slice.scala 94:16]
  wire  abc_mshr_6_io_tasks_sink_c_bits_save; // @[Slice.scala 94:16]
  wire  abc_mshr_6_io_tasks_sink_c_bits_drop; // @[Slice.scala 94:16]
  wire  abc_mshr_6_io_tasks_sink_c_bits_release; // @[Slice.scala 94:16]
  wire  abc_mshr_6_io_tasks_sink_c_bits_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_6_io_tasks_source_d_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_6_io_tasks_source_d_valid; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_6_io_tasks_source_d_bits_sourceId; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_6_io_tasks_source_d_bits_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_6_io_tasks_source_d_bits_tag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_6_io_tasks_source_d_bits_channel; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_6_io_tasks_source_d_bits_opcode; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_6_io_tasks_source_d_bits_param; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_6_io_tasks_source_d_bits_size; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_6_io_tasks_source_d_bits_way; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_6_io_tasks_source_d_bits_off; // @[Slice.scala 94:16]
  wire  abc_mshr_6_io_tasks_source_d_bits_useBypass; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_6_io_tasks_source_d_bits_bufIdx; // @[Slice.scala 94:16]
  wire  abc_mshr_6_io_tasks_source_d_bits_denied; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_6_io_tasks_source_d_bits_sinkId; // @[Slice.scala 94:16]
  wire  abc_mshr_6_io_tasks_source_d_bits_bypassPut; // @[Slice.scala 94:16]
  wire  abc_mshr_6_io_tasks_source_d_bits_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_6_io_tasks_source_a_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_6_io_tasks_source_a_valid; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_6_io_tasks_source_a_bits_tag; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_6_io_tasks_source_a_bits_set; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_6_io_tasks_source_a_bits_off; // @[Slice.scala 94:16]
  wire [31:0] abc_mshr_6_io_tasks_source_a_bits_mask; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_6_io_tasks_source_a_bits_opcode; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_6_io_tasks_source_a_bits_param; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_6_io_tasks_source_a_bits_source; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_6_io_tasks_source_a_bits_bufIdx; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_6_io_tasks_source_a_bits_size; // @[Slice.scala 94:16]
  wire  abc_mshr_6_io_tasks_source_a_bits_needData; // @[Slice.scala 94:16]
  wire  abc_mshr_6_io_tasks_source_a_bits_putData; // @[Slice.scala 94:16]
  wire  abc_mshr_6_io_tasks_source_c_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_6_io_tasks_source_c_valid; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_6_io_tasks_source_c_bits_opcode; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_6_io_tasks_source_c_bits_tag; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_6_io_tasks_source_c_bits_set; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_6_io_tasks_source_c_bits_param; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_6_io_tasks_source_c_bits_source; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_6_io_tasks_source_c_bits_way; // @[Slice.scala 94:16]
  wire  abc_mshr_6_io_tasks_source_c_bits_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_6_io_tasks_source_e_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_6_io_tasks_source_e_valid; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_6_io_tasks_source_e_bits_sink; // @[Slice.scala 94:16]
  wire  abc_mshr_6_io_tasks_dir_write_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_6_io_tasks_dir_write_valid; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_6_io_tasks_dir_write_bits_set; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_6_io_tasks_dir_write_bits_way; // @[Slice.scala 94:16]
  wire  abc_mshr_6_io_tasks_dir_write_bits_data_dirty; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_6_io_tasks_dir_write_bits_data_state; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_6_io_tasks_dir_write_bits_data_clientStates_0; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_6_io_tasks_dir_write_bits_data_clientStates_1; // @[Slice.scala 94:16]
  wire  abc_mshr_6_io_tasks_tag_write_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_6_io_tasks_tag_write_valid; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_6_io_tasks_tag_write_bits_set; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_6_io_tasks_tag_write_bits_way; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_6_io_tasks_tag_write_bits_tag; // @[Slice.scala 94:16]
  wire  abc_mshr_6_io_tasks_client_dir_write_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_6_io_tasks_client_dir_write_valid; // @[Slice.scala 94:16]
  wire [6:0] abc_mshr_6_io_tasks_client_dir_write_bits_set; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_6_io_tasks_client_dir_write_bits_way; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_6_io_tasks_client_dir_write_bits_data_0_state; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_6_io_tasks_client_dir_write_bits_data_1_state; // @[Slice.scala 94:16]
  wire  abc_mshr_6_io_tasks_client_tag_write_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_6_io_tasks_client_tag_write_valid; // @[Slice.scala 94:16]
  wire [6:0] abc_mshr_6_io_tasks_client_tag_write_bits_set; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_6_io_tasks_client_tag_write_bits_way; // @[Slice.scala 94:16]
  wire [22:0] abc_mshr_6_io_tasks_client_tag_write_bits_tag; // @[Slice.scala 94:16]
  wire  abc_mshr_6_io_dirResult_valid; // @[Slice.scala 94:16]
  wire  abc_mshr_6_io_dirResult_bits_self_dirty; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_6_io_dirResult_bits_self_state; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_6_io_dirResult_bits_self_clientStates_0; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_6_io_dirResult_bits_self_clientStates_1; // @[Slice.scala 94:16]
  wire  abc_mshr_6_io_dirResult_bits_self_hit; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_6_io_dirResult_bits_self_way; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_6_io_dirResult_bits_self_tag; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_6_io_dirResult_bits_clients_states_0_state; // @[Slice.scala 94:16]
  wire  abc_mshr_6_io_dirResult_bits_clients_states_0_hit; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_6_io_dirResult_bits_clients_states_1_state; // @[Slice.scala 94:16]
  wire  abc_mshr_6_io_dirResult_bits_clients_states_1_hit; // @[Slice.scala 94:16]
  wire [22:0] abc_mshr_6_io_dirResult_bits_clients_tag; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_6_io_dirResult_bits_clients_way; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_6_io_c_status_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_6_io_c_status_tag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_6_io_c_status_way; // @[Slice.scala 94:16]
  wire  abc_mshr_6_io_c_status_nestedReleaseData; // @[Slice.scala 94:16]
  wire  abc_mshr_6_io_c_status_releaseThrough; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_6_io_bstatus_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_6_io_bstatus_tag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_6_io_bstatus_way; // @[Slice.scala 94:16]
  wire  abc_mshr_6_io_bstatus_nestedProbeAckData; // @[Slice.scala 94:16]
  wire  abc_mshr_6_io_bstatus_probeHelperFinish; // @[Slice.scala 94:16]
  wire  abc_mshr_6_io_bstatus_probeAckDataThrough; // @[Slice.scala 94:16]
  wire  abc_mshr_6_io_releaseThrough; // @[Slice.scala 94:16]
  wire  abc_mshr_6_io_probeAckDataThrough; // @[Slice.scala 94:16]
  wire  abc_mshr_6_io_is_nestedReleaseData; // @[Slice.scala 94:16]
  wire  abc_mshr_6_io_is_nestedProbeAckData; // @[Slice.scala 94:16]
  wire  abc_mshr_6_io_probeHelperFinish; // @[Slice.scala 94:16]
  wire  abc_mshr_7_clock; // @[Slice.scala 94:16]
  wire  abc_mshr_7_reset; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_7_io_id; // @[Slice.scala 94:16]
  wire  abc_mshr_7_io_enable; // @[Slice.scala 94:16]
  wire  abc_mshr_7_io_alloc_valid; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_7_io_alloc_bits_channel; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_7_io_alloc_bits_opcode; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_7_io_alloc_bits_param; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_7_io_alloc_bits_size; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_7_io_alloc_bits_source; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_7_io_alloc_bits_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_7_io_alloc_bits_tag; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_7_io_alloc_bits_off; // @[Slice.scala 94:16]
  wire [31:0] abc_mshr_7_io_alloc_bits_mask; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_7_io_alloc_bits_bufIdx; // @[Slice.scala 94:16]
  wire  abc_mshr_7_io_alloc_bits_preferCache; // @[Slice.scala 94:16]
  wire  abc_mshr_7_io_alloc_bits_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_7_io_alloc_bits_fromProbeHelper; // @[Slice.scala 94:16]
  wire  abc_mshr_7_io_alloc_bits_fromCmoHelper; // @[Slice.scala 94:16]
  wire  abc_mshr_7_io_alloc_bits_needProbeAckData; // @[Slice.scala 94:16]
  wire  abc_mshr_7_io_status_valid; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_7_io_status_bits_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_7_io_status_bits_tag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_7_io_status_bits_way; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_7_io_status_bits_way_reg; // @[Slice.scala 94:16]
  wire  abc_mshr_7_io_status_bits_nestB; // @[Slice.scala 94:16]
  wire  abc_mshr_7_io_status_bits_nestC; // @[Slice.scala 94:16]
  wire  abc_mshr_7_io_status_bits_will_grant_data; // @[Slice.scala 94:16]
  wire  abc_mshr_7_io_status_bits_will_save_data; // @[Slice.scala 94:16]
  wire  abc_mshr_7_io_status_bits_will_free; // @[Slice.scala 94:16]
  wire  abc_mshr_7_io_resps_sink_c_valid; // @[Slice.scala 94:16]
  wire  abc_mshr_7_io_resps_sink_c_bits_hasData; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_7_io_resps_sink_c_bits_param; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_7_io_resps_sink_c_bits_source; // @[Slice.scala 94:16]
  wire  abc_mshr_7_io_resps_sink_c_bits_last; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_7_io_resps_sink_c_bits_bufIdx; // @[Slice.scala 94:16]
  wire  abc_mshr_7_io_resps_sink_d_valid; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_7_io_resps_sink_d_bits_opcode; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_7_io_resps_sink_d_bits_param; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_7_io_resps_sink_d_bits_sink; // @[Slice.scala 94:16]
  wire  abc_mshr_7_io_resps_sink_d_bits_last; // @[Slice.scala 94:16]
  wire  abc_mshr_7_io_resps_sink_d_bits_denied; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_7_io_resps_sink_d_bits_bufIdx; // @[Slice.scala 94:16]
  wire  abc_mshr_7_io_resps_sink_e_valid; // @[Slice.scala 94:16]
  wire  abc_mshr_7_io_resps_source_d_valid; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_7_io_nestedwb_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_7_io_nestedwb_tag; // @[Slice.scala 94:16]
  wire  abc_mshr_7_io_nestedwb_btoN; // @[Slice.scala 94:16]
  wire  abc_mshr_7_io_nestedwb_btoB; // @[Slice.scala 94:16]
  wire  abc_mshr_7_io_nestedwb_bclr_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_7_io_nestedwb_bset_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_7_io_nestedwb_c_set_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_7_io_nestedwb_c_set_hit; // @[Slice.scala 94:16]
  wire  abc_mshr_7_io_nestedwb_clients_0_isToN; // @[Slice.scala 94:16]
  wire  abc_mshr_7_io_nestedwb_clients_1_isToN; // @[Slice.scala 94:16]
  wire  abc_mshr_7_io_tasks_sink_a_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_7_io_tasks_sink_a_valid; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_7_io_tasks_sink_a_bits_sourceId; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_7_io_tasks_sink_a_bits_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_7_io_tasks_sink_a_bits_tag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_7_io_tasks_sink_a_bits_size; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_7_io_tasks_sink_a_bits_off; // @[Slice.scala 94:16]
  wire  abc_mshr_7_io_tasks_source_bready; // @[Slice.scala 94:16]
  wire  abc_mshr_7_io_tasks_source_bvalid; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_7_io_tasks_source_bset; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_7_io_tasks_source_btag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_7_io_tasks_source_bparam; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_7_io_tasks_source_bclients; // @[Slice.scala 94:16]
  wire  abc_mshr_7_io_tasks_source_bneedData; // @[Slice.scala 94:16]
  wire  abc_mshr_7_io_tasks_sink_c_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_7_io_tasks_sink_c_valid; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_7_io_tasks_sink_c_bits_sourceId; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_7_io_tasks_sink_c_bits_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_7_io_tasks_sink_c_bits_tag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_7_io_tasks_sink_c_bits_size; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_7_io_tasks_sink_c_bits_way; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_7_io_tasks_sink_c_bits_off; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_7_io_tasks_sink_c_bits_bufIdx; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_7_io_tasks_sink_c_bits_opcode; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_7_io_tasks_sink_c_bits_param; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_7_io_tasks_sink_c_bits_source; // @[Slice.scala 94:16]
  wire  abc_mshr_7_io_tasks_sink_c_bits_save; // @[Slice.scala 94:16]
  wire  abc_mshr_7_io_tasks_sink_c_bits_drop; // @[Slice.scala 94:16]
  wire  abc_mshr_7_io_tasks_sink_c_bits_release; // @[Slice.scala 94:16]
  wire  abc_mshr_7_io_tasks_sink_c_bits_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_7_io_tasks_source_d_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_7_io_tasks_source_d_valid; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_7_io_tasks_source_d_bits_sourceId; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_7_io_tasks_source_d_bits_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_7_io_tasks_source_d_bits_tag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_7_io_tasks_source_d_bits_channel; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_7_io_tasks_source_d_bits_opcode; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_7_io_tasks_source_d_bits_param; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_7_io_tasks_source_d_bits_size; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_7_io_tasks_source_d_bits_way; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_7_io_tasks_source_d_bits_off; // @[Slice.scala 94:16]
  wire  abc_mshr_7_io_tasks_source_d_bits_useBypass; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_7_io_tasks_source_d_bits_bufIdx; // @[Slice.scala 94:16]
  wire  abc_mshr_7_io_tasks_source_d_bits_denied; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_7_io_tasks_source_d_bits_sinkId; // @[Slice.scala 94:16]
  wire  abc_mshr_7_io_tasks_source_d_bits_bypassPut; // @[Slice.scala 94:16]
  wire  abc_mshr_7_io_tasks_source_d_bits_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_7_io_tasks_source_a_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_7_io_tasks_source_a_valid; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_7_io_tasks_source_a_bits_tag; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_7_io_tasks_source_a_bits_set; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_7_io_tasks_source_a_bits_off; // @[Slice.scala 94:16]
  wire [31:0] abc_mshr_7_io_tasks_source_a_bits_mask; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_7_io_tasks_source_a_bits_opcode; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_7_io_tasks_source_a_bits_param; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_7_io_tasks_source_a_bits_source; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_7_io_tasks_source_a_bits_bufIdx; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_7_io_tasks_source_a_bits_size; // @[Slice.scala 94:16]
  wire  abc_mshr_7_io_tasks_source_a_bits_needData; // @[Slice.scala 94:16]
  wire  abc_mshr_7_io_tasks_source_a_bits_putData; // @[Slice.scala 94:16]
  wire  abc_mshr_7_io_tasks_source_c_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_7_io_tasks_source_c_valid; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_7_io_tasks_source_c_bits_opcode; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_7_io_tasks_source_c_bits_tag; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_7_io_tasks_source_c_bits_set; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_7_io_tasks_source_c_bits_param; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_7_io_tasks_source_c_bits_source; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_7_io_tasks_source_c_bits_way; // @[Slice.scala 94:16]
  wire  abc_mshr_7_io_tasks_source_c_bits_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_7_io_tasks_source_e_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_7_io_tasks_source_e_valid; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_7_io_tasks_source_e_bits_sink; // @[Slice.scala 94:16]
  wire  abc_mshr_7_io_tasks_dir_write_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_7_io_tasks_dir_write_valid; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_7_io_tasks_dir_write_bits_set; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_7_io_tasks_dir_write_bits_way; // @[Slice.scala 94:16]
  wire  abc_mshr_7_io_tasks_dir_write_bits_data_dirty; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_7_io_tasks_dir_write_bits_data_state; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_7_io_tasks_dir_write_bits_data_clientStates_0; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_7_io_tasks_dir_write_bits_data_clientStates_1; // @[Slice.scala 94:16]
  wire  abc_mshr_7_io_tasks_tag_write_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_7_io_tasks_tag_write_valid; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_7_io_tasks_tag_write_bits_set; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_7_io_tasks_tag_write_bits_way; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_7_io_tasks_tag_write_bits_tag; // @[Slice.scala 94:16]
  wire  abc_mshr_7_io_tasks_client_dir_write_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_7_io_tasks_client_dir_write_valid; // @[Slice.scala 94:16]
  wire [6:0] abc_mshr_7_io_tasks_client_dir_write_bits_set; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_7_io_tasks_client_dir_write_bits_way; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_7_io_tasks_client_dir_write_bits_data_0_state; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_7_io_tasks_client_dir_write_bits_data_1_state; // @[Slice.scala 94:16]
  wire  abc_mshr_7_io_tasks_client_tag_write_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_7_io_tasks_client_tag_write_valid; // @[Slice.scala 94:16]
  wire [6:0] abc_mshr_7_io_tasks_client_tag_write_bits_set; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_7_io_tasks_client_tag_write_bits_way; // @[Slice.scala 94:16]
  wire [22:0] abc_mshr_7_io_tasks_client_tag_write_bits_tag; // @[Slice.scala 94:16]
  wire  abc_mshr_7_io_dirResult_valid; // @[Slice.scala 94:16]
  wire  abc_mshr_7_io_dirResult_bits_self_dirty; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_7_io_dirResult_bits_self_state; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_7_io_dirResult_bits_self_clientStates_0; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_7_io_dirResult_bits_self_clientStates_1; // @[Slice.scala 94:16]
  wire  abc_mshr_7_io_dirResult_bits_self_hit; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_7_io_dirResult_bits_self_way; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_7_io_dirResult_bits_self_tag; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_7_io_dirResult_bits_clients_states_0_state; // @[Slice.scala 94:16]
  wire  abc_mshr_7_io_dirResult_bits_clients_states_0_hit; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_7_io_dirResult_bits_clients_states_1_state; // @[Slice.scala 94:16]
  wire  abc_mshr_7_io_dirResult_bits_clients_states_1_hit; // @[Slice.scala 94:16]
  wire [22:0] abc_mshr_7_io_dirResult_bits_clients_tag; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_7_io_dirResult_bits_clients_way; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_7_io_c_status_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_7_io_c_status_tag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_7_io_c_status_way; // @[Slice.scala 94:16]
  wire  abc_mshr_7_io_c_status_nestedReleaseData; // @[Slice.scala 94:16]
  wire  abc_mshr_7_io_c_status_releaseThrough; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_7_io_bstatus_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_7_io_bstatus_tag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_7_io_bstatus_way; // @[Slice.scala 94:16]
  wire  abc_mshr_7_io_bstatus_nestedProbeAckData; // @[Slice.scala 94:16]
  wire  abc_mshr_7_io_bstatus_probeHelperFinish; // @[Slice.scala 94:16]
  wire  abc_mshr_7_io_bstatus_probeAckDataThrough; // @[Slice.scala 94:16]
  wire  abc_mshr_7_io_releaseThrough; // @[Slice.scala 94:16]
  wire  abc_mshr_7_io_probeAckDataThrough; // @[Slice.scala 94:16]
  wire  abc_mshr_7_io_is_nestedReleaseData; // @[Slice.scala 94:16]
  wire  abc_mshr_7_io_is_nestedProbeAckData; // @[Slice.scala 94:16]
  wire  abc_mshr_7_io_probeHelperFinish; // @[Slice.scala 94:16]
  wire  abc_mshr_8_clock; // @[Slice.scala 94:16]
  wire  abc_mshr_8_reset; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_8_io_id; // @[Slice.scala 94:16]
  wire  abc_mshr_8_io_enable; // @[Slice.scala 94:16]
  wire  abc_mshr_8_io_alloc_valid; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_8_io_alloc_bits_channel; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_8_io_alloc_bits_opcode; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_8_io_alloc_bits_param; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_8_io_alloc_bits_size; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_8_io_alloc_bits_source; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_8_io_alloc_bits_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_8_io_alloc_bits_tag; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_8_io_alloc_bits_off; // @[Slice.scala 94:16]
  wire [31:0] abc_mshr_8_io_alloc_bits_mask; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_8_io_alloc_bits_bufIdx; // @[Slice.scala 94:16]
  wire  abc_mshr_8_io_alloc_bits_preferCache; // @[Slice.scala 94:16]
  wire  abc_mshr_8_io_alloc_bits_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_8_io_alloc_bits_fromProbeHelper; // @[Slice.scala 94:16]
  wire  abc_mshr_8_io_alloc_bits_fromCmoHelper; // @[Slice.scala 94:16]
  wire  abc_mshr_8_io_alloc_bits_needProbeAckData; // @[Slice.scala 94:16]
  wire  abc_mshr_8_io_status_valid; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_8_io_status_bits_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_8_io_status_bits_tag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_8_io_status_bits_way; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_8_io_status_bits_way_reg; // @[Slice.scala 94:16]
  wire  abc_mshr_8_io_status_bits_nestB; // @[Slice.scala 94:16]
  wire  abc_mshr_8_io_status_bits_nestC; // @[Slice.scala 94:16]
  wire  abc_mshr_8_io_status_bits_will_grant_data; // @[Slice.scala 94:16]
  wire  abc_mshr_8_io_status_bits_will_save_data; // @[Slice.scala 94:16]
  wire  abc_mshr_8_io_status_bits_will_free; // @[Slice.scala 94:16]
  wire  abc_mshr_8_io_resps_sink_c_valid; // @[Slice.scala 94:16]
  wire  abc_mshr_8_io_resps_sink_c_bits_hasData; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_8_io_resps_sink_c_bits_param; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_8_io_resps_sink_c_bits_source; // @[Slice.scala 94:16]
  wire  abc_mshr_8_io_resps_sink_c_bits_last; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_8_io_resps_sink_c_bits_bufIdx; // @[Slice.scala 94:16]
  wire  abc_mshr_8_io_resps_sink_d_valid; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_8_io_resps_sink_d_bits_opcode; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_8_io_resps_sink_d_bits_param; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_8_io_resps_sink_d_bits_sink; // @[Slice.scala 94:16]
  wire  abc_mshr_8_io_resps_sink_d_bits_last; // @[Slice.scala 94:16]
  wire  abc_mshr_8_io_resps_sink_d_bits_denied; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_8_io_resps_sink_d_bits_bufIdx; // @[Slice.scala 94:16]
  wire  abc_mshr_8_io_resps_sink_e_valid; // @[Slice.scala 94:16]
  wire  abc_mshr_8_io_resps_source_d_valid; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_8_io_nestedwb_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_8_io_nestedwb_tag; // @[Slice.scala 94:16]
  wire  abc_mshr_8_io_nestedwb_btoN; // @[Slice.scala 94:16]
  wire  abc_mshr_8_io_nestedwb_btoB; // @[Slice.scala 94:16]
  wire  abc_mshr_8_io_nestedwb_bclr_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_8_io_nestedwb_bset_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_8_io_nestedwb_c_set_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_8_io_nestedwb_c_set_hit; // @[Slice.scala 94:16]
  wire  abc_mshr_8_io_nestedwb_clients_0_isToN; // @[Slice.scala 94:16]
  wire  abc_mshr_8_io_nestedwb_clients_1_isToN; // @[Slice.scala 94:16]
  wire  abc_mshr_8_io_tasks_sink_a_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_8_io_tasks_sink_a_valid; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_8_io_tasks_sink_a_bits_sourceId; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_8_io_tasks_sink_a_bits_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_8_io_tasks_sink_a_bits_tag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_8_io_tasks_sink_a_bits_size; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_8_io_tasks_sink_a_bits_off; // @[Slice.scala 94:16]
  wire  abc_mshr_8_io_tasks_source_bready; // @[Slice.scala 94:16]
  wire  abc_mshr_8_io_tasks_source_bvalid; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_8_io_tasks_source_bset; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_8_io_tasks_source_btag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_8_io_tasks_source_bparam; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_8_io_tasks_source_bclients; // @[Slice.scala 94:16]
  wire  abc_mshr_8_io_tasks_source_bneedData; // @[Slice.scala 94:16]
  wire  abc_mshr_8_io_tasks_sink_c_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_8_io_tasks_sink_c_valid; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_8_io_tasks_sink_c_bits_sourceId; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_8_io_tasks_sink_c_bits_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_8_io_tasks_sink_c_bits_tag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_8_io_tasks_sink_c_bits_size; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_8_io_tasks_sink_c_bits_way; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_8_io_tasks_sink_c_bits_off; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_8_io_tasks_sink_c_bits_bufIdx; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_8_io_tasks_sink_c_bits_opcode; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_8_io_tasks_sink_c_bits_param; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_8_io_tasks_sink_c_bits_source; // @[Slice.scala 94:16]
  wire  abc_mshr_8_io_tasks_sink_c_bits_save; // @[Slice.scala 94:16]
  wire  abc_mshr_8_io_tasks_sink_c_bits_drop; // @[Slice.scala 94:16]
  wire  abc_mshr_8_io_tasks_sink_c_bits_release; // @[Slice.scala 94:16]
  wire  abc_mshr_8_io_tasks_sink_c_bits_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_8_io_tasks_source_d_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_8_io_tasks_source_d_valid; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_8_io_tasks_source_d_bits_sourceId; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_8_io_tasks_source_d_bits_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_8_io_tasks_source_d_bits_tag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_8_io_tasks_source_d_bits_channel; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_8_io_tasks_source_d_bits_opcode; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_8_io_tasks_source_d_bits_param; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_8_io_tasks_source_d_bits_size; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_8_io_tasks_source_d_bits_way; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_8_io_tasks_source_d_bits_off; // @[Slice.scala 94:16]
  wire  abc_mshr_8_io_tasks_source_d_bits_useBypass; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_8_io_tasks_source_d_bits_bufIdx; // @[Slice.scala 94:16]
  wire  abc_mshr_8_io_tasks_source_d_bits_denied; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_8_io_tasks_source_d_bits_sinkId; // @[Slice.scala 94:16]
  wire  abc_mshr_8_io_tasks_source_d_bits_bypassPut; // @[Slice.scala 94:16]
  wire  abc_mshr_8_io_tasks_source_d_bits_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_8_io_tasks_source_a_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_8_io_tasks_source_a_valid; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_8_io_tasks_source_a_bits_tag; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_8_io_tasks_source_a_bits_set; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_8_io_tasks_source_a_bits_off; // @[Slice.scala 94:16]
  wire [31:0] abc_mshr_8_io_tasks_source_a_bits_mask; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_8_io_tasks_source_a_bits_opcode; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_8_io_tasks_source_a_bits_param; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_8_io_tasks_source_a_bits_source; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_8_io_tasks_source_a_bits_bufIdx; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_8_io_tasks_source_a_bits_size; // @[Slice.scala 94:16]
  wire  abc_mshr_8_io_tasks_source_a_bits_needData; // @[Slice.scala 94:16]
  wire  abc_mshr_8_io_tasks_source_a_bits_putData; // @[Slice.scala 94:16]
  wire  abc_mshr_8_io_tasks_source_c_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_8_io_tasks_source_c_valid; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_8_io_tasks_source_c_bits_opcode; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_8_io_tasks_source_c_bits_tag; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_8_io_tasks_source_c_bits_set; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_8_io_tasks_source_c_bits_param; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_8_io_tasks_source_c_bits_source; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_8_io_tasks_source_c_bits_way; // @[Slice.scala 94:16]
  wire  abc_mshr_8_io_tasks_source_c_bits_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_8_io_tasks_source_e_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_8_io_tasks_source_e_valid; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_8_io_tasks_source_e_bits_sink; // @[Slice.scala 94:16]
  wire  abc_mshr_8_io_tasks_dir_write_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_8_io_tasks_dir_write_valid; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_8_io_tasks_dir_write_bits_set; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_8_io_tasks_dir_write_bits_way; // @[Slice.scala 94:16]
  wire  abc_mshr_8_io_tasks_dir_write_bits_data_dirty; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_8_io_tasks_dir_write_bits_data_state; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_8_io_tasks_dir_write_bits_data_clientStates_0; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_8_io_tasks_dir_write_bits_data_clientStates_1; // @[Slice.scala 94:16]
  wire  abc_mshr_8_io_tasks_tag_write_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_8_io_tasks_tag_write_valid; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_8_io_tasks_tag_write_bits_set; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_8_io_tasks_tag_write_bits_way; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_8_io_tasks_tag_write_bits_tag; // @[Slice.scala 94:16]
  wire  abc_mshr_8_io_tasks_client_dir_write_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_8_io_tasks_client_dir_write_valid; // @[Slice.scala 94:16]
  wire [6:0] abc_mshr_8_io_tasks_client_dir_write_bits_set; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_8_io_tasks_client_dir_write_bits_way; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_8_io_tasks_client_dir_write_bits_data_0_state; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_8_io_tasks_client_dir_write_bits_data_1_state; // @[Slice.scala 94:16]
  wire  abc_mshr_8_io_tasks_client_tag_write_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_8_io_tasks_client_tag_write_valid; // @[Slice.scala 94:16]
  wire [6:0] abc_mshr_8_io_tasks_client_tag_write_bits_set; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_8_io_tasks_client_tag_write_bits_way; // @[Slice.scala 94:16]
  wire [22:0] abc_mshr_8_io_tasks_client_tag_write_bits_tag; // @[Slice.scala 94:16]
  wire  abc_mshr_8_io_dirResult_valid; // @[Slice.scala 94:16]
  wire  abc_mshr_8_io_dirResult_bits_self_dirty; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_8_io_dirResult_bits_self_state; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_8_io_dirResult_bits_self_clientStates_0; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_8_io_dirResult_bits_self_clientStates_1; // @[Slice.scala 94:16]
  wire  abc_mshr_8_io_dirResult_bits_self_hit; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_8_io_dirResult_bits_self_way; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_8_io_dirResult_bits_self_tag; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_8_io_dirResult_bits_clients_states_0_state; // @[Slice.scala 94:16]
  wire  abc_mshr_8_io_dirResult_bits_clients_states_0_hit; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_8_io_dirResult_bits_clients_states_1_state; // @[Slice.scala 94:16]
  wire  abc_mshr_8_io_dirResult_bits_clients_states_1_hit; // @[Slice.scala 94:16]
  wire [22:0] abc_mshr_8_io_dirResult_bits_clients_tag; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_8_io_dirResult_bits_clients_way; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_8_io_c_status_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_8_io_c_status_tag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_8_io_c_status_way; // @[Slice.scala 94:16]
  wire  abc_mshr_8_io_c_status_nestedReleaseData; // @[Slice.scala 94:16]
  wire  abc_mshr_8_io_c_status_releaseThrough; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_8_io_bstatus_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_8_io_bstatus_tag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_8_io_bstatus_way; // @[Slice.scala 94:16]
  wire  abc_mshr_8_io_bstatus_nestedProbeAckData; // @[Slice.scala 94:16]
  wire  abc_mshr_8_io_bstatus_probeHelperFinish; // @[Slice.scala 94:16]
  wire  abc_mshr_8_io_bstatus_probeAckDataThrough; // @[Slice.scala 94:16]
  wire  abc_mshr_8_io_releaseThrough; // @[Slice.scala 94:16]
  wire  abc_mshr_8_io_probeAckDataThrough; // @[Slice.scala 94:16]
  wire  abc_mshr_8_io_is_nestedReleaseData; // @[Slice.scala 94:16]
  wire  abc_mshr_8_io_is_nestedProbeAckData; // @[Slice.scala 94:16]
  wire  abc_mshr_8_io_probeHelperFinish; // @[Slice.scala 94:16]
  wire  abc_mshr_9_clock; // @[Slice.scala 94:16]
  wire  abc_mshr_9_reset; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_9_io_id; // @[Slice.scala 94:16]
  wire  abc_mshr_9_io_enable; // @[Slice.scala 94:16]
  wire  abc_mshr_9_io_alloc_valid; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_9_io_alloc_bits_channel; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_9_io_alloc_bits_opcode; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_9_io_alloc_bits_param; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_9_io_alloc_bits_size; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_9_io_alloc_bits_source; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_9_io_alloc_bits_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_9_io_alloc_bits_tag; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_9_io_alloc_bits_off; // @[Slice.scala 94:16]
  wire [31:0] abc_mshr_9_io_alloc_bits_mask; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_9_io_alloc_bits_bufIdx; // @[Slice.scala 94:16]
  wire  abc_mshr_9_io_alloc_bits_preferCache; // @[Slice.scala 94:16]
  wire  abc_mshr_9_io_alloc_bits_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_9_io_alloc_bits_fromProbeHelper; // @[Slice.scala 94:16]
  wire  abc_mshr_9_io_alloc_bits_fromCmoHelper; // @[Slice.scala 94:16]
  wire  abc_mshr_9_io_alloc_bits_needProbeAckData; // @[Slice.scala 94:16]
  wire  abc_mshr_9_io_status_valid; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_9_io_status_bits_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_9_io_status_bits_tag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_9_io_status_bits_way; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_9_io_status_bits_way_reg; // @[Slice.scala 94:16]
  wire  abc_mshr_9_io_status_bits_nestB; // @[Slice.scala 94:16]
  wire  abc_mshr_9_io_status_bits_nestC; // @[Slice.scala 94:16]
  wire  abc_mshr_9_io_status_bits_will_grant_data; // @[Slice.scala 94:16]
  wire  abc_mshr_9_io_status_bits_will_save_data; // @[Slice.scala 94:16]
  wire  abc_mshr_9_io_status_bits_will_free; // @[Slice.scala 94:16]
  wire  abc_mshr_9_io_resps_sink_c_valid; // @[Slice.scala 94:16]
  wire  abc_mshr_9_io_resps_sink_c_bits_hasData; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_9_io_resps_sink_c_bits_param; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_9_io_resps_sink_c_bits_source; // @[Slice.scala 94:16]
  wire  abc_mshr_9_io_resps_sink_c_bits_last; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_9_io_resps_sink_c_bits_bufIdx; // @[Slice.scala 94:16]
  wire  abc_mshr_9_io_resps_sink_d_valid; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_9_io_resps_sink_d_bits_opcode; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_9_io_resps_sink_d_bits_param; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_9_io_resps_sink_d_bits_sink; // @[Slice.scala 94:16]
  wire  abc_mshr_9_io_resps_sink_d_bits_last; // @[Slice.scala 94:16]
  wire  abc_mshr_9_io_resps_sink_d_bits_denied; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_9_io_resps_sink_d_bits_bufIdx; // @[Slice.scala 94:16]
  wire  abc_mshr_9_io_resps_sink_e_valid; // @[Slice.scala 94:16]
  wire  abc_mshr_9_io_resps_source_d_valid; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_9_io_nestedwb_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_9_io_nestedwb_tag; // @[Slice.scala 94:16]
  wire  abc_mshr_9_io_nestedwb_btoN; // @[Slice.scala 94:16]
  wire  abc_mshr_9_io_nestedwb_btoB; // @[Slice.scala 94:16]
  wire  abc_mshr_9_io_nestedwb_bclr_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_9_io_nestedwb_bset_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_9_io_nestedwb_c_set_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_9_io_nestedwb_c_set_hit; // @[Slice.scala 94:16]
  wire  abc_mshr_9_io_nestedwb_clients_0_isToN; // @[Slice.scala 94:16]
  wire  abc_mshr_9_io_nestedwb_clients_1_isToN; // @[Slice.scala 94:16]
  wire  abc_mshr_9_io_tasks_sink_a_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_9_io_tasks_sink_a_valid; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_9_io_tasks_sink_a_bits_sourceId; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_9_io_tasks_sink_a_bits_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_9_io_tasks_sink_a_bits_tag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_9_io_tasks_sink_a_bits_size; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_9_io_tasks_sink_a_bits_off; // @[Slice.scala 94:16]
  wire  abc_mshr_9_io_tasks_source_bready; // @[Slice.scala 94:16]
  wire  abc_mshr_9_io_tasks_source_bvalid; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_9_io_tasks_source_bset; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_9_io_tasks_source_btag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_9_io_tasks_source_bparam; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_9_io_tasks_source_bclients; // @[Slice.scala 94:16]
  wire  abc_mshr_9_io_tasks_source_bneedData; // @[Slice.scala 94:16]
  wire  abc_mshr_9_io_tasks_sink_c_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_9_io_tasks_sink_c_valid; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_9_io_tasks_sink_c_bits_sourceId; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_9_io_tasks_sink_c_bits_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_9_io_tasks_sink_c_bits_tag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_9_io_tasks_sink_c_bits_size; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_9_io_tasks_sink_c_bits_way; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_9_io_tasks_sink_c_bits_off; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_9_io_tasks_sink_c_bits_bufIdx; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_9_io_tasks_sink_c_bits_opcode; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_9_io_tasks_sink_c_bits_param; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_9_io_tasks_sink_c_bits_source; // @[Slice.scala 94:16]
  wire  abc_mshr_9_io_tasks_sink_c_bits_save; // @[Slice.scala 94:16]
  wire  abc_mshr_9_io_tasks_sink_c_bits_drop; // @[Slice.scala 94:16]
  wire  abc_mshr_9_io_tasks_sink_c_bits_release; // @[Slice.scala 94:16]
  wire  abc_mshr_9_io_tasks_sink_c_bits_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_9_io_tasks_source_d_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_9_io_tasks_source_d_valid; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_9_io_tasks_source_d_bits_sourceId; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_9_io_tasks_source_d_bits_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_9_io_tasks_source_d_bits_tag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_9_io_tasks_source_d_bits_channel; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_9_io_tasks_source_d_bits_opcode; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_9_io_tasks_source_d_bits_param; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_9_io_tasks_source_d_bits_size; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_9_io_tasks_source_d_bits_way; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_9_io_tasks_source_d_bits_off; // @[Slice.scala 94:16]
  wire  abc_mshr_9_io_tasks_source_d_bits_useBypass; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_9_io_tasks_source_d_bits_bufIdx; // @[Slice.scala 94:16]
  wire  abc_mshr_9_io_tasks_source_d_bits_denied; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_9_io_tasks_source_d_bits_sinkId; // @[Slice.scala 94:16]
  wire  abc_mshr_9_io_tasks_source_d_bits_bypassPut; // @[Slice.scala 94:16]
  wire  abc_mshr_9_io_tasks_source_d_bits_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_9_io_tasks_source_a_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_9_io_tasks_source_a_valid; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_9_io_tasks_source_a_bits_tag; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_9_io_tasks_source_a_bits_set; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_9_io_tasks_source_a_bits_off; // @[Slice.scala 94:16]
  wire [31:0] abc_mshr_9_io_tasks_source_a_bits_mask; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_9_io_tasks_source_a_bits_opcode; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_9_io_tasks_source_a_bits_param; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_9_io_tasks_source_a_bits_source; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_9_io_tasks_source_a_bits_bufIdx; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_9_io_tasks_source_a_bits_size; // @[Slice.scala 94:16]
  wire  abc_mshr_9_io_tasks_source_a_bits_needData; // @[Slice.scala 94:16]
  wire  abc_mshr_9_io_tasks_source_a_bits_putData; // @[Slice.scala 94:16]
  wire  abc_mshr_9_io_tasks_source_c_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_9_io_tasks_source_c_valid; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_9_io_tasks_source_c_bits_opcode; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_9_io_tasks_source_c_bits_tag; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_9_io_tasks_source_c_bits_set; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_9_io_tasks_source_c_bits_param; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_9_io_tasks_source_c_bits_source; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_9_io_tasks_source_c_bits_way; // @[Slice.scala 94:16]
  wire  abc_mshr_9_io_tasks_source_c_bits_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_9_io_tasks_source_e_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_9_io_tasks_source_e_valid; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_9_io_tasks_source_e_bits_sink; // @[Slice.scala 94:16]
  wire  abc_mshr_9_io_tasks_dir_write_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_9_io_tasks_dir_write_valid; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_9_io_tasks_dir_write_bits_set; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_9_io_tasks_dir_write_bits_way; // @[Slice.scala 94:16]
  wire  abc_mshr_9_io_tasks_dir_write_bits_data_dirty; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_9_io_tasks_dir_write_bits_data_state; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_9_io_tasks_dir_write_bits_data_clientStates_0; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_9_io_tasks_dir_write_bits_data_clientStates_1; // @[Slice.scala 94:16]
  wire  abc_mshr_9_io_tasks_tag_write_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_9_io_tasks_tag_write_valid; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_9_io_tasks_tag_write_bits_set; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_9_io_tasks_tag_write_bits_way; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_9_io_tasks_tag_write_bits_tag; // @[Slice.scala 94:16]
  wire  abc_mshr_9_io_tasks_client_dir_write_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_9_io_tasks_client_dir_write_valid; // @[Slice.scala 94:16]
  wire [6:0] abc_mshr_9_io_tasks_client_dir_write_bits_set; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_9_io_tasks_client_dir_write_bits_way; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_9_io_tasks_client_dir_write_bits_data_0_state; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_9_io_tasks_client_dir_write_bits_data_1_state; // @[Slice.scala 94:16]
  wire  abc_mshr_9_io_tasks_client_tag_write_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_9_io_tasks_client_tag_write_valid; // @[Slice.scala 94:16]
  wire [6:0] abc_mshr_9_io_tasks_client_tag_write_bits_set; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_9_io_tasks_client_tag_write_bits_way; // @[Slice.scala 94:16]
  wire [22:0] abc_mshr_9_io_tasks_client_tag_write_bits_tag; // @[Slice.scala 94:16]
  wire  abc_mshr_9_io_dirResult_valid; // @[Slice.scala 94:16]
  wire  abc_mshr_9_io_dirResult_bits_self_dirty; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_9_io_dirResult_bits_self_state; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_9_io_dirResult_bits_self_clientStates_0; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_9_io_dirResult_bits_self_clientStates_1; // @[Slice.scala 94:16]
  wire  abc_mshr_9_io_dirResult_bits_self_hit; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_9_io_dirResult_bits_self_way; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_9_io_dirResult_bits_self_tag; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_9_io_dirResult_bits_clients_states_0_state; // @[Slice.scala 94:16]
  wire  abc_mshr_9_io_dirResult_bits_clients_states_0_hit; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_9_io_dirResult_bits_clients_states_1_state; // @[Slice.scala 94:16]
  wire  abc_mshr_9_io_dirResult_bits_clients_states_1_hit; // @[Slice.scala 94:16]
  wire [22:0] abc_mshr_9_io_dirResult_bits_clients_tag; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_9_io_dirResult_bits_clients_way; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_9_io_c_status_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_9_io_c_status_tag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_9_io_c_status_way; // @[Slice.scala 94:16]
  wire  abc_mshr_9_io_c_status_nestedReleaseData; // @[Slice.scala 94:16]
  wire  abc_mshr_9_io_c_status_releaseThrough; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_9_io_bstatus_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_9_io_bstatus_tag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_9_io_bstatus_way; // @[Slice.scala 94:16]
  wire  abc_mshr_9_io_bstatus_nestedProbeAckData; // @[Slice.scala 94:16]
  wire  abc_mshr_9_io_bstatus_probeHelperFinish; // @[Slice.scala 94:16]
  wire  abc_mshr_9_io_bstatus_probeAckDataThrough; // @[Slice.scala 94:16]
  wire  abc_mshr_9_io_releaseThrough; // @[Slice.scala 94:16]
  wire  abc_mshr_9_io_probeAckDataThrough; // @[Slice.scala 94:16]
  wire  abc_mshr_9_io_is_nestedReleaseData; // @[Slice.scala 94:16]
  wire  abc_mshr_9_io_is_nestedProbeAckData; // @[Slice.scala 94:16]
  wire  abc_mshr_9_io_probeHelperFinish; // @[Slice.scala 94:16]
  wire  abc_mshr_10_clock; // @[Slice.scala 94:16]
  wire  abc_mshr_10_reset; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_10_io_id; // @[Slice.scala 94:16]
  wire  abc_mshr_10_io_enable; // @[Slice.scala 94:16]
  wire  abc_mshr_10_io_alloc_valid; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_10_io_alloc_bits_channel; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_10_io_alloc_bits_opcode; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_10_io_alloc_bits_param; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_10_io_alloc_bits_size; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_10_io_alloc_bits_source; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_10_io_alloc_bits_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_10_io_alloc_bits_tag; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_10_io_alloc_bits_off; // @[Slice.scala 94:16]
  wire [31:0] abc_mshr_10_io_alloc_bits_mask; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_10_io_alloc_bits_bufIdx; // @[Slice.scala 94:16]
  wire  abc_mshr_10_io_alloc_bits_preferCache; // @[Slice.scala 94:16]
  wire  abc_mshr_10_io_alloc_bits_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_10_io_alloc_bits_fromProbeHelper; // @[Slice.scala 94:16]
  wire  abc_mshr_10_io_alloc_bits_fromCmoHelper; // @[Slice.scala 94:16]
  wire  abc_mshr_10_io_alloc_bits_needProbeAckData; // @[Slice.scala 94:16]
  wire  abc_mshr_10_io_status_valid; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_10_io_status_bits_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_10_io_status_bits_tag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_10_io_status_bits_way; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_10_io_status_bits_way_reg; // @[Slice.scala 94:16]
  wire  abc_mshr_10_io_status_bits_nestB; // @[Slice.scala 94:16]
  wire  abc_mshr_10_io_status_bits_nestC; // @[Slice.scala 94:16]
  wire  abc_mshr_10_io_status_bits_will_grant_data; // @[Slice.scala 94:16]
  wire  abc_mshr_10_io_status_bits_will_save_data; // @[Slice.scala 94:16]
  wire  abc_mshr_10_io_status_bits_will_free; // @[Slice.scala 94:16]
  wire  abc_mshr_10_io_resps_sink_c_valid; // @[Slice.scala 94:16]
  wire  abc_mshr_10_io_resps_sink_c_bits_hasData; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_10_io_resps_sink_c_bits_param; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_10_io_resps_sink_c_bits_source; // @[Slice.scala 94:16]
  wire  abc_mshr_10_io_resps_sink_c_bits_last; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_10_io_resps_sink_c_bits_bufIdx; // @[Slice.scala 94:16]
  wire  abc_mshr_10_io_resps_sink_d_valid; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_10_io_resps_sink_d_bits_opcode; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_10_io_resps_sink_d_bits_param; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_10_io_resps_sink_d_bits_sink; // @[Slice.scala 94:16]
  wire  abc_mshr_10_io_resps_sink_d_bits_last; // @[Slice.scala 94:16]
  wire  abc_mshr_10_io_resps_sink_d_bits_denied; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_10_io_resps_sink_d_bits_bufIdx; // @[Slice.scala 94:16]
  wire  abc_mshr_10_io_resps_sink_e_valid; // @[Slice.scala 94:16]
  wire  abc_mshr_10_io_resps_source_d_valid; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_10_io_nestedwb_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_10_io_nestedwb_tag; // @[Slice.scala 94:16]
  wire  abc_mshr_10_io_nestedwb_btoN; // @[Slice.scala 94:16]
  wire  abc_mshr_10_io_nestedwb_btoB; // @[Slice.scala 94:16]
  wire  abc_mshr_10_io_nestedwb_bclr_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_10_io_nestedwb_bset_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_10_io_nestedwb_c_set_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_10_io_nestedwb_c_set_hit; // @[Slice.scala 94:16]
  wire  abc_mshr_10_io_nestedwb_clients_0_isToN; // @[Slice.scala 94:16]
  wire  abc_mshr_10_io_nestedwb_clients_1_isToN; // @[Slice.scala 94:16]
  wire  abc_mshr_10_io_tasks_sink_a_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_10_io_tasks_sink_a_valid; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_10_io_tasks_sink_a_bits_sourceId; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_10_io_tasks_sink_a_bits_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_10_io_tasks_sink_a_bits_tag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_10_io_tasks_sink_a_bits_size; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_10_io_tasks_sink_a_bits_off; // @[Slice.scala 94:16]
  wire  abc_mshr_10_io_tasks_source_bready; // @[Slice.scala 94:16]
  wire  abc_mshr_10_io_tasks_source_bvalid; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_10_io_tasks_source_bset; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_10_io_tasks_source_btag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_10_io_tasks_source_bparam; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_10_io_tasks_source_bclients; // @[Slice.scala 94:16]
  wire  abc_mshr_10_io_tasks_source_bneedData; // @[Slice.scala 94:16]
  wire  abc_mshr_10_io_tasks_sink_c_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_10_io_tasks_sink_c_valid; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_10_io_tasks_sink_c_bits_sourceId; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_10_io_tasks_sink_c_bits_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_10_io_tasks_sink_c_bits_tag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_10_io_tasks_sink_c_bits_size; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_10_io_tasks_sink_c_bits_way; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_10_io_tasks_sink_c_bits_off; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_10_io_tasks_sink_c_bits_bufIdx; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_10_io_tasks_sink_c_bits_opcode; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_10_io_tasks_sink_c_bits_param; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_10_io_tasks_sink_c_bits_source; // @[Slice.scala 94:16]
  wire  abc_mshr_10_io_tasks_sink_c_bits_save; // @[Slice.scala 94:16]
  wire  abc_mshr_10_io_tasks_sink_c_bits_drop; // @[Slice.scala 94:16]
  wire  abc_mshr_10_io_tasks_sink_c_bits_release; // @[Slice.scala 94:16]
  wire  abc_mshr_10_io_tasks_sink_c_bits_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_10_io_tasks_source_d_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_10_io_tasks_source_d_valid; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_10_io_tasks_source_d_bits_sourceId; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_10_io_tasks_source_d_bits_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_10_io_tasks_source_d_bits_tag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_10_io_tasks_source_d_bits_channel; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_10_io_tasks_source_d_bits_opcode; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_10_io_tasks_source_d_bits_param; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_10_io_tasks_source_d_bits_size; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_10_io_tasks_source_d_bits_way; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_10_io_tasks_source_d_bits_off; // @[Slice.scala 94:16]
  wire  abc_mshr_10_io_tasks_source_d_bits_useBypass; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_10_io_tasks_source_d_bits_bufIdx; // @[Slice.scala 94:16]
  wire  abc_mshr_10_io_tasks_source_d_bits_denied; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_10_io_tasks_source_d_bits_sinkId; // @[Slice.scala 94:16]
  wire  abc_mshr_10_io_tasks_source_d_bits_bypassPut; // @[Slice.scala 94:16]
  wire  abc_mshr_10_io_tasks_source_d_bits_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_10_io_tasks_source_a_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_10_io_tasks_source_a_valid; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_10_io_tasks_source_a_bits_tag; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_10_io_tasks_source_a_bits_set; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_10_io_tasks_source_a_bits_off; // @[Slice.scala 94:16]
  wire [31:0] abc_mshr_10_io_tasks_source_a_bits_mask; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_10_io_tasks_source_a_bits_opcode; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_10_io_tasks_source_a_bits_param; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_10_io_tasks_source_a_bits_source; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_10_io_tasks_source_a_bits_bufIdx; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_10_io_tasks_source_a_bits_size; // @[Slice.scala 94:16]
  wire  abc_mshr_10_io_tasks_source_a_bits_needData; // @[Slice.scala 94:16]
  wire  abc_mshr_10_io_tasks_source_a_bits_putData; // @[Slice.scala 94:16]
  wire  abc_mshr_10_io_tasks_source_c_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_10_io_tasks_source_c_valid; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_10_io_tasks_source_c_bits_opcode; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_10_io_tasks_source_c_bits_tag; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_10_io_tasks_source_c_bits_set; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_10_io_tasks_source_c_bits_param; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_10_io_tasks_source_c_bits_source; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_10_io_tasks_source_c_bits_way; // @[Slice.scala 94:16]
  wire  abc_mshr_10_io_tasks_source_c_bits_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_10_io_tasks_source_e_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_10_io_tasks_source_e_valid; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_10_io_tasks_source_e_bits_sink; // @[Slice.scala 94:16]
  wire  abc_mshr_10_io_tasks_dir_write_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_10_io_tasks_dir_write_valid; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_10_io_tasks_dir_write_bits_set; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_10_io_tasks_dir_write_bits_way; // @[Slice.scala 94:16]
  wire  abc_mshr_10_io_tasks_dir_write_bits_data_dirty; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_10_io_tasks_dir_write_bits_data_state; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_10_io_tasks_dir_write_bits_data_clientStates_0; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_10_io_tasks_dir_write_bits_data_clientStates_1; // @[Slice.scala 94:16]
  wire  abc_mshr_10_io_tasks_tag_write_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_10_io_tasks_tag_write_valid; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_10_io_tasks_tag_write_bits_set; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_10_io_tasks_tag_write_bits_way; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_10_io_tasks_tag_write_bits_tag; // @[Slice.scala 94:16]
  wire  abc_mshr_10_io_tasks_client_dir_write_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_10_io_tasks_client_dir_write_valid; // @[Slice.scala 94:16]
  wire [6:0] abc_mshr_10_io_tasks_client_dir_write_bits_set; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_10_io_tasks_client_dir_write_bits_way; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_10_io_tasks_client_dir_write_bits_data_0_state; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_10_io_tasks_client_dir_write_bits_data_1_state; // @[Slice.scala 94:16]
  wire  abc_mshr_10_io_tasks_client_tag_write_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_10_io_tasks_client_tag_write_valid; // @[Slice.scala 94:16]
  wire [6:0] abc_mshr_10_io_tasks_client_tag_write_bits_set; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_10_io_tasks_client_tag_write_bits_way; // @[Slice.scala 94:16]
  wire [22:0] abc_mshr_10_io_tasks_client_tag_write_bits_tag; // @[Slice.scala 94:16]
  wire  abc_mshr_10_io_dirResult_valid; // @[Slice.scala 94:16]
  wire  abc_mshr_10_io_dirResult_bits_self_dirty; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_10_io_dirResult_bits_self_state; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_10_io_dirResult_bits_self_clientStates_0; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_10_io_dirResult_bits_self_clientStates_1; // @[Slice.scala 94:16]
  wire  abc_mshr_10_io_dirResult_bits_self_hit; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_10_io_dirResult_bits_self_way; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_10_io_dirResult_bits_self_tag; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_10_io_dirResult_bits_clients_states_0_state; // @[Slice.scala 94:16]
  wire  abc_mshr_10_io_dirResult_bits_clients_states_0_hit; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_10_io_dirResult_bits_clients_states_1_state; // @[Slice.scala 94:16]
  wire  abc_mshr_10_io_dirResult_bits_clients_states_1_hit; // @[Slice.scala 94:16]
  wire [22:0] abc_mshr_10_io_dirResult_bits_clients_tag; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_10_io_dirResult_bits_clients_way; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_10_io_c_status_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_10_io_c_status_tag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_10_io_c_status_way; // @[Slice.scala 94:16]
  wire  abc_mshr_10_io_c_status_nestedReleaseData; // @[Slice.scala 94:16]
  wire  abc_mshr_10_io_c_status_releaseThrough; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_10_io_bstatus_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_10_io_bstatus_tag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_10_io_bstatus_way; // @[Slice.scala 94:16]
  wire  abc_mshr_10_io_bstatus_nestedProbeAckData; // @[Slice.scala 94:16]
  wire  abc_mshr_10_io_bstatus_probeHelperFinish; // @[Slice.scala 94:16]
  wire  abc_mshr_10_io_bstatus_probeAckDataThrough; // @[Slice.scala 94:16]
  wire  abc_mshr_10_io_releaseThrough; // @[Slice.scala 94:16]
  wire  abc_mshr_10_io_probeAckDataThrough; // @[Slice.scala 94:16]
  wire  abc_mshr_10_io_is_nestedReleaseData; // @[Slice.scala 94:16]
  wire  abc_mshr_10_io_is_nestedProbeAckData; // @[Slice.scala 94:16]
  wire  abc_mshr_10_io_probeHelperFinish; // @[Slice.scala 94:16]
  wire  abc_mshr_11_clock; // @[Slice.scala 94:16]
  wire  abc_mshr_11_reset; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_11_io_id; // @[Slice.scala 94:16]
  wire  abc_mshr_11_io_enable; // @[Slice.scala 94:16]
  wire  abc_mshr_11_io_alloc_valid; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_11_io_alloc_bits_channel; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_11_io_alloc_bits_opcode; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_11_io_alloc_bits_param; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_11_io_alloc_bits_size; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_11_io_alloc_bits_source; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_11_io_alloc_bits_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_11_io_alloc_bits_tag; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_11_io_alloc_bits_off; // @[Slice.scala 94:16]
  wire [31:0] abc_mshr_11_io_alloc_bits_mask; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_11_io_alloc_bits_bufIdx; // @[Slice.scala 94:16]
  wire  abc_mshr_11_io_alloc_bits_preferCache; // @[Slice.scala 94:16]
  wire  abc_mshr_11_io_alloc_bits_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_11_io_alloc_bits_fromProbeHelper; // @[Slice.scala 94:16]
  wire  abc_mshr_11_io_alloc_bits_fromCmoHelper; // @[Slice.scala 94:16]
  wire  abc_mshr_11_io_alloc_bits_needProbeAckData; // @[Slice.scala 94:16]
  wire  abc_mshr_11_io_status_valid; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_11_io_status_bits_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_11_io_status_bits_tag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_11_io_status_bits_way; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_11_io_status_bits_way_reg; // @[Slice.scala 94:16]
  wire  abc_mshr_11_io_status_bits_nestB; // @[Slice.scala 94:16]
  wire  abc_mshr_11_io_status_bits_nestC; // @[Slice.scala 94:16]
  wire  abc_mshr_11_io_status_bits_will_grant_data; // @[Slice.scala 94:16]
  wire  abc_mshr_11_io_status_bits_will_save_data; // @[Slice.scala 94:16]
  wire  abc_mshr_11_io_status_bits_will_free; // @[Slice.scala 94:16]
  wire  abc_mshr_11_io_resps_sink_c_valid; // @[Slice.scala 94:16]
  wire  abc_mshr_11_io_resps_sink_c_bits_hasData; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_11_io_resps_sink_c_bits_param; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_11_io_resps_sink_c_bits_source; // @[Slice.scala 94:16]
  wire  abc_mshr_11_io_resps_sink_c_bits_last; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_11_io_resps_sink_c_bits_bufIdx; // @[Slice.scala 94:16]
  wire  abc_mshr_11_io_resps_sink_d_valid; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_11_io_resps_sink_d_bits_opcode; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_11_io_resps_sink_d_bits_param; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_11_io_resps_sink_d_bits_sink; // @[Slice.scala 94:16]
  wire  abc_mshr_11_io_resps_sink_d_bits_last; // @[Slice.scala 94:16]
  wire  abc_mshr_11_io_resps_sink_d_bits_denied; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_11_io_resps_sink_d_bits_bufIdx; // @[Slice.scala 94:16]
  wire  abc_mshr_11_io_resps_sink_e_valid; // @[Slice.scala 94:16]
  wire  abc_mshr_11_io_resps_source_d_valid; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_11_io_nestedwb_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_11_io_nestedwb_tag; // @[Slice.scala 94:16]
  wire  abc_mshr_11_io_nestedwb_btoN; // @[Slice.scala 94:16]
  wire  abc_mshr_11_io_nestedwb_btoB; // @[Slice.scala 94:16]
  wire  abc_mshr_11_io_nestedwb_bclr_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_11_io_nestedwb_bset_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_11_io_nestedwb_c_set_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_11_io_nestedwb_c_set_hit; // @[Slice.scala 94:16]
  wire  abc_mshr_11_io_nestedwb_clients_0_isToN; // @[Slice.scala 94:16]
  wire  abc_mshr_11_io_nestedwb_clients_1_isToN; // @[Slice.scala 94:16]
  wire  abc_mshr_11_io_tasks_sink_a_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_11_io_tasks_sink_a_valid; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_11_io_tasks_sink_a_bits_sourceId; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_11_io_tasks_sink_a_bits_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_11_io_tasks_sink_a_bits_tag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_11_io_tasks_sink_a_bits_size; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_11_io_tasks_sink_a_bits_off; // @[Slice.scala 94:16]
  wire  abc_mshr_11_io_tasks_source_bready; // @[Slice.scala 94:16]
  wire  abc_mshr_11_io_tasks_source_bvalid; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_11_io_tasks_source_bset; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_11_io_tasks_source_btag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_11_io_tasks_source_bparam; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_11_io_tasks_source_bclients; // @[Slice.scala 94:16]
  wire  abc_mshr_11_io_tasks_source_bneedData; // @[Slice.scala 94:16]
  wire  abc_mshr_11_io_tasks_sink_c_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_11_io_tasks_sink_c_valid; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_11_io_tasks_sink_c_bits_sourceId; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_11_io_tasks_sink_c_bits_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_11_io_tasks_sink_c_bits_tag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_11_io_tasks_sink_c_bits_size; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_11_io_tasks_sink_c_bits_way; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_11_io_tasks_sink_c_bits_off; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_11_io_tasks_sink_c_bits_bufIdx; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_11_io_tasks_sink_c_bits_opcode; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_11_io_tasks_sink_c_bits_param; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_11_io_tasks_sink_c_bits_source; // @[Slice.scala 94:16]
  wire  abc_mshr_11_io_tasks_sink_c_bits_save; // @[Slice.scala 94:16]
  wire  abc_mshr_11_io_tasks_sink_c_bits_drop; // @[Slice.scala 94:16]
  wire  abc_mshr_11_io_tasks_sink_c_bits_release; // @[Slice.scala 94:16]
  wire  abc_mshr_11_io_tasks_sink_c_bits_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_11_io_tasks_source_d_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_11_io_tasks_source_d_valid; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_11_io_tasks_source_d_bits_sourceId; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_11_io_tasks_source_d_bits_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_11_io_tasks_source_d_bits_tag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_11_io_tasks_source_d_bits_channel; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_11_io_tasks_source_d_bits_opcode; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_11_io_tasks_source_d_bits_param; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_11_io_tasks_source_d_bits_size; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_11_io_tasks_source_d_bits_way; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_11_io_tasks_source_d_bits_off; // @[Slice.scala 94:16]
  wire  abc_mshr_11_io_tasks_source_d_bits_useBypass; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_11_io_tasks_source_d_bits_bufIdx; // @[Slice.scala 94:16]
  wire  abc_mshr_11_io_tasks_source_d_bits_denied; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_11_io_tasks_source_d_bits_sinkId; // @[Slice.scala 94:16]
  wire  abc_mshr_11_io_tasks_source_d_bits_bypassPut; // @[Slice.scala 94:16]
  wire  abc_mshr_11_io_tasks_source_d_bits_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_11_io_tasks_source_a_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_11_io_tasks_source_a_valid; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_11_io_tasks_source_a_bits_tag; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_11_io_tasks_source_a_bits_set; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_11_io_tasks_source_a_bits_off; // @[Slice.scala 94:16]
  wire [31:0] abc_mshr_11_io_tasks_source_a_bits_mask; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_11_io_tasks_source_a_bits_opcode; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_11_io_tasks_source_a_bits_param; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_11_io_tasks_source_a_bits_source; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_11_io_tasks_source_a_bits_bufIdx; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_11_io_tasks_source_a_bits_size; // @[Slice.scala 94:16]
  wire  abc_mshr_11_io_tasks_source_a_bits_needData; // @[Slice.scala 94:16]
  wire  abc_mshr_11_io_tasks_source_a_bits_putData; // @[Slice.scala 94:16]
  wire  abc_mshr_11_io_tasks_source_c_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_11_io_tasks_source_c_valid; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_11_io_tasks_source_c_bits_opcode; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_11_io_tasks_source_c_bits_tag; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_11_io_tasks_source_c_bits_set; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_11_io_tasks_source_c_bits_param; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_11_io_tasks_source_c_bits_source; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_11_io_tasks_source_c_bits_way; // @[Slice.scala 94:16]
  wire  abc_mshr_11_io_tasks_source_c_bits_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_11_io_tasks_source_e_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_11_io_tasks_source_e_valid; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_11_io_tasks_source_e_bits_sink; // @[Slice.scala 94:16]
  wire  abc_mshr_11_io_tasks_dir_write_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_11_io_tasks_dir_write_valid; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_11_io_tasks_dir_write_bits_set; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_11_io_tasks_dir_write_bits_way; // @[Slice.scala 94:16]
  wire  abc_mshr_11_io_tasks_dir_write_bits_data_dirty; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_11_io_tasks_dir_write_bits_data_state; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_11_io_tasks_dir_write_bits_data_clientStates_0; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_11_io_tasks_dir_write_bits_data_clientStates_1; // @[Slice.scala 94:16]
  wire  abc_mshr_11_io_tasks_tag_write_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_11_io_tasks_tag_write_valid; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_11_io_tasks_tag_write_bits_set; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_11_io_tasks_tag_write_bits_way; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_11_io_tasks_tag_write_bits_tag; // @[Slice.scala 94:16]
  wire  abc_mshr_11_io_tasks_client_dir_write_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_11_io_tasks_client_dir_write_valid; // @[Slice.scala 94:16]
  wire [6:0] abc_mshr_11_io_tasks_client_dir_write_bits_set; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_11_io_tasks_client_dir_write_bits_way; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_11_io_tasks_client_dir_write_bits_data_0_state; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_11_io_tasks_client_dir_write_bits_data_1_state; // @[Slice.scala 94:16]
  wire  abc_mshr_11_io_tasks_client_tag_write_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_11_io_tasks_client_tag_write_valid; // @[Slice.scala 94:16]
  wire [6:0] abc_mshr_11_io_tasks_client_tag_write_bits_set; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_11_io_tasks_client_tag_write_bits_way; // @[Slice.scala 94:16]
  wire [22:0] abc_mshr_11_io_tasks_client_tag_write_bits_tag; // @[Slice.scala 94:16]
  wire  abc_mshr_11_io_dirResult_valid; // @[Slice.scala 94:16]
  wire  abc_mshr_11_io_dirResult_bits_self_dirty; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_11_io_dirResult_bits_self_state; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_11_io_dirResult_bits_self_clientStates_0; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_11_io_dirResult_bits_self_clientStates_1; // @[Slice.scala 94:16]
  wire  abc_mshr_11_io_dirResult_bits_self_hit; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_11_io_dirResult_bits_self_way; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_11_io_dirResult_bits_self_tag; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_11_io_dirResult_bits_clients_states_0_state; // @[Slice.scala 94:16]
  wire  abc_mshr_11_io_dirResult_bits_clients_states_0_hit; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_11_io_dirResult_bits_clients_states_1_state; // @[Slice.scala 94:16]
  wire  abc_mshr_11_io_dirResult_bits_clients_states_1_hit; // @[Slice.scala 94:16]
  wire [22:0] abc_mshr_11_io_dirResult_bits_clients_tag; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_11_io_dirResult_bits_clients_way; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_11_io_c_status_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_11_io_c_status_tag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_11_io_c_status_way; // @[Slice.scala 94:16]
  wire  abc_mshr_11_io_c_status_nestedReleaseData; // @[Slice.scala 94:16]
  wire  abc_mshr_11_io_c_status_releaseThrough; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_11_io_bstatus_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_11_io_bstatus_tag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_11_io_bstatus_way; // @[Slice.scala 94:16]
  wire  abc_mshr_11_io_bstatus_nestedProbeAckData; // @[Slice.scala 94:16]
  wire  abc_mshr_11_io_bstatus_probeHelperFinish; // @[Slice.scala 94:16]
  wire  abc_mshr_11_io_bstatus_probeAckDataThrough; // @[Slice.scala 94:16]
  wire  abc_mshr_11_io_releaseThrough; // @[Slice.scala 94:16]
  wire  abc_mshr_11_io_probeAckDataThrough; // @[Slice.scala 94:16]
  wire  abc_mshr_11_io_is_nestedReleaseData; // @[Slice.scala 94:16]
  wire  abc_mshr_11_io_is_nestedProbeAckData; // @[Slice.scala 94:16]
  wire  abc_mshr_11_io_probeHelperFinish; // @[Slice.scala 94:16]
  wire  abc_mshr_12_clock; // @[Slice.scala 94:16]
  wire  abc_mshr_12_reset; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_12_io_id; // @[Slice.scala 94:16]
  wire  abc_mshr_12_io_enable; // @[Slice.scala 94:16]
  wire  abc_mshr_12_io_alloc_valid; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_12_io_alloc_bits_channel; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_12_io_alloc_bits_opcode; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_12_io_alloc_bits_param; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_12_io_alloc_bits_size; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_12_io_alloc_bits_source; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_12_io_alloc_bits_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_12_io_alloc_bits_tag; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_12_io_alloc_bits_off; // @[Slice.scala 94:16]
  wire [31:0] abc_mshr_12_io_alloc_bits_mask; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_12_io_alloc_bits_bufIdx; // @[Slice.scala 94:16]
  wire  abc_mshr_12_io_alloc_bits_preferCache; // @[Slice.scala 94:16]
  wire  abc_mshr_12_io_alloc_bits_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_12_io_alloc_bits_fromProbeHelper; // @[Slice.scala 94:16]
  wire  abc_mshr_12_io_alloc_bits_fromCmoHelper; // @[Slice.scala 94:16]
  wire  abc_mshr_12_io_alloc_bits_needProbeAckData; // @[Slice.scala 94:16]
  wire  abc_mshr_12_io_status_valid; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_12_io_status_bits_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_12_io_status_bits_tag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_12_io_status_bits_way; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_12_io_status_bits_way_reg; // @[Slice.scala 94:16]
  wire  abc_mshr_12_io_status_bits_nestB; // @[Slice.scala 94:16]
  wire  abc_mshr_12_io_status_bits_nestC; // @[Slice.scala 94:16]
  wire  abc_mshr_12_io_status_bits_will_grant_data; // @[Slice.scala 94:16]
  wire  abc_mshr_12_io_status_bits_will_save_data; // @[Slice.scala 94:16]
  wire  abc_mshr_12_io_status_bits_will_free; // @[Slice.scala 94:16]
  wire  abc_mshr_12_io_resps_sink_c_valid; // @[Slice.scala 94:16]
  wire  abc_mshr_12_io_resps_sink_c_bits_hasData; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_12_io_resps_sink_c_bits_param; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_12_io_resps_sink_c_bits_source; // @[Slice.scala 94:16]
  wire  abc_mshr_12_io_resps_sink_c_bits_last; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_12_io_resps_sink_c_bits_bufIdx; // @[Slice.scala 94:16]
  wire  abc_mshr_12_io_resps_sink_d_valid; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_12_io_resps_sink_d_bits_opcode; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_12_io_resps_sink_d_bits_param; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_12_io_resps_sink_d_bits_sink; // @[Slice.scala 94:16]
  wire  abc_mshr_12_io_resps_sink_d_bits_last; // @[Slice.scala 94:16]
  wire  abc_mshr_12_io_resps_sink_d_bits_denied; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_12_io_resps_sink_d_bits_bufIdx; // @[Slice.scala 94:16]
  wire  abc_mshr_12_io_resps_sink_e_valid; // @[Slice.scala 94:16]
  wire  abc_mshr_12_io_resps_source_d_valid; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_12_io_nestedwb_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_12_io_nestedwb_tag; // @[Slice.scala 94:16]
  wire  abc_mshr_12_io_nestedwb_btoN; // @[Slice.scala 94:16]
  wire  abc_mshr_12_io_nestedwb_btoB; // @[Slice.scala 94:16]
  wire  abc_mshr_12_io_nestedwb_bclr_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_12_io_nestedwb_bset_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_12_io_nestedwb_c_set_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_12_io_nestedwb_c_set_hit; // @[Slice.scala 94:16]
  wire  abc_mshr_12_io_nestedwb_clients_0_isToN; // @[Slice.scala 94:16]
  wire  abc_mshr_12_io_nestedwb_clients_1_isToN; // @[Slice.scala 94:16]
  wire  abc_mshr_12_io_tasks_sink_a_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_12_io_tasks_sink_a_valid; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_12_io_tasks_sink_a_bits_sourceId; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_12_io_tasks_sink_a_bits_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_12_io_tasks_sink_a_bits_tag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_12_io_tasks_sink_a_bits_size; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_12_io_tasks_sink_a_bits_off; // @[Slice.scala 94:16]
  wire  abc_mshr_12_io_tasks_source_bready; // @[Slice.scala 94:16]
  wire  abc_mshr_12_io_tasks_source_bvalid; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_12_io_tasks_source_bset; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_12_io_tasks_source_btag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_12_io_tasks_source_bparam; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_12_io_tasks_source_bclients; // @[Slice.scala 94:16]
  wire  abc_mshr_12_io_tasks_source_bneedData; // @[Slice.scala 94:16]
  wire  abc_mshr_12_io_tasks_sink_c_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_12_io_tasks_sink_c_valid; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_12_io_tasks_sink_c_bits_sourceId; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_12_io_tasks_sink_c_bits_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_12_io_tasks_sink_c_bits_tag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_12_io_tasks_sink_c_bits_size; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_12_io_tasks_sink_c_bits_way; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_12_io_tasks_sink_c_bits_off; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_12_io_tasks_sink_c_bits_bufIdx; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_12_io_tasks_sink_c_bits_opcode; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_12_io_tasks_sink_c_bits_param; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_12_io_tasks_sink_c_bits_source; // @[Slice.scala 94:16]
  wire  abc_mshr_12_io_tasks_sink_c_bits_save; // @[Slice.scala 94:16]
  wire  abc_mshr_12_io_tasks_sink_c_bits_drop; // @[Slice.scala 94:16]
  wire  abc_mshr_12_io_tasks_sink_c_bits_release; // @[Slice.scala 94:16]
  wire  abc_mshr_12_io_tasks_sink_c_bits_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_12_io_tasks_source_d_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_12_io_tasks_source_d_valid; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_12_io_tasks_source_d_bits_sourceId; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_12_io_tasks_source_d_bits_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_12_io_tasks_source_d_bits_tag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_12_io_tasks_source_d_bits_channel; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_12_io_tasks_source_d_bits_opcode; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_12_io_tasks_source_d_bits_param; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_12_io_tasks_source_d_bits_size; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_12_io_tasks_source_d_bits_way; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_12_io_tasks_source_d_bits_off; // @[Slice.scala 94:16]
  wire  abc_mshr_12_io_tasks_source_d_bits_useBypass; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_12_io_tasks_source_d_bits_bufIdx; // @[Slice.scala 94:16]
  wire  abc_mshr_12_io_tasks_source_d_bits_denied; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_12_io_tasks_source_d_bits_sinkId; // @[Slice.scala 94:16]
  wire  abc_mshr_12_io_tasks_source_d_bits_bypassPut; // @[Slice.scala 94:16]
  wire  abc_mshr_12_io_tasks_source_d_bits_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_12_io_tasks_source_a_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_12_io_tasks_source_a_valid; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_12_io_tasks_source_a_bits_tag; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_12_io_tasks_source_a_bits_set; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_12_io_tasks_source_a_bits_off; // @[Slice.scala 94:16]
  wire [31:0] abc_mshr_12_io_tasks_source_a_bits_mask; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_12_io_tasks_source_a_bits_opcode; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_12_io_tasks_source_a_bits_param; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_12_io_tasks_source_a_bits_source; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_12_io_tasks_source_a_bits_bufIdx; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_12_io_tasks_source_a_bits_size; // @[Slice.scala 94:16]
  wire  abc_mshr_12_io_tasks_source_a_bits_needData; // @[Slice.scala 94:16]
  wire  abc_mshr_12_io_tasks_source_a_bits_putData; // @[Slice.scala 94:16]
  wire  abc_mshr_12_io_tasks_source_c_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_12_io_tasks_source_c_valid; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_12_io_tasks_source_c_bits_opcode; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_12_io_tasks_source_c_bits_tag; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_12_io_tasks_source_c_bits_set; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_12_io_tasks_source_c_bits_param; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_12_io_tasks_source_c_bits_source; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_12_io_tasks_source_c_bits_way; // @[Slice.scala 94:16]
  wire  abc_mshr_12_io_tasks_source_c_bits_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_12_io_tasks_source_e_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_12_io_tasks_source_e_valid; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_12_io_tasks_source_e_bits_sink; // @[Slice.scala 94:16]
  wire  abc_mshr_12_io_tasks_dir_write_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_12_io_tasks_dir_write_valid; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_12_io_tasks_dir_write_bits_set; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_12_io_tasks_dir_write_bits_way; // @[Slice.scala 94:16]
  wire  abc_mshr_12_io_tasks_dir_write_bits_data_dirty; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_12_io_tasks_dir_write_bits_data_state; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_12_io_tasks_dir_write_bits_data_clientStates_0; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_12_io_tasks_dir_write_bits_data_clientStates_1; // @[Slice.scala 94:16]
  wire  abc_mshr_12_io_tasks_tag_write_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_12_io_tasks_tag_write_valid; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_12_io_tasks_tag_write_bits_set; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_12_io_tasks_tag_write_bits_way; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_12_io_tasks_tag_write_bits_tag; // @[Slice.scala 94:16]
  wire  abc_mshr_12_io_tasks_client_dir_write_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_12_io_tasks_client_dir_write_valid; // @[Slice.scala 94:16]
  wire [6:0] abc_mshr_12_io_tasks_client_dir_write_bits_set; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_12_io_tasks_client_dir_write_bits_way; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_12_io_tasks_client_dir_write_bits_data_0_state; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_12_io_tasks_client_dir_write_bits_data_1_state; // @[Slice.scala 94:16]
  wire  abc_mshr_12_io_tasks_client_tag_write_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_12_io_tasks_client_tag_write_valid; // @[Slice.scala 94:16]
  wire [6:0] abc_mshr_12_io_tasks_client_tag_write_bits_set; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_12_io_tasks_client_tag_write_bits_way; // @[Slice.scala 94:16]
  wire [22:0] abc_mshr_12_io_tasks_client_tag_write_bits_tag; // @[Slice.scala 94:16]
  wire  abc_mshr_12_io_dirResult_valid; // @[Slice.scala 94:16]
  wire  abc_mshr_12_io_dirResult_bits_self_dirty; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_12_io_dirResult_bits_self_state; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_12_io_dirResult_bits_self_clientStates_0; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_12_io_dirResult_bits_self_clientStates_1; // @[Slice.scala 94:16]
  wire  abc_mshr_12_io_dirResult_bits_self_hit; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_12_io_dirResult_bits_self_way; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_12_io_dirResult_bits_self_tag; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_12_io_dirResult_bits_clients_states_0_state; // @[Slice.scala 94:16]
  wire  abc_mshr_12_io_dirResult_bits_clients_states_0_hit; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_12_io_dirResult_bits_clients_states_1_state; // @[Slice.scala 94:16]
  wire  abc_mshr_12_io_dirResult_bits_clients_states_1_hit; // @[Slice.scala 94:16]
  wire [22:0] abc_mshr_12_io_dirResult_bits_clients_tag; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_12_io_dirResult_bits_clients_way; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_12_io_c_status_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_12_io_c_status_tag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_12_io_c_status_way; // @[Slice.scala 94:16]
  wire  abc_mshr_12_io_c_status_nestedReleaseData; // @[Slice.scala 94:16]
  wire  abc_mshr_12_io_c_status_releaseThrough; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_12_io_bstatus_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_12_io_bstatus_tag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_12_io_bstatus_way; // @[Slice.scala 94:16]
  wire  abc_mshr_12_io_bstatus_nestedProbeAckData; // @[Slice.scala 94:16]
  wire  abc_mshr_12_io_bstatus_probeHelperFinish; // @[Slice.scala 94:16]
  wire  abc_mshr_12_io_bstatus_probeAckDataThrough; // @[Slice.scala 94:16]
  wire  abc_mshr_12_io_releaseThrough; // @[Slice.scala 94:16]
  wire  abc_mshr_12_io_probeAckDataThrough; // @[Slice.scala 94:16]
  wire  abc_mshr_12_io_is_nestedReleaseData; // @[Slice.scala 94:16]
  wire  abc_mshr_12_io_is_nestedProbeAckData; // @[Slice.scala 94:16]
  wire  abc_mshr_12_io_probeHelperFinish; // @[Slice.scala 94:16]
  wire  abc_mshr_13_clock; // @[Slice.scala 94:16]
  wire  abc_mshr_13_reset; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_13_io_id; // @[Slice.scala 94:16]
  wire  abc_mshr_13_io_enable; // @[Slice.scala 94:16]
  wire  abc_mshr_13_io_alloc_valid; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_13_io_alloc_bits_channel; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_13_io_alloc_bits_opcode; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_13_io_alloc_bits_param; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_13_io_alloc_bits_size; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_13_io_alloc_bits_source; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_13_io_alloc_bits_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_13_io_alloc_bits_tag; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_13_io_alloc_bits_off; // @[Slice.scala 94:16]
  wire [31:0] abc_mshr_13_io_alloc_bits_mask; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_13_io_alloc_bits_bufIdx; // @[Slice.scala 94:16]
  wire  abc_mshr_13_io_alloc_bits_preferCache; // @[Slice.scala 94:16]
  wire  abc_mshr_13_io_alloc_bits_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_13_io_alloc_bits_fromProbeHelper; // @[Slice.scala 94:16]
  wire  abc_mshr_13_io_alloc_bits_fromCmoHelper; // @[Slice.scala 94:16]
  wire  abc_mshr_13_io_alloc_bits_needProbeAckData; // @[Slice.scala 94:16]
  wire  abc_mshr_13_io_status_valid; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_13_io_status_bits_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_13_io_status_bits_tag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_13_io_status_bits_way; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_13_io_status_bits_way_reg; // @[Slice.scala 94:16]
  wire  abc_mshr_13_io_status_bits_nestB; // @[Slice.scala 94:16]
  wire  abc_mshr_13_io_status_bits_nestC; // @[Slice.scala 94:16]
  wire  abc_mshr_13_io_status_bits_will_grant_data; // @[Slice.scala 94:16]
  wire  abc_mshr_13_io_status_bits_will_save_data; // @[Slice.scala 94:16]
  wire  abc_mshr_13_io_status_bits_will_free; // @[Slice.scala 94:16]
  wire  abc_mshr_13_io_resps_sink_c_valid; // @[Slice.scala 94:16]
  wire  abc_mshr_13_io_resps_sink_c_bits_hasData; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_13_io_resps_sink_c_bits_param; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_13_io_resps_sink_c_bits_source; // @[Slice.scala 94:16]
  wire  abc_mshr_13_io_resps_sink_c_bits_last; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_13_io_resps_sink_c_bits_bufIdx; // @[Slice.scala 94:16]
  wire  abc_mshr_13_io_resps_sink_d_valid; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_13_io_resps_sink_d_bits_opcode; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_13_io_resps_sink_d_bits_param; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_13_io_resps_sink_d_bits_sink; // @[Slice.scala 94:16]
  wire  abc_mshr_13_io_resps_sink_d_bits_last; // @[Slice.scala 94:16]
  wire  abc_mshr_13_io_resps_sink_d_bits_denied; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_13_io_resps_sink_d_bits_bufIdx; // @[Slice.scala 94:16]
  wire  abc_mshr_13_io_resps_sink_e_valid; // @[Slice.scala 94:16]
  wire  abc_mshr_13_io_resps_source_d_valid; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_13_io_nestedwb_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_13_io_nestedwb_tag; // @[Slice.scala 94:16]
  wire  abc_mshr_13_io_nestedwb_btoN; // @[Slice.scala 94:16]
  wire  abc_mshr_13_io_nestedwb_btoB; // @[Slice.scala 94:16]
  wire  abc_mshr_13_io_nestedwb_bclr_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_13_io_nestedwb_bset_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_13_io_nestedwb_c_set_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_13_io_nestedwb_c_set_hit; // @[Slice.scala 94:16]
  wire  abc_mshr_13_io_nestedwb_clients_0_isToN; // @[Slice.scala 94:16]
  wire  abc_mshr_13_io_nestedwb_clients_1_isToN; // @[Slice.scala 94:16]
  wire  abc_mshr_13_io_tasks_sink_a_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_13_io_tasks_sink_a_valid; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_13_io_tasks_sink_a_bits_sourceId; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_13_io_tasks_sink_a_bits_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_13_io_tasks_sink_a_bits_tag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_13_io_tasks_sink_a_bits_size; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_13_io_tasks_sink_a_bits_off; // @[Slice.scala 94:16]
  wire  abc_mshr_13_io_tasks_source_bready; // @[Slice.scala 94:16]
  wire  abc_mshr_13_io_tasks_source_bvalid; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_13_io_tasks_source_bset; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_13_io_tasks_source_btag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_13_io_tasks_source_bparam; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_13_io_tasks_source_bclients; // @[Slice.scala 94:16]
  wire  abc_mshr_13_io_tasks_source_bneedData; // @[Slice.scala 94:16]
  wire  abc_mshr_13_io_tasks_sink_c_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_13_io_tasks_sink_c_valid; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_13_io_tasks_sink_c_bits_sourceId; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_13_io_tasks_sink_c_bits_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_13_io_tasks_sink_c_bits_tag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_13_io_tasks_sink_c_bits_size; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_13_io_tasks_sink_c_bits_way; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_13_io_tasks_sink_c_bits_off; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_13_io_tasks_sink_c_bits_bufIdx; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_13_io_tasks_sink_c_bits_opcode; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_13_io_tasks_sink_c_bits_param; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_13_io_tasks_sink_c_bits_source; // @[Slice.scala 94:16]
  wire  abc_mshr_13_io_tasks_sink_c_bits_save; // @[Slice.scala 94:16]
  wire  abc_mshr_13_io_tasks_sink_c_bits_drop; // @[Slice.scala 94:16]
  wire  abc_mshr_13_io_tasks_sink_c_bits_release; // @[Slice.scala 94:16]
  wire  abc_mshr_13_io_tasks_sink_c_bits_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_13_io_tasks_source_d_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_13_io_tasks_source_d_valid; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_13_io_tasks_source_d_bits_sourceId; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_13_io_tasks_source_d_bits_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_13_io_tasks_source_d_bits_tag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_13_io_tasks_source_d_bits_channel; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_13_io_tasks_source_d_bits_opcode; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_13_io_tasks_source_d_bits_param; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_13_io_tasks_source_d_bits_size; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_13_io_tasks_source_d_bits_way; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_13_io_tasks_source_d_bits_off; // @[Slice.scala 94:16]
  wire  abc_mshr_13_io_tasks_source_d_bits_useBypass; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_13_io_tasks_source_d_bits_bufIdx; // @[Slice.scala 94:16]
  wire  abc_mshr_13_io_tasks_source_d_bits_denied; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_13_io_tasks_source_d_bits_sinkId; // @[Slice.scala 94:16]
  wire  abc_mshr_13_io_tasks_source_d_bits_bypassPut; // @[Slice.scala 94:16]
  wire  abc_mshr_13_io_tasks_source_d_bits_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_13_io_tasks_source_a_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_13_io_tasks_source_a_valid; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_13_io_tasks_source_a_bits_tag; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_13_io_tasks_source_a_bits_set; // @[Slice.scala 94:16]
  wire [5:0] abc_mshr_13_io_tasks_source_a_bits_off; // @[Slice.scala 94:16]
  wire [31:0] abc_mshr_13_io_tasks_source_a_bits_mask; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_13_io_tasks_source_a_bits_opcode; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_13_io_tasks_source_a_bits_param; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_13_io_tasks_source_a_bits_source; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_13_io_tasks_source_a_bits_bufIdx; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_13_io_tasks_source_a_bits_size; // @[Slice.scala 94:16]
  wire  abc_mshr_13_io_tasks_source_a_bits_needData; // @[Slice.scala 94:16]
  wire  abc_mshr_13_io_tasks_source_a_bits_putData; // @[Slice.scala 94:16]
  wire  abc_mshr_13_io_tasks_source_c_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_13_io_tasks_source_c_valid; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_13_io_tasks_source_c_bits_opcode; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_13_io_tasks_source_c_bits_tag; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_13_io_tasks_source_c_bits_set; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_13_io_tasks_source_c_bits_param; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_13_io_tasks_source_c_bits_source; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_13_io_tasks_source_c_bits_way; // @[Slice.scala 94:16]
  wire  abc_mshr_13_io_tasks_source_c_bits_dirty; // @[Slice.scala 94:16]
  wire  abc_mshr_13_io_tasks_source_e_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_13_io_tasks_source_e_valid; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_13_io_tasks_source_e_bits_sink; // @[Slice.scala 94:16]
  wire  abc_mshr_13_io_tasks_dir_write_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_13_io_tasks_dir_write_valid; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_13_io_tasks_dir_write_bits_set; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_13_io_tasks_dir_write_bits_way; // @[Slice.scala 94:16]
  wire  abc_mshr_13_io_tasks_dir_write_bits_data_dirty; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_13_io_tasks_dir_write_bits_data_state; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_13_io_tasks_dir_write_bits_data_clientStates_0; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_13_io_tasks_dir_write_bits_data_clientStates_1; // @[Slice.scala 94:16]
  wire  abc_mshr_13_io_tasks_tag_write_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_13_io_tasks_tag_write_valid; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_13_io_tasks_tag_write_bits_set; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_13_io_tasks_tag_write_bits_way; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_13_io_tasks_tag_write_bits_tag; // @[Slice.scala 94:16]
  wire  abc_mshr_13_io_tasks_client_dir_write_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_13_io_tasks_client_dir_write_valid; // @[Slice.scala 94:16]
  wire [6:0] abc_mshr_13_io_tasks_client_dir_write_bits_set; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_13_io_tasks_client_dir_write_bits_way; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_13_io_tasks_client_dir_write_bits_data_0_state; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_13_io_tasks_client_dir_write_bits_data_1_state; // @[Slice.scala 94:16]
  wire  abc_mshr_13_io_tasks_client_tag_write_ready; // @[Slice.scala 94:16]
  wire  abc_mshr_13_io_tasks_client_tag_write_valid; // @[Slice.scala 94:16]
  wire [6:0] abc_mshr_13_io_tasks_client_tag_write_bits_set; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_13_io_tasks_client_tag_write_bits_way; // @[Slice.scala 94:16]
  wire [22:0] abc_mshr_13_io_tasks_client_tag_write_bits_tag; // @[Slice.scala 94:16]
  wire  abc_mshr_13_io_dirResult_valid; // @[Slice.scala 94:16]
  wire  abc_mshr_13_io_dirResult_bits_self_dirty; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_13_io_dirResult_bits_self_state; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_13_io_dirResult_bits_self_clientStates_0; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_13_io_dirResult_bits_self_clientStates_1; // @[Slice.scala 94:16]
  wire  abc_mshr_13_io_dirResult_bits_self_hit; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_13_io_dirResult_bits_self_way; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_13_io_dirResult_bits_self_tag; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_13_io_dirResult_bits_clients_states_0_state; // @[Slice.scala 94:16]
  wire  abc_mshr_13_io_dirResult_bits_clients_states_0_hit; // @[Slice.scala 94:16]
  wire [1:0] abc_mshr_13_io_dirResult_bits_clients_states_1_state; // @[Slice.scala 94:16]
  wire  abc_mshr_13_io_dirResult_bits_clients_states_1_hit; // @[Slice.scala 94:16]
  wire [22:0] abc_mshr_13_io_dirResult_bits_clients_tag; // @[Slice.scala 94:16]
  wire [3:0] abc_mshr_13_io_dirResult_bits_clients_way; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_13_io_c_status_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_13_io_c_status_tag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_13_io_c_status_way; // @[Slice.scala 94:16]
  wire  abc_mshr_13_io_c_status_nestedReleaseData; // @[Slice.scala 94:16]
  wire  abc_mshr_13_io_c_status_releaseThrough; // @[Slice.scala 94:16]
  wire [9:0] abc_mshr_13_io_bstatus_set; // @[Slice.scala 94:16]
  wire [19:0] abc_mshr_13_io_bstatus_tag; // @[Slice.scala 94:16]
  wire [2:0] abc_mshr_13_io_bstatus_way; // @[Slice.scala 94:16]
  wire  abc_mshr_13_io_bstatus_nestedProbeAckData; // @[Slice.scala 94:16]
  wire  abc_mshr_13_io_bstatus_probeHelperFinish; // @[Slice.scala 94:16]
  wire  abc_mshr_13_io_bstatus_probeAckDataThrough; // @[Slice.scala 94:16]
  wire  abc_mshr_13_io_releaseThrough; // @[Slice.scala 94:16]
  wire  abc_mshr_13_io_probeAckDataThrough; // @[Slice.scala 94:16]
  wire  abc_mshr_13_io_is_nestedReleaseData; // @[Slice.scala 94:16]
  wire  abc_mshr_13_io_is_nestedProbeAckData; // @[Slice.scala 94:16]
  wire  abc_mshr_13_io_probeHelperFinish; // @[Slice.scala 94:16]
  wire  bc_mshr_clock; // @[Slice.scala 94:16]
  wire  bc_mshr_reset; // @[Slice.scala 94:16]
  wire [3:0] bc_mshr_io_id; // @[Slice.scala 94:16]
  wire  bc_mshr_io_enable; // @[Slice.scala 94:16]
  wire  bc_mshr_io_alloc_valid; // @[Slice.scala 94:16]
  wire [2:0] bc_mshr_io_alloc_bits_channel; // @[Slice.scala 94:16]
  wire [2:0] bc_mshr_io_alloc_bits_opcode; // @[Slice.scala 94:16]
  wire [2:0] bc_mshr_io_alloc_bits_param; // @[Slice.scala 94:16]
  wire [2:0] bc_mshr_io_alloc_bits_size; // @[Slice.scala 94:16]
  wire [5:0] bc_mshr_io_alloc_bits_source; // @[Slice.scala 94:16]
  wire [9:0] bc_mshr_io_alloc_bits_set; // @[Slice.scala 94:16]
  wire [19:0] bc_mshr_io_alloc_bits_tag; // @[Slice.scala 94:16]
  wire [5:0] bc_mshr_io_alloc_bits_off; // @[Slice.scala 94:16]
  wire [31:0] bc_mshr_io_alloc_bits_mask; // @[Slice.scala 94:16]
  wire [2:0] bc_mshr_io_alloc_bits_bufIdx; // @[Slice.scala 94:16]
  wire  bc_mshr_io_alloc_bits_preferCache; // @[Slice.scala 94:16]
  wire  bc_mshr_io_alloc_bits_dirty; // @[Slice.scala 94:16]
  wire  bc_mshr_io_alloc_bits_fromProbeHelper; // @[Slice.scala 94:16]
  wire  bc_mshr_io_alloc_bits_fromCmoHelper; // @[Slice.scala 94:16]
  wire  bc_mshr_io_alloc_bits_needProbeAckData; // @[Slice.scala 94:16]
  wire  bc_mshr_io_status_valid; // @[Slice.scala 94:16]
  wire [9:0] bc_mshr_io_status_bits_set; // @[Slice.scala 94:16]
  wire [19:0] bc_mshr_io_status_bits_tag; // @[Slice.scala 94:16]
  wire [2:0] bc_mshr_io_status_bits_way; // @[Slice.scala 94:16]
  wire [2:0] bc_mshr_io_status_bits_way_reg; // @[Slice.scala 94:16]
  wire  bc_mshr_io_status_bits_nestB; // @[Slice.scala 94:16]
  wire  bc_mshr_io_status_bits_nestC; // @[Slice.scala 94:16]
  wire  bc_mshr_io_status_bits_will_grant_data; // @[Slice.scala 94:16]
  wire  bc_mshr_io_status_bits_will_save_data; // @[Slice.scala 94:16]
  wire  bc_mshr_io_status_bits_will_free; // @[Slice.scala 94:16]
  wire  bc_mshr_io_resps_sink_c_valid; // @[Slice.scala 94:16]
  wire  bc_mshr_io_resps_sink_c_bits_hasData; // @[Slice.scala 94:16]
  wire [2:0] bc_mshr_io_resps_sink_c_bits_param; // @[Slice.scala 94:16]
  wire [5:0] bc_mshr_io_resps_sink_c_bits_source; // @[Slice.scala 94:16]
  wire  bc_mshr_io_resps_sink_c_bits_last; // @[Slice.scala 94:16]
  wire [2:0] bc_mshr_io_resps_sink_c_bits_bufIdx; // @[Slice.scala 94:16]
  wire  bc_mshr_io_resps_sink_d_valid; // @[Slice.scala 94:16]
  wire [2:0] bc_mshr_io_resps_sink_d_bits_opcode; // @[Slice.scala 94:16]
  wire [2:0] bc_mshr_io_resps_sink_d_bits_param; // @[Slice.scala 94:16]
  wire [2:0] bc_mshr_io_resps_sink_d_bits_sink; // @[Slice.scala 94:16]
  wire  bc_mshr_io_resps_sink_d_bits_last; // @[Slice.scala 94:16]
  wire  bc_mshr_io_resps_sink_d_bits_denied; // @[Slice.scala 94:16]
  wire [2:0] bc_mshr_io_resps_sink_d_bits_bufIdx; // @[Slice.scala 94:16]
  wire  bc_mshr_io_resps_sink_e_valid; // @[Slice.scala 94:16]
  wire  bc_mshr_io_resps_source_d_valid; // @[Slice.scala 94:16]
  wire [9:0] bc_mshr_io_nestedwb_set; // @[Slice.scala 94:16]
  wire [19:0] bc_mshr_io_nestedwb_tag; // @[Slice.scala 94:16]
  wire  bc_mshr_io_nestedwb_btoN; // @[Slice.scala 94:16]
  wire  bc_mshr_io_nestedwb_btoB; // @[Slice.scala 94:16]
  wire  bc_mshr_io_nestedwb_bclr_dirty; // @[Slice.scala 94:16]
  wire  bc_mshr_io_nestedwb_bset_dirty; // @[Slice.scala 94:16]
  wire  bc_mshr_io_nestedwb_c_set_dirty; // @[Slice.scala 94:16]
  wire  bc_mshr_io_nestedwb_c_set_hit; // @[Slice.scala 94:16]
  wire  bc_mshr_io_nestedwb_clients_0_isToN; // @[Slice.scala 94:16]
  wire  bc_mshr_io_nestedwb_clients_1_isToN; // @[Slice.scala 94:16]
  wire  bc_mshr_io_tasks_sink_a_ready; // @[Slice.scala 94:16]
  wire  bc_mshr_io_tasks_sink_a_valid; // @[Slice.scala 94:16]
  wire [5:0] bc_mshr_io_tasks_sink_a_bits_sourceId; // @[Slice.scala 94:16]
  wire [9:0] bc_mshr_io_tasks_sink_a_bits_set; // @[Slice.scala 94:16]
  wire [19:0] bc_mshr_io_tasks_sink_a_bits_tag; // @[Slice.scala 94:16]
  wire [2:0] bc_mshr_io_tasks_sink_a_bits_size; // @[Slice.scala 94:16]
  wire [5:0] bc_mshr_io_tasks_sink_a_bits_off; // @[Slice.scala 94:16]
  wire  bc_mshr_io_tasks_source_bready; // @[Slice.scala 94:16]
  wire  bc_mshr_io_tasks_source_bvalid; // @[Slice.scala 94:16]
  wire [9:0] bc_mshr_io_tasks_source_bset; // @[Slice.scala 94:16]
  wire [19:0] bc_mshr_io_tasks_source_btag; // @[Slice.scala 94:16]
  wire [2:0] bc_mshr_io_tasks_source_bparam; // @[Slice.scala 94:16]
  wire [1:0] bc_mshr_io_tasks_source_bclients; // @[Slice.scala 94:16]
  wire  bc_mshr_io_tasks_source_bneedData; // @[Slice.scala 94:16]
  wire  bc_mshr_io_tasks_sink_c_ready; // @[Slice.scala 94:16]
  wire  bc_mshr_io_tasks_sink_c_valid; // @[Slice.scala 94:16]
  wire [5:0] bc_mshr_io_tasks_sink_c_bits_sourceId; // @[Slice.scala 94:16]
  wire [9:0] bc_mshr_io_tasks_sink_c_bits_set; // @[Slice.scala 94:16]
  wire [19:0] bc_mshr_io_tasks_sink_c_bits_tag; // @[Slice.scala 94:16]
  wire [2:0] bc_mshr_io_tasks_sink_c_bits_size; // @[Slice.scala 94:16]
  wire [2:0] bc_mshr_io_tasks_sink_c_bits_way; // @[Slice.scala 94:16]
  wire [5:0] bc_mshr_io_tasks_sink_c_bits_off; // @[Slice.scala 94:16]
  wire [2:0] bc_mshr_io_tasks_sink_c_bits_bufIdx; // @[Slice.scala 94:16]
  wire [2:0] bc_mshr_io_tasks_sink_c_bits_opcode; // @[Slice.scala 94:16]
  wire [2:0] bc_mshr_io_tasks_sink_c_bits_param; // @[Slice.scala 94:16]
  wire [3:0] bc_mshr_io_tasks_sink_c_bits_source; // @[Slice.scala 94:16]
  wire  bc_mshr_io_tasks_sink_c_bits_save; // @[Slice.scala 94:16]
  wire  bc_mshr_io_tasks_sink_c_bits_drop; // @[Slice.scala 94:16]
  wire  bc_mshr_io_tasks_sink_c_bits_release; // @[Slice.scala 94:16]
  wire  bc_mshr_io_tasks_sink_c_bits_dirty; // @[Slice.scala 94:16]
  wire  bc_mshr_io_tasks_source_d_ready; // @[Slice.scala 94:16]
  wire  bc_mshr_io_tasks_source_d_valid; // @[Slice.scala 94:16]
  wire [5:0] bc_mshr_io_tasks_source_d_bits_sourceId; // @[Slice.scala 94:16]
  wire [9:0] bc_mshr_io_tasks_source_d_bits_set; // @[Slice.scala 94:16]
  wire [19:0] bc_mshr_io_tasks_source_d_bits_tag; // @[Slice.scala 94:16]
  wire [2:0] bc_mshr_io_tasks_source_d_bits_channel; // @[Slice.scala 94:16]
  wire [2:0] bc_mshr_io_tasks_source_d_bits_opcode; // @[Slice.scala 94:16]
  wire [2:0] bc_mshr_io_tasks_source_d_bits_param; // @[Slice.scala 94:16]
  wire [2:0] bc_mshr_io_tasks_source_d_bits_size; // @[Slice.scala 94:16]
  wire [2:0] bc_mshr_io_tasks_source_d_bits_way; // @[Slice.scala 94:16]
  wire [5:0] bc_mshr_io_tasks_source_d_bits_off; // @[Slice.scala 94:16]
  wire  bc_mshr_io_tasks_source_d_bits_useBypass; // @[Slice.scala 94:16]
  wire [2:0] bc_mshr_io_tasks_source_d_bits_bufIdx; // @[Slice.scala 94:16]
  wire  bc_mshr_io_tasks_source_d_bits_denied; // @[Slice.scala 94:16]
  wire [3:0] bc_mshr_io_tasks_source_d_bits_sinkId; // @[Slice.scala 94:16]
  wire  bc_mshr_io_tasks_source_d_bits_bypassPut; // @[Slice.scala 94:16]
  wire  bc_mshr_io_tasks_source_d_bits_dirty; // @[Slice.scala 94:16]
  wire  bc_mshr_io_tasks_source_a_ready; // @[Slice.scala 94:16]
  wire  bc_mshr_io_tasks_source_a_valid; // @[Slice.scala 94:16]
  wire [19:0] bc_mshr_io_tasks_source_a_bits_tag; // @[Slice.scala 94:16]
  wire [9:0] bc_mshr_io_tasks_source_a_bits_set; // @[Slice.scala 94:16]
  wire [5:0] bc_mshr_io_tasks_source_a_bits_off; // @[Slice.scala 94:16]
  wire [31:0] bc_mshr_io_tasks_source_a_bits_mask; // @[Slice.scala 94:16]
  wire [2:0] bc_mshr_io_tasks_source_a_bits_opcode; // @[Slice.scala 94:16]
  wire [2:0] bc_mshr_io_tasks_source_a_bits_param; // @[Slice.scala 94:16]
  wire [3:0] bc_mshr_io_tasks_source_a_bits_source; // @[Slice.scala 94:16]
  wire [2:0] bc_mshr_io_tasks_source_a_bits_bufIdx; // @[Slice.scala 94:16]
  wire [2:0] bc_mshr_io_tasks_source_a_bits_size; // @[Slice.scala 94:16]
  wire  bc_mshr_io_tasks_source_a_bits_needData; // @[Slice.scala 94:16]
  wire  bc_mshr_io_tasks_source_a_bits_putData; // @[Slice.scala 94:16]
  wire  bc_mshr_io_tasks_source_c_ready; // @[Slice.scala 94:16]
  wire  bc_mshr_io_tasks_source_c_valid; // @[Slice.scala 94:16]
  wire [2:0] bc_mshr_io_tasks_source_c_bits_opcode; // @[Slice.scala 94:16]
  wire [19:0] bc_mshr_io_tasks_source_c_bits_tag; // @[Slice.scala 94:16]
  wire [9:0] bc_mshr_io_tasks_source_c_bits_set; // @[Slice.scala 94:16]
  wire [2:0] bc_mshr_io_tasks_source_c_bits_param; // @[Slice.scala 94:16]
  wire [3:0] bc_mshr_io_tasks_source_c_bits_source; // @[Slice.scala 94:16]
  wire [2:0] bc_mshr_io_tasks_source_c_bits_way; // @[Slice.scala 94:16]
  wire  bc_mshr_io_tasks_source_c_bits_dirty; // @[Slice.scala 94:16]
  wire  bc_mshr_io_tasks_source_e_ready; // @[Slice.scala 94:16]
  wire  bc_mshr_io_tasks_source_e_valid; // @[Slice.scala 94:16]
  wire [2:0] bc_mshr_io_tasks_source_e_bits_sink; // @[Slice.scala 94:16]
  wire  bc_mshr_io_tasks_dir_write_ready; // @[Slice.scala 94:16]
  wire  bc_mshr_io_tasks_dir_write_valid; // @[Slice.scala 94:16]
  wire [9:0] bc_mshr_io_tasks_dir_write_bits_set; // @[Slice.scala 94:16]
  wire [2:0] bc_mshr_io_tasks_dir_write_bits_way; // @[Slice.scala 94:16]
  wire  bc_mshr_io_tasks_dir_write_bits_data_dirty; // @[Slice.scala 94:16]
  wire [1:0] bc_mshr_io_tasks_dir_write_bits_data_state; // @[Slice.scala 94:16]
  wire [1:0] bc_mshr_io_tasks_dir_write_bits_data_clientStates_0; // @[Slice.scala 94:16]
  wire [1:0] bc_mshr_io_tasks_dir_write_bits_data_clientStates_1; // @[Slice.scala 94:16]
  wire  bc_mshr_io_tasks_tag_write_ready; // @[Slice.scala 94:16]
  wire  bc_mshr_io_tasks_tag_write_valid; // @[Slice.scala 94:16]
  wire [9:0] bc_mshr_io_tasks_tag_write_bits_set; // @[Slice.scala 94:16]
  wire [2:0] bc_mshr_io_tasks_tag_write_bits_way; // @[Slice.scala 94:16]
  wire [19:0] bc_mshr_io_tasks_tag_write_bits_tag; // @[Slice.scala 94:16]
  wire  bc_mshr_io_tasks_client_dir_write_ready; // @[Slice.scala 94:16]
  wire  bc_mshr_io_tasks_client_dir_write_valid; // @[Slice.scala 94:16]
  wire [6:0] bc_mshr_io_tasks_client_dir_write_bits_set; // @[Slice.scala 94:16]
  wire [3:0] bc_mshr_io_tasks_client_dir_write_bits_way; // @[Slice.scala 94:16]
  wire [1:0] bc_mshr_io_tasks_client_dir_write_bits_data_0_state; // @[Slice.scala 94:16]
  wire [1:0] bc_mshr_io_tasks_client_dir_write_bits_data_1_state; // @[Slice.scala 94:16]
  wire  bc_mshr_io_tasks_client_tag_write_ready; // @[Slice.scala 94:16]
  wire  bc_mshr_io_tasks_client_tag_write_valid; // @[Slice.scala 94:16]
  wire [6:0] bc_mshr_io_tasks_client_tag_write_bits_set; // @[Slice.scala 94:16]
  wire [3:0] bc_mshr_io_tasks_client_tag_write_bits_way; // @[Slice.scala 94:16]
  wire [22:0] bc_mshr_io_tasks_client_tag_write_bits_tag; // @[Slice.scala 94:16]
  wire  bc_mshr_io_dirResult_valid; // @[Slice.scala 94:16]
  wire  bc_mshr_io_dirResult_bits_self_dirty; // @[Slice.scala 94:16]
  wire [1:0] bc_mshr_io_dirResult_bits_self_state; // @[Slice.scala 94:16]
  wire [1:0] bc_mshr_io_dirResult_bits_self_clientStates_0; // @[Slice.scala 94:16]
  wire [1:0] bc_mshr_io_dirResult_bits_self_clientStates_1; // @[Slice.scala 94:16]
  wire  bc_mshr_io_dirResult_bits_self_hit; // @[Slice.scala 94:16]
  wire [2:0] bc_mshr_io_dirResult_bits_self_way; // @[Slice.scala 94:16]
  wire [19:0] bc_mshr_io_dirResult_bits_self_tag; // @[Slice.scala 94:16]
  wire [1:0] bc_mshr_io_dirResult_bits_clients_states_0_state; // @[Slice.scala 94:16]
  wire  bc_mshr_io_dirResult_bits_clients_states_0_hit; // @[Slice.scala 94:16]
  wire [1:0] bc_mshr_io_dirResult_bits_clients_states_1_state; // @[Slice.scala 94:16]
  wire  bc_mshr_io_dirResult_bits_clients_states_1_hit; // @[Slice.scala 94:16]
  wire [22:0] bc_mshr_io_dirResult_bits_clients_tag; // @[Slice.scala 94:16]
  wire [3:0] bc_mshr_io_dirResult_bits_clients_way; // @[Slice.scala 94:16]
  wire [9:0] bc_mshr_io_c_status_set; // @[Slice.scala 94:16]
  wire [19:0] bc_mshr_io_c_status_tag; // @[Slice.scala 94:16]
  wire [2:0] bc_mshr_io_c_status_way; // @[Slice.scala 94:16]
  wire  bc_mshr_io_c_status_nestedReleaseData; // @[Slice.scala 94:16]
  wire  bc_mshr_io_c_status_releaseThrough; // @[Slice.scala 94:16]
  wire [9:0] bc_mshr_io_bstatus_set; // @[Slice.scala 94:16]
  wire [19:0] bc_mshr_io_bstatus_tag; // @[Slice.scala 94:16]
  wire [2:0] bc_mshr_io_bstatus_way; // @[Slice.scala 94:16]
  wire  bc_mshr_io_bstatus_nestedProbeAckData; // @[Slice.scala 94:16]
  wire  bc_mshr_io_bstatus_probeHelperFinish; // @[Slice.scala 94:16]
  wire  bc_mshr_io_bstatus_probeAckDataThrough; // @[Slice.scala 94:16]
  wire  bc_mshr_io_releaseThrough; // @[Slice.scala 94:16]
  wire  bc_mshr_io_probeAckDataThrough; // @[Slice.scala 94:16]
  wire  bc_mshr_io_is_nestedReleaseData; // @[Slice.scala 94:16]
  wire  bc_mshr_io_is_nestedProbeAckData; // @[Slice.scala 94:16]
  wire  bc_mshr_io_probeHelperFinish; // @[Slice.scala 94:16]
  wire  c_mshr_clock; // @[Slice.scala 94:16]
  wire  c_mshr_reset; // @[Slice.scala 94:16]
  wire [3:0] c_mshr_io_id; // @[Slice.scala 94:16]
  wire  c_mshr_io_enable; // @[Slice.scala 94:16]
  wire  c_mshr_io_alloc_valid; // @[Slice.scala 94:16]
  wire [2:0] c_mshr_io_alloc_bits_channel; // @[Slice.scala 94:16]
  wire [2:0] c_mshr_io_alloc_bits_opcode; // @[Slice.scala 94:16]
  wire [2:0] c_mshr_io_alloc_bits_param; // @[Slice.scala 94:16]
  wire [2:0] c_mshr_io_alloc_bits_size; // @[Slice.scala 94:16]
  wire [5:0] c_mshr_io_alloc_bits_source; // @[Slice.scala 94:16]
  wire [9:0] c_mshr_io_alloc_bits_set; // @[Slice.scala 94:16]
  wire [19:0] c_mshr_io_alloc_bits_tag; // @[Slice.scala 94:16]
  wire [5:0] c_mshr_io_alloc_bits_off; // @[Slice.scala 94:16]
  wire [31:0] c_mshr_io_alloc_bits_mask; // @[Slice.scala 94:16]
  wire [2:0] c_mshr_io_alloc_bits_bufIdx; // @[Slice.scala 94:16]
  wire  c_mshr_io_alloc_bits_preferCache; // @[Slice.scala 94:16]
  wire  c_mshr_io_alloc_bits_dirty; // @[Slice.scala 94:16]
  wire  c_mshr_io_alloc_bits_fromProbeHelper; // @[Slice.scala 94:16]
  wire  c_mshr_io_alloc_bits_fromCmoHelper; // @[Slice.scala 94:16]
  wire  c_mshr_io_alloc_bits_needProbeAckData; // @[Slice.scala 94:16]
  wire  c_mshr_io_status_valid; // @[Slice.scala 94:16]
  wire [9:0] c_mshr_io_status_bits_set; // @[Slice.scala 94:16]
  wire [19:0] c_mshr_io_status_bits_tag; // @[Slice.scala 94:16]
  wire [2:0] c_mshr_io_status_bits_way; // @[Slice.scala 94:16]
  wire [2:0] c_mshr_io_status_bits_way_reg; // @[Slice.scala 94:16]
  wire  c_mshr_io_status_bits_nestB; // @[Slice.scala 94:16]
  wire  c_mshr_io_status_bits_nestC; // @[Slice.scala 94:16]
  wire  c_mshr_io_status_bits_will_grant_data; // @[Slice.scala 94:16]
  wire  c_mshr_io_status_bits_will_save_data; // @[Slice.scala 94:16]
  wire  c_mshr_io_status_bits_will_free; // @[Slice.scala 94:16]
  wire  c_mshr_io_resps_sink_c_valid; // @[Slice.scala 94:16]
  wire  c_mshr_io_resps_sink_c_bits_hasData; // @[Slice.scala 94:16]
  wire [2:0] c_mshr_io_resps_sink_c_bits_param; // @[Slice.scala 94:16]
  wire [5:0] c_mshr_io_resps_sink_c_bits_source; // @[Slice.scala 94:16]
  wire  c_mshr_io_resps_sink_c_bits_last; // @[Slice.scala 94:16]
  wire [2:0] c_mshr_io_resps_sink_c_bits_bufIdx; // @[Slice.scala 94:16]
  wire  c_mshr_io_resps_sink_d_valid; // @[Slice.scala 94:16]
  wire [2:0] c_mshr_io_resps_sink_d_bits_opcode; // @[Slice.scala 94:16]
  wire [2:0] c_mshr_io_resps_sink_d_bits_param; // @[Slice.scala 94:16]
  wire [2:0] c_mshr_io_resps_sink_d_bits_sink; // @[Slice.scala 94:16]
  wire  c_mshr_io_resps_sink_d_bits_last; // @[Slice.scala 94:16]
  wire  c_mshr_io_resps_sink_d_bits_denied; // @[Slice.scala 94:16]
  wire [2:0] c_mshr_io_resps_sink_d_bits_bufIdx; // @[Slice.scala 94:16]
  wire  c_mshr_io_resps_sink_e_valid; // @[Slice.scala 94:16]
  wire  c_mshr_io_resps_source_d_valid; // @[Slice.scala 94:16]
  wire [9:0] c_mshr_io_nestedwb_set; // @[Slice.scala 94:16]
  wire [19:0] c_mshr_io_nestedwb_tag; // @[Slice.scala 94:16]
  wire  c_mshr_io_nestedwb_btoN; // @[Slice.scala 94:16]
  wire  c_mshr_io_nestedwb_btoB; // @[Slice.scala 94:16]
  wire  c_mshr_io_nestedwb_bclr_dirty; // @[Slice.scala 94:16]
  wire  c_mshr_io_nestedwb_bset_dirty; // @[Slice.scala 94:16]
  wire  c_mshr_io_nestedwb_c_set_dirty; // @[Slice.scala 94:16]
  wire  c_mshr_io_nestedwb_c_set_hit; // @[Slice.scala 94:16]
  wire  c_mshr_io_nestedwb_clients_0_isToN; // @[Slice.scala 94:16]
  wire  c_mshr_io_nestedwb_clients_1_isToN; // @[Slice.scala 94:16]
  wire  c_mshr_io_tasks_sink_a_ready; // @[Slice.scala 94:16]
  wire  c_mshr_io_tasks_sink_a_valid; // @[Slice.scala 94:16]
  wire [5:0] c_mshr_io_tasks_sink_a_bits_sourceId; // @[Slice.scala 94:16]
  wire [9:0] c_mshr_io_tasks_sink_a_bits_set; // @[Slice.scala 94:16]
  wire [19:0] c_mshr_io_tasks_sink_a_bits_tag; // @[Slice.scala 94:16]
  wire [2:0] c_mshr_io_tasks_sink_a_bits_size; // @[Slice.scala 94:16]
  wire [5:0] c_mshr_io_tasks_sink_a_bits_off; // @[Slice.scala 94:16]
  wire  c_mshr_io_tasks_source_bready; // @[Slice.scala 94:16]
  wire  c_mshr_io_tasks_source_bvalid; // @[Slice.scala 94:16]
  wire [9:0] c_mshr_io_tasks_source_bset; // @[Slice.scala 94:16]
  wire [19:0] c_mshr_io_tasks_source_btag; // @[Slice.scala 94:16]
  wire [2:0] c_mshr_io_tasks_source_bparam; // @[Slice.scala 94:16]
  wire [1:0] c_mshr_io_tasks_source_bclients; // @[Slice.scala 94:16]
  wire  c_mshr_io_tasks_source_bneedData; // @[Slice.scala 94:16]
  wire  c_mshr_io_tasks_sink_c_ready; // @[Slice.scala 94:16]
  wire  c_mshr_io_tasks_sink_c_valid; // @[Slice.scala 94:16]
  wire [5:0] c_mshr_io_tasks_sink_c_bits_sourceId; // @[Slice.scala 94:16]
  wire [9:0] c_mshr_io_tasks_sink_c_bits_set; // @[Slice.scala 94:16]
  wire [19:0] c_mshr_io_tasks_sink_c_bits_tag; // @[Slice.scala 94:16]
  wire [2:0] c_mshr_io_tasks_sink_c_bits_size; // @[Slice.scala 94:16]
  wire [2:0] c_mshr_io_tasks_sink_c_bits_way; // @[Slice.scala 94:16]
  wire [5:0] c_mshr_io_tasks_sink_c_bits_off; // @[Slice.scala 94:16]
  wire [2:0] c_mshr_io_tasks_sink_c_bits_bufIdx; // @[Slice.scala 94:16]
  wire [2:0] c_mshr_io_tasks_sink_c_bits_opcode; // @[Slice.scala 94:16]
  wire [2:0] c_mshr_io_tasks_sink_c_bits_param; // @[Slice.scala 94:16]
  wire [3:0] c_mshr_io_tasks_sink_c_bits_source; // @[Slice.scala 94:16]
  wire  c_mshr_io_tasks_sink_c_bits_save; // @[Slice.scala 94:16]
  wire  c_mshr_io_tasks_sink_c_bits_drop; // @[Slice.scala 94:16]
  wire  c_mshr_io_tasks_sink_c_bits_release; // @[Slice.scala 94:16]
  wire  c_mshr_io_tasks_sink_c_bits_dirty; // @[Slice.scala 94:16]
  wire  c_mshr_io_tasks_source_d_ready; // @[Slice.scala 94:16]
  wire  c_mshr_io_tasks_source_d_valid; // @[Slice.scala 94:16]
  wire [5:0] c_mshr_io_tasks_source_d_bits_sourceId; // @[Slice.scala 94:16]
  wire [9:0] c_mshr_io_tasks_source_d_bits_set; // @[Slice.scala 94:16]
  wire [19:0] c_mshr_io_tasks_source_d_bits_tag; // @[Slice.scala 94:16]
  wire [2:0] c_mshr_io_tasks_source_d_bits_channel; // @[Slice.scala 94:16]
  wire [2:0] c_mshr_io_tasks_source_d_bits_opcode; // @[Slice.scala 94:16]
  wire [2:0] c_mshr_io_tasks_source_d_bits_param; // @[Slice.scala 94:16]
  wire [2:0] c_mshr_io_tasks_source_d_bits_size; // @[Slice.scala 94:16]
  wire [2:0] c_mshr_io_tasks_source_d_bits_way; // @[Slice.scala 94:16]
  wire [5:0] c_mshr_io_tasks_source_d_bits_off; // @[Slice.scala 94:16]
  wire  c_mshr_io_tasks_source_d_bits_useBypass; // @[Slice.scala 94:16]
  wire [2:0] c_mshr_io_tasks_source_d_bits_bufIdx; // @[Slice.scala 94:16]
  wire  c_mshr_io_tasks_source_d_bits_denied; // @[Slice.scala 94:16]
  wire [3:0] c_mshr_io_tasks_source_d_bits_sinkId; // @[Slice.scala 94:16]
  wire  c_mshr_io_tasks_source_d_bits_bypassPut; // @[Slice.scala 94:16]
  wire  c_mshr_io_tasks_source_d_bits_dirty; // @[Slice.scala 94:16]
  wire  c_mshr_io_tasks_source_a_ready; // @[Slice.scala 94:16]
  wire  c_mshr_io_tasks_source_a_valid; // @[Slice.scala 94:16]
  wire [19:0] c_mshr_io_tasks_source_a_bits_tag; // @[Slice.scala 94:16]
  wire [9:0] c_mshr_io_tasks_source_a_bits_set; // @[Slice.scala 94:16]
  wire [5:0] c_mshr_io_tasks_source_a_bits_off; // @[Slice.scala 94:16]
  wire [31:0] c_mshr_io_tasks_source_a_bits_mask; // @[Slice.scala 94:16]
  wire [2:0] c_mshr_io_tasks_source_a_bits_opcode; // @[Slice.scala 94:16]
  wire [2:0] c_mshr_io_tasks_source_a_bits_param; // @[Slice.scala 94:16]
  wire [3:0] c_mshr_io_tasks_source_a_bits_source; // @[Slice.scala 94:16]
  wire [2:0] c_mshr_io_tasks_source_a_bits_bufIdx; // @[Slice.scala 94:16]
  wire [2:0] c_mshr_io_tasks_source_a_bits_size; // @[Slice.scala 94:16]
  wire  c_mshr_io_tasks_source_a_bits_needData; // @[Slice.scala 94:16]
  wire  c_mshr_io_tasks_source_a_bits_putData; // @[Slice.scala 94:16]
  wire  c_mshr_io_tasks_source_c_ready; // @[Slice.scala 94:16]
  wire  c_mshr_io_tasks_source_c_valid; // @[Slice.scala 94:16]
  wire [2:0] c_mshr_io_tasks_source_c_bits_opcode; // @[Slice.scala 94:16]
  wire [19:0] c_mshr_io_tasks_source_c_bits_tag; // @[Slice.scala 94:16]
  wire [9:0] c_mshr_io_tasks_source_c_bits_set; // @[Slice.scala 94:16]
  wire [2:0] c_mshr_io_tasks_source_c_bits_param; // @[Slice.scala 94:16]
  wire [3:0] c_mshr_io_tasks_source_c_bits_source; // @[Slice.scala 94:16]
  wire [2:0] c_mshr_io_tasks_source_c_bits_way; // @[Slice.scala 94:16]
  wire  c_mshr_io_tasks_source_c_bits_dirty; // @[Slice.scala 94:16]
  wire  c_mshr_io_tasks_source_e_ready; // @[Slice.scala 94:16]
  wire  c_mshr_io_tasks_source_e_valid; // @[Slice.scala 94:16]
  wire [2:0] c_mshr_io_tasks_source_e_bits_sink; // @[Slice.scala 94:16]
  wire  c_mshr_io_tasks_dir_write_ready; // @[Slice.scala 94:16]
  wire  c_mshr_io_tasks_dir_write_valid; // @[Slice.scala 94:16]
  wire [9:0] c_mshr_io_tasks_dir_write_bits_set; // @[Slice.scala 94:16]
  wire [2:0] c_mshr_io_tasks_dir_write_bits_way; // @[Slice.scala 94:16]
  wire  c_mshr_io_tasks_dir_write_bits_data_dirty; // @[Slice.scala 94:16]
  wire [1:0] c_mshr_io_tasks_dir_write_bits_data_state; // @[Slice.scala 94:16]
  wire [1:0] c_mshr_io_tasks_dir_write_bits_data_clientStates_0; // @[Slice.scala 94:16]
  wire [1:0] c_mshr_io_tasks_dir_write_bits_data_clientStates_1; // @[Slice.scala 94:16]
  wire  c_mshr_io_tasks_tag_write_ready; // @[Slice.scala 94:16]
  wire  c_mshr_io_tasks_tag_write_valid; // @[Slice.scala 94:16]
  wire [9:0] c_mshr_io_tasks_tag_write_bits_set; // @[Slice.scala 94:16]
  wire [2:0] c_mshr_io_tasks_tag_write_bits_way; // @[Slice.scala 94:16]
  wire [19:0] c_mshr_io_tasks_tag_write_bits_tag; // @[Slice.scala 94:16]
  wire  c_mshr_io_tasks_client_dir_write_ready; // @[Slice.scala 94:16]
  wire  c_mshr_io_tasks_client_dir_write_valid; // @[Slice.scala 94:16]
  wire [6:0] c_mshr_io_tasks_client_dir_write_bits_set; // @[Slice.scala 94:16]
  wire [3:0] c_mshr_io_tasks_client_dir_write_bits_way; // @[Slice.scala 94:16]
  wire [1:0] c_mshr_io_tasks_client_dir_write_bits_data_0_state; // @[Slice.scala 94:16]
  wire [1:0] c_mshr_io_tasks_client_dir_write_bits_data_1_state; // @[Slice.scala 94:16]
  wire  c_mshr_io_tasks_client_tag_write_ready; // @[Slice.scala 94:16]
  wire  c_mshr_io_tasks_client_tag_write_valid; // @[Slice.scala 94:16]
  wire [6:0] c_mshr_io_tasks_client_tag_write_bits_set; // @[Slice.scala 94:16]
  wire [3:0] c_mshr_io_tasks_client_tag_write_bits_way; // @[Slice.scala 94:16]
  wire [22:0] c_mshr_io_tasks_client_tag_write_bits_tag; // @[Slice.scala 94:16]
  wire  c_mshr_io_dirResult_valid; // @[Slice.scala 94:16]
  wire  c_mshr_io_dirResult_bits_self_dirty; // @[Slice.scala 94:16]
  wire [1:0] c_mshr_io_dirResult_bits_self_state; // @[Slice.scala 94:16]
  wire [1:0] c_mshr_io_dirResult_bits_self_clientStates_0; // @[Slice.scala 94:16]
  wire [1:0] c_mshr_io_dirResult_bits_self_clientStates_1; // @[Slice.scala 94:16]
  wire  c_mshr_io_dirResult_bits_self_hit; // @[Slice.scala 94:16]
  wire [2:0] c_mshr_io_dirResult_bits_self_way; // @[Slice.scala 94:16]
  wire [19:0] c_mshr_io_dirResult_bits_self_tag; // @[Slice.scala 94:16]
  wire [1:0] c_mshr_io_dirResult_bits_clients_states_0_state; // @[Slice.scala 94:16]
  wire  c_mshr_io_dirResult_bits_clients_states_0_hit; // @[Slice.scala 94:16]
  wire [1:0] c_mshr_io_dirResult_bits_clients_states_1_state; // @[Slice.scala 94:16]
  wire  c_mshr_io_dirResult_bits_clients_states_1_hit; // @[Slice.scala 94:16]
  wire [22:0] c_mshr_io_dirResult_bits_clients_tag; // @[Slice.scala 94:16]
  wire [3:0] c_mshr_io_dirResult_bits_clients_way; // @[Slice.scala 94:16]
  wire [9:0] c_mshr_io_c_status_set; // @[Slice.scala 94:16]
  wire [19:0] c_mshr_io_c_status_tag; // @[Slice.scala 94:16]
  wire [2:0] c_mshr_io_c_status_way; // @[Slice.scala 94:16]
  wire  c_mshr_io_c_status_nestedReleaseData; // @[Slice.scala 94:16]
  wire  c_mshr_io_c_status_releaseThrough; // @[Slice.scala 94:16]
  wire [9:0] c_mshr_io_bstatus_set; // @[Slice.scala 94:16]
  wire [19:0] c_mshr_io_bstatus_tag; // @[Slice.scala 94:16]
  wire [2:0] c_mshr_io_bstatus_way; // @[Slice.scala 94:16]
  wire  c_mshr_io_bstatus_nestedProbeAckData; // @[Slice.scala 94:16]
  wire  c_mshr_io_bstatus_probeHelperFinish; // @[Slice.scala 94:16]
  wire  c_mshr_io_bstatus_probeAckDataThrough; // @[Slice.scala 94:16]
  wire  c_mshr_io_releaseThrough; // @[Slice.scala 94:16]
  wire  c_mshr_io_probeAckDataThrough; // @[Slice.scala 94:16]
  wire  c_mshr_io_is_nestedReleaseData; // @[Slice.scala 94:16]
  wire  c_mshr_io_is_nestedProbeAckData; // @[Slice.scala 94:16]
  wire  c_mshr_io_probeHelperFinish; // @[Slice.scala 94:16]
  wire  dataStorage_clock; // @[Slice.scala 101:27]
  wire  dataStorage_reset; // @[Slice.scala 101:27]
  wire  dataStorage_io_sourceC_raddr_ready; // @[Slice.scala 101:27]
  wire  dataStorage_io_sourceC_raddr_valid; // @[Slice.scala 101:27]
  wire [2:0] dataStorage_io_sourceC_raddr_bits_way; // @[Slice.scala 101:27]
  wire [9:0] dataStorage_io_sourceC_raddr_bits_set; // @[Slice.scala 101:27]
  wire  dataStorage_io_sourceC_raddr_bits_beat; // @[Slice.scala 101:27]
  wire [255:0] dataStorage_io_sourceC_rdata_data; // @[Slice.scala 101:27]
  wire  dataStorage_io_sinkD_waddr_ready; // @[Slice.scala 101:27]
  wire  dataStorage_io_sinkD_waddr_valid; // @[Slice.scala 101:27]
  wire [2:0] dataStorage_io_sinkD_waddr_bits_way; // @[Slice.scala 101:27]
  wire [9:0] dataStorage_io_sinkD_waddr_bits_set; // @[Slice.scala 101:27]
  wire  dataStorage_io_sinkD_waddr_bits_beat; // @[Slice.scala 101:27]
  wire  dataStorage_io_sinkD_waddr_bits_noop; // @[Slice.scala 101:27]
  wire [255:0] dataStorage_io_sinkD_wdata_data; // @[Slice.scala 101:27]
  wire  dataStorage_io_sourceD_raddr_ready; // @[Slice.scala 101:27]
  wire  dataStorage_io_sourceD_raddr_valid; // @[Slice.scala 101:27]
  wire [2:0] dataStorage_io_sourceD_raddr_bits_way; // @[Slice.scala 101:27]
  wire [9:0] dataStorage_io_sourceD_raddr_bits_set; // @[Slice.scala 101:27]
  wire  dataStorage_io_sourceD_raddr_bits_beat; // @[Slice.scala 101:27]
  wire [255:0] dataStorage_io_sourceD_rdata_data; // @[Slice.scala 101:27]
  wire  dataStorage_io_sourceD_waddr_ready; // @[Slice.scala 101:27]
  wire  dataStorage_io_sourceD_waddr_valid; // @[Slice.scala 101:27]
  wire [2:0] dataStorage_io_sourceD_waddr_bits_way; // @[Slice.scala 101:27]
  wire [9:0] dataStorage_io_sourceD_waddr_bits_set; // @[Slice.scala 101:27]
  wire  dataStorage_io_sourceD_waddr_bits_beat; // @[Slice.scala 101:27]
  wire [255:0] dataStorage_io_sourceD_wdata_data; // @[Slice.scala 101:27]
  wire  dataStorage_io_sinkC_waddr_ready; // @[Slice.scala 101:27]
  wire  dataStorage_io_sinkC_waddr_valid; // @[Slice.scala 101:27]
  wire [2:0] dataStorage_io_sinkC_waddr_bits_way; // @[Slice.scala 101:27]
  wire [9:0] dataStorage_io_sinkC_waddr_bits_set; // @[Slice.scala 101:27]
  wire  dataStorage_io_sinkC_waddr_bits_beat; // @[Slice.scala 101:27]
  wire  dataStorage_io_sinkC_waddr_bits_noop; // @[Slice.scala 101:27]
  wire [255:0] dataStorage_io_sinkC_wdata_data; // @[Slice.scala 101:27]
  wire  mshrAlloc_io_a_req_ready; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_a_req_valid; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_a_req_bits_channel; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_a_req_bits_opcode; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_a_req_bits_param; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_a_req_bits_size; // @[Slice.scala 123:25]
  wire [5:0] mshrAlloc_io_a_req_bits_source; // @[Slice.scala 123:25]
  wire [9:0] mshrAlloc_io_a_req_bits_set; // @[Slice.scala 123:25]
  wire [19:0] mshrAlloc_io_a_req_bits_tag; // @[Slice.scala 123:25]
  wire [5:0] mshrAlloc_io_a_req_bits_off; // @[Slice.scala 123:25]
  wire [31:0] mshrAlloc_io_a_req_bits_mask; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_a_req_bits_bufIdx; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_a_req_bits_preferCache; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_a_req_bits_dirty; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_a_req_bits_fromProbeHelper; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_a_req_bits_fromCmoHelper; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_a_req_bits_needProbeAckData; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_breq_ready; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_breq_valid; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_breq_bits_channel; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_breq_bits_opcode; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_breq_bits_param; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_breq_bits_size; // @[Slice.scala 123:25]
  wire [5:0] mshrAlloc_io_breq_bits_source; // @[Slice.scala 123:25]
  wire [9:0] mshrAlloc_io_breq_bits_set; // @[Slice.scala 123:25]
  wire [19:0] mshrAlloc_io_breq_bits_tag; // @[Slice.scala 123:25]
  wire [5:0] mshrAlloc_io_breq_bits_off; // @[Slice.scala 123:25]
  wire [31:0] mshrAlloc_io_breq_bits_mask; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_breq_bits_bufIdx; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_breq_bits_preferCache; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_breq_bits_dirty; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_breq_bits_fromProbeHelper; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_breq_bits_fromCmoHelper; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_breq_bits_needProbeAckData; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_c_req_ready; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_c_req_valid; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_c_req_bits_opcode; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_c_req_bits_param; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_c_req_bits_size; // @[Slice.scala 123:25]
  wire [5:0] mshrAlloc_io_c_req_bits_source; // @[Slice.scala 123:25]
  wire [9:0] mshrAlloc_io_c_req_bits_set; // @[Slice.scala 123:25]
  wire [19:0] mshrAlloc_io_c_req_bits_tag; // @[Slice.scala 123:25]
  wire [5:0] mshrAlloc_io_c_req_bits_off; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_c_req_bits_bufIdx; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_c_req_bits_dirty; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_status_0_valid; // @[Slice.scala 123:25]
  wire [9:0] mshrAlloc_io_status_0_bits_set; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_status_0_bits_nestB; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_status_0_bits_nestC; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_status_1_valid; // @[Slice.scala 123:25]
  wire [9:0] mshrAlloc_io_status_1_bits_set; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_status_1_bits_nestB; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_status_1_bits_nestC; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_status_2_valid; // @[Slice.scala 123:25]
  wire [9:0] mshrAlloc_io_status_2_bits_set; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_status_2_bits_nestB; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_status_2_bits_nestC; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_status_3_valid; // @[Slice.scala 123:25]
  wire [9:0] mshrAlloc_io_status_3_bits_set; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_status_3_bits_nestB; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_status_3_bits_nestC; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_status_4_valid; // @[Slice.scala 123:25]
  wire [9:0] mshrAlloc_io_status_4_bits_set; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_status_4_bits_nestB; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_status_4_bits_nestC; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_status_5_valid; // @[Slice.scala 123:25]
  wire [9:0] mshrAlloc_io_status_5_bits_set; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_status_5_bits_nestB; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_status_5_bits_nestC; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_status_6_valid; // @[Slice.scala 123:25]
  wire [9:0] mshrAlloc_io_status_6_bits_set; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_status_6_bits_nestB; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_status_6_bits_nestC; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_status_7_valid; // @[Slice.scala 123:25]
  wire [9:0] mshrAlloc_io_status_7_bits_set; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_status_7_bits_nestB; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_status_7_bits_nestC; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_status_8_valid; // @[Slice.scala 123:25]
  wire [9:0] mshrAlloc_io_status_8_bits_set; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_status_8_bits_nestB; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_status_8_bits_nestC; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_status_9_valid; // @[Slice.scala 123:25]
  wire [9:0] mshrAlloc_io_status_9_bits_set; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_status_9_bits_nestB; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_status_9_bits_nestC; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_status_10_valid; // @[Slice.scala 123:25]
  wire [9:0] mshrAlloc_io_status_10_bits_set; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_status_10_bits_nestB; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_status_10_bits_nestC; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_status_11_valid; // @[Slice.scala 123:25]
  wire [9:0] mshrAlloc_io_status_11_bits_set; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_status_11_bits_nestB; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_status_11_bits_nestC; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_status_12_valid; // @[Slice.scala 123:25]
  wire [9:0] mshrAlloc_io_status_12_bits_set; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_status_12_bits_nestB; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_status_12_bits_nestC; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_status_13_valid; // @[Slice.scala 123:25]
  wire [9:0] mshrAlloc_io_status_13_bits_set; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_status_13_bits_nestB; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_status_13_bits_nestC; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_status_14_valid; // @[Slice.scala 123:25]
  wire [9:0] mshrAlloc_io_status_14_bits_set; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_status_14_bits_nestC; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_status_15_valid; // @[Slice.scala 123:25]
  wire [9:0] mshrAlloc_io_status_15_bits_set; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_0_valid; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_alloc_0_bits_channel; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_alloc_0_bits_opcode; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_alloc_0_bits_param; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_alloc_0_bits_size; // @[Slice.scala 123:25]
  wire [5:0] mshrAlloc_io_alloc_0_bits_source; // @[Slice.scala 123:25]
  wire [9:0] mshrAlloc_io_alloc_0_bits_set; // @[Slice.scala 123:25]
  wire [19:0] mshrAlloc_io_alloc_0_bits_tag; // @[Slice.scala 123:25]
  wire [5:0] mshrAlloc_io_alloc_0_bits_off; // @[Slice.scala 123:25]
  wire [31:0] mshrAlloc_io_alloc_0_bits_mask; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_alloc_0_bits_bufIdx; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_0_bits_preferCache; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_0_bits_dirty; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_0_bits_fromProbeHelper; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_0_bits_fromCmoHelper; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_0_bits_needProbeAckData; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_1_valid; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_alloc_1_bits_channel; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_alloc_1_bits_opcode; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_alloc_1_bits_param; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_alloc_1_bits_size; // @[Slice.scala 123:25]
  wire [5:0] mshrAlloc_io_alloc_1_bits_source; // @[Slice.scala 123:25]
  wire [9:0] mshrAlloc_io_alloc_1_bits_set; // @[Slice.scala 123:25]
  wire [19:0] mshrAlloc_io_alloc_1_bits_tag; // @[Slice.scala 123:25]
  wire [5:0] mshrAlloc_io_alloc_1_bits_off; // @[Slice.scala 123:25]
  wire [31:0] mshrAlloc_io_alloc_1_bits_mask; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_alloc_1_bits_bufIdx; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_1_bits_preferCache; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_1_bits_dirty; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_1_bits_fromProbeHelper; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_1_bits_fromCmoHelper; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_1_bits_needProbeAckData; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_2_valid; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_alloc_2_bits_channel; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_alloc_2_bits_opcode; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_alloc_2_bits_param; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_alloc_2_bits_size; // @[Slice.scala 123:25]
  wire [5:0] mshrAlloc_io_alloc_2_bits_source; // @[Slice.scala 123:25]
  wire [9:0] mshrAlloc_io_alloc_2_bits_set; // @[Slice.scala 123:25]
  wire [19:0] mshrAlloc_io_alloc_2_bits_tag; // @[Slice.scala 123:25]
  wire [5:0] mshrAlloc_io_alloc_2_bits_off; // @[Slice.scala 123:25]
  wire [31:0] mshrAlloc_io_alloc_2_bits_mask; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_alloc_2_bits_bufIdx; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_2_bits_preferCache; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_2_bits_dirty; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_2_bits_fromProbeHelper; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_2_bits_fromCmoHelper; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_2_bits_needProbeAckData; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_3_valid; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_alloc_3_bits_channel; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_alloc_3_bits_opcode; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_alloc_3_bits_param; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_alloc_3_bits_size; // @[Slice.scala 123:25]
  wire [5:0] mshrAlloc_io_alloc_3_bits_source; // @[Slice.scala 123:25]
  wire [9:0] mshrAlloc_io_alloc_3_bits_set; // @[Slice.scala 123:25]
  wire [19:0] mshrAlloc_io_alloc_3_bits_tag; // @[Slice.scala 123:25]
  wire [5:0] mshrAlloc_io_alloc_3_bits_off; // @[Slice.scala 123:25]
  wire [31:0] mshrAlloc_io_alloc_3_bits_mask; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_alloc_3_bits_bufIdx; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_3_bits_preferCache; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_3_bits_dirty; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_3_bits_fromProbeHelper; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_3_bits_fromCmoHelper; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_3_bits_needProbeAckData; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_4_valid; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_alloc_4_bits_channel; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_alloc_4_bits_opcode; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_alloc_4_bits_param; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_alloc_4_bits_size; // @[Slice.scala 123:25]
  wire [5:0] mshrAlloc_io_alloc_4_bits_source; // @[Slice.scala 123:25]
  wire [9:0] mshrAlloc_io_alloc_4_bits_set; // @[Slice.scala 123:25]
  wire [19:0] mshrAlloc_io_alloc_4_bits_tag; // @[Slice.scala 123:25]
  wire [5:0] mshrAlloc_io_alloc_4_bits_off; // @[Slice.scala 123:25]
  wire [31:0] mshrAlloc_io_alloc_4_bits_mask; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_alloc_4_bits_bufIdx; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_4_bits_preferCache; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_4_bits_dirty; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_4_bits_fromProbeHelper; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_4_bits_fromCmoHelper; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_4_bits_needProbeAckData; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_5_valid; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_alloc_5_bits_channel; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_alloc_5_bits_opcode; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_alloc_5_bits_param; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_alloc_5_bits_size; // @[Slice.scala 123:25]
  wire [5:0] mshrAlloc_io_alloc_5_bits_source; // @[Slice.scala 123:25]
  wire [9:0] mshrAlloc_io_alloc_5_bits_set; // @[Slice.scala 123:25]
  wire [19:0] mshrAlloc_io_alloc_5_bits_tag; // @[Slice.scala 123:25]
  wire [5:0] mshrAlloc_io_alloc_5_bits_off; // @[Slice.scala 123:25]
  wire [31:0] mshrAlloc_io_alloc_5_bits_mask; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_alloc_5_bits_bufIdx; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_5_bits_preferCache; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_5_bits_dirty; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_5_bits_fromProbeHelper; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_5_bits_fromCmoHelper; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_5_bits_needProbeAckData; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_6_valid; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_alloc_6_bits_channel; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_alloc_6_bits_opcode; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_alloc_6_bits_param; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_alloc_6_bits_size; // @[Slice.scala 123:25]
  wire [5:0] mshrAlloc_io_alloc_6_bits_source; // @[Slice.scala 123:25]
  wire [9:0] mshrAlloc_io_alloc_6_bits_set; // @[Slice.scala 123:25]
  wire [19:0] mshrAlloc_io_alloc_6_bits_tag; // @[Slice.scala 123:25]
  wire [5:0] mshrAlloc_io_alloc_6_bits_off; // @[Slice.scala 123:25]
  wire [31:0] mshrAlloc_io_alloc_6_bits_mask; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_alloc_6_bits_bufIdx; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_6_bits_preferCache; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_6_bits_dirty; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_6_bits_fromProbeHelper; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_6_bits_fromCmoHelper; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_6_bits_needProbeAckData; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_7_valid; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_alloc_7_bits_channel; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_alloc_7_bits_opcode; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_alloc_7_bits_param; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_alloc_7_bits_size; // @[Slice.scala 123:25]
  wire [5:0] mshrAlloc_io_alloc_7_bits_source; // @[Slice.scala 123:25]
  wire [9:0] mshrAlloc_io_alloc_7_bits_set; // @[Slice.scala 123:25]
  wire [19:0] mshrAlloc_io_alloc_7_bits_tag; // @[Slice.scala 123:25]
  wire [5:0] mshrAlloc_io_alloc_7_bits_off; // @[Slice.scala 123:25]
  wire [31:0] mshrAlloc_io_alloc_7_bits_mask; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_alloc_7_bits_bufIdx; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_7_bits_preferCache; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_7_bits_dirty; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_7_bits_fromProbeHelper; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_7_bits_fromCmoHelper; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_7_bits_needProbeAckData; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_8_valid; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_alloc_8_bits_channel; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_alloc_8_bits_opcode; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_alloc_8_bits_param; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_alloc_8_bits_size; // @[Slice.scala 123:25]
  wire [5:0] mshrAlloc_io_alloc_8_bits_source; // @[Slice.scala 123:25]
  wire [9:0] mshrAlloc_io_alloc_8_bits_set; // @[Slice.scala 123:25]
  wire [19:0] mshrAlloc_io_alloc_8_bits_tag; // @[Slice.scala 123:25]
  wire [5:0] mshrAlloc_io_alloc_8_bits_off; // @[Slice.scala 123:25]
  wire [31:0] mshrAlloc_io_alloc_8_bits_mask; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_alloc_8_bits_bufIdx; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_8_bits_preferCache; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_8_bits_dirty; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_8_bits_fromProbeHelper; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_8_bits_fromCmoHelper; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_8_bits_needProbeAckData; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_9_valid; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_alloc_9_bits_channel; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_alloc_9_bits_opcode; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_alloc_9_bits_param; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_alloc_9_bits_size; // @[Slice.scala 123:25]
  wire [5:0] mshrAlloc_io_alloc_9_bits_source; // @[Slice.scala 123:25]
  wire [9:0] mshrAlloc_io_alloc_9_bits_set; // @[Slice.scala 123:25]
  wire [19:0] mshrAlloc_io_alloc_9_bits_tag; // @[Slice.scala 123:25]
  wire [5:0] mshrAlloc_io_alloc_9_bits_off; // @[Slice.scala 123:25]
  wire [31:0] mshrAlloc_io_alloc_9_bits_mask; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_alloc_9_bits_bufIdx; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_9_bits_preferCache; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_9_bits_dirty; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_9_bits_fromProbeHelper; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_9_bits_fromCmoHelper; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_9_bits_needProbeAckData; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_10_valid; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_alloc_10_bits_channel; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_alloc_10_bits_opcode; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_alloc_10_bits_param; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_alloc_10_bits_size; // @[Slice.scala 123:25]
  wire [5:0] mshrAlloc_io_alloc_10_bits_source; // @[Slice.scala 123:25]
  wire [9:0] mshrAlloc_io_alloc_10_bits_set; // @[Slice.scala 123:25]
  wire [19:0] mshrAlloc_io_alloc_10_bits_tag; // @[Slice.scala 123:25]
  wire [5:0] mshrAlloc_io_alloc_10_bits_off; // @[Slice.scala 123:25]
  wire [31:0] mshrAlloc_io_alloc_10_bits_mask; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_alloc_10_bits_bufIdx; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_10_bits_preferCache; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_10_bits_dirty; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_10_bits_fromProbeHelper; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_10_bits_fromCmoHelper; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_10_bits_needProbeAckData; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_11_valid; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_alloc_11_bits_channel; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_alloc_11_bits_opcode; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_alloc_11_bits_param; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_alloc_11_bits_size; // @[Slice.scala 123:25]
  wire [5:0] mshrAlloc_io_alloc_11_bits_source; // @[Slice.scala 123:25]
  wire [9:0] mshrAlloc_io_alloc_11_bits_set; // @[Slice.scala 123:25]
  wire [19:0] mshrAlloc_io_alloc_11_bits_tag; // @[Slice.scala 123:25]
  wire [5:0] mshrAlloc_io_alloc_11_bits_off; // @[Slice.scala 123:25]
  wire [31:0] mshrAlloc_io_alloc_11_bits_mask; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_alloc_11_bits_bufIdx; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_11_bits_preferCache; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_11_bits_dirty; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_11_bits_fromProbeHelper; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_11_bits_fromCmoHelper; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_11_bits_needProbeAckData; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_12_valid; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_alloc_12_bits_channel; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_alloc_12_bits_opcode; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_alloc_12_bits_param; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_alloc_12_bits_size; // @[Slice.scala 123:25]
  wire [5:0] mshrAlloc_io_alloc_12_bits_source; // @[Slice.scala 123:25]
  wire [9:0] mshrAlloc_io_alloc_12_bits_set; // @[Slice.scala 123:25]
  wire [19:0] mshrAlloc_io_alloc_12_bits_tag; // @[Slice.scala 123:25]
  wire [5:0] mshrAlloc_io_alloc_12_bits_off; // @[Slice.scala 123:25]
  wire [31:0] mshrAlloc_io_alloc_12_bits_mask; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_alloc_12_bits_bufIdx; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_12_bits_preferCache; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_12_bits_dirty; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_12_bits_fromProbeHelper; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_12_bits_fromCmoHelper; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_12_bits_needProbeAckData; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_13_valid; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_alloc_13_bits_channel; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_alloc_13_bits_opcode; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_alloc_13_bits_param; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_alloc_13_bits_size; // @[Slice.scala 123:25]
  wire [5:0] mshrAlloc_io_alloc_13_bits_source; // @[Slice.scala 123:25]
  wire [9:0] mshrAlloc_io_alloc_13_bits_set; // @[Slice.scala 123:25]
  wire [19:0] mshrAlloc_io_alloc_13_bits_tag; // @[Slice.scala 123:25]
  wire [5:0] mshrAlloc_io_alloc_13_bits_off; // @[Slice.scala 123:25]
  wire [31:0] mshrAlloc_io_alloc_13_bits_mask; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_alloc_13_bits_bufIdx; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_13_bits_preferCache; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_13_bits_dirty; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_13_bits_fromProbeHelper; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_13_bits_fromCmoHelper; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_13_bits_needProbeAckData; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_14_valid; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_alloc_14_bits_channel; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_alloc_14_bits_opcode; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_alloc_14_bits_param; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_alloc_14_bits_size; // @[Slice.scala 123:25]
  wire [5:0] mshrAlloc_io_alloc_14_bits_source; // @[Slice.scala 123:25]
  wire [9:0] mshrAlloc_io_alloc_14_bits_set; // @[Slice.scala 123:25]
  wire [19:0] mshrAlloc_io_alloc_14_bits_tag; // @[Slice.scala 123:25]
  wire [5:0] mshrAlloc_io_alloc_14_bits_off; // @[Slice.scala 123:25]
  wire [31:0] mshrAlloc_io_alloc_14_bits_mask; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_alloc_14_bits_bufIdx; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_14_bits_preferCache; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_14_bits_dirty; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_14_bits_fromProbeHelper; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_14_bits_fromCmoHelper; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_14_bits_needProbeAckData; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_15_valid; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_alloc_15_bits_opcode; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_alloc_15_bits_param; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_alloc_15_bits_size; // @[Slice.scala 123:25]
  wire [5:0] mshrAlloc_io_alloc_15_bits_source; // @[Slice.scala 123:25]
  wire [9:0] mshrAlloc_io_alloc_15_bits_set; // @[Slice.scala 123:25]
  wire [19:0] mshrAlloc_io_alloc_15_bits_tag; // @[Slice.scala 123:25]
  wire [5:0] mshrAlloc_io_alloc_15_bits_off; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_alloc_15_bits_bufIdx; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_alloc_15_bits_dirty; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_dirRead_ready; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_dirRead_valid; // @[Slice.scala 123:25]
  wire [15:0] mshrAlloc_io_dirRead_bits_idOH; // @[Slice.scala 123:25]
  wire [19:0] mshrAlloc_io_dirRead_bits_tag; // @[Slice.scala 123:25]
  wire [9:0] mshrAlloc_io_dirRead_bits_set; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_dirRead_bits_replacerInfo_channel; // @[Slice.scala 123:25]
  wire [2:0] mshrAlloc_io_dirRead_bits_replacerInfo_opcode; // @[Slice.scala 123:25]
  wire [5:0] mshrAlloc_io_dirRead_bits_source; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_bc_mask_valid; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_bc_mask_bits_0; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_bc_mask_bits_1; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_bc_mask_bits_2; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_bc_mask_bits_3; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_bc_mask_bits_4; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_bc_mask_bits_5; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_bc_mask_bits_6; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_bc_mask_bits_7; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_bc_mask_bits_8; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_bc_mask_bits_9; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_bc_mask_bits_10; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_bc_mask_bits_11; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_bc_mask_bits_12; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_bc_mask_bits_13; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_c_mask_valid; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_c_mask_bits_0; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_c_mask_bits_1; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_c_mask_bits_2; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_c_mask_bits_3; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_c_mask_bits_4; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_c_mask_bits_5; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_c_mask_bits_6; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_c_mask_bits_7; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_c_mask_bits_8; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_c_mask_bits_9; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_c_mask_bits_10; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_c_mask_bits_11; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_c_mask_bits_12; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_c_mask_bits_13; // @[Slice.scala 123:25]
  wire  mshrAlloc_io_c_mask_bits_14; // @[Slice.scala 123:25]
  wire  a_req_buffer_clock; // @[Slice.scala 124:28]
  wire  a_req_buffer_reset; // @[Slice.scala 124:28]
  wire  a_req_buffer_io_in_ready; // @[Slice.scala 124:28]
  wire  a_req_buffer_io_in_valid; // @[Slice.scala 124:28]
  wire [2:0] a_req_buffer_io_in_bits_opcode; // @[Slice.scala 124:28]
  wire [2:0] a_req_buffer_io_in_bits_param; // @[Slice.scala 124:28]
  wire [2:0] a_req_buffer_io_in_bits_size; // @[Slice.scala 124:28]
  wire [5:0] a_req_buffer_io_in_bits_source; // @[Slice.scala 124:28]
  wire [9:0] a_req_buffer_io_in_bits_set; // @[Slice.scala 124:28]
  wire [19:0] a_req_buffer_io_in_bits_tag; // @[Slice.scala 124:28]
  wire [5:0] a_req_buffer_io_in_bits_off; // @[Slice.scala 124:28]
  wire [31:0] a_req_buffer_io_in_bits_mask; // @[Slice.scala 124:28]
  wire [2:0] a_req_buffer_io_in_bits_bufIdx; // @[Slice.scala 124:28]
  wire  a_req_buffer_io_in_bits_preferCache; // @[Slice.scala 124:28]
  wire  a_req_buffer_io_out_ready; // @[Slice.scala 124:28]
  wire  a_req_buffer_io_out_valid; // @[Slice.scala 124:28]
  wire [2:0] a_req_buffer_io_out_bits_channel; // @[Slice.scala 124:28]
  wire [2:0] a_req_buffer_io_out_bits_opcode; // @[Slice.scala 124:28]
  wire [2:0] a_req_buffer_io_out_bits_param; // @[Slice.scala 124:28]
  wire [2:0] a_req_buffer_io_out_bits_size; // @[Slice.scala 124:28]
  wire [5:0] a_req_buffer_io_out_bits_source; // @[Slice.scala 124:28]
  wire [9:0] a_req_buffer_io_out_bits_set; // @[Slice.scala 124:28]
  wire [19:0] a_req_buffer_io_out_bits_tag; // @[Slice.scala 124:28]
  wire [5:0] a_req_buffer_io_out_bits_off; // @[Slice.scala 124:28]
  wire [31:0] a_req_buffer_io_out_bits_mask; // @[Slice.scala 124:28]
  wire [2:0] a_req_buffer_io_out_bits_bufIdx; // @[Slice.scala 124:28]
  wire  a_req_buffer_io_out_bits_preferCache; // @[Slice.scala 124:28]
  wire  a_req_buffer_io_out_bits_dirty; // @[Slice.scala 124:28]
  wire  a_req_buffer_io_out_bits_fromProbeHelper; // @[Slice.scala 124:28]
  wire  a_req_buffer_io_out_bits_fromCmoHelper; // @[Slice.scala 124:28]
  wire  a_req_buffer_io_out_bits_needProbeAckData; // @[Slice.scala 124:28]
  wire  a_req_buffer_io_mshr_status_0_valid; // @[Slice.scala 124:28]
  wire [9:0] a_req_buffer_io_mshr_status_0_bits_set; // @[Slice.scala 124:28]
  wire  a_req_buffer_io_mshr_status_0_bits_will_free; // @[Slice.scala 124:28]
  wire  a_req_buffer_io_mshr_status_1_valid; // @[Slice.scala 124:28]
  wire [9:0] a_req_buffer_io_mshr_status_1_bits_set; // @[Slice.scala 124:28]
  wire  a_req_buffer_io_mshr_status_1_bits_will_free; // @[Slice.scala 124:28]
  wire  a_req_buffer_io_mshr_status_2_valid; // @[Slice.scala 124:28]
  wire [9:0] a_req_buffer_io_mshr_status_2_bits_set; // @[Slice.scala 124:28]
  wire  a_req_buffer_io_mshr_status_2_bits_will_free; // @[Slice.scala 124:28]
  wire  a_req_buffer_io_mshr_status_3_valid; // @[Slice.scala 124:28]
  wire [9:0] a_req_buffer_io_mshr_status_3_bits_set; // @[Slice.scala 124:28]
  wire  a_req_buffer_io_mshr_status_3_bits_will_free; // @[Slice.scala 124:28]
  wire  a_req_buffer_io_mshr_status_4_valid; // @[Slice.scala 124:28]
  wire [9:0] a_req_buffer_io_mshr_status_4_bits_set; // @[Slice.scala 124:28]
  wire  a_req_buffer_io_mshr_status_4_bits_will_free; // @[Slice.scala 124:28]
  wire  a_req_buffer_io_mshr_status_5_valid; // @[Slice.scala 124:28]
  wire [9:0] a_req_buffer_io_mshr_status_5_bits_set; // @[Slice.scala 124:28]
  wire  a_req_buffer_io_mshr_status_5_bits_will_free; // @[Slice.scala 124:28]
  wire  a_req_buffer_io_mshr_status_6_valid; // @[Slice.scala 124:28]
  wire [9:0] a_req_buffer_io_mshr_status_6_bits_set; // @[Slice.scala 124:28]
  wire  a_req_buffer_io_mshr_status_6_bits_will_free; // @[Slice.scala 124:28]
  wire  a_req_buffer_io_mshr_status_7_valid; // @[Slice.scala 124:28]
  wire [9:0] a_req_buffer_io_mshr_status_7_bits_set; // @[Slice.scala 124:28]
  wire  a_req_buffer_io_mshr_status_7_bits_will_free; // @[Slice.scala 124:28]
  wire  a_req_buffer_io_mshr_status_8_valid; // @[Slice.scala 124:28]
  wire [9:0] a_req_buffer_io_mshr_status_8_bits_set; // @[Slice.scala 124:28]
  wire  a_req_buffer_io_mshr_status_8_bits_will_free; // @[Slice.scala 124:28]
  wire  a_req_buffer_io_mshr_status_9_valid; // @[Slice.scala 124:28]
  wire [9:0] a_req_buffer_io_mshr_status_9_bits_set; // @[Slice.scala 124:28]
  wire  a_req_buffer_io_mshr_status_9_bits_will_free; // @[Slice.scala 124:28]
  wire  a_req_buffer_io_mshr_status_10_valid; // @[Slice.scala 124:28]
  wire [9:0] a_req_buffer_io_mshr_status_10_bits_set; // @[Slice.scala 124:28]
  wire  a_req_buffer_io_mshr_status_10_bits_will_free; // @[Slice.scala 124:28]
  wire  a_req_buffer_io_mshr_status_11_valid; // @[Slice.scala 124:28]
  wire [9:0] a_req_buffer_io_mshr_status_11_bits_set; // @[Slice.scala 124:28]
  wire  a_req_buffer_io_mshr_status_11_bits_will_free; // @[Slice.scala 124:28]
  wire  a_req_buffer_io_mshr_status_12_valid; // @[Slice.scala 124:28]
  wire [9:0] a_req_buffer_io_mshr_status_12_bits_set; // @[Slice.scala 124:28]
  wire  a_req_buffer_io_mshr_status_12_bits_will_free; // @[Slice.scala 124:28]
  wire  a_req_buffer_io_mshr_status_13_valid; // @[Slice.scala 124:28]
  wire [9:0] a_req_buffer_io_mshr_status_13_bits_set; // @[Slice.scala 124:28]
  wire  a_req_buffer_io_mshr_status_13_bits_will_free; // @[Slice.scala 124:28]
  wire  probeHelperOpt_clock; // @[Slice.scala 126:16]
  wire  probeHelperOpt_reset; // @[Slice.scala 126:16]
  wire  probeHelperOpt_io_dirResult_valid; // @[Slice.scala 126:16]
  wire [1:0] probeHelperOpt_io_dirResult_bits_clients_states_0_state; // @[Slice.scala 126:16]
  wire  probeHelperOpt_io_dirResult_bits_clients_states_0_hit; // @[Slice.scala 126:16]
  wire [1:0] probeHelperOpt_io_dirResult_bits_clients_states_1_state; // @[Slice.scala 126:16]
  wire  probeHelperOpt_io_dirResult_bits_clients_states_1_hit; // @[Slice.scala 126:16]
  wire  probeHelperOpt_io_dirResult_bits_clients_tag_match; // @[Slice.scala 126:16]
  wire [22:0] probeHelperOpt_io_dirResult_bits_clients_tag; // @[Slice.scala 126:16]
  wire [5:0] probeHelperOpt_io_dirResult_bits_sourceId; // @[Slice.scala 126:16]
  wire [9:0] probeHelperOpt_io_dirResult_bits_set; // @[Slice.scala 126:16]
  wire [2:0] probeHelperOpt_io_dirResult_bits_replacerInfo_channel; // @[Slice.scala 126:16]
  wire [2:0] probeHelperOpt_io_dirResult_bits_replacerInfo_opcode; // @[Slice.scala 126:16]
  wire  probeHelperOpt_io_probe_ready; // @[Slice.scala 126:16]
  wire  probeHelperOpt_io_probe_valid; // @[Slice.scala 126:16]
  wire [2:0] probeHelperOpt_io_probe_bits_channel; // @[Slice.scala 126:16]
  wire [2:0] probeHelperOpt_io_probe_bits_opcode; // @[Slice.scala 126:16]
  wire [2:0] probeHelperOpt_io_probe_bits_param; // @[Slice.scala 126:16]
  wire [2:0] probeHelperOpt_io_probe_bits_size; // @[Slice.scala 126:16]
  wire [5:0] probeHelperOpt_io_probe_bits_source; // @[Slice.scala 126:16]
  wire [9:0] probeHelperOpt_io_probe_bits_set; // @[Slice.scala 126:16]
  wire [19:0] probeHelperOpt_io_probe_bits_tag; // @[Slice.scala 126:16]
  wire [5:0] probeHelperOpt_io_probe_bits_off; // @[Slice.scala 126:16]
  wire [31:0] probeHelperOpt_io_probe_bits_mask; // @[Slice.scala 126:16]
  wire [2:0] probeHelperOpt_io_probe_bits_bufIdx; // @[Slice.scala 126:16]
  wire  probeHelperOpt_io_probe_bits_preferCache; // @[Slice.scala 126:16]
  wire  probeHelperOpt_io_probe_bits_dirty; // @[Slice.scala 126:16]
  wire  probeHelperOpt_io_probe_bits_fromProbeHelper; // @[Slice.scala 126:16]
  wire  probeHelperOpt_io_probe_bits_fromCmoHelper; // @[Slice.scala 126:16]
  wire  probeHelperOpt_io_probe_bits_needProbeAckData; // @[Slice.scala 126:16]
  wire  probeHelperOpt_io_full; // @[Slice.scala 126:16]
  wire  b_arb_io_in_0_ready; // @[Slice.scala 136:23]
  wire  b_arb_io_in_0_valid; // @[Slice.scala 136:23]
  wire [2:0] b_arb_io_in_0_bits_channel; // @[Slice.scala 136:23]
  wire [2:0] b_arb_io_in_0_bits_opcode; // @[Slice.scala 136:23]
  wire [2:0] b_arb_io_in_0_bits_param; // @[Slice.scala 136:23]
  wire [2:0] b_arb_io_in_0_bits_size; // @[Slice.scala 136:23]
  wire [5:0] b_arb_io_in_0_bits_source; // @[Slice.scala 136:23]
  wire [9:0] b_arb_io_in_0_bits_set; // @[Slice.scala 136:23]
  wire [19:0] b_arb_io_in_0_bits_tag; // @[Slice.scala 136:23]
  wire [5:0] b_arb_io_in_0_bits_off; // @[Slice.scala 136:23]
  wire [31:0] b_arb_io_in_0_bits_mask; // @[Slice.scala 136:23]
  wire [2:0] b_arb_io_in_0_bits_bufIdx; // @[Slice.scala 136:23]
  wire  b_arb_io_in_0_bits_preferCache; // @[Slice.scala 136:23]
  wire  b_arb_io_in_0_bits_dirty; // @[Slice.scala 136:23]
  wire  b_arb_io_in_0_bits_fromProbeHelper; // @[Slice.scala 136:23]
  wire  b_arb_io_in_0_bits_fromCmoHelper; // @[Slice.scala 136:23]
  wire  b_arb_io_in_0_bits_needProbeAckData; // @[Slice.scala 136:23]
  wire  b_arb_io_in_1_ready; // @[Slice.scala 136:23]
  wire  b_arb_io_in_1_valid; // @[Slice.scala 136:23]
  wire [2:0] b_arb_io_in_1_bits_opcode; // @[Slice.scala 136:23]
  wire [2:0] b_arb_io_in_1_bits_param; // @[Slice.scala 136:23]
  wire [2:0] b_arb_io_in_1_bits_size; // @[Slice.scala 136:23]
  wire [5:0] b_arb_io_in_1_bits_source; // @[Slice.scala 136:23]
  wire [9:0] b_arb_io_in_1_bits_set; // @[Slice.scala 136:23]
  wire [19:0] b_arb_io_in_1_bits_tag; // @[Slice.scala 136:23]
  wire [5:0] b_arb_io_in_1_bits_off; // @[Slice.scala 136:23]
  wire [31:0] b_arb_io_in_1_bits_mask; // @[Slice.scala 136:23]
  wire  b_arb_io_in_1_bits_needProbeAckData; // @[Slice.scala 136:23]
  wire  b_arb_io_out_ready; // @[Slice.scala 136:23]
  wire  b_arb_io_out_valid; // @[Slice.scala 136:23]
  wire [2:0] b_arb_io_out_bits_channel; // @[Slice.scala 136:23]
  wire [2:0] b_arb_io_out_bits_opcode; // @[Slice.scala 136:23]
  wire [2:0] b_arb_io_out_bits_param; // @[Slice.scala 136:23]
  wire [2:0] b_arb_io_out_bits_size; // @[Slice.scala 136:23]
  wire [5:0] b_arb_io_out_bits_source; // @[Slice.scala 136:23]
  wire [9:0] b_arb_io_out_bits_set; // @[Slice.scala 136:23]
  wire [19:0] b_arb_io_out_bits_tag; // @[Slice.scala 136:23]
  wire [5:0] b_arb_io_out_bits_off; // @[Slice.scala 136:23]
  wire [31:0] b_arb_io_out_bits_mask; // @[Slice.scala 136:23]
  wire [2:0] b_arb_io_out_bits_bufIdx; // @[Slice.scala 136:23]
  wire  b_arb_io_out_bits_preferCache; // @[Slice.scala 136:23]
  wire  b_arb_io_out_bits_dirty; // @[Slice.scala 136:23]
  wire  b_arb_io_out_bits_fromProbeHelper; // @[Slice.scala 136:23]
  wire  b_arb_io_out_bits_fromCmoHelper; // @[Slice.scala 136:23]
  wire  b_arb_io_out_bits_needProbeAckData; // @[Slice.scala 136:23]
  wire  directory_clock; // @[Slice.scala 372:25]
  wire  directory_reset; // @[Slice.scala 372:25]
  wire  directory_io_read_ready; // @[Slice.scala 372:25]
  wire  directory_io_read_valid; // @[Slice.scala 372:25]
  wire [15:0] directory_io_read_bits_idOH; // @[Slice.scala 372:25]
  wire [19:0] directory_io_read_bits_tag; // @[Slice.scala 372:25]
  wire [9:0] directory_io_read_bits_set; // @[Slice.scala 372:25]
  wire [2:0] directory_io_read_bits_replacerInfo_channel; // @[Slice.scala 372:25]
  wire [2:0] directory_io_read_bits_replacerInfo_opcode; // @[Slice.scala 372:25]
  wire [5:0] directory_io_read_bits_source; // @[Slice.scala 372:25]
  wire  directory_io_result_valid; // @[Slice.scala 372:25]
  wire [15:0] directory_io_result_bits_idOH; // @[Slice.scala 372:25]
  wire  directory_io_result_bits_self_dirty; // @[Slice.scala 372:25]
  wire [1:0] directory_io_result_bits_self_state; // @[Slice.scala 372:25]
  wire [1:0] directory_io_result_bits_self_clientStates_0; // @[Slice.scala 372:25]
  wire [1:0] directory_io_result_bits_self_clientStates_1; // @[Slice.scala 372:25]
  wire  directory_io_result_bits_self_hit; // @[Slice.scala 372:25]
  wire [2:0] directory_io_result_bits_self_way; // @[Slice.scala 372:25]
  wire [19:0] directory_io_result_bits_self_tag; // @[Slice.scala 372:25]
  wire [1:0] directory_io_result_bits_clients_states_0_state; // @[Slice.scala 372:25]
  wire  directory_io_result_bits_clients_states_0_hit; // @[Slice.scala 372:25]
  wire [1:0] directory_io_result_bits_clients_states_1_state; // @[Slice.scala 372:25]
  wire  directory_io_result_bits_clients_states_1_hit; // @[Slice.scala 372:25]
  wire  directory_io_result_bits_clients_tag_match; // @[Slice.scala 372:25]
  wire [22:0] directory_io_result_bits_clients_tag; // @[Slice.scala 372:25]
  wire [3:0] directory_io_result_bits_clients_way; // @[Slice.scala 372:25]
  wire [5:0] directory_io_result_bits_sourceId; // @[Slice.scala 372:25]
  wire [9:0] directory_io_result_bits_set; // @[Slice.scala 372:25]
  wire [2:0] directory_io_result_bits_replacerInfo_channel; // @[Slice.scala 372:25]
  wire [2:0] directory_io_result_bits_replacerInfo_opcode; // @[Slice.scala 372:25]
  wire  directory_io_dirWReq_valid; // @[Slice.scala 372:25]
  wire [9:0] directory_io_dirWReq_bits_set; // @[Slice.scala 372:25]
  wire [2:0] directory_io_dirWReq_bits_way; // @[Slice.scala 372:25]
  wire  directory_io_dirWReq_bits_data_dirty; // @[Slice.scala 372:25]
  wire [1:0] directory_io_dirWReq_bits_data_state; // @[Slice.scala 372:25]
  wire [1:0] directory_io_dirWReq_bits_data_clientStates_0; // @[Slice.scala 372:25]
  wire [1:0] directory_io_dirWReq_bits_data_clientStates_1; // @[Slice.scala 372:25]
  wire  directory_io_tagWReq_valid; // @[Slice.scala 372:25]
  wire [9:0] directory_io_tagWReq_bits_set; // @[Slice.scala 372:25]
  wire [2:0] directory_io_tagWReq_bits_way; // @[Slice.scala 372:25]
  wire [19:0] directory_io_tagWReq_bits_tag; // @[Slice.scala 372:25]
  wire  directory_io_clientDirWReq_valid; // @[Slice.scala 372:25]
  wire [6:0] directory_io_clientDirWReq_bits_set; // @[Slice.scala 372:25]
  wire [3:0] directory_io_clientDirWReq_bits_way; // @[Slice.scala 372:25]
  wire [1:0] directory_io_clientDirWReq_bits_data_0_state; // @[Slice.scala 372:25]
  wire [1:0] directory_io_clientDirWReq_bits_data_1_state; // @[Slice.scala 372:25]
  wire  directory_io_clientTagWreq_valid; // @[Slice.scala 372:25]
  wire [6:0] directory_io_clientTagWreq_bits_set; // @[Slice.scala 372:25]
  wire [3:0] directory_io_clientTagWreq_bits_way; // @[Slice.scala 372:25]
  wire [22:0] directory_io_clientTagWreq_bits_tag; // @[Slice.scala 372:25]
  wire  pipeline_clock; // @[Pipeline.scala 39:26]
  wire  pipeline_reset; // @[Pipeline.scala 39:26]
  wire  pipeline_io_in_valid; // @[Pipeline.scala 39:26]
  wire [9:0] pipeline_io_in_bits_set; // @[Pipeline.scala 39:26]
  wire [2:0] pipeline_io_in_bits_way; // @[Pipeline.scala 39:26]
  wire  pipeline_io_in_bits_data_dirty; // @[Pipeline.scala 39:26]
  wire [1:0] pipeline_io_in_bits_data_state; // @[Pipeline.scala 39:26]
  wire [1:0] pipeline_io_in_bits_data_clientStates_0; // @[Pipeline.scala 39:26]
  wire [1:0] pipeline_io_in_bits_data_clientStates_1; // @[Pipeline.scala 39:26]
  wire  pipeline_io_out_valid; // @[Pipeline.scala 39:26]
  wire [9:0] pipeline_io_out_bits_set; // @[Pipeline.scala 39:26]
  wire [2:0] pipeline_io_out_bits_way; // @[Pipeline.scala 39:26]
  wire  pipeline_io_out_bits_data_dirty; // @[Pipeline.scala 39:26]
  wire [1:0] pipeline_io_out_bits_data_state; // @[Pipeline.scala 39:26]
  wire [1:0] pipeline_io_out_bits_data_clientStates_0; // @[Pipeline.scala 39:26]
  wire [1:0] pipeline_io_out_bits_data_clientStates_1; // @[Pipeline.scala 39:26]
  wire  arbiter_clock; // @[Slice.scala 405:25]
  wire  arbiter_reset; // @[Slice.scala 405:25]
  wire  arbiter_io_in_0_ready; // @[Slice.scala 405:25]
  wire  arbiter_io_in_0_valid; // @[Slice.scala 405:25]
  wire [9:0] arbiter_io_in_0_bits_set; // @[Slice.scala 405:25]
  wire [2:0] arbiter_io_in_0_bits_way; // @[Slice.scala 405:25]
  wire  arbiter_io_in_0_bits_data_dirty; // @[Slice.scala 405:25]
  wire [1:0] arbiter_io_in_0_bits_data_state; // @[Slice.scala 405:25]
  wire [1:0] arbiter_io_in_0_bits_data_clientStates_0; // @[Slice.scala 405:25]
  wire [1:0] arbiter_io_in_0_bits_data_clientStates_1; // @[Slice.scala 405:25]
  wire  arbiter_io_in_1_ready; // @[Slice.scala 405:25]
  wire  arbiter_io_in_1_valid; // @[Slice.scala 405:25]
  wire [9:0] arbiter_io_in_1_bits_set; // @[Slice.scala 405:25]
  wire [2:0] arbiter_io_in_1_bits_way; // @[Slice.scala 405:25]
  wire  arbiter_io_in_1_bits_data_dirty; // @[Slice.scala 405:25]
  wire [1:0] arbiter_io_in_1_bits_data_state; // @[Slice.scala 405:25]
  wire [1:0] arbiter_io_in_1_bits_data_clientStates_0; // @[Slice.scala 405:25]
  wire [1:0] arbiter_io_in_1_bits_data_clientStates_1; // @[Slice.scala 405:25]
  wire  arbiter_io_in_2_ready; // @[Slice.scala 405:25]
  wire  arbiter_io_in_2_valid; // @[Slice.scala 405:25]
  wire [9:0] arbiter_io_in_2_bits_set; // @[Slice.scala 405:25]
  wire [2:0] arbiter_io_in_2_bits_way; // @[Slice.scala 405:25]
  wire  arbiter_io_in_2_bits_data_dirty; // @[Slice.scala 405:25]
  wire [1:0] arbiter_io_in_2_bits_data_state; // @[Slice.scala 405:25]
  wire [1:0] arbiter_io_in_2_bits_data_clientStates_0; // @[Slice.scala 405:25]
  wire [1:0] arbiter_io_in_2_bits_data_clientStates_1; // @[Slice.scala 405:25]
  wire  arbiter_io_in_3_ready; // @[Slice.scala 405:25]
  wire  arbiter_io_in_3_valid; // @[Slice.scala 405:25]
  wire [9:0] arbiter_io_in_3_bits_set; // @[Slice.scala 405:25]
  wire [2:0] arbiter_io_in_3_bits_way; // @[Slice.scala 405:25]
  wire  arbiter_io_in_3_bits_data_dirty; // @[Slice.scala 405:25]
  wire [1:0] arbiter_io_in_3_bits_data_state; // @[Slice.scala 405:25]
  wire [1:0] arbiter_io_in_3_bits_data_clientStates_0; // @[Slice.scala 405:25]
  wire [1:0] arbiter_io_in_3_bits_data_clientStates_1; // @[Slice.scala 405:25]
  wire  arbiter_io_in_4_ready; // @[Slice.scala 405:25]
  wire  arbiter_io_in_4_valid; // @[Slice.scala 405:25]
  wire [9:0] arbiter_io_in_4_bits_set; // @[Slice.scala 405:25]
  wire [2:0] arbiter_io_in_4_bits_way; // @[Slice.scala 405:25]
  wire  arbiter_io_in_4_bits_data_dirty; // @[Slice.scala 405:25]
  wire [1:0] arbiter_io_in_4_bits_data_state; // @[Slice.scala 405:25]
  wire [1:0] arbiter_io_in_4_bits_data_clientStates_0; // @[Slice.scala 405:25]
  wire [1:0] arbiter_io_in_4_bits_data_clientStates_1; // @[Slice.scala 405:25]
  wire  arbiter_io_in_5_ready; // @[Slice.scala 405:25]
  wire  arbiter_io_in_5_valid; // @[Slice.scala 405:25]
  wire [9:0] arbiter_io_in_5_bits_set; // @[Slice.scala 405:25]
  wire [2:0] arbiter_io_in_5_bits_way; // @[Slice.scala 405:25]
  wire  arbiter_io_in_5_bits_data_dirty; // @[Slice.scala 405:25]
  wire [1:0] arbiter_io_in_5_bits_data_state; // @[Slice.scala 405:25]
  wire [1:0] arbiter_io_in_5_bits_data_clientStates_0; // @[Slice.scala 405:25]
  wire [1:0] arbiter_io_in_5_bits_data_clientStates_1; // @[Slice.scala 405:25]
  wire  arbiter_io_in_6_ready; // @[Slice.scala 405:25]
  wire  arbiter_io_in_6_valid; // @[Slice.scala 405:25]
  wire [9:0] arbiter_io_in_6_bits_set; // @[Slice.scala 405:25]
  wire [2:0] arbiter_io_in_6_bits_way; // @[Slice.scala 405:25]
  wire  arbiter_io_in_6_bits_data_dirty; // @[Slice.scala 405:25]
  wire [1:0] arbiter_io_in_6_bits_data_state; // @[Slice.scala 405:25]
  wire [1:0] arbiter_io_in_6_bits_data_clientStates_0; // @[Slice.scala 405:25]
  wire [1:0] arbiter_io_in_6_bits_data_clientStates_1; // @[Slice.scala 405:25]
  wire  arbiter_io_in_7_ready; // @[Slice.scala 405:25]
  wire  arbiter_io_in_7_valid; // @[Slice.scala 405:25]
  wire [9:0] arbiter_io_in_7_bits_set; // @[Slice.scala 405:25]
  wire [2:0] arbiter_io_in_7_bits_way; // @[Slice.scala 405:25]
  wire  arbiter_io_in_7_bits_data_dirty; // @[Slice.scala 405:25]
  wire [1:0] arbiter_io_in_7_bits_data_state; // @[Slice.scala 405:25]
  wire [1:0] arbiter_io_in_7_bits_data_clientStates_0; // @[Slice.scala 405:25]
  wire [1:0] arbiter_io_in_7_bits_data_clientStates_1; // @[Slice.scala 405:25]
  wire  arbiter_io_in_8_ready; // @[Slice.scala 405:25]
  wire  arbiter_io_in_8_valid; // @[Slice.scala 405:25]
  wire [9:0] arbiter_io_in_8_bits_set; // @[Slice.scala 405:25]
  wire [2:0] arbiter_io_in_8_bits_way; // @[Slice.scala 405:25]
  wire  arbiter_io_in_8_bits_data_dirty; // @[Slice.scala 405:25]
  wire [1:0] arbiter_io_in_8_bits_data_state; // @[Slice.scala 405:25]
  wire [1:0] arbiter_io_in_8_bits_data_clientStates_0; // @[Slice.scala 405:25]
  wire [1:0] arbiter_io_in_8_bits_data_clientStates_1; // @[Slice.scala 405:25]
  wire  arbiter_io_in_9_ready; // @[Slice.scala 405:25]
  wire  arbiter_io_in_9_valid; // @[Slice.scala 405:25]
  wire [9:0] arbiter_io_in_9_bits_set; // @[Slice.scala 405:25]
  wire [2:0] arbiter_io_in_9_bits_way; // @[Slice.scala 405:25]
  wire  arbiter_io_in_9_bits_data_dirty; // @[Slice.scala 405:25]
  wire [1:0] arbiter_io_in_9_bits_data_state; // @[Slice.scala 405:25]
  wire [1:0] arbiter_io_in_9_bits_data_clientStates_0; // @[Slice.scala 405:25]
  wire [1:0] arbiter_io_in_9_bits_data_clientStates_1; // @[Slice.scala 405:25]
  wire  arbiter_io_in_10_ready; // @[Slice.scala 405:25]
  wire  arbiter_io_in_10_valid; // @[Slice.scala 405:25]
  wire [9:0] arbiter_io_in_10_bits_set; // @[Slice.scala 405:25]
  wire [2:0] arbiter_io_in_10_bits_way; // @[Slice.scala 405:25]
  wire  arbiter_io_in_10_bits_data_dirty; // @[Slice.scala 405:25]
  wire [1:0] arbiter_io_in_10_bits_data_state; // @[Slice.scala 405:25]
  wire [1:0] arbiter_io_in_10_bits_data_clientStates_0; // @[Slice.scala 405:25]
  wire [1:0] arbiter_io_in_10_bits_data_clientStates_1; // @[Slice.scala 405:25]
  wire  arbiter_io_in_11_ready; // @[Slice.scala 405:25]
  wire  arbiter_io_in_11_valid; // @[Slice.scala 405:25]
  wire [9:0] arbiter_io_in_11_bits_set; // @[Slice.scala 405:25]
  wire [2:0] arbiter_io_in_11_bits_way; // @[Slice.scala 405:25]
  wire  arbiter_io_in_11_bits_data_dirty; // @[Slice.scala 405:25]
  wire [1:0] arbiter_io_in_11_bits_data_state; // @[Slice.scala 405:25]
  wire [1:0] arbiter_io_in_11_bits_data_clientStates_0; // @[Slice.scala 405:25]
  wire [1:0] arbiter_io_in_11_bits_data_clientStates_1; // @[Slice.scala 405:25]
  wire  arbiter_io_in_12_ready; // @[Slice.scala 405:25]
  wire  arbiter_io_in_12_valid; // @[Slice.scala 405:25]
  wire [9:0] arbiter_io_in_12_bits_set; // @[Slice.scala 405:25]
  wire [2:0] arbiter_io_in_12_bits_way; // @[Slice.scala 405:25]
  wire  arbiter_io_in_12_bits_data_dirty; // @[Slice.scala 405:25]
  wire [1:0] arbiter_io_in_12_bits_data_state; // @[Slice.scala 405:25]
  wire [1:0] arbiter_io_in_12_bits_data_clientStates_0; // @[Slice.scala 405:25]
  wire [1:0] arbiter_io_in_12_bits_data_clientStates_1; // @[Slice.scala 405:25]
  wire  arbiter_io_in_13_ready; // @[Slice.scala 405:25]
  wire  arbiter_io_in_13_valid; // @[Slice.scala 405:25]
  wire [9:0] arbiter_io_in_13_bits_set; // @[Slice.scala 405:25]
  wire [2:0] arbiter_io_in_13_bits_way; // @[Slice.scala 405:25]
  wire  arbiter_io_in_13_bits_data_dirty; // @[Slice.scala 405:25]
  wire [1:0] arbiter_io_in_13_bits_data_state; // @[Slice.scala 405:25]
  wire [1:0] arbiter_io_in_13_bits_data_clientStates_0; // @[Slice.scala 405:25]
  wire [1:0] arbiter_io_in_13_bits_data_clientStates_1; // @[Slice.scala 405:25]
  wire  arbiter_io_in_14_ready; // @[Slice.scala 405:25]
  wire  arbiter_io_in_14_valid; // @[Slice.scala 405:25]
  wire [9:0] arbiter_io_in_14_bits_set; // @[Slice.scala 405:25]
  wire [2:0] arbiter_io_in_14_bits_way; // @[Slice.scala 405:25]
  wire  arbiter_io_in_14_bits_data_dirty; // @[Slice.scala 405:25]
  wire [1:0] arbiter_io_in_14_bits_data_state; // @[Slice.scala 405:25]
  wire [1:0] arbiter_io_in_14_bits_data_clientStates_0; // @[Slice.scala 405:25]
  wire [1:0] arbiter_io_in_14_bits_data_clientStates_1; // @[Slice.scala 405:25]
  wire  arbiter_io_in_15_ready; // @[Slice.scala 405:25]
  wire  arbiter_io_in_15_valid; // @[Slice.scala 405:25]
  wire [9:0] arbiter_io_in_15_bits_set; // @[Slice.scala 405:25]
  wire [2:0] arbiter_io_in_15_bits_way; // @[Slice.scala 405:25]
  wire  arbiter_io_in_15_bits_data_dirty; // @[Slice.scala 405:25]
  wire [1:0] arbiter_io_in_15_bits_data_state; // @[Slice.scala 405:25]
  wire [1:0] arbiter_io_in_15_bits_data_clientStates_0; // @[Slice.scala 405:25]
  wire [1:0] arbiter_io_in_15_bits_data_clientStates_1; // @[Slice.scala 405:25]
  wire  arbiter_io_out_valid; // @[Slice.scala 405:25]
  wire [9:0] arbiter_io_out_bits_set; // @[Slice.scala 405:25]
  wire [2:0] arbiter_io_out_bits_way; // @[Slice.scala 405:25]
  wire  arbiter_io_out_bits_data_dirty; // @[Slice.scala 405:25]
  wire [1:0] arbiter_io_out_bits_data_state; // @[Slice.scala 405:25]
  wire [1:0] arbiter_io_out_bits_data_clientStates_0; // @[Slice.scala 405:25]
  wire [1:0] arbiter_io_out_bits_data_clientStates_1; // @[Slice.scala 405:25]
  wire  sourceA_task_arb_clock; // @[Slice.scala 468:27]
  wire  sourceA_task_arb_reset; // @[Slice.scala 468:27]
  wire  sourceA_task_arb_io_in_0_ready; // @[Slice.scala 468:27]
  wire  sourceA_task_arb_io_in_0_valid; // @[Slice.scala 468:27]
  wire [19:0] sourceA_task_arb_io_in_0_bits_tag; // @[Slice.scala 468:27]
  wire [9:0] sourceA_task_arb_io_in_0_bits_set; // @[Slice.scala 468:27]
  wire [5:0] sourceA_task_arb_io_in_0_bits_off; // @[Slice.scala 468:27]
  wire [2:0] sourceA_task_arb_io_in_0_bits_opcode; // @[Slice.scala 468:27]
  wire [2:0] sourceA_task_arb_io_in_0_bits_param; // @[Slice.scala 468:27]
  wire [3:0] sourceA_task_arb_io_in_0_bits_source; // @[Slice.scala 468:27]
  wire [2:0] sourceA_task_arb_io_in_0_bits_bufIdx; // @[Slice.scala 468:27]
  wire [2:0] sourceA_task_arb_io_in_0_bits_size; // @[Slice.scala 468:27]
  wire  sourceA_task_arb_io_in_0_bits_putData; // @[Slice.scala 468:27]
  wire  sourceA_task_arb_io_in_1_ready; // @[Slice.scala 468:27]
  wire  sourceA_task_arb_io_in_1_valid; // @[Slice.scala 468:27]
  wire [19:0] sourceA_task_arb_io_in_1_bits_tag; // @[Slice.scala 468:27]
  wire [9:0] sourceA_task_arb_io_in_1_bits_set; // @[Slice.scala 468:27]
  wire [5:0] sourceA_task_arb_io_in_1_bits_off; // @[Slice.scala 468:27]
  wire [2:0] sourceA_task_arb_io_in_1_bits_opcode; // @[Slice.scala 468:27]
  wire [2:0] sourceA_task_arb_io_in_1_bits_param; // @[Slice.scala 468:27]
  wire [3:0] sourceA_task_arb_io_in_1_bits_source; // @[Slice.scala 468:27]
  wire [2:0] sourceA_task_arb_io_in_1_bits_bufIdx; // @[Slice.scala 468:27]
  wire [2:0] sourceA_task_arb_io_in_1_bits_size; // @[Slice.scala 468:27]
  wire  sourceA_task_arb_io_in_1_bits_putData; // @[Slice.scala 468:27]
  wire  sourceA_task_arb_io_in_2_ready; // @[Slice.scala 468:27]
  wire  sourceA_task_arb_io_in_2_valid; // @[Slice.scala 468:27]
  wire [19:0] sourceA_task_arb_io_in_2_bits_tag; // @[Slice.scala 468:27]
  wire [9:0] sourceA_task_arb_io_in_2_bits_set; // @[Slice.scala 468:27]
  wire [5:0] sourceA_task_arb_io_in_2_bits_off; // @[Slice.scala 468:27]
  wire [2:0] sourceA_task_arb_io_in_2_bits_opcode; // @[Slice.scala 468:27]
  wire [2:0] sourceA_task_arb_io_in_2_bits_param; // @[Slice.scala 468:27]
  wire [3:0] sourceA_task_arb_io_in_2_bits_source; // @[Slice.scala 468:27]
  wire [2:0] sourceA_task_arb_io_in_2_bits_bufIdx; // @[Slice.scala 468:27]
  wire [2:0] sourceA_task_arb_io_in_2_bits_size; // @[Slice.scala 468:27]
  wire  sourceA_task_arb_io_in_2_bits_putData; // @[Slice.scala 468:27]
  wire  sourceA_task_arb_io_in_3_ready; // @[Slice.scala 468:27]
  wire  sourceA_task_arb_io_in_3_valid; // @[Slice.scala 468:27]
  wire [19:0] sourceA_task_arb_io_in_3_bits_tag; // @[Slice.scala 468:27]
  wire [9:0] sourceA_task_arb_io_in_3_bits_set; // @[Slice.scala 468:27]
  wire [5:0] sourceA_task_arb_io_in_3_bits_off; // @[Slice.scala 468:27]
  wire [2:0] sourceA_task_arb_io_in_3_bits_opcode; // @[Slice.scala 468:27]
  wire [2:0] sourceA_task_arb_io_in_3_bits_param; // @[Slice.scala 468:27]
  wire [3:0] sourceA_task_arb_io_in_3_bits_source; // @[Slice.scala 468:27]
  wire [2:0] sourceA_task_arb_io_in_3_bits_bufIdx; // @[Slice.scala 468:27]
  wire [2:0] sourceA_task_arb_io_in_3_bits_size; // @[Slice.scala 468:27]
  wire  sourceA_task_arb_io_in_3_bits_putData; // @[Slice.scala 468:27]
  wire  sourceA_task_arb_io_in_4_ready; // @[Slice.scala 468:27]
  wire  sourceA_task_arb_io_in_4_valid; // @[Slice.scala 468:27]
  wire [19:0] sourceA_task_arb_io_in_4_bits_tag; // @[Slice.scala 468:27]
  wire [9:0] sourceA_task_arb_io_in_4_bits_set; // @[Slice.scala 468:27]
  wire [5:0] sourceA_task_arb_io_in_4_bits_off; // @[Slice.scala 468:27]
  wire [2:0] sourceA_task_arb_io_in_4_bits_opcode; // @[Slice.scala 468:27]
  wire [2:0] sourceA_task_arb_io_in_4_bits_param; // @[Slice.scala 468:27]
  wire [3:0] sourceA_task_arb_io_in_4_bits_source; // @[Slice.scala 468:27]
  wire [2:0] sourceA_task_arb_io_in_4_bits_bufIdx; // @[Slice.scala 468:27]
  wire [2:0] sourceA_task_arb_io_in_4_bits_size; // @[Slice.scala 468:27]
  wire  sourceA_task_arb_io_in_4_bits_putData; // @[Slice.scala 468:27]
  wire  sourceA_task_arb_io_in_5_ready; // @[Slice.scala 468:27]
  wire  sourceA_task_arb_io_in_5_valid; // @[Slice.scala 468:27]
  wire [19:0] sourceA_task_arb_io_in_5_bits_tag; // @[Slice.scala 468:27]
  wire [9:0] sourceA_task_arb_io_in_5_bits_set; // @[Slice.scala 468:27]
  wire [5:0] sourceA_task_arb_io_in_5_bits_off; // @[Slice.scala 468:27]
  wire [2:0] sourceA_task_arb_io_in_5_bits_opcode; // @[Slice.scala 468:27]
  wire [2:0] sourceA_task_arb_io_in_5_bits_param; // @[Slice.scala 468:27]
  wire [3:0] sourceA_task_arb_io_in_5_bits_source; // @[Slice.scala 468:27]
  wire [2:0] sourceA_task_arb_io_in_5_bits_bufIdx; // @[Slice.scala 468:27]
  wire [2:0] sourceA_task_arb_io_in_5_bits_size; // @[Slice.scala 468:27]
  wire  sourceA_task_arb_io_in_5_bits_putData; // @[Slice.scala 468:27]
  wire  sourceA_task_arb_io_in_6_ready; // @[Slice.scala 468:27]
  wire  sourceA_task_arb_io_in_6_valid; // @[Slice.scala 468:27]
  wire [19:0] sourceA_task_arb_io_in_6_bits_tag; // @[Slice.scala 468:27]
  wire [9:0] sourceA_task_arb_io_in_6_bits_set; // @[Slice.scala 468:27]
  wire [5:0] sourceA_task_arb_io_in_6_bits_off; // @[Slice.scala 468:27]
  wire [2:0] sourceA_task_arb_io_in_6_bits_opcode; // @[Slice.scala 468:27]
  wire [2:0] sourceA_task_arb_io_in_6_bits_param; // @[Slice.scala 468:27]
  wire [3:0] sourceA_task_arb_io_in_6_bits_source; // @[Slice.scala 468:27]
  wire [2:0] sourceA_task_arb_io_in_6_bits_bufIdx; // @[Slice.scala 468:27]
  wire [2:0] sourceA_task_arb_io_in_6_bits_size; // @[Slice.scala 468:27]
  wire  sourceA_task_arb_io_in_6_bits_putData; // @[Slice.scala 468:27]
  wire  sourceA_task_arb_io_in_7_ready; // @[Slice.scala 468:27]
  wire  sourceA_task_arb_io_in_7_valid; // @[Slice.scala 468:27]
  wire [19:0] sourceA_task_arb_io_in_7_bits_tag; // @[Slice.scala 468:27]
  wire [9:0] sourceA_task_arb_io_in_7_bits_set; // @[Slice.scala 468:27]
  wire [5:0] sourceA_task_arb_io_in_7_bits_off; // @[Slice.scala 468:27]
  wire [2:0] sourceA_task_arb_io_in_7_bits_opcode; // @[Slice.scala 468:27]
  wire [2:0] sourceA_task_arb_io_in_7_bits_param; // @[Slice.scala 468:27]
  wire [3:0] sourceA_task_arb_io_in_7_bits_source; // @[Slice.scala 468:27]
  wire [2:0] sourceA_task_arb_io_in_7_bits_bufIdx; // @[Slice.scala 468:27]
  wire [2:0] sourceA_task_arb_io_in_7_bits_size; // @[Slice.scala 468:27]
  wire  sourceA_task_arb_io_in_7_bits_putData; // @[Slice.scala 468:27]
  wire  sourceA_task_arb_io_in_8_ready; // @[Slice.scala 468:27]
  wire  sourceA_task_arb_io_in_8_valid; // @[Slice.scala 468:27]
  wire [19:0] sourceA_task_arb_io_in_8_bits_tag; // @[Slice.scala 468:27]
  wire [9:0] sourceA_task_arb_io_in_8_bits_set; // @[Slice.scala 468:27]
  wire [5:0] sourceA_task_arb_io_in_8_bits_off; // @[Slice.scala 468:27]
  wire [2:0] sourceA_task_arb_io_in_8_bits_opcode; // @[Slice.scala 468:27]
  wire [2:0] sourceA_task_arb_io_in_8_bits_param; // @[Slice.scala 468:27]
  wire [3:0] sourceA_task_arb_io_in_8_bits_source; // @[Slice.scala 468:27]
  wire [2:0] sourceA_task_arb_io_in_8_bits_bufIdx; // @[Slice.scala 468:27]
  wire [2:0] sourceA_task_arb_io_in_8_bits_size; // @[Slice.scala 468:27]
  wire  sourceA_task_arb_io_in_8_bits_putData; // @[Slice.scala 468:27]
  wire  sourceA_task_arb_io_in_9_ready; // @[Slice.scala 468:27]
  wire  sourceA_task_arb_io_in_9_valid; // @[Slice.scala 468:27]
  wire [19:0] sourceA_task_arb_io_in_9_bits_tag; // @[Slice.scala 468:27]
  wire [9:0] sourceA_task_arb_io_in_9_bits_set; // @[Slice.scala 468:27]
  wire [5:0] sourceA_task_arb_io_in_9_bits_off; // @[Slice.scala 468:27]
  wire [2:0] sourceA_task_arb_io_in_9_bits_opcode; // @[Slice.scala 468:27]
  wire [2:0] sourceA_task_arb_io_in_9_bits_param; // @[Slice.scala 468:27]
  wire [3:0] sourceA_task_arb_io_in_9_bits_source; // @[Slice.scala 468:27]
  wire [2:0] sourceA_task_arb_io_in_9_bits_bufIdx; // @[Slice.scala 468:27]
  wire [2:0] sourceA_task_arb_io_in_9_bits_size; // @[Slice.scala 468:27]
  wire  sourceA_task_arb_io_in_9_bits_putData; // @[Slice.scala 468:27]
  wire  sourceA_task_arb_io_in_10_ready; // @[Slice.scala 468:27]
  wire  sourceA_task_arb_io_in_10_valid; // @[Slice.scala 468:27]
  wire [19:0] sourceA_task_arb_io_in_10_bits_tag; // @[Slice.scala 468:27]
  wire [9:0] sourceA_task_arb_io_in_10_bits_set; // @[Slice.scala 468:27]
  wire [5:0] sourceA_task_arb_io_in_10_bits_off; // @[Slice.scala 468:27]
  wire [2:0] sourceA_task_arb_io_in_10_bits_opcode; // @[Slice.scala 468:27]
  wire [2:0] sourceA_task_arb_io_in_10_bits_param; // @[Slice.scala 468:27]
  wire [3:0] sourceA_task_arb_io_in_10_bits_source; // @[Slice.scala 468:27]
  wire [2:0] sourceA_task_arb_io_in_10_bits_bufIdx; // @[Slice.scala 468:27]
  wire [2:0] sourceA_task_arb_io_in_10_bits_size; // @[Slice.scala 468:27]
  wire  sourceA_task_arb_io_in_10_bits_putData; // @[Slice.scala 468:27]
  wire  sourceA_task_arb_io_in_11_ready; // @[Slice.scala 468:27]
  wire  sourceA_task_arb_io_in_11_valid; // @[Slice.scala 468:27]
  wire [19:0] sourceA_task_arb_io_in_11_bits_tag; // @[Slice.scala 468:27]
  wire [9:0] sourceA_task_arb_io_in_11_bits_set; // @[Slice.scala 468:27]
  wire [5:0] sourceA_task_arb_io_in_11_bits_off; // @[Slice.scala 468:27]
  wire [2:0] sourceA_task_arb_io_in_11_bits_opcode; // @[Slice.scala 468:27]
  wire [2:0] sourceA_task_arb_io_in_11_bits_param; // @[Slice.scala 468:27]
  wire [3:0] sourceA_task_arb_io_in_11_bits_source; // @[Slice.scala 468:27]
  wire [2:0] sourceA_task_arb_io_in_11_bits_bufIdx; // @[Slice.scala 468:27]
  wire [2:0] sourceA_task_arb_io_in_11_bits_size; // @[Slice.scala 468:27]
  wire  sourceA_task_arb_io_in_11_bits_putData; // @[Slice.scala 468:27]
  wire  sourceA_task_arb_io_in_12_ready; // @[Slice.scala 468:27]
  wire  sourceA_task_arb_io_in_12_valid; // @[Slice.scala 468:27]
  wire [19:0] sourceA_task_arb_io_in_12_bits_tag; // @[Slice.scala 468:27]
  wire [9:0] sourceA_task_arb_io_in_12_bits_set; // @[Slice.scala 468:27]
  wire [5:0] sourceA_task_arb_io_in_12_bits_off; // @[Slice.scala 468:27]
  wire [2:0] sourceA_task_arb_io_in_12_bits_opcode; // @[Slice.scala 468:27]
  wire [2:0] sourceA_task_arb_io_in_12_bits_param; // @[Slice.scala 468:27]
  wire [3:0] sourceA_task_arb_io_in_12_bits_source; // @[Slice.scala 468:27]
  wire [2:0] sourceA_task_arb_io_in_12_bits_bufIdx; // @[Slice.scala 468:27]
  wire [2:0] sourceA_task_arb_io_in_12_bits_size; // @[Slice.scala 468:27]
  wire  sourceA_task_arb_io_in_12_bits_putData; // @[Slice.scala 468:27]
  wire  sourceA_task_arb_io_in_13_ready; // @[Slice.scala 468:27]
  wire  sourceA_task_arb_io_in_13_valid; // @[Slice.scala 468:27]
  wire [19:0] sourceA_task_arb_io_in_13_bits_tag; // @[Slice.scala 468:27]
  wire [9:0] sourceA_task_arb_io_in_13_bits_set; // @[Slice.scala 468:27]
  wire [5:0] sourceA_task_arb_io_in_13_bits_off; // @[Slice.scala 468:27]
  wire [2:0] sourceA_task_arb_io_in_13_bits_opcode; // @[Slice.scala 468:27]
  wire [2:0] sourceA_task_arb_io_in_13_bits_param; // @[Slice.scala 468:27]
  wire [3:0] sourceA_task_arb_io_in_13_bits_source; // @[Slice.scala 468:27]
  wire [2:0] sourceA_task_arb_io_in_13_bits_bufIdx; // @[Slice.scala 468:27]
  wire [2:0] sourceA_task_arb_io_in_13_bits_size; // @[Slice.scala 468:27]
  wire  sourceA_task_arb_io_in_13_bits_putData; // @[Slice.scala 468:27]
  wire  sourceA_task_arb_io_out_ready; // @[Slice.scala 468:27]
  wire  sourceA_task_arb_io_out_valid; // @[Slice.scala 468:27]
  wire [19:0] sourceA_task_arb_io_out_bits_tag; // @[Slice.scala 468:27]
  wire [9:0] sourceA_task_arb_io_out_bits_set; // @[Slice.scala 468:27]
  wire [5:0] sourceA_task_arb_io_out_bits_off; // @[Slice.scala 468:27]
  wire [2:0] sourceA_task_arb_io_out_bits_opcode; // @[Slice.scala 468:27]
  wire [2:0] sourceA_task_arb_io_out_bits_param; // @[Slice.scala 468:27]
  wire [3:0] sourceA_task_arb_io_out_bits_source; // @[Slice.scala 468:27]
  wire [2:0] sourceA_task_arb_io_out_bits_bufIdx; // @[Slice.scala 468:27]
  wire [2:0] sourceA_task_arb_io_out_bits_size; // @[Slice.scala 468:27]
  wire  sourceA_task_arb_io_out_bits_putData; // @[Slice.scala 468:27]
  wire  sourceB_task_arb_clock; // @[Slice.scala 468:27]
  wire  sourceB_task_arb_reset; // @[Slice.scala 468:27]
  wire  sourceB_task_arb_io_in_0_ready; // @[Slice.scala 468:27]
  wire  sourceB_task_arb_io_in_0_valid; // @[Slice.scala 468:27]
  wire [9:0] sourceB_task_arb_io_in_0_bits_set; // @[Slice.scala 468:27]
  wire [19:0] sourceB_task_arb_io_in_0_bits_tag; // @[Slice.scala 468:27]
  wire [2:0] sourceB_task_arb_io_in_0_bits_param; // @[Slice.scala 468:27]
  wire [1:0] sourceB_task_arb_io_in_0_bits_clients; // @[Slice.scala 468:27]
  wire  sourceB_task_arb_io_in_0_bits_needData; // @[Slice.scala 468:27]
  wire  sourceB_task_arb_io_in_1_ready; // @[Slice.scala 468:27]
  wire  sourceB_task_arb_io_in_1_valid; // @[Slice.scala 468:27]
  wire [9:0] sourceB_task_arb_io_in_1_bits_set; // @[Slice.scala 468:27]
  wire [19:0] sourceB_task_arb_io_in_1_bits_tag; // @[Slice.scala 468:27]
  wire [2:0] sourceB_task_arb_io_in_1_bits_param; // @[Slice.scala 468:27]
  wire [1:0] sourceB_task_arb_io_in_1_bits_clients; // @[Slice.scala 468:27]
  wire  sourceB_task_arb_io_in_1_bits_needData; // @[Slice.scala 468:27]
  wire  sourceB_task_arb_io_in_2_ready; // @[Slice.scala 468:27]
  wire  sourceB_task_arb_io_in_2_valid; // @[Slice.scala 468:27]
  wire [9:0] sourceB_task_arb_io_in_2_bits_set; // @[Slice.scala 468:27]
  wire [19:0] sourceB_task_arb_io_in_2_bits_tag; // @[Slice.scala 468:27]
  wire [2:0] sourceB_task_arb_io_in_2_bits_param; // @[Slice.scala 468:27]
  wire [1:0] sourceB_task_arb_io_in_2_bits_clients; // @[Slice.scala 468:27]
  wire  sourceB_task_arb_io_in_2_bits_needData; // @[Slice.scala 468:27]
  wire  sourceB_task_arb_io_in_3_ready; // @[Slice.scala 468:27]
  wire  sourceB_task_arb_io_in_3_valid; // @[Slice.scala 468:27]
  wire [9:0] sourceB_task_arb_io_in_3_bits_set; // @[Slice.scala 468:27]
  wire [19:0] sourceB_task_arb_io_in_3_bits_tag; // @[Slice.scala 468:27]
  wire [2:0] sourceB_task_arb_io_in_3_bits_param; // @[Slice.scala 468:27]
  wire [1:0] sourceB_task_arb_io_in_3_bits_clients; // @[Slice.scala 468:27]
  wire  sourceB_task_arb_io_in_3_bits_needData; // @[Slice.scala 468:27]
  wire  sourceB_task_arb_io_in_4_ready; // @[Slice.scala 468:27]
  wire  sourceB_task_arb_io_in_4_valid; // @[Slice.scala 468:27]
  wire [9:0] sourceB_task_arb_io_in_4_bits_set; // @[Slice.scala 468:27]
  wire [19:0] sourceB_task_arb_io_in_4_bits_tag; // @[Slice.scala 468:27]
  wire [2:0] sourceB_task_arb_io_in_4_bits_param; // @[Slice.scala 468:27]
  wire [1:0] sourceB_task_arb_io_in_4_bits_clients; // @[Slice.scala 468:27]
  wire  sourceB_task_arb_io_in_4_bits_needData; // @[Slice.scala 468:27]
  wire  sourceB_task_arb_io_in_5_ready; // @[Slice.scala 468:27]
  wire  sourceB_task_arb_io_in_5_valid; // @[Slice.scala 468:27]
  wire [9:0] sourceB_task_arb_io_in_5_bits_set; // @[Slice.scala 468:27]
  wire [19:0] sourceB_task_arb_io_in_5_bits_tag; // @[Slice.scala 468:27]
  wire [2:0] sourceB_task_arb_io_in_5_bits_param; // @[Slice.scala 468:27]
  wire [1:0] sourceB_task_arb_io_in_5_bits_clients; // @[Slice.scala 468:27]
  wire  sourceB_task_arb_io_in_5_bits_needData; // @[Slice.scala 468:27]
  wire  sourceB_task_arb_io_in_6_ready; // @[Slice.scala 468:27]
  wire  sourceB_task_arb_io_in_6_valid; // @[Slice.scala 468:27]
  wire [9:0] sourceB_task_arb_io_in_6_bits_set; // @[Slice.scala 468:27]
  wire [19:0] sourceB_task_arb_io_in_6_bits_tag; // @[Slice.scala 468:27]
  wire [2:0] sourceB_task_arb_io_in_6_bits_param; // @[Slice.scala 468:27]
  wire [1:0] sourceB_task_arb_io_in_6_bits_clients; // @[Slice.scala 468:27]
  wire  sourceB_task_arb_io_in_6_bits_needData; // @[Slice.scala 468:27]
  wire  sourceB_task_arb_io_in_7_ready; // @[Slice.scala 468:27]
  wire  sourceB_task_arb_io_in_7_valid; // @[Slice.scala 468:27]
  wire [9:0] sourceB_task_arb_io_in_7_bits_set; // @[Slice.scala 468:27]
  wire [19:0] sourceB_task_arb_io_in_7_bits_tag; // @[Slice.scala 468:27]
  wire [2:0] sourceB_task_arb_io_in_7_bits_param; // @[Slice.scala 468:27]
  wire [1:0] sourceB_task_arb_io_in_7_bits_clients; // @[Slice.scala 468:27]
  wire  sourceB_task_arb_io_in_7_bits_needData; // @[Slice.scala 468:27]
  wire  sourceB_task_arb_io_in_8_ready; // @[Slice.scala 468:27]
  wire  sourceB_task_arb_io_in_8_valid; // @[Slice.scala 468:27]
  wire [9:0] sourceB_task_arb_io_in_8_bits_set; // @[Slice.scala 468:27]
  wire [19:0] sourceB_task_arb_io_in_8_bits_tag; // @[Slice.scala 468:27]
  wire [2:0] sourceB_task_arb_io_in_8_bits_param; // @[Slice.scala 468:27]
  wire [1:0] sourceB_task_arb_io_in_8_bits_clients; // @[Slice.scala 468:27]
  wire  sourceB_task_arb_io_in_8_bits_needData; // @[Slice.scala 468:27]
  wire  sourceB_task_arb_io_in_9_ready; // @[Slice.scala 468:27]
  wire  sourceB_task_arb_io_in_9_valid; // @[Slice.scala 468:27]
  wire [9:0] sourceB_task_arb_io_in_9_bits_set; // @[Slice.scala 468:27]
  wire [19:0] sourceB_task_arb_io_in_9_bits_tag; // @[Slice.scala 468:27]
  wire [2:0] sourceB_task_arb_io_in_9_bits_param; // @[Slice.scala 468:27]
  wire [1:0] sourceB_task_arb_io_in_9_bits_clients; // @[Slice.scala 468:27]
  wire  sourceB_task_arb_io_in_9_bits_needData; // @[Slice.scala 468:27]
  wire  sourceB_task_arb_io_in_10_ready; // @[Slice.scala 468:27]
  wire  sourceB_task_arb_io_in_10_valid; // @[Slice.scala 468:27]
  wire [9:0] sourceB_task_arb_io_in_10_bits_set; // @[Slice.scala 468:27]
  wire [19:0] sourceB_task_arb_io_in_10_bits_tag; // @[Slice.scala 468:27]
  wire [2:0] sourceB_task_arb_io_in_10_bits_param; // @[Slice.scala 468:27]
  wire [1:0] sourceB_task_arb_io_in_10_bits_clients; // @[Slice.scala 468:27]
  wire  sourceB_task_arb_io_in_10_bits_needData; // @[Slice.scala 468:27]
  wire  sourceB_task_arb_io_in_11_ready; // @[Slice.scala 468:27]
  wire  sourceB_task_arb_io_in_11_valid; // @[Slice.scala 468:27]
  wire [9:0] sourceB_task_arb_io_in_11_bits_set; // @[Slice.scala 468:27]
  wire [19:0] sourceB_task_arb_io_in_11_bits_tag; // @[Slice.scala 468:27]
  wire [2:0] sourceB_task_arb_io_in_11_bits_param; // @[Slice.scala 468:27]
  wire [1:0] sourceB_task_arb_io_in_11_bits_clients; // @[Slice.scala 468:27]
  wire  sourceB_task_arb_io_in_11_bits_needData; // @[Slice.scala 468:27]
  wire  sourceB_task_arb_io_in_12_ready; // @[Slice.scala 468:27]
  wire  sourceB_task_arb_io_in_12_valid; // @[Slice.scala 468:27]
  wire [9:0] sourceB_task_arb_io_in_12_bits_set; // @[Slice.scala 468:27]
  wire [19:0] sourceB_task_arb_io_in_12_bits_tag; // @[Slice.scala 468:27]
  wire [2:0] sourceB_task_arb_io_in_12_bits_param; // @[Slice.scala 468:27]
  wire [1:0] sourceB_task_arb_io_in_12_bits_clients; // @[Slice.scala 468:27]
  wire  sourceB_task_arb_io_in_12_bits_needData; // @[Slice.scala 468:27]
  wire  sourceB_task_arb_io_in_13_ready; // @[Slice.scala 468:27]
  wire  sourceB_task_arb_io_in_13_valid; // @[Slice.scala 468:27]
  wire [9:0] sourceB_task_arb_io_in_13_bits_set; // @[Slice.scala 468:27]
  wire [19:0] sourceB_task_arb_io_in_13_bits_tag; // @[Slice.scala 468:27]
  wire [2:0] sourceB_task_arb_io_in_13_bits_param; // @[Slice.scala 468:27]
  wire [1:0] sourceB_task_arb_io_in_13_bits_clients; // @[Slice.scala 468:27]
  wire  sourceB_task_arb_io_in_13_bits_needData; // @[Slice.scala 468:27]
  wire  sourceB_task_arb_io_out_ready; // @[Slice.scala 468:27]
  wire  sourceB_task_arb_io_out_valid; // @[Slice.scala 468:27]
  wire [9:0] sourceB_task_arb_io_out_bits_set; // @[Slice.scala 468:27]
  wire [19:0] sourceB_task_arb_io_out_bits_tag; // @[Slice.scala 468:27]
  wire [2:0] sourceB_task_arb_io_out_bits_param; // @[Slice.scala 468:27]
  wire [1:0] sourceB_task_arb_io_out_bits_clients; // @[Slice.scala 468:27]
  wire  sourceB_task_arb_io_out_bits_needData; // @[Slice.scala 468:27]
  wire  sourceC_task_arb_clock; // @[Slice.scala 468:27]
  wire  sourceC_task_arb_reset; // @[Slice.scala 468:27]
  wire  sourceC_task_arb_io_in_0_ready; // @[Slice.scala 468:27]
  wire  sourceC_task_arb_io_in_0_valid; // @[Slice.scala 468:27]
  wire [2:0] sourceC_task_arb_io_in_0_bits_opcode; // @[Slice.scala 468:27]
  wire [19:0] sourceC_task_arb_io_in_0_bits_tag; // @[Slice.scala 468:27]
  wire [9:0] sourceC_task_arb_io_in_0_bits_set; // @[Slice.scala 468:27]
  wire [3:0] sourceC_task_arb_io_in_0_bits_source; // @[Slice.scala 468:27]
  wire [2:0] sourceC_task_arb_io_in_0_bits_way; // @[Slice.scala 468:27]
  wire  sourceC_task_arb_io_in_1_ready; // @[Slice.scala 468:27]
  wire  sourceC_task_arb_io_in_1_valid; // @[Slice.scala 468:27]
  wire [2:0] sourceC_task_arb_io_in_1_bits_opcode; // @[Slice.scala 468:27]
  wire [19:0] sourceC_task_arb_io_in_1_bits_tag; // @[Slice.scala 468:27]
  wire [9:0] sourceC_task_arb_io_in_1_bits_set; // @[Slice.scala 468:27]
  wire [3:0] sourceC_task_arb_io_in_1_bits_source; // @[Slice.scala 468:27]
  wire [2:0] sourceC_task_arb_io_in_1_bits_way; // @[Slice.scala 468:27]
  wire  sourceC_task_arb_io_in_2_ready; // @[Slice.scala 468:27]
  wire  sourceC_task_arb_io_in_2_valid; // @[Slice.scala 468:27]
  wire [2:0] sourceC_task_arb_io_in_2_bits_opcode; // @[Slice.scala 468:27]
  wire [19:0] sourceC_task_arb_io_in_2_bits_tag; // @[Slice.scala 468:27]
  wire [9:0] sourceC_task_arb_io_in_2_bits_set; // @[Slice.scala 468:27]
  wire [3:0] sourceC_task_arb_io_in_2_bits_source; // @[Slice.scala 468:27]
  wire [2:0] sourceC_task_arb_io_in_2_bits_way; // @[Slice.scala 468:27]
  wire  sourceC_task_arb_io_in_3_ready; // @[Slice.scala 468:27]
  wire  sourceC_task_arb_io_in_3_valid; // @[Slice.scala 468:27]
  wire [2:0] sourceC_task_arb_io_in_3_bits_opcode; // @[Slice.scala 468:27]
  wire [19:0] sourceC_task_arb_io_in_3_bits_tag; // @[Slice.scala 468:27]
  wire [9:0] sourceC_task_arb_io_in_3_bits_set; // @[Slice.scala 468:27]
  wire [3:0] sourceC_task_arb_io_in_3_bits_source; // @[Slice.scala 468:27]
  wire [2:0] sourceC_task_arb_io_in_3_bits_way; // @[Slice.scala 468:27]
  wire  sourceC_task_arb_io_in_4_ready; // @[Slice.scala 468:27]
  wire  sourceC_task_arb_io_in_4_valid; // @[Slice.scala 468:27]
  wire [2:0] sourceC_task_arb_io_in_4_bits_opcode; // @[Slice.scala 468:27]
  wire [19:0] sourceC_task_arb_io_in_4_bits_tag; // @[Slice.scala 468:27]
  wire [9:0] sourceC_task_arb_io_in_4_bits_set; // @[Slice.scala 468:27]
  wire [3:0] sourceC_task_arb_io_in_4_bits_source; // @[Slice.scala 468:27]
  wire [2:0] sourceC_task_arb_io_in_4_bits_way; // @[Slice.scala 468:27]
  wire  sourceC_task_arb_io_in_5_ready; // @[Slice.scala 468:27]
  wire  sourceC_task_arb_io_in_5_valid; // @[Slice.scala 468:27]
  wire [2:0] sourceC_task_arb_io_in_5_bits_opcode; // @[Slice.scala 468:27]
  wire [19:0] sourceC_task_arb_io_in_5_bits_tag; // @[Slice.scala 468:27]
  wire [9:0] sourceC_task_arb_io_in_5_bits_set; // @[Slice.scala 468:27]
  wire [3:0] sourceC_task_arb_io_in_5_bits_source; // @[Slice.scala 468:27]
  wire [2:0] sourceC_task_arb_io_in_5_bits_way; // @[Slice.scala 468:27]
  wire  sourceC_task_arb_io_in_6_ready; // @[Slice.scala 468:27]
  wire  sourceC_task_arb_io_in_6_valid; // @[Slice.scala 468:27]
  wire [2:0] sourceC_task_arb_io_in_6_bits_opcode; // @[Slice.scala 468:27]
  wire [19:0] sourceC_task_arb_io_in_6_bits_tag; // @[Slice.scala 468:27]
  wire [9:0] sourceC_task_arb_io_in_6_bits_set; // @[Slice.scala 468:27]
  wire [3:0] sourceC_task_arb_io_in_6_bits_source; // @[Slice.scala 468:27]
  wire [2:0] sourceC_task_arb_io_in_6_bits_way; // @[Slice.scala 468:27]
  wire  sourceC_task_arb_io_in_7_ready; // @[Slice.scala 468:27]
  wire  sourceC_task_arb_io_in_7_valid; // @[Slice.scala 468:27]
  wire [2:0] sourceC_task_arb_io_in_7_bits_opcode; // @[Slice.scala 468:27]
  wire [19:0] sourceC_task_arb_io_in_7_bits_tag; // @[Slice.scala 468:27]
  wire [9:0] sourceC_task_arb_io_in_7_bits_set; // @[Slice.scala 468:27]
  wire [3:0] sourceC_task_arb_io_in_7_bits_source; // @[Slice.scala 468:27]
  wire [2:0] sourceC_task_arb_io_in_7_bits_way; // @[Slice.scala 468:27]
  wire  sourceC_task_arb_io_in_8_ready; // @[Slice.scala 468:27]
  wire  sourceC_task_arb_io_in_8_valid; // @[Slice.scala 468:27]
  wire [2:0] sourceC_task_arb_io_in_8_bits_opcode; // @[Slice.scala 468:27]
  wire [19:0] sourceC_task_arb_io_in_8_bits_tag; // @[Slice.scala 468:27]
  wire [9:0] sourceC_task_arb_io_in_8_bits_set; // @[Slice.scala 468:27]
  wire [3:0] sourceC_task_arb_io_in_8_bits_source; // @[Slice.scala 468:27]
  wire [2:0] sourceC_task_arb_io_in_8_bits_way; // @[Slice.scala 468:27]
  wire  sourceC_task_arb_io_in_9_ready; // @[Slice.scala 468:27]
  wire  sourceC_task_arb_io_in_9_valid; // @[Slice.scala 468:27]
  wire [2:0] sourceC_task_arb_io_in_9_bits_opcode; // @[Slice.scala 468:27]
  wire [19:0] sourceC_task_arb_io_in_9_bits_tag; // @[Slice.scala 468:27]
  wire [9:0] sourceC_task_arb_io_in_9_bits_set; // @[Slice.scala 468:27]
  wire [3:0] sourceC_task_arb_io_in_9_bits_source; // @[Slice.scala 468:27]
  wire [2:0] sourceC_task_arb_io_in_9_bits_way; // @[Slice.scala 468:27]
  wire  sourceC_task_arb_io_in_10_ready; // @[Slice.scala 468:27]
  wire  sourceC_task_arb_io_in_10_valid; // @[Slice.scala 468:27]
  wire [2:0] sourceC_task_arb_io_in_10_bits_opcode; // @[Slice.scala 468:27]
  wire [19:0] sourceC_task_arb_io_in_10_bits_tag; // @[Slice.scala 468:27]
  wire [9:0] sourceC_task_arb_io_in_10_bits_set; // @[Slice.scala 468:27]
  wire [3:0] sourceC_task_arb_io_in_10_bits_source; // @[Slice.scala 468:27]
  wire [2:0] sourceC_task_arb_io_in_10_bits_way; // @[Slice.scala 468:27]
  wire  sourceC_task_arb_io_in_11_ready; // @[Slice.scala 468:27]
  wire  sourceC_task_arb_io_in_11_valid; // @[Slice.scala 468:27]
  wire [2:0] sourceC_task_arb_io_in_11_bits_opcode; // @[Slice.scala 468:27]
  wire [19:0] sourceC_task_arb_io_in_11_bits_tag; // @[Slice.scala 468:27]
  wire [9:0] sourceC_task_arb_io_in_11_bits_set; // @[Slice.scala 468:27]
  wire [3:0] sourceC_task_arb_io_in_11_bits_source; // @[Slice.scala 468:27]
  wire [2:0] sourceC_task_arb_io_in_11_bits_way; // @[Slice.scala 468:27]
  wire  sourceC_task_arb_io_in_12_ready; // @[Slice.scala 468:27]
  wire  sourceC_task_arb_io_in_12_valid; // @[Slice.scala 468:27]
  wire [2:0] sourceC_task_arb_io_in_12_bits_opcode; // @[Slice.scala 468:27]
  wire [19:0] sourceC_task_arb_io_in_12_bits_tag; // @[Slice.scala 468:27]
  wire [9:0] sourceC_task_arb_io_in_12_bits_set; // @[Slice.scala 468:27]
  wire [3:0] sourceC_task_arb_io_in_12_bits_source; // @[Slice.scala 468:27]
  wire [2:0] sourceC_task_arb_io_in_12_bits_way; // @[Slice.scala 468:27]
  wire  sourceC_task_arb_io_in_13_ready; // @[Slice.scala 468:27]
  wire  sourceC_task_arb_io_in_13_valid; // @[Slice.scala 468:27]
  wire [2:0] sourceC_task_arb_io_in_13_bits_opcode; // @[Slice.scala 468:27]
  wire [19:0] sourceC_task_arb_io_in_13_bits_tag; // @[Slice.scala 468:27]
  wire [9:0] sourceC_task_arb_io_in_13_bits_set; // @[Slice.scala 468:27]
  wire [3:0] sourceC_task_arb_io_in_13_bits_source; // @[Slice.scala 468:27]
  wire [2:0] sourceC_task_arb_io_in_13_bits_way; // @[Slice.scala 468:27]
  wire  sourceC_task_arb_io_out_ready; // @[Slice.scala 468:27]
  wire  sourceC_task_arb_io_out_valid; // @[Slice.scala 468:27]
  wire [2:0] sourceC_task_arb_io_out_bits_opcode; // @[Slice.scala 468:27]
  wire [19:0] sourceC_task_arb_io_out_bits_tag; // @[Slice.scala 468:27]
  wire [9:0] sourceC_task_arb_io_out_bits_set; // @[Slice.scala 468:27]
  wire [3:0] sourceC_task_arb_io_out_bits_source; // @[Slice.scala 468:27]
  wire [2:0] sourceC_task_arb_io_out_bits_way; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_clock; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_reset; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_in_0_ready; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_in_0_valid; // @[Slice.scala 468:27]
  wire [5:0] sourceD_task_arb_io_in_0_bits_sourceId; // @[Slice.scala 468:27]
  wire [9:0] sourceD_task_arb_io_in_0_bits_set; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_in_0_bits_channel; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_in_0_bits_opcode; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_in_0_bits_param; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_in_0_bits_size; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_in_0_bits_way; // @[Slice.scala 468:27]
  wire [5:0] sourceD_task_arb_io_in_0_bits_off; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_in_0_bits_useBypass; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_in_0_bits_bufIdx; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_in_0_bits_denied; // @[Slice.scala 468:27]
  wire [3:0] sourceD_task_arb_io_in_0_bits_sinkId; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_in_0_bits_bypassPut; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_in_0_bits_dirty; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_in_1_ready; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_in_1_valid; // @[Slice.scala 468:27]
  wire [5:0] sourceD_task_arb_io_in_1_bits_sourceId; // @[Slice.scala 468:27]
  wire [9:0] sourceD_task_arb_io_in_1_bits_set; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_in_1_bits_channel; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_in_1_bits_opcode; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_in_1_bits_param; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_in_1_bits_size; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_in_1_bits_way; // @[Slice.scala 468:27]
  wire [5:0] sourceD_task_arb_io_in_1_bits_off; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_in_1_bits_useBypass; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_in_1_bits_bufIdx; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_in_1_bits_denied; // @[Slice.scala 468:27]
  wire [3:0] sourceD_task_arb_io_in_1_bits_sinkId; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_in_1_bits_bypassPut; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_in_1_bits_dirty; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_in_2_ready; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_in_2_valid; // @[Slice.scala 468:27]
  wire [5:0] sourceD_task_arb_io_in_2_bits_sourceId; // @[Slice.scala 468:27]
  wire [9:0] sourceD_task_arb_io_in_2_bits_set; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_in_2_bits_channel; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_in_2_bits_opcode; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_in_2_bits_param; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_in_2_bits_size; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_in_2_bits_way; // @[Slice.scala 468:27]
  wire [5:0] sourceD_task_arb_io_in_2_bits_off; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_in_2_bits_useBypass; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_in_2_bits_bufIdx; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_in_2_bits_denied; // @[Slice.scala 468:27]
  wire [3:0] sourceD_task_arb_io_in_2_bits_sinkId; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_in_2_bits_bypassPut; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_in_2_bits_dirty; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_in_3_ready; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_in_3_valid; // @[Slice.scala 468:27]
  wire [5:0] sourceD_task_arb_io_in_3_bits_sourceId; // @[Slice.scala 468:27]
  wire [9:0] sourceD_task_arb_io_in_3_bits_set; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_in_3_bits_channel; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_in_3_bits_opcode; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_in_3_bits_param; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_in_3_bits_size; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_in_3_bits_way; // @[Slice.scala 468:27]
  wire [5:0] sourceD_task_arb_io_in_3_bits_off; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_in_3_bits_useBypass; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_in_3_bits_bufIdx; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_in_3_bits_denied; // @[Slice.scala 468:27]
  wire [3:0] sourceD_task_arb_io_in_3_bits_sinkId; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_in_3_bits_bypassPut; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_in_3_bits_dirty; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_in_4_ready; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_in_4_valid; // @[Slice.scala 468:27]
  wire [5:0] sourceD_task_arb_io_in_4_bits_sourceId; // @[Slice.scala 468:27]
  wire [9:0] sourceD_task_arb_io_in_4_bits_set; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_in_4_bits_channel; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_in_4_bits_opcode; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_in_4_bits_param; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_in_4_bits_size; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_in_4_bits_way; // @[Slice.scala 468:27]
  wire [5:0] sourceD_task_arb_io_in_4_bits_off; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_in_4_bits_useBypass; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_in_4_bits_bufIdx; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_in_4_bits_denied; // @[Slice.scala 468:27]
  wire [3:0] sourceD_task_arb_io_in_4_bits_sinkId; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_in_4_bits_bypassPut; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_in_4_bits_dirty; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_in_5_ready; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_in_5_valid; // @[Slice.scala 468:27]
  wire [5:0] sourceD_task_arb_io_in_5_bits_sourceId; // @[Slice.scala 468:27]
  wire [9:0] sourceD_task_arb_io_in_5_bits_set; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_in_5_bits_channel; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_in_5_bits_opcode; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_in_5_bits_param; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_in_5_bits_size; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_in_5_bits_way; // @[Slice.scala 468:27]
  wire [5:0] sourceD_task_arb_io_in_5_bits_off; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_in_5_bits_useBypass; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_in_5_bits_bufIdx; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_in_5_bits_denied; // @[Slice.scala 468:27]
  wire [3:0] sourceD_task_arb_io_in_5_bits_sinkId; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_in_5_bits_bypassPut; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_in_5_bits_dirty; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_in_6_ready; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_in_6_valid; // @[Slice.scala 468:27]
  wire [5:0] sourceD_task_arb_io_in_6_bits_sourceId; // @[Slice.scala 468:27]
  wire [9:0] sourceD_task_arb_io_in_6_bits_set; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_in_6_bits_channel; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_in_6_bits_opcode; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_in_6_bits_param; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_in_6_bits_size; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_in_6_bits_way; // @[Slice.scala 468:27]
  wire [5:0] sourceD_task_arb_io_in_6_bits_off; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_in_6_bits_useBypass; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_in_6_bits_bufIdx; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_in_6_bits_denied; // @[Slice.scala 468:27]
  wire [3:0] sourceD_task_arb_io_in_6_bits_sinkId; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_in_6_bits_bypassPut; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_in_6_bits_dirty; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_in_7_ready; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_in_7_valid; // @[Slice.scala 468:27]
  wire [5:0] sourceD_task_arb_io_in_7_bits_sourceId; // @[Slice.scala 468:27]
  wire [9:0] sourceD_task_arb_io_in_7_bits_set; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_in_7_bits_channel; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_in_7_bits_opcode; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_in_7_bits_param; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_in_7_bits_size; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_in_7_bits_way; // @[Slice.scala 468:27]
  wire [5:0] sourceD_task_arb_io_in_7_bits_off; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_in_7_bits_useBypass; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_in_7_bits_bufIdx; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_in_7_bits_denied; // @[Slice.scala 468:27]
  wire [3:0] sourceD_task_arb_io_in_7_bits_sinkId; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_in_7_bits_bypassPut; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_in_7_bits_dirty; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_in_8_ready; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_in_8_valid; // @[Slice.scala 468:27]
  wire [5:0] sourceD_task_arb_io_in_8_bits_sourceId; // @[Slice.scala 468:27]
  wire [9:0] sourceD_task_arb_io_in_8_bits_set; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_in_8_bits_channel; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_in_8_bits_opcode; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_in_8_bits_param; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_in_8_bits_size; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_in_8_bits_way; // @[Slice.scala 468:27]
  wire [5:0] sourceD_task_arb_io_in_8_bits_off; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_in_8_bits_useBypass; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_in_8_bits_bufIdx; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_in_8_bits_denied; // @[Slice.scala 468:27]
  wire [3:0] sourceD_task_arb_io_in_8_bits_sinkId; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_in_8_bits_bypassPut; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_in_8_bits_dirty; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_in_9_ready; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_in_9_valid; // @[Slice.scala 468:27]
  wire [5:0] sourceD_task_arb_io_in_9_bits_sourceId; // @[Slice.scala 468:27]
  wire [9:0] sourceD_task_arb_io_in_9_bits_set; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_in_9_bits_channel; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_in_9_bits_opcode; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_in_9_bits_param; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_in_9_bits_size; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_in_9_bits_way; // @[Slice.scala 468:27]
  wire [5:0] sourceD_task_arb_io_in_9_bits_off; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_in_9_bits_useBypass; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_in_9_bits_bufIdx; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_in_9_bits_denied; // @[Slice.scala 468:27]
  wire [3:0] sourceD_task_arb_io_in_9_bits_sinkId; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_in_9_bits_bypassPut; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_in_9_bits_dirty; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_in_10_ready; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_in_10_valid; // @[Slice.scala 468:27]
  wire [5:0] sourceD_task_arb_io_in_10_bits_sourceId; // @[Slice.scala 468:27]
  wire [9:0] sourceD_task_arb_io_in_10_bits_set; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_in_10_bits_channel; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_in_10_bits_opcode; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_in_10_bits_param; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_in_10_bits_size; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_in_10_bits_way; // @[Slice.scala 468:27]
  wire [5:0] sourceD_task_arb_io_in_10_bits_off; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_in_10_bits_useBypass; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_in_10_bits_bufIdx; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_in_10_bits_denied; // @[Slice.scala 468:27]
  wire [3:0] sourceD_task_arb_io_in_10_bits_sinkId; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_in_10_bits_bypassPut; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_in_10_bits_dirty; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_in_11_ready; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_in_11_valid; // @[Slice.scala 468:27]
  wire [5:0] sourceD_task_arb_io_in_11_bits_sourceId; // @[Slice.scala 468:27]
  wire [9:0] sourceD_task_arb_io_in_11_bits_set; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_in_11_bits_channel; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_in_11_bits_opcode; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_in_11_bits_param; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_in_11_bits_size; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_in_11_bits_way; // @[Slice.scala 468:27]
  wire [5:0] sourceD_task_arb_io_in_11_bits_off; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_in_11_bits_useBypass; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_in_11_bits_bufIdx; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_in_11_bits_denied; // @[Slice.scala 468:27]
  wire [3:0] sourceD_task_arb_io_in_11_bits_sinkId; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_in_11_bits_bypassPut; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_in_11_bits_dirty; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_in_12_ready; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_in_12_valid; // @[Slice.scala 468:27]
  wire [5:0] sourceD_task_arb_io_in_12_bits_sourceId; // @[Slice.scala 468:27]
  wire [9:0] sourceD_task_arb_io_in_12_bits_set; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_in_12_bits_channel; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_in_12_bits_opcode; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_in_12_bits_param; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_in_12_bits_size; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_in_12_bits_way; // @[Slice.scala 468:27]
  wire [5:0] sourceD_task_arb_io_in_12_bits_off; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_in_12_bits_useBypass; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_in_12_bits_bufIdx; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_in_12_bits_denied; // @[Slice.scala 468:27]
  wire [3:0] sourceD_task_arb_io_in_12_bits_sinkId; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_in_12_bits_bypassPut; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_in_12_bits_dirty; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_in_13_ready; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_in_13_valid; // @[Slice.scala 468:27]
  wire [5:0] sourceD_task_arb_io_in_13_bits_sourceId; // @[Slice.scala 468:27]
  wire [9:0] sourceD_task_arb_io_in_13_bits_set; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_in_13_bits_channel; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_in_13_bits_opcode; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_in_13_bits_param; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_in_13_bits_size; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_in_13_bits_way; // @[Slice.scala 468:27]
  wire [5:0] sourceD_task_arb_io_in_13_bits_off; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_in_13_bits_useBypass; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_in_13_bits_bufIdx; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_in_13_bits_denied; // @[Slice.scala 468:27]
  wire [3:0] sourceD_task_arb_io_in_13_bits_sinkId; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_in_13_bits_bypassPut; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_in_13_bits_dirty; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_out_ready; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_out_valid; // @[Slice.scala 468:27]
  wire [5:0] sourceD_task_arb_io_out_bits_sourceId; // @[Slice.scala 468:27]
  wire [9:0] sourceD_task_arb_io_out_bits_set; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_out_bits_channel; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_out_bits_opcode; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_out_bits_param; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_out_bits_size; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_out_bits_way; // @[Slice.scala 468:27]
  wire [5:0] sourceD_task_arb_io_out_bits_off; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_out_bits_useBypass; // @[Slice.scala 468:27]
  wire [2:0] sourceD_task_arb_io_out_bits_bufIdx; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_out_bits_denied; // @[Slice.scala 468:27]
  wire [3:0] sourceD_task_arb_io_out_bits_sinkId; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_out_bits_bypassPut; // @[Slice.scala 468:27]
  wire  sourceD_task_arb_io_out_bits_dirty; // @[Slice.scala 468:27]
  wire  sourceE_task_arb_clock; // @[Slice.scala 468:27]
  wire  sourceE_task_arb_reset; // @[Slice.scala 468:27]
  wire  sourceE_task_arb_io_in_0_ready; // @[Slice.scala 468:27]
  wire  sourceE_task_arb_io_in_0_valid; // @[Slice.scala 468:27]
  wire [2:0] sourceE_task_arb_io_in_0_bits_sink; // @[Slice.scala 468:27]
  wire  sourceE_task_arb_io_in_1_ready; // @[Slice.scala 468:27]
  wire  sourceE_task_arb_io_in_1_valid; // @[Slice.scala 468:27]
  wire [2:0] sourceE_task_arb_io_in_1_bits_sink; // @[Slice.scala 468:27]
  wire  sourceE_task_arb_io_in_2_ready; // @[Slice.scala 468:27]
  wire  sourceE_task_arb_io_in_2_valid; // @[Slice.scala 468:27]
  wire [2:0] sourceE_task_arb_io_in_2_bits_sink; // @[Slice.scala 468:27]
  wire  sourceE_task_arb_io_in_3_ready; // @[Slice.scala 468:27]
  wire  sourceE_task_arb_io_in_3_valid; // @[Slice.scala 468:27]
  wire [2:0] sourceE_task_arb_io_in_3_bits_sink; // @[Slice.scala 468:27]
  wire  sourceE_task_arb_io_in_4_ready; // @[Slice.scala 468:27]
  wire  sourceE_task_arb_io_in_4_valid; // @[Slice.scala 468:27]
  wire [2:0] sourceE_task_arb_io_in_4_bits_sink; // @[Slice.scala 468:27]
  wire  sourceE_task_arb_io_in_5_ready; // @[Slice.scala 468:27]
  wire  sourceE_task_arb_io_in_5_valid; // @[Slice.scala 468:27]
  wire [2:0] sourceE_task_arb_io_in_5_bits_sink; // @[Slice.scala 468:27]
  wire  sourceE_task_arb_io_in_6_ready; // @[Slice.scala 468:27]
  wire  sourceE_task_arb_io_in_6_valid; // @[Slice.scala 468:27]
  wire [2:0] sourceE_task_arb_io_in_6_bits_sink; // @[Slice.scala 468:27]
  wire  sourceE_task_arb_io_in_7_ready; // @[Slice.scala 468:27]
  wire  sourceE_task_arb_io_in_7_valid; // @[Slice.scala 468:27]
  wire [2:0] sourceE_task_arb_io_in_7_bits_sink; // @[Slice.scala 468:27]
  wire  sourceE_task_arb_io_in_8_ready; // @[Slice.scala 468:27]
  wire  sourceE_task_arb_io_in_8_valid; // @[Slice.scala 468:27]
  wire [2:0] sourceE_task_arb_io_in_8_bits_sink; // @[Slice.scala 468:27]
  wire  sourceE_task_arb_io_in_9_ready; // @[Slice.scala 468:27]
  wire  sourceE_task_arb_io_in_9_valid; // @[Slice.scala 468:27]
  wire [2:0] sourceE_task_arb_io_in_9_bits_sink; // @[Slice.scala 468:27]
  wire  sourceE_task_arb_io_in_10_ready; // @[Slice.scala 468:27]
  wire  sourceE_task_arb_io_in_10_valid; // @[Slice.scala 468:27]
  wire [2:0] sourceE_task_arb_io_in_10_bits_sink; // @[Slice.scala 468:27]
  wire  sourceE_task_arb_io_in_11_ready; // @[Slice.scala 468:27]
  wire  sourceE_task_arb_io_in_11_valid; // @[Slice.scala 468:27]
  wire [2:0] sourceE_task_arb_io_in_11_bits_sink; // @[Slice.scala 468:27]
  wire  sourceE_task_arb_io_in_12_ready; // @[Slice.scala 468:27]
  wire  sourceE_task_arb_io_in_12_valid; // @[Slice.scala 468:27]
  wire [2:0] sourceE_task_arb_io_in_12_bits_sink; // @[Slice.scala 468:27]
  wire  sourceE_task_arb_io_in_13_ready; // @[Slice.scala 468:27]
  wire  sourceE_task_arb_io_in_13_valid; // @[Slice.scala 468:27]
  wire [2:0] sourceE_task_arb_io_in_13_bits_sink; // @[Slice.scala 468:27]
  wire  sourceE_task_arb_io_out_ready; // @[Slice.scala 468:27]
  wire  sourceE_task_arb_io_out_valid; // @[Slice.scala 468:27]
  wire [2:0] sourceE_task_arb_io_out_bits_sink; // @[Slice.scala 468:27]
  wire  sinkC_task_arb_clock; // @[Slice.scala 468:27]
  wire  sinkC_task_arb_reset; // @[Slice.scala 468:27]
  wire  sinkC_task_arb_io_in_0_ready; // @[Slice.scala 468:27]
  wire  sinkC_task_arb_io_in_0_valid; // @[Slice.scala 468:27]
  wire [9:0] sinkC_task_arb_io_in_0_bits_set; // @[Slice.scala 468:27]
  wire [19:0] sinkC_task_arb_io_in_0_bits_tag; // @[Slice.scala 468:27]
  wire [2:0] sinkC_task_arb_io_in_0_bits_way; // @[Slice.scala 468:27]
  wire [2:0] sinkC_task_arb_io_in_0_bits_bufIdx; // @[Slice.scala 468:27]
  wire [2:0] sinkC_task_arb_io_in_0_bits_opcode; // @[Slice.scala 468:27]
  wire [3:0] sinkC_task_arb_io_in_0_bits_source; // @[Slice.scala 468:27]
  wire  sinkC_task_arb_io_in_0_bits_save; // @[Slice.scala 468:27]
  wire  sinkC_task_arb_io_in_0_bits_drop; // @[Slice.scala 468:27]
  wire  sinkC_task_arb_io_in_0_bits_release; // @[Slice.scala 468:27]
  wire  sinkC_task_arb_io_in_1_ready; // @[Slice.scala 468:27]
  wire  sinkC_task_arb_io_in_1_valid; // @[Slice.scala 468:27]
  wire [9:0] sinkC_task_arb_io_in_1_bits_set; // @[Slice.scala 468:27]
  wire [19:0] sinkC_task_arb_io_in_1_bits_tag; // @[Slice.scala 468:27]
  wire [2:0] sinkC_task_arb_io_in_1_bits_way; // @[Slice.scala 468:27]
  wire [2:0] sinkC_task_arb_io_in_1_bits_bufIdx; // @[Slice.scala 468:27]
  wire [2:0] sinkC_task_arb_io_in_1_bits_opcode; // @[Slice.scala 468:27]
  wire [3:0] sinkC_task_arb_io_in_1_bits_source; // @[Slice.scala 468:27]
  wire  sinkC_task_arb_io_in_1_bits_save; // @[Slice.scala 468:27]
  wire  sinkC_task_arb_io_in_1_bits_drop; // @[Slice.scala 468:27]
  wire  sinkC_task_arb_io_in_1_bits_release; // @[Slice.scala 468:27]
  wire  sinkC_task_arb_io_in_2_ready; // @[Slice.scala 468:27]
  wire  sinkC_task_arb_io_in_2_valid; // @[Slice.scala 468:27]
  wire [9:0] sinkC_task_arb_io_in_2_bits_set; // @[Slice.scala 468:27]
  wire [19:0] sinkC_task_arb_io_in_2_bits_tag; // @[Slice.scala 468:27]
  wire [2:0] sinkC_task_arb_io_in_2_bits_way; // @[Slice.scala 468:27]
  wire [2:0] sinkC_task_arb_io_in_2_bits_bufIdx; // @[Slice.scala 468:27]
  wire [2:0] sinkC_task_arb_io_in_2_bits_opcode; // @[Slice.scala 468:27]
  wire [3:0] sinkC_task_arb_io_in_2_bits_source; // @[Slice.scala 468:27]
  wire  sinkC_task_arb_io_in_2_bits_save; // @[Slice.scala 468:27]
  wire  sinkC_task_arb_io_in_2_bits_drop; // @[Slice.scala 468:27]
  wire  sinkC_task_arb_io_in_2_bits_release; // @[Slice.scala 468:27]
  wire  sinkC_task_arb_io_in_3_ready; // @[Slice.scala 468:27]
  wire  sinkC_task_arb_io_in_3_valid; // @[Slice.scala 468:27]
  wire [9:0] sinkC_task_arb_io_in_3_bits_set; // @[Slice.scala 468:27]
  wire [19:0] sinkC_task_arb_io_in_3_bits_tag; // @[Slice.scala 468:27]
  wire [2:0] sinkC_task_arb_io_in_3_bits_way; // @[Slice.scala 468:27]
  wire [2:0] sinkC_task_arb_io_in_3_bits_bufIdx; // @[Slice.scala 468:27]
  wire [2:0] sinkC_task_arb_io_in_3_bits_opcode; // @[Slice.scala 468:27]
  wire [3:0] sinkC_task_arb_io_in_3_bits_source; // @[Slice.scala 468:27]
  wire  sinkC_task_arb_io_in_3_bits_save; // @[Slice.scala 468:27]
  wire  sinkC_task_arb_io_in_3_bits_drop; // @[Slice.scala 468:27]
  wire  sinkC_task_arb_io_in_3_bits_release; // @[Slice.scala 468:27]
  wire  sinkC_task_arb_io_in_4_ready; // @[Slice.scala 468:27]
  wire  sinkC_task_arb_io_in_4_valid; // @[Slice.scala 468:27]
  wire [9:0] sinkC_task_arb_io_in_4_bits_set; // @[Slice.scala 468:27]
  wire [19:0] sinkC_task_arb_io_in_4_bits_tag; // @[Slice.scala 468:27]
  wire [2:0] sinkC_task_arb_io_in_4_bits_way; // @[Slice.scala 468:27]
  wire [2:0] sinkC_task_arb_io_in_4_bits_bufIdx; // @[Slice.scala 468:27]
  wire [2:0] sinkC_task_arb_io_in_4_bits_opcode; // @[Slice.scala 468:27]
  wire [3:0] sinkC_task_arb_io_in_4_bits_source; // @[Slice.scala 468:27]
  wire  sinkC_task_arb_io_in_4_bits_save; // @[Slice.scala 468:27]
  wire  sinkC_task_arb_io_in_4_bits_drop; // @[Slice.scala 468:27]
  wire  sinkC_task_arb_io_in_4_bits_release; // @[Slice.scala 468:27]
  wire  sinkC_task_arb_io_in_5_ready; // @[Slice.scala 468:27]
  wire  sinkC_task_arb_io_in_5_valid; // @[Slice.scala 468:27]
  wire [9:0] sinkC_task_arb_io_in_5_bits_set; // @[Slice.scala 468:27]
  wire [19:0] sinkC_task_arb_io_in_5_bits_tag; // @[Slice.scala 468:27]
  wire [2:0] sinkC_task_arb_io_in_5_bits_way; // @[Slice.scala 468:27]
  wire [2:0] sinkC_task_arb_io_in_5_bits_bufIdx; // @[Slice.scala 468:27]
  wire [2:0] sinkC_task_arb_io_in_5_bits_opcode; // @[Slice.scala 468:27]
  wire [3:0] sinkC_task_arb_io_in_5_bits_source; // @[Slice.scala 468:27]
  wire  sinkC_task_arb_io_in_5_bits_save; // @[Slice.scala 468:27]
  wire  sinkC_task_arb_io_in_5_bits_drop; // @[Slice.scala 468:27]
  wire  sinkC_task_arb_io_in_5_bits_release; // @[Slice.scala 468:27]
  wire  sinkC_task_arb_io_in_6_ready; // @[Slice.scala 468:27]
  wire  sinkC_task_arb_io_in_6_valid; // @[Slice.scala 468:27]
  wire [9:0] sinkC_task_arb_io_in_6_bits_set; // @[Slice.scala 468:27]
  wire [19:0] sinkC_task_arb_io_in_6_bits_tag; // @[Slice.scala 468:27]
  wire [2:0] sinkC_task_arb_io_in_6_bits_way; // @[Slice.scala 468:27]
  wire [2:0] sinkC_task_arb_io_in_6_bits_bufIdx; // @[Slice.scala 468:27]
  wire [2:0] sinkC_task_arb_io_in_6_bits_opcode; // @[Slice.scala 468:27]
  wire [3:0] sinkC_task_arb_io_in_6_bits_source; // @[Slice.scala 468:27]
  wire  sinkC_task_arb_io_in_6_bits_save; // @[Slice.scala 468:27]
  wire  sinkC_task_arb_io_in_6_bits_drop; // @[Slice.scala 468:27]
  wire  sinkC_task_arb_io_in_6_bits_release; // @[Slice.scala 468:27]
  wire  sinkC_task_arb_io_in_7_ready; // @[Slice.scala 468:27]
  wire  sinkC_task_arb_io_in_7_valid; // @[Slice.scala 468:27]
  wire [9:0] sinkC_task_arb_io_in_7_bits_set; // @[Slice.scala 468:27]
  wire [19:0] sinkC_task_arb_io_in_7_bits_tag; // @[Slice.scala 468:27]
  wire [2:0] sinkC_task_arb_io_in_7_bits_way; // @[Slice.scala 468:27]
  wire [2:0] sinkC_task_arb_io_in_7_bits_bufIdx; // @[Slice.scala 468:27]
  wire [2:0] sinkC_task_arb_io_in_7_bits_opcode; // @[Slice.scala 468:27]
  wire [3:0] sinkC_task_arb_io_in_7_bits_source; // @[Slice.scala 468:27]
  wire  sinkC_task_arb_io_in_7_bits_save; // @[Slice.scala 468:27]
  wire  sinkC_task_arb_io_in_7_bits_drop; // @[Slice.scala 468:27]
  wire  sinkC_task_arb_io_in_7_bits_release; // @[Slice.scala 468:27]
  wire  sinkC_task_arb_io_in_8_ready; // @[Slice.scala 468:27]
  wire  sinkC_task_arb_io_in_8_valid; // @[Slice.scala 468:27]
  wire [9:0] sinkC_task_arb_io_in_8_bits_set; // @[Slice.scala 468:27]
  wire [19:0] sinkC_task_arb_io_in_8_bits_tag; // @[Slice.scala 468:27]
  wire [2:0] sinkC_task_arb_io_in_8_bits_way; // @[Slice.scala 468:27]
  wire [2:0] sinkC_task_arb_io_in_8_bits_bufIdx; // @[Slice.scala 468:27]
  wire [2:0] sinkC_task_arb_io_in_8_bits_opcode; // @[Slice.scala 468:27]
  wire [3:0] sinkC_task_arb_io_in_8_bits_source; // @[Slice.scala 468:27]
  wire  sinkC_task_arb_io_in_8_bits_save; // @[Slice.scala 468:27]
  wire  sinkC_task_arb_io_in_8_bits_drop; // @[Slice.scala 468:27]
  wire  sinkC_task_arb_io_in_8_bits_release; // @[Slice.scala 468:27]
  wire  sinkC_task_arb_io_in_9_ready; // @[Slice.scala 468:27]
  wire  sinkC_task_arb_io_in_9_valid; // @[Slice.scala 468:27]
  wire [9:0] sinkC_task_arb_io_in_9_bits_set; // @[Slice.scala 468:27]
  wire [19:0] sinkC_task_arb_io_in_9_bits_tag; // @[Slice.scala 468:27]
  wire [2:0] sinkC_task_arb_io_in_9_bits_way; // @[Slice.scala 468:27]
  wire [2:0] sinkC_task_arb_io_in_9_bits_bufIdx; // @[Slice.scala 468:27]
  wire [2:0] sinkC_task_arb_io_in_9_bits_opcode; // @[Slice.scala 468:27]
  wire [3:0] sinkC_task_arb_io_in_9_bits_source; // @[Slice.scala 468:27]
  wire  sinkC_task_arb_io_in_9_bits_save; // @[Slice.scala 468:27]
  wire  sinkC_task_arb_io_in_9_bits_drop; // @[Slice.scala 468:27]
  wire  sinkC_task_arb_io_in_9_bits_release; // @[Slice.scala 468:27]
  wire  sinkC_task_arb_io_in_10_ready; // @[Slice.scala 468:27]
  wire  sinkC_task_arb_io_in_10_valid; // @[Slice.scala 468:27]
  wire [9:0] sinkC_task_arb_io_in_10_bits_set; // @[Slice.scala 468:27]
  wire [19:0] sinkC_task_arb_io_in_10_bits_tag; // @[Slice.scala 468:27]
  wire [2:0] sinkC_task_arb_io_in_10_bits_way; // @[Slice.scala 468:27]
  wire [2:0] sinkC_task_arb_io_in_10_bits_bufIdx; // @[Slice.scala 468:27]
  wire [2:0] sinkC_task_arb_io_in_10_bits_opcode; // @[Slice.scala 468:27]
  wire [3:0] sinkC_task_arb_io_in_10_bits_source; // @[Slice.scala 468:27]
  wire  sinkC_task_arb_io_in_10_bits_save; // @[Slice.scala 468:27]
  wire  sinkC_task_arb_io_in_10_bits_drop; // @[Slice.scala 468:27]
  wire  sinkC_task_arb_io_in_10_bits_release; // @[Slice.scala 468:27]
  wire  sinkC_task_arb_io_in_11_ready; // @[Slice.scala 468:27]
  wire  sinkC_task_arb_io_in_11_valid; // @[Slice.scala 468:27]
  wire [9:0] sinkC_task_arb_io_in_11_bits_set; // @[Slice.scala 468:27]
  wire [19:0] sinkC_task_arb_io_in_11_bits_tag; // @[Slice.scala 468:27]
  wire [2:0] sinkC_task_arb_io_in_11_bits_way; // @[Slice.scala 468:27]
  wire [2:0] sinkC_task_arb_io_in_11_bits_bufIdx; // @[Slice.scala 468:27]
  wire [2:0] sinkC_task_arb_io_in_11_bits_opcode; // @[Slice.scala 468:27]
  wire [3:0] sinkC_task_arb_io_in_11_bits_source; // @[Slice.scala 468:27]
  wire  sinkC_task_arb_io_in_11_bits_save; // @[Slice.scala 468:27]
  wire  sinkC_task_arb_io_in_11_bits_drop; // @[Slice.scala 468:27]
  wire  sinkC_task_arb_io_in_11_bits_release; // @[Slice.scala 468:27]
  wire  sinkC_task_arb_io_in_12_ready; // @[Slice.scala 468:27]
  wire  sinkC_task_arb_io_in_12_valid; // @[Slice.scala 468:27]
  wire [9:0] sinkC_task_arb_io_in_12_bits_set; // @[Slice.scala 468:27]
  wire [19:0] sinkC_task_arb_io_in_12_bits_tag; // @[Slice.scala 468:27]
  wire [2:0] sinkC_task_arb_io_in_12_bits_way; // @[Slice.scala 468:27]
  wire [2:0] sinkC_task_arb_io_in_12_bits_bufIdx; // @[Slice.scala 468:27]
  wire [2:0] sinkC_task_arb_io_in_12_bits_opcode; // @[Slice.scala 468:27]
  wire [3:0] sinkC_task_arb_io_in_12_bits_source; // @[Slice.scala 468:27]
  wire  sinkC_task_arb_io_in_12_bits_save; // @[Slice.scala 468:27]
  wire  sinkC_task_arb_io_in_12_bits_drop; // @[Slice.scala 468:27]
  wire  sinkC_task_arb_io_in_12_bits_release; // @[Slice.scala 468:27]
  wire  sinkC_task_arb_io_in_13_ready; // @[Slice.scala 468:27]
  wire  sinkC_task_arb_io_in_13_valid; // @[Slice.scala 468:27]
  wire [9:0] sinkC_task_arb_io_in_13_bits_set; // @[Slice.scala 468:27]
  wire [19:0] sinkC_task_arb_io_in_13_bits_tag; // @[Slice.scala 468:27]
  wire [2:0] sinkC_task_arb_io_in_13_bits_way; // @[Slice.scala 468:27]
  wire [2:0] sinkC_task_arb_io_in_13_bits_bufIdx; // @[Slice.scala 468:27]
  wire [2:0] sinkC_task_arb_io_in_13_bits_opcode; // @[Slice.scala 468:27]
  wire [3:0] sinkC_task_arb_io_in_13_bits_source; // @[Slice.scala 468:27]
  wire  sinkC_task_arb_io_in_13_bits_save; // @[Slice.scala 468:27]
  wire  sinkC_task_arb_io_in_13_bits_drop; // @[Slice.scala 468:27]
  wire  sinkC_task_arb_io_in_13_bits_release; // @[Slice.scala 468:27]
  wire  sinkC_task_arb_io_out_ready; // @[Slice.scala 468:27]
  wire  sinkC_task_arb_io_out_valid; // @[Slice.scala 468:27]
  wire [9:0] sinkC_task_arb_io_out_bits_set; // @[Slice.scala 468:27]
  wire [19:0] sinkC_task_arb_io_out_bits_tag; // @[Slice.scala 468:27]
  wire [2:0] sinkC_task_arb_io_out_bits_way; // @[Slice.scala 468:27]
  wire [2:0] sinkC_task_arb_io_out_bits_bufIdx; // @[Slice.scala 468:27]
  wire [2:0] sinkC_task_arb_io_out_bits_opcode; // @[Slice.scala 468:27]
  wire [3:0] sinkC_task_arb_io_out_bits_source; // @[Slice.scala 468:27]
  wire  sinkC_task_arb_io_out_bits_save; // @[Slice.scala 468:27]
  wire  sinkC_task_arb_io_out_bits_drop; // @[Slice.scala 468:27]
  wire  sinkC_task_arb_io_out_bits_release; // @[Slice.scala 468:27]
  wire  pipeline_1_clock; // @[Pipeline.scala 39:26]
  wire  pipeline_1_reset; // @[Pipeline.scala 39:26]
  wire  pipeline_1_io_in_valid; // @[Pipeline.scala 39:26]
  wire [9:0] pipeline_1_io_in_bits_set; // @[Pipeline.scala 39:26]
  wire [2:0] pipeline_1_io_in_bits_way; // @[Pipeline.scala 39:26]
  wire [19:0] pipeline_1_io_in_bits_tag; // @[Pipeline.scala 39:26]
  wire  pipeline_1_io_out_valid; // @[Pipeline.scala 39:26]
  wire [9:0] pipeline_1_io_out_bits_set; // @[Pipeline.scala 39:26]
  wire [2:0] pipeline_1_io_out_bits_way; // @[Pipeline.scala 39:26]
  wire [19:0] pipeline_1_io_out_bits_tag; // @[Pipeline.scala 39:26]
  wire  tagWrite_task_arb_clock; // @[Slice.scala 468:27]
  wire  tagWrite_task_arb_reset; // @[Slice.scala 468:27]
  wire  tagWrite_task_arb_io_in_0_ready; // @[Slice.scala 468:27]
  wire  tagWrite_task_arb_io_in_0_valid; // @[Slice.scala 468:27]
  wire [9:0] tagWrite_task_arb_io_in_0_bits_set; // @[Slice.scala 468:27]
  wire [2:0] tagWrite_task_arb_io_in_0_bits_way; // @[Slice.scala 468:27]
  wire [19:0] tagWrite_task_arb_io_in_0_bits_tag; // @[Slice.scala 468:27]
  wire  tagWrite_task_arb_io_in_1_ready; // @[Slice.scala 468:27]
  wire  tagWrite_task_arb_io_in_1_valid; // @[Slice.scala 468:27]
  wire [9:0] tagWrite_task_arb_io_in_1_bits_set; // @[Slice.scala 468:27]
  wire [2:0] tagWrite_task_arb_io_in_1_bits_way; // @[Slice.scala 468:27]
  wire [19:0] tagWrite_task_arb_io_in_1_bits_tag; // @[Slice.scala 468:27]
  wire  tagWrite_task_arb_io_in_2_ready; // @[Slice.scala 468:27]
  wire  tagWrite_task_arb_io_in_2_valid; // @[Slice.scala 468:27]
  wire [9:0] tagWrite_task_arb_io_in_2_bits_set; // @[Slice.scala 468:27]
  wire [2:0] tagWrite_task_arb_io_in_2_bits_way; // @[Slice.scala 468:27]
  wire [19:0] tagWrite_task_arb_io_in_2_bits_tag; // @[Slice.scala 468:27]
  wire  tagWrite_task_arb_io_in_3_ready; // @[Slice.scala 468:27]
  wire  tagWrite_task_arb_io_in_3_valid; // @[Slice.scala 468:27]
  wire [9:0] tagWrite_task_arb_io_in_3_bits_set; // @[Slice.scala 468:27]
  wire [2:0] tagWrite_task_arb_io_in_3_bits_way; // @[Slice.scala 468:27]
  wire [19:0] tagWrite_task_arb_io_in_3_bits_tag; // @[Slice.scala 468:27]
  wire  tagWrite_task_arb_io_in_4_ready; // @[Slice.scala 468:27]
  wire  tagWrite_task_arb_io_in_4_valid; // @[Slice.scala 468:27]
  wire [9:0] tagWrite_task_arb_io_in_4_bits_set; // @[Slice.scala 468:27]
  wire [2:0] tagWrite_task_arb_io_in_4_bits_way; // @[Slice.scala 468:27]
  wire [19:0] tagWrite_task_arb_io_in_4_bits_tag; // @[Slice.scala 468:27]
  wire  tagWrite_task_arb_io_in_5_ready; // @[Slice.scala 468:27]
  wire  tagWrite_task_arb_io_in_5_valid; // @[Slice.scala 468:27]
  wire [9:0] tagWrite_task_arb_io_in_5_bits_set; // @[Slice.scala 468:27]
  wire [2:0] tagWrite_task_arb_io_in_5_bits_way; // @[Slice.scala 468:27]
  wire [19:0] tagWrite_task_arb_io_in_5_bits_tag; // @[Slice.scala 468:27]
  wire  tagWrite_task_arb_io_in_6_ready; // @[Slice.scala 468:27]
  wire  tagWrite_task_arb_io_in_6_valid; // @[Slice.scala 468:27]
  wire [9:0] tagWrite_task_arb_io_in_6_bits_set; // @[Slice.scala 468:27]
  wire [2:0] tagWrite_task_arb_io_in_6_bits_way; // @[Slice.scala 468:27]
  wire [19:0] tagWrite_task_arb_io_in_6_bits_tag; // @[Slice.scala 468:27]
  wire  tagWrite_task_arb_io_in_7_ready; // @[Slice.scala 468:27]
  wire  tagWrite_task_arb_io_in_7_valid; // @[Slice.scala 468:27]
  wire [9:0] tagWrite_task_arb_io_in_7_bits_set; // @[Slice.scala 468:27]
  wire [2:0] tagWrite_task_arb_io_in_7_bits_way; // @[Slice.scala 468:27]
  wire [19:0] tagWrite_task_arb_io_in_7_bits_tag; // @[Slice.scala 468:27]
  wire  tagWrite_task_arb_io_in_8_ready; // @[Slice.scala 468:27]
  wire  tagWrite_task_arb_io_in_8_valid; // @[Slice.scala 468:27]
  wire [9:0] tagWrite_task_arb_io_in_8_bits_set; // @[Slice.scala 468:27]
  wire [2:0] tagWrite_task_arb_io_in_8_bits_way; // @[Slice.scala 468:27]
  wire [19:0] tagWrite_task_arb_io_in_8_bits_tag; // @[Slice.scala 468:27]
  wire  tagWrite_task_arb_io_in_9_ready; // @[Slice.scala 468:27]
  wire  tagWrite_task_arb_io_in_9_valid; // @[Slice.scala 468:27]
  wire [9:0] tagWrite_task_arb_io_in_9_bits_set; // @[Slice.scala 468:27]
  wire [2:0] tagWrite_task_arb_io_in_9_bits_way; // @[Slice.scala 468:27]
  wire [19:0] tagWrite_task_arb_io_in_9_bits_tag; // @[Slice.scala 468:27]
  wire  tagWrite_task_arb_io_in_10_ready; // @[Slice.scala 468:27]
  wire  tagWrite_task_arb_io_in_10_valid; // @[Slice.scala 468:27]
  wire [9:0] tagWrite_task_arb_io_in_10_bits_set; // @[Slice.scala 468:27]
  wire [2:0] tagWrite_task_arb_io_in_10_bits_way; // @[Slice.scala 468:27]
  wire [19:0] tagWrite_task_arb_io_in_10_bits_tag; // @[Slice.scala 468:27]
  wire  tagWrite_task_arb_io_in_11_ready; // @[Slice.scala 468:27]
  wire  tagWrite_task_arb_io_in_11_valid; // @[Slice.scala 468:27]
  wire [9:0] tagWrite_task_arb_io_in_11_bits_set; // @[Slice.scala 468:27]
  wire [2:0] tagWrite_task_arb_io_in_11_bits_way; // @[Slice.scala 468:27]
  wire [19:0] tagWrite_task_arb_io_in_11_bits_tag; // @[Slice.scala 468:27]
  wire  tagWrite_task_arb_io_in_12_ready; // @[Slice.scala 468:27]
  wire  tagWrite_task_arb_io_in_12_valid; // @[Slice.scala 468:27]
  wire [9:0] tagWrite_task_arb_io_in_12_bits_set; // @[Slice.scala 468:27]
  wire [2:0] tagWrite_task_arb_io_in_12_bits_way; // @[Slice.scala 468:27]
  wire [19:0] tagWrite_task_arb_io_in_12_bits_tag; // @[Slice.scala 468:27]
  wire  tagWrite_task_arb_io_in_13_ready; // @[Slice.scala 468:27]
  wire  tagWrite_task_arb_io_in_13_valid; // @[Slice.scala 468:27]
  wire [9:0] tagWrite_task_arb_io_in_13_bits_set; // @[Slice.scala 468:27]
  wire [2:0] tagWrite_task_arb_io_in_13_bits_way; // @[Slice.scala 468:27]
  wire [19:0] tagWrite_task_arb_io_in_13_bits_tag; // @[Slice.scala 468:27]
  wire  tagWrite_task_arb_io_out_ready; // @[Slice.scala 468:27]
  wire  tagWrite_task_arb_io_out_valid; // @[Slice.scala 468:27]
  wire [9:0] tagWrite_task_arb_io_out_bits_set; // @[Slice.scala 468:27]
  wire [2:0] tagWrite_task_arb_io_out_bits_way; // @[Slice.scala 468:27]
  wire [19:0] tagWrite_task_arb_io_out_bits_tag; // @[Slice.scala 468:27]
  wire  pipeline_2_clock; // @[Pipeline.scala 39:26]
  wire  pipeline_2_reset; // @[Pipeline.scala 39:26]
  wire  pipeline_2_io_in_valid; // @[Pipeline.scala 39:26]
  wire [6:0] pipeline_2_io_in_bits_set; // @[Pipeline.scala 39:26]
  wire [3:0] pipeline_2_io_in_bits_way; // @[Pipeline.scala 39:26]
  wire [1:0] pipeline_2_io_in_bits_data_0_state; // @[Pipeline.scala 39:26]
  wire [1:0] pipeline_2_io_in_bits_data_1_state; // @[Pipeline.scala 39:26]
  wire  pipeline_2_io_out_valid; // @[Pipeline.scala 39:26]
  wire [6:0] pipeline_2_io_out_bits_set; // @[Pipeline.scala 39:26]
  wire [3:0] pipeline_2_io_out_bits_way; // @[Pipeline.scala 39:26]
  wire [1:0] pipeline_2_io_out_bits_data_0_state; // @[Pipeline.scala 39:26]
  wire [1:0] pipeline_2_io_out_bits_data_1_state; // @[Pipeline.scala 39:26]
  wire  arbiter_1_clock; // @[Slice.scala 405:25]
  wire  arbiter_1_reset; // @[Slice.scala 405:25]
  wire  arbiter_1_io_in_0_ready; // @[Slice.scala 405:25]
  wire  arbiter_1_io_in_0_valid; // @[Slice.scala 405:25]
  wire [6:0] arbiter_1_io_in_0_bits_set; // @[Slice.scala 405:25]
  wire [3:0] arbiter_1_io_in_0_bits_way; // @[Slice.scala 405:25]
  wire [1:0] arbiter_1_io_in_0_bits_data_0_state; // @[Slice.scala 405:25]
  wire [1:0] arbiter_1_io_in_0_bits_data_1_state; // @[Slice.scala 405:25]
  wire  arbiter_1_io_in_1_ready; // @[Slice.scala 405:25]
  wire  arbiter_1_io_in_1_valid; // @[Slice.scala 405:25]
  wire [6:0] arbiter_1_io_in_1_bits_set; // @[Slice.scala 405:25]
  wire [3:0] arbiter_1_io_in_1_bits_way; // @[Slice.scala 405:25]
  wire [1:0] arbiter_1_io_in_1_bits_data_0_state; // @[Slice.scala 405:25]
  wire [1:0] arbiter_1_io_in_1_bits_data_1_state; // @[Slice.scala 405:25]
  wire  arbiter_1_io_in_2_ready; // @[Slice.scala 405:25]
  wire  arbiter_1_io_in_2_valid; // @[Slice.scala 405:25]
  wire [6:0] arbiter_1_io_in_2_bits_set; // @[Slice.scala 405:25]
  wire [3:0] arbiter_1_io_in_2_bits_way; // @[Slice.scala 405:25]
  wire [1:0] arbiter_1_io_in_2_bits_data_0_state; // @[Slice.scala 405:25]
  wire [1:0] arbiter_1_io_in_2_bits_data_1_state; // @[Slice.scala 405:25]
  wire  arbiter_1_io_in_3_ready; // @[Slice.scala 405:25]
  wire  arbiter_1_io_in_3_valid; // @[Slice.scala 405:25]
  wire [6:0] arbiter_1_io_in_3_bits_set; // @[Slice.scala 405:25]
  wire [3:0] arbiter_1_io_in_3_bits_way; // @[Slice.scala 405:25]
  wire [1:0] arbiter_1_io_in_3_bits_data_0_state; // @[Slice.scala 405:25]
  wire [1:0] arbiter_1_io_in_3_bits_data_1_state; // @[Slice.scala 405:25]
  wire  arbiter_1_io_in_4_ready; // @[Slice.scala 405:25]
  wire  arbiter_1_io_in_4_valid; // @[Slice.scala 405:25]
  wire [6:0] arbiter_1_io_in_4_bits_set; // @[Slice.scala 405:25]
  wire [3:0] arbiter_1_io_in_4_bits_way; // @[Slice.scala 405:25]
  wire [1:0] arbiter_1_io_in_4_bits_data_0_state; // @[Slice.scala 405:25]
  wire [1:0] arbiter_1_io_in_4_bits_data_1_state; // @[Slice.scala 405:25]
  wire  arbiter_1_io_in_5_ready; // @[Slice.scala 405:25]
  wire  arbiter_1_io_in_5_valid; // @[Slice.scala 405:25]
  wire [6:0] arbiter_1_io_in_5_bits_set; // @[Slice.scala 405:25]
  wire [3:0] arbiter_1_io_in_5_bits_way; // @[Slice.scala 405:25]
  wire [1:0] arbiter_1_io_in_5_bits_data_0_state; // @[Slice.scala 405:25]
  wire [1:0] arbiter_1_io_in_5_bits_data_1_state; // @[Slice.scala 405:25]
  wire  arbiter_1_io_in_6_ready; // @[Slice.scala 405:25]
  wire  arbiter_1_io_in_6_valid; // @[Slice.scala 405:25]
  wire [6:0] arbiter_1_io_in_6_bits_set; // @[Slice.scala 405:25]
  wire [3:0] arbiter_1_io_in_6_bits_way; // @[Slice.scala 405:25]
  wire [1:0] arbiter_1_io_in_6_bits_data_0_state; // @[Slice.scala 405:25]
  wire [1:0] arbiter_1_io_in_6_bits_data_1_state; // @[Slice.scala 405:25]
  wire  arbiter_1_io_in_7_ready; // @[Slice.scala 405:25]
  wire  arbiter_1_io_in_7_valid; // @[Slice.scala 405:25]
  wire [6:0] arbiter_1_io_in_7_bits_set; // @[Slice.scala 405:25]
  wire [3:0] arbiter_1_io_in_7_bits_way; // @[Slice.scala 405:25]
  wire [1:0] arbiter_1_io_in_7_bits_data_0_state; // @[Slice.scala 405:25]
  wire [1:0] arbiter_1_io_in_7_bits_data_1_state; // @[Slice.scala 405:25]
  wire  arbiter_1_io_in_8_ready; // @[Slice.scala 405:25]
  wire  arbiter_1_io_in_8_valid; // @[Slice.scala 405:25]
  wire [6:0] arbiter_1_io_in_8_bits_set; // @[Slice.scala 405:25]
  wire [3:0] arbiter_1_io_in_8_bits_way; // @[Slice.scala 405:25]
  wire [1:0] arbiter_1_io_in_8_bits_data_0_state; // @[Slice.scala 405:25]
  wire [1:0] arbiter_1_io_in_8_bits_data_1_state; // @[Slice.scala 405:25]
  wire  arbiter_1_io_in_9_ready; // @[Slice.scala 405:25]
  wire  arbiter_1_io_in_9_valid; // @[Slice.scala 405:25]
  wire [6:0] arbiter_1_io_in_9_bits_set; // @[Slice.scala 405:25]
  wire [3:0] arbiter_1_io_in_9_bits_way; // @[Slice.scala 405:25]
  wire [1:0] arbiter_1_io_in_9_bits_data_0_state; // @[Slice.scala 405:25]
  wire [1:0] arbiter_1_io_in_9_bits_data_1_state; // @[Slice.scala 405:25]
  wire  arbiter_1_io_in_10_ready; // @[Slice.scala 405:25]
  wire  arbiter_1_io_in_10_valid; // @[Slice.scala 405:25]
  wire [6:0] arbiter_1_io_in_10_bits_set; // @[Slice.scala 405:25]
  wire [3:0] arbiter_1_io_in_10_bits_way; // @[Slice.scala 405:25]
  wire [1:0] arbiter_1_io_in_10_bits_data_0_state; // @[Slice.scala 405:25]
  wire [1:0] arbiter_1_io_in_10_bits_data_1_state; // @[Slice.scala 405:25]
  wire  arbiter_1_io_in_11_ready; // @[Slice.scala 405:25]
  wire  arbiter_1_io_in_11_valid; // @[Slice.scala 405:25]
  wire [6:0] arbiter_1_io_in_11_bits_set; // @[Slice.scala 405:25]
  wire [3:0] arbiter_1_io_in_11_bits_way; // @[Slice.scala 405:25]
  wire [1:0] arbiter_1_io_in_11_bits_data_0_state; // @[Slice.scala 405:25]
  wire [1:0] arbiter_1_io_in_11_bits_data_1_state; // @[Slice.scala 405:25]
  wire  arbiter_1_io_in_12_ready; // @[Slice.scala 405:25]
  wire  arbiter_1_io_in_12_valid; // @[Slice.scala 405:25]
  wire [6:0] arbiter_1_io_in_12_bits_set; // @[Slice.scala 405:25]
  wire [3:0] arbiter_1_io_in_12_bits_way; // @[Slice.scala 405:25]
  wire [1:0] arbiter_1_io_in_12_bits_data_0_state; // @[Slice.scala 405:25]
  wire [1:0] arbiter_1_io_in_12_bits_data_1_state; // @[Slice.scala 405:25]
  wire  arbiter_1_io_in_13_ready; // @[Slice.scala 405:25]
  wire  arbiter_1_io_in_13_valid; // @[Slice.scala 405:25]
  wire [6:0] arbiter_1_io_in_13_bits_set; // @[Slice.scala 405:25]
  wire [3:0] arbiter_1_io_in_13_bits_way; // @[Slice.scala 405:25]
  wire [1:0] arbiter_1_io_in_13_bits_data_0_state; // @[Slice.scala 405:25]
  wire [1:0] arbiter_1_io_in_13_bits_data_1_state; // @[Slice.scala 405:25]
  wire  arbiter_1_io_in_14_ready; // @[Slice.scala 405:25]
  wire  arbiter_1_io_in_14_valid; // @[Slice.scala 405:25]
  wire [6:0] arbiter_1_io_in_14_bits_set; // @[Slice.scala 405:25]
  wire [3:0] arbiter_1_io_in_14_bits_way; // @[Slice.scala 405:25]
  wire [1:0] arbiter_1_io_in_14_bits_data_0_state; // @[Slice.scala 405:25]
  wire [1:0] arbiter_1_io_in_14_bits_data_1_state; // @[Slice.scala 405:25]
  wire  arbiter_1_io_in_15_ready; // @[Slice.scala 405:25]
  wire  arbiter_1_io_in_15_valid; // @[Slice.scala 405:25]
  wire [6:0] arbiter_1_io_in_15_bits_set; // @[Slice.scala 405:25]
  wire [3:0] arbiter_1_io_in_15_bits_way; // @[Slice.scala 405:25]
  wire [1:0] arbiter_1_io_in_15_bits_data_0_state; // @[Slice.scala 405:25]
  wire [1:0] arbiter_1_io_in_15_bits_data_1_state; // @[Slice.scala 405:25]
  wire  arbiter_1_io_out_valid; // @[Slice.scala 405:25]
  wire [6:0] arbiter_1_io_out_bits_set; // @[Slice.scala 405:25]
  wire [3:0] arbiter_1_io_out_bits_way; // @[Slice.scala 405:25]
  wire [1:0] arbiter_1_io_out_bits_data_0_state; // @[Slice.scala 405:25]
  wire [1:0] arbiter_1_io_out_bits_data_1_state; // @[Slice.scala 405:25]
  wire  pipeline_3_clock; // @[Pipeline.scala 39:26]
  wire  pipeline_3_reset; // @[Pipeline.scala 39:26]
  wire  pipeline_3_io_in_valid; // @[Pipeline.scala 39:26]
  wire [6:0] pipeline_3_io_in_bits_set; // @[Pipeline.scala 39:26]
  wire [3:0] pipeline_3_io_in_bits_way; // @[Pipeline.scala 39:26]
  wire [22:0] pipeline_3_io_in_bits_tag; // @[Pipeline.scala 39:26]
  wire  pipeline_3_io_out_valid; // @[Pipeline.scala 39:26]
  wire [6:0] pipeline_3_io_out_bits_set; // @[Pipeline.scala 39:26]
  wire [3:0] pipeline_3_io_out_bits_way; // @[Pipeline.scala 39:26]
  wire [22:0] pipeline_3_io_out_bits_tag; // @[Pipeline.scala 39:26]
  wire  arbiter_2_clock; // @[Slice.scala 468:27]
  wire  arbiter_2_reset; // @[Slice.scala 468:27]
  wire  arbiter_2_io_in_0_ready; // @[Slice.scala 468:27]
  wire  arbiter_2_io_in_0_valid; // @[Slice.scala 468:27]
  wire [6:0] arbiter_2_io_in_0_bits_set; // @[Slice.scala 468:27]
  wire [3:0] arbiter_2_io_in_0_bits_way; // @[Slice.scala 468:27]
  wire [22:0] arbiter_2_io_in_0_bits_tag; // @[Slice.scala 468:27]
  wire  arbiter_2_io_in_1_ready; // @[Slice.scala 468:27]
  wire  arbiter_2_io_in_1_valid; // @[Slice.scala 468:27]
  wire [6:0] arbiter_2_io_in_1_bits_set; // @[Slice.scala 468:27]
  wire [3:0] arbiter_2_io_in_1_bits_way; // @[Slice.scala 468:27]
  wire [22:0] arbiter_2_io_in_1_bits_tag; // @[Slice.scala 468:27]
  wire  arbiter_2_io_in_2_ready; // @[Slice.scala 468:27]
  wire  arbiter_2_io_in_2_valid; // @[Slice.scala 468:27]
  wire [6:0] arbiter_2_io_in_2_bits_set; // @[Slice.scala 468:27]
  wire [3:0] arbiter_2_io_in_2_bits_way; // @[Slice.scala 468:27]
  wire [22:0] arbiter_2_io_in_2_bits_tag; // @[Slice.scala 468:27]
  wire  arbiter_2_io_in_3_ready; // @[Slice.scala 468:27]
  wire  arbiter_2_io_in_3_valid; // @[Slice.scala 468:27]
  wire [6:0] arbiter_2_io_in_3_bits_set; // @[Slice.scala 468:27]
  wire [3:0] arbiter_2_io_in_3_bits_way; // @[Slice.scala 468:27]
  wire [22:0] arbiter_2_io_in_3_bits_tag; // @[Slice.scala 468:27]
  wire  arbiter_2_io_in_4_ready; // @[Slice.scala 468:27]
  wire  arbiter_2_io_in_4_valid; // @[Slice.scala 468:27]
  wire [6:0] arbiter_2_io_in_4_bits_set; // @[Slice.scala 468:27]
  wire [3:0] arbiter_2_io_in_4_bits_way; // @[Slice.scala 468:27]
  wire [22:0] arbiter_2_io_in_4_bits_tag; // @[Slice.scala 468:27]
  wire  arbiter_2_io_in_5_ready; // @[Slice.scala 468:27]
  wire  arbiter_2_io_in_5_valid; // @[Slice.scala 468:27]
  wire [6:0] arbiter_2_io_in_5_bits_set; // @[Slice.scala 468:27]
  wire [3:0] arbiter_2_io_in_5_bits_way; // @[Slice.scala 468:27]
  wire [22:0] arbiter_2_io_in_5_bits_tag; // @[Slice.scala 468:27]
  wire  arbiter_2_io_in_6_ready; // @[Slice.scala 468:27]
  wire  arbiter_2_io_in_6_valid; // @[Slice.scala 468:27]
  wire [6:0] arbiter_2_io_in_6_bits_set; // @[Slice.scala 468:27]
  wire [3:0] arbiter_2_io_in_6_bits_way; // @[Slice.scala 468:27]
  wire [22:0] arbiter_2_io_in_6_bits_tag; // @[Slice.scala 468:27]
  wire  arbiter_2_io_in_7_ready; // @[Slice.scala 468:27]
  wire  arbiter_2_io_in_7_valid; // @[Slice.scala 468:27]
  wire [6:0] arbiter_2_io_in_7_bits_set; // @[Slice.scala 468:27]
  wire [3:0] arbiter_2_io_in_7_bits_way; // @[Slice.scala 468:27]
  wire [22:0] arbiter_2_io_in_7_bits_tag; // @[Slice.scala 468:27]
  wire  arbiter_2_io_in_8_ready; // @[Slice.scala 468:27]
  wire  arbiter_2_io_in_8_valid; // @[Slice.scala 468:27]
  wire [6:0] arbiter_2_io_in_8_bits_set; // @[Slice.scala 468:27]
  wire [3:0] arbiter_2_io_in_8_bits_way; // @[Slice.scala 468:27]
  wire [22:0] arbiter_2_io_in_8_bits_tag; // @[Slice.scala 468:27]
  wire  arbiter_2_io_in_9_ready; // @[Slice.scala 468:27]
  wire  arbiter_2_io_in_9_valid; // @[Slice.scala 468:27]
  wire [6:0] arbiter_2_io_in_9_bits_set; // @[Slice.scala 468:27]
  wire [3:0] arbiter_2_io_in_9_bits_way; // @[Slice.scala 468:27]
  wire [22:0] arbiter_2_io_in_9_bits_tag; // @[Slice.scala 468:27]
  wire  arbiter_2_io_in_10_ready; // @[Slice.scala 468:27]
  wire  arbiter_2_io_in_10_valid; // @[Slice.scala 468:27]
  wire [6:0] arbiter_2_io_in_10_bits_set; // @[Slice.scala 468:27]
  wire [3:0] arbiter_2_io_in_10_bits_way; // @[Slice.scala 468:27]
  wire [22:0] arbiter_2_io_in_10_bits_tag; // @[Slice.scala 468:27]
  wire  arbiter_2_io_in_11_ready; // @[Slice.scala 468:27]
  wire  arbiter_2_io_in_11_valid; // @[Slice.scala 468:27]
  wire [6:0] arbiter_2_io_in_11_bits_set; // @[Slice.scala 468:27]
  wire [3:0] arbiter_2_io_in_11_bits_way; // @[Slice.scala 468:27]
  wire [22:0] arbiter_2_io_in_11_bits_tag; // @[Slice.scala 468:27]
  wire  arbiter_2_io_in_12_ready; // @[Slice.scala 468:27]
  wire  arbiter_2_io_in_12_valid; // @[Slice.scala 468:27]
  wire [6:0] arbiter_2_io_in_12_bits_set; // @[Slice.scala 468:27]
  wire [3:0] arbiter_2_io_in_12_bits_way; // @[Slice.scala 468:27]
  wire [22:0] arbiter_2_io_in_12_bits_tag; // @[Slice.scala 468:27]
  wire  arbiter_2_io_in_13_ready; // @[Slice.scala 468:27]
  wire  arbiter_2_io_in_13_valid; // @[Slice.scala 468:27]
  wire [6:0] arbiter_2_io_in_13_bits_set; // @[Slice.scala 468:27]
  wire [3:0] arbiter_2_io_in_13_bits_way; // @[Slice.scala 468:27]
  wire [22:0] arbiter_2_io_in_13_bits_tag; // @[Slice.scala 468:27]
  wire  arbiter_2_io_out_ready; // @[Slice.scala 468:27]
  wire  arbiter_2_io_out_valid; // @[Slice.scala 468:27]
  wire [6:0] arbiter_2_io_out_bits_set; // @[Slice.scala 468:27]
  wire [3:0] arbiter_2_io_out_bits_way; // @[Slice.scala 468:27]
  wire [22:0] arbiter_2_io_out_bits_tag; // @[Slice.scala 468:27]
  wire  opdata = sinkC_io_release_bits_opcode[0]; // @[Edges.scala 101:36]
  wire [12:0] _decode_T_5 = 13'h3f << sourceC_io_c_bits_size; // @[package.scala 234:77]
  wire [5:0] _decode_T_7 = ~_decode_T_5[5:0]; // @[package.scala 234:46]
  wire  decode_1 = _decode_T_7[5]; // @[Edges.scala 219:59]
  wire  opdata_1 = sourceC_io_c_bits_opcode[0]; // @[Edges.scala 101:36]
  wire  _T_1 = opdata_1 & decode_1; // @[Edges.scala 220:14]
  reg  beatsLeft; // @[Arbiter.scala 87:30]
  wire  idle = ~beatsLeft; // @[Arbiter.scala 88:28]
  wire  out_c_ready = io_out_c_q_io_enq_ready; // @[Decoupled.scala 365:17 Slice.scala 84:19]
  wire  latch = idle & out_c_ready; // @[Arbiter.scala 89:24]
  wire  out_earlyValid = sinkC_io_release_valid; // @[ReadyValidCancel.scala 68:19 69:20]
  wire  out_1_earlyValid = sourceC_io_c_valid; // @[ReadyValidCancel.scala 68:19 69:20]
  wire [1:0] _readys_T = {out_1_earlyValid,out_earlyValid}; // @[Cat.scala 31:58]
  wire [2:0] _readys_T_1 = {_readys_T, 1'h0}; // @[package.scala 244:48]
  wire [1:0] _readys_T_3 = _readys_T | _readys_T_1[1:0]; // @[package.scala 244:43]
  wire [2:0] _readys_T_5 = {_readys_T_3, 1'h0}; // @[Arbiter.scala 16:78]
  wire [1:0] _readys_T_7 = ~_readys_T_5[1:0]; // @[Arbiter.scala 16:61]
  wire  readys_0 = _readys_T_7[0]; // @[Arbiter.scala 95:86]
  wire  readys_1 = _readys_T_7[1]; // @[Arbiter.scala 95:86]
  wire  earlyWinner_0 = readys_0 & out_earlyValid; // @[Arbiter.scala 97:79]
  wire  earlyWinner_1 = readys_1 & out_1_earlyValid; // @[Arbiter.scala 97:79]
  wire  _T_12 = out_earlyValid | out_1_earlyValid; // @[Arbiter.scala 107:36]
  wire  maskedBeats_0 = earlyWinner_0 & opdata; // @[Arbiter.scala 111:73]
  wire  maskedBeats_1 = earlyWinner_1 & _T_1; // @[Arbiter.scala 111:73]
  wire  initBeats = maskedBeats_0 | maskedBeats_1; // @[Arbiter.scala 112:44]
  reg  state_0; // @[Arbiter.scala 116:26]
  wire  muxStateEarly_0 = idle ? earlyWinner_0 : state_0; // @[Arbiter.scala 117:30]
  reg  state_1; // @[Arbiter.scala 116:26]
  wire  muxStateEarly_1 = idle ? earlyWinner_1 : state_1; // @[Arbiter.scala 117:30]
  wire  _sink_ACancel_earlyValid_T_3 = state_0 & out_earlyValid | state_1 & out_1_earlyValid; // @[Mux.scala 27:73]
  wire  sink_ACancel_earlyValid = idle ? _T_12 : _sink_ACancel_earlyValid_T_3; // @[Arbiter.scala 125:29]
  wire  _beatsLeft_T_2 = out_c_ready & sink_ACancel_earlyValid; // @[ReadyValidCancel.scala 49:33]
  wire  allowed_0 = idle ? readys_0 : state_0; // @[Arbiter.scala 121:24]
  wire  allowed_1 = idle ? readys_1 : state_1; // @[Arbiter.scala 121:24]
  wire [255:0] out_bits_data = sinkC_io_release_bits_data; // @[ReadyValidCancel.scala 68:19 71:14]
  wire [255:0] _T_29 = muxStateEarly_0 ? out_bits_data : 256'h0; // @[Mux.scala 27:73]
  wire [255:0] out_1_bits_data = sourceC_io_c_bits_data; // @[ReadyValidCancel.scala 68:19 71:14]
  wire [255:0] _T_30 = muxStateEarly_1 ? out_1_bits_data : 256'h0; // @[Mux.scala 27:73]
  wire [35:0] out_bits_address = sinkC_io_release_bits_address; // @[ReadyValidCancel.scala 68:19 71:14]
  wire [35:0] _T_32 = muxStateEarly_0 ? out_bits_address : 36'h0; // @[Mux.scala 27:73]
  wire [35:0] out_1_bits_address = sourceC_io_c_bits_address; // @[ReadyValidCancel.scala 68:19 71:14]
  wire [35:0] _T_33 = muxStateEarly_1 ? out_1_bits_address : 36'h0; // @[Mux.scala 27:73]
  wire [3:0] out_bits_source = sinkC_io_release_bits_source; // @[ReadyValidCancel.scala 68:19 71:14]
  wire [3:0] _T_35 = muxStateEarly_0 ? out_bits_source : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] out_1_bits_source = sourceC_io_c_bits_source; // @[ReadyValidCancel.scala 68:19 71:14]
  wire [3:0] _T_36 = muxStateEarly_1 ? out_1_bits_source : 4'h0; // @[Mux.scala 27:73]
  wire [2:0] _T_38 = muxStateEarly_0 ? 3'h6 : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] out_1_bits_size = sourceC_io_c_bits_size; // @[ReadyValidCancel.scala 68:19 71:14]
  wire [2:0] _T_39 = muxStateEarly_1 ? out_1_bits_size : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] out_bits_opcode = sinkC_io_release_bits_opcode; // @[ReadyValidCancel.scala 68:19 71:14]
  wire [2:0] _T_44 = muxStateEarly_0 ? out_bits_opcode : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] out_1_bits_opcode = sourceC_io_c_bits_opcode; // @[ReadyValidCancel.scala 68:19 71:14]
  wire [2:0] _T_45 = muxStateEarly_1 ? out_1_bits_opcode : 3'h0; // @[Mux.scala 27:73]
  wire  _a_req_valid_T = ~probeHelperOpt_io_full; // @[Slice.scala 389:19]
  wire  a_req_ready = a_req_buffer_io_in_ready; // @[Slice.scala 129:19 148:24]
  reg  bc_mask_latch_0; // @[Slice.scala 186:30]
  reg  bc_mask_latch_1; // @[Slice.scala 186:30]
  reg  bc_mask_latch_2; // @[Slice.scala 186:30]
  reg  bc_mask_latch_3; // @[Slice.scala 186:30]
  reg  bc_mask_latch_4; // @[Slice.scala 186:30]
  reg  bc_mask_latch_5; // @[Slice.scala 186:30]
  reg  bc_mask_latch_6; // @[Slice.scala 186:30]
  reg  bc_mask_latch_7; // @[Slice.scala 186:30]
  reg  bc_mask_latch_8; // @[Slice.scala 186:30]
  reg  bc_mask_latch_9; // @[Slice.scala 186:30]
  reg  bc_mask_latch_10; // @[Slice.scala 186:30]
  reg  bc_mask_latch_11; // @[Slice.scala 186:30]
  reg  bc_mask_latch_12; // @[Slice.scala 186:30]
  reg  bc_mask_latch_13; // @[Slice.scala 186:30]
  reg  c_mask_latch_0; // @[Slice.scala 187:29]
  reg  c_mask_latch_1; // @[Slice.scala 187:29]
  reg  c_mask_latch_2; // @[Slice.scala 187:29]
  reg  c_mask_latch_3; // @[Slice.scala 187:29]
  reg  c_mask_latch_4; // @[Slice.scala 187:29]
  reg  c_mask_latch_5; // @[Slice.scala 187:29]
  reg  c_mask_latch_6; // @[Slice.scala 187:29]
  reg  c_mask_latch_7; // @[Slice.scala 187:29]
  reg  c_mask_latch_8; // @[Slice.scala 187:29]
  reg  c_mask_latch_9; // @[Slice.scala 187:29]
  reg  c_mask_latch_10; // @[Slice.scala 187:29]
  reg  c_mask_latch_11; // @[Slice.scala 187:29]
  reg  c_mask_latch_12; // @[Slice.scala 187:29]
  reg  c_mask_latch_13; // @[Slice.scala 187:29]
  reg  c_mask_latch_14; // @[Slice.scala 187:29]
  wire  bc_disable = bc_mask_latch_0 & bc_mshr_io_status_valid; // @[Slice.scala 196:41]
  wire  c_disable = c_mask_latch_0 & c_mshr_io_status_valid; // @[Slice.scala 197:39]
  wire  bc_disable_1 = bc_mask_latch_1 & bc_mshr_io_status_valid; // @[Slice.scala 196:41]
  wire  c_disable_1 = c_mask_latch_1 & c_mshr_io_status_valid; // @[Slice.scala 197:39]
  wire  bc_disable_2 = bc_mask_latch_2 & bc_mshr_io_status_valid; // @[Slice.scala 196:41]
  wire  c_disable_2 = c_mask_latch_2 & c_mshr_io_status_valid; // @[Slice.scala 197:39]
  wire  bc_disable_3 = bc_mask_latch_3 & bc_mshr_io_status_valid; // @[Slice.scala 196:41]
  wire  c_disable_3 = c_mask_latch_3 & c_mshr_io_status_valid; // @[Slice.scala 197:39]
  wire  bc_disable_4 = bc_mask_latch_4 & bc_mshr_io_status_valid; // @[Slice.scala 196:41]
  wire  c_disable_4 = c_mask_latch_4 & c_mshr_io_status_valid; // @[Slice.scala 197:39]
  wire  bc_disable_5 = bc_mask_latch_5 & bc_mshr_io_status_valid; // @[Slice.scala 196:41]
  wire  c_disable_5 = c_mask_latch_5 & c_mshr_io_status_valid; // @[Slice.scala 197:39]
  wire  bc_disable_6 = bc_mask_latch_6 & bc_mshr_io_status_valid; // @[Slice.scala 196:41]
  wire  c_disable_6 = c_mask_latch_6 & c_mshr_io_status_valid; // @[Slice.scala 197:39]
  wire  bc_disable_7 = bc_mask_latch_7 & bc_mshr_io_status_valid; // @[Slice.scala 196:41]
  wire  c_disable_7 = c_mask_latch_7 & c_mshr_io_status_valid; // @[Slice.scala 197:39]
  wire  bc_disable_8 = bc_mask_latch_8 & bc_mshr_io_status_valid; // @[Slice.scala 196:41]
  wire  c_disable_8 = c_mask_latch_8 & c_mshr_io_status_valid; // @[Slice.scala 197:39]
  wire  bc_disable_9 = bc_mask_latch_9 & bc_mshr_io_status_valid; // @[Slice.scala 196:41]
  wire  c_disable_9 = c_mask_latch_9 & c_mshr_io_status_valid; // @[Slice.scala 197:39]
  wire  bc_disable_10 = bc_mask_latch_10 & bc_mshr_io_status_valid; // @[Slice.scala 196:41]
  wire  c_disable_10 = c_mask_latch_10 & c_mshr_io_status_valid; // @[Slice.scala 197:39]
  wire  bc_disable_11 = bc_mask_latch_11 & bc_mshr_io_status_valid; // @[Slice.scala 196:41]
  wire  c_disable_11 = c_mask_latch_11 & c_mshr_io_status_valid; // @[Slice.scala 197:39]
  wire  bc_disable_12 = bc_mask_latch_12 & bc_mshr_io_status_valid; // @[Slice.scala 196:41]
  wire  c_disable_12 = c_mask_latch_12 & c_mshr_io_status_valid; // @[Slice.scala 197:39]
  wire  bc_disable_13 = bc_mask_latch_13 & bc_mshr_io_status_valid; // @[Slice.scala 196:41]
  wire  c_disable_13 = c_mask_latch_13 & c_mshr_io_status_valid; // @[Slice.scala 197:39]
  wire  _nestedWb_btoN_T = ~c_mshr_io_status_valid; // @[Slice.scala 279:34]
  wire  _nestedWb_btoN_T_2 = bc_mshr_io_status_valid & ~c_mshr_io_status_valid & bc_mshr_io_tasks_dir_write_valid; // @[Slice.scala 279:44]
  wire  _nestedWb_btoN_T_3 = bc_mshr_io_tasks_dir_write_bits_data_state == 2'h0; // @[Slice.scala 281:17]
  wire  _nestedWb_btoB_T_3 = bc_mshr_io_tasks_dir_write_bits_data_state == 2'h1; // @[Slice.scala 284:17]
  wire  _nestedWb_bclr_dirty_T_4 = ~bc_mshr_io_tasks_dir_write_bits_data_state[1]; // @[Slice.scala 287:5]
  wire  _nestedWb_c_set_dirty_T = c_mshr_io_status_valid & c_mshr_io_tasks_dir_write_valid; // @[Slice.scala 291:36]
  wire  _nestedWb_c_set_hit_T_1 = c_mshr_io_tasks_tag_write_bits_tag == abc_mshr_0_io_status_bits_tag; // @[Slice.scala 305:43]
  wire  _nestedWb_c_set_hit_T_3 = c_mshr_io_tasks_tag_write_bits_tag == abc_mshr_1_io_status_bits_tag; // @[Slice.scala 305:43]
  wire  _nestedWb_c_set_hit_T_5 = c_mshr_io_tasks_tag_write_bits_tag == abc_mshr_2_io_status_bits_tag; // @[Slice.scala 305:43]
  wire  _nestedWb_c_set_hit_T_7 = c_mshr_io_tasks_tag_write_bits_tag == abc_mshr_3_io_status_bits_tag; // @[Slice.scala 305:43]
  wire  _nestedWb_c_set_hit_T_9 = c_mshr_io_tasks_tag_write_bits_tag == abc_mshr_4_io_status_bits_tag; // @[Slice.scala 305:43]
  wire  _nestedWb_c_set_hit_T_11 = c_mshr_io_tasks_tag_write_bits_tag == abc_mshr_5_io_status_bits_tag; // @[Slice.scala 305:43]
  wire  _nestedWb_c_set_hit_T_13 = c_mshr_io_tasks_tag_write_bits_tag == abc_mshr_6_io_status_bits_tag; // @[Slice.scala 305:43]
  wire  _nestedWb_c_set_hit_T_15 = c_mshr_io_tasks_tag_write_bits_tag == abc_mshr_7_io_status_bits_tag; // @[Slice.scala 305:43]
  wire  _nestedWb_c_set_hit_T_17 = c_mshr_io_tasks_tag_write_bits_tag == abc_mshr_8_io_status_bits_tag; // @[Slice.scala 305:43]
  wire  _nestedWb_c_set_hit_T_19 = c_mshr_io_tasks_tag_write_bits_tag == abc_mshr_9_io_status_bits_tag; // @[Slice.scala 305:43]
  wire  _nestedWb_c_set_hit_T_21 = c_mshr_io_tasks_tag_write_bits_tag == abc_mshr_10_io_status_bits_tag; // @[Slice.scala 305:43]
  wire  _nestedWb_c_set_hit_T_23 = c_mshr_io_tasks_tag_write_bits_tag == abc_mshr_11_io_status_bits_tag; // @[Slice.scala 305:43]
  wire  _nestedWb_c_set_hit_T_25 = c_mshr_io_tasks_tag_write_bits_tag == abc_mshr_12_io_status_bits_tag; // @[Slice.scala 305:43]
  wire  _nestedWb_c_set_hit_T_27 = c_mshr_io_tasks_tag_write_bits_tag == abc_mshr_13_io_status_bits_tag; // @[Slice.scala 305:43]
  wire  _nestedWb_c_set_hit_T_29 = c_mshr_io_tasks_tag_write_bits_tag == bc_mshr_io_status_bits_tag; // @[Slice.scala 305:43]
  wire  _nestedWb_clients_0_isToN_T = c_mshr_io_tasks_client_dir_write_bits_data_0_state == 2'h0; // @[Slice.scala 317:67]
  wire  _nestedWb_clients_0_isToN_T_1 = c_mshr_io_tasks_client_dir_write_valid & _nestedWb_clients_0_isToN_T; // @[Slice.scala 316:52]
  wire  _nestedWb_clients_0_isToN_T_2 = bc_mshr_io_tasks_client_dir_write_bits_data_0_state == 2'h0; // @[Slice.scala 319:68]
  wire  _nestedWb_clients_0_isToN_T_3 = bc_mshr_io_tasks_client_dir_write_valid & _nestedWb_clients_0_isToN_T_2; // @[Slice.scala 318:53]
  wire  nestedWb_clients_0_isToN = c_mshr_io_status_valid ? _nestedWb_clients_0_isToN_T_1 :
    _nestedWb_clients_0_isToN_T_3; // @[Slice.scala 314:25]
  wire  _nestedWb_clients_1_isToN_T = c_mshr_io_tasks_client_dir_write_bits_data_1_state == 2'h0; // @[Slice.scala 317:67]
  wire  _nestedWb_clients_1_isToN_T_1 = c_mshr_io_tasks_client_dir_write_valid & _nestedWb_clients_1_isToN_T; // @[Slice.scala 316:52]
  wire  _nestedWb_clients_1_isToN_T_2 = bc_mshr_io_tasks_client_dir_write_bits_data_1_state == 2'h0; // @[Slice.scala 319:68]
  wire  _nestedWb_clients_1_isToN_T_3 = bc_mshr_io_tasks_client_dir_write_valid & _nestedWb_clients_1_isToN_T_2; // @[Slice.scala 318:53]
  wire  nestedWb_clients_1_isToN = c_mshr_io_status_valid ? _nestedWb_clients_1_isToN_T_1 :
    _nestedWb_clients_1_isToN_T_3; // @[Slice.scala 314:25]
  wire [6:0] ms_14_io_probeAckDataThrough_lo = {abc_mshr_7_io_bstatus_probeAckDataThrough,
    abc_mshr_8_io_bstatus_probeAckDataThrough,abc_mshr_9_io_bstatus_probeAckDataThrough,
    abc_mshr_10_io_bstatus_probeAckDataThrough,abc_mshr_11_io_bstatus_probeAckDataThrough,
    abc_mshr_12_io_bstatus_probeAckDataThrough,abc_mshr_13_io_bstatus_probeAckDataThrough}; // @[Cat.scala 31:58]
  wire [13:0] _ms_14_io_probeAckDataThrough_T = {abc_mshr_0_io_bstatus_probeAckDataThrough,
    abc_mshr_1_io_bstatus_probeAckDataThrough,abc_mshr_2_io_bstatus_probeAckDataThrough,
    abc_mshr_3_io_bstatus_probeAckDataThrough,abc_mshr_4_io_bstatus_probeAckDataThrough,
    abc_mshr_5_io_bstatus_probeAckDataThrough,abc_mshr_6_io_bstatus_probeAckDataThrough,
    ms_14_io_probeAckDataThrough_lo}; // @[Cat.scala 31:58]
  wire [6:0] ms_15_io_releaseThrough_lo = {abc_mshr_8_io_c_status_releaseThrough,abc_mshr_9_io_c_status_releaseThrough,
    abc_mshr_10_io_c_status_releaseThrough,abc_mshr_11_io_c_status_releaseThrough,abc_mshr_12_io_c_status_releaseThrough
    ,abc_mshr_13_io_c_status_releaseThrough,bc_mshr_io_c_status_releaseThrough}; // @[Cat.scala 31:58]
  wire [14:0] _ms_15_io_releaseThrough_T = {abc_mshr_0_io_c_status_releaseThrough,abc_mshr_1_io_c_status_releaseThrough,
    abc_mshr_2_io_c_status_releaseThrough,abc_mshr_3_io_c_status_releaseThrough,abc_mshr_4_io_c_status_releaseThrough,
    abc_mshr_5_io_c_status_releaseThrough,abc_mshr_6_io_c_status_releaseThrough,abc_mshr_7_io_c_status_releaseThrough,
    ms_15_io_releaseThrough_lo}; // @[Cat.scala 31:58]
  reg [19:0] bc_bits_latch_tag; // @[Reg.scala 16:16]
  reg [9:0] bc_bits_latch_set; // @[Reg.scala 16:16]
  reg [5:0] bc_bits_latch_off; // @[Reg.scala 16:16]
  reg [2:0] bc_bits_latch_opcode; // @[Reg.scala 16:16]
  reg [2:0] bc_bits_latch_param; // @[Reg.scala 16:16]
  reg [3:0] bc_bits_latch_source; // @[Reg.scala 16:16]
  reg [2:0] bc_bits_latch_bufIdx; // @[Reg.scala 16:16]
  reg [2:0] bc_bits_latch_size; // @[Reg.scala 16:16]
  reg  bc_bits_latch_putData; // @[Reg.scala 16:16]
  reg  bc_valid_latch; // @[Slice.scala 484:37]
  reg [19:0] c_bits_latch_tag; // @[Reg.scala 16:16]
  reg [9:0] c_bits_latch_set; // @[Reg.scala 16:16]
  reg [5:0] c_bits_latch_off; // @[Reg.scala 16:16]
  reg [2:0] c_bits_latch_opcode; // @[Reg.scala 16:16]
  reg [2:0] c_bits_latch_param; // @[Reg.scala 16:16]
  reg [3:0] c_bits_latch_source; // @[Reg.scala 16:16]
  reg [2:0] c_bits_latch_bufIdx; // @[Reg.scala 16:16]
  reg [2:0] c_bits_latch_size; // @[Reg.scala 16:16]
  reg  c_bits_latch_putData; // @[Reg.scala 16:16]
  reg  c_valid_latch; // @[Slice.scala 486:36]
  wire  bc_real_valid = bc_mshr_io_tasks_source_a_valid & bc_valid_latch; // @[Slice.scala 487:38]
  wire  c_real_valid = c_mshr_io_tasks_source_a_valid & c_valid_latch; // @[Slice.scala 488:36]
  wire [19:0] _sourceA_io_task_bits_T_tag = bc_real_valid ? bc_bits_latch_tag : sourceA_task_arb_io_out_bits_tag; // @[Slice.scala 490:56]
  wire [9:0] _sourceA_io_task_bits_T_set = bc_real_valid ? bc_bits_latch_set : sourceA_task_arb_io_out_bits_set; // @[Slice.scala 490:56]
  wire [5:0] _sourceA_io_task_bits_T_off = bc_real_valid ? bc_bits_latch_off : sourceA_task_arb_io_out_bits_off; // @[Slice.scala 490:56]
  wire [2:0] _sourceA_io_task_bits_T_opcode = bc_real_valid ? bc_bits_latch_opcode : sourceA_task_arb_io_out_bits_opcode
    ; // @[Slice.scala 490:56]
  wire [2:0] _sourceA_io_task_bits_T_param = bc_real_valid ? bc_bits_latch_param : sourceA_task_arb_io_out_bits_param; // @[Slice.scala 490:56]
  wire [3:0] _sourceA_io_task_bits_T_source = bc_real_valid ? bc_bits_latch_source : sourceA_task_arb_io_out_bits_source
    ; // @[Slice.scala 490:56]
  wire [2:0] _sourceA_io_task_bits_T_bufIdx = bc_real_valid ? bc_bits_latch_bufIdx : sourceA_task_arb_io_out_bits_bufIdx
    ; // @[Slice.scala 490:56]
  wire [2:0] _sourceA_io_task_bits_T_size = bc_real_valid ? bc_bits_latch_size : sourceA_task_arb_io_out_bits_size; // @[Slice.scala 490:56]
  wire  _sourceA_io_task_bits_T_putData = bc_real_valid ? bc_bits_latch_putData : sourceA_task_arb_io_out_bits_putData; // @[Slice.scala 490:56]
  wire  _ms_14_io_tasks_source_a_ready_T_1 = ~c_real_valid; // @[Slice.scala 492:52]
  reg [9:0] bc_bits_latch_1_set; // @[Reg.scala 16:16]
  reg [19:0] bc_bits_latch_1_tag; // @[Reg.scala 16:16]
  reg [2:0] bc_bits_latch_1_param; // @[Reg.scala 16:16]
  reg [1:0] bc_bits_latch_1_clients; // @[Reg.scala 16:16]
  reg  bc_bits_latch_1_needData; // @[Reg.scala 16:16]
  reg  bc_valid_latch_1; // @[Slice.scala 484:37]
  reg [9:0] c_bits_latch_1_set; // @[Reg.scala 16:16]
  reg [19:0] c_bits_latch_1_tag; // @[Reg.scala 16:16]
  reg [2:0] c_bits_latch_1_param; // @[Reg.scala 16:16]
  reg [1:0] c_bits_latch_1_clients; // @[Reg.scala 16:16]
  reg  c_bits_latch_1_needData; // @[Reg.scala 16:16]
  reg  c_valid_latch_1; // @[Slice.scala 486:36]
  wire  bc_real_valid_1 = bc_mshr_io_tasks_source_bvalid & bc_valid_latch_1; // @[Slice.scala 487:38]
  wire  c_real_valid_1 = c_mshr_io_tasks_source_bvalid & c_valid_latch_1; // @[Slice.scala 488:36]
  wire [9:0] _sourceB_io_task_bits_T_set = bc_real_valid_1 ? bc_bits_latch_1_set : sourceB_task_arb_io_out_bits_set; // @[Slice.scala 490:56]
  wire [19:0] _sourceB_io_task_bits_T_tag = bc_real_valid_1 ? bc_bits_latch_1_tag : sourceB_task_arb_io_out_bits_tag; // @[Slice.scala 490:56]
  wire [2:0] _sourceB_io_task_bits_T_param = bc_real_valid_1 ? bc_bits_latch_1_param :
    sourceB_task_arb_io_out_bits_param; // @[Slice.scala 490:56]
  wire [1:0] _sourceB_io_task_bits_T_clients = bc_real_valid_1 ? bc_bits_latch_1_clients :
    sourceB_task_arb_io_out_bits_clients; // @[Slice.scala 490:56]
  wire  _sourceB_io_task_bits_T_needData = bc_real_valid_1 ? bc_bits_latch_1_needData :
    sourceB_task_arb_io_out_bits_needData; // @[Slice.scala 490:56]
  wire  _ms_14_io_tasks_source_bready_T_1 = ~c_real_valid_1; // @[Slice.scala 492:52]
  reg [2:0] bc_bits_latch_2_opcode; // @[Reg.scala 16:16]
  reg [19:0] bc_bits_latch_2_tag; // @[Reg.scala 16:16]
  reg [9:0] bc_bits_latch_2_set; // @[Reg.scala 16:16]
  reg [3:0] bc_bits_latch_2_source; // @[Reg.scala 16:16]
  reg [2:0] bc_bits_latch_2_way; // @[Reg.scala 16:16]
  reg  bc_valid_latch_2; // @[Slice.scala 484:37]
  reg [2:0] c_bits_latch_2_opcode; // @[Reg.scala 16:16]
  reg [19:0] c_bits_latch_2_tag; // @[Reg.scala 16:16]
  reg [9:0] c_bits_latch_2_set; // @[Reg.scala 16:16]
  reg [3:0] c_bits_latch_2_source; // @[Reg.scala 16:16]
  reg [2:0] c_bits_latch_2_way; // @[Reg.scala 16:16]
  reg  c_valid_latch_2; // @[Slice.scala 486:36]
  wire  bc_real_valid_2 = bc_mshr_io_tasks_source_c_valid & bc_valid_latch_2; // @[Slice.scala 487:38]
  wire  c_real_valid_2 = c_mshr_io_tasks_source_c_valid & c_valid_latch_2; // @[Slice.scala 488:36]
  wire [2:0] _sourceC_io_task_bits_T_opcode = bc_real_valid_2 ? bc_bits_latch_2_opcode :
    sourceC_task_arb_io_out_bits_opcode; // @[Slice.scala 490:56]
  wire [19:0] _sourceC_io_task_bits_T_tag = bc_real_valid_2 ? bc_bits_latch_2_tag : sourceC_task_arb_io_out_bits_tag; // @[Slice.scala 490:56]
  wire [9:0] _sourceC_io_task_bits_T_set = bc_real_valid_2 ? bc_bits_latch_2_set : sourceC_task_arb_io_out_bits_set; // @[Slice.scala 490:56]
  wire [3:0] _sourceC_io_task_bits_T_source = bc_real_valid_2 ? bc_bits_latch_2_source :
    sourceC_task_arb_io_out_bits_source; // @[Slice.scala 490:56]
  wire [2:0] _sourceC_io_task_bits_T_way = bc_real_valid_2 ? bc_bits_latch_2_way : sourceC_task_arb_io_out_bits_way; // @[Slice.scala 490:56]
  wire  _ms_14_io_tasks_source_c_ready_T_1 = ~c_real_valid_2; // @[Slice.scala 492:52]
  reg [5:0] bc_bits_latch_3_sourceId; // @[Reg.scala 16:16]
  reg [9:0] bc_bits_latch_3_set; // @[Reg.scala 16:16]
  reg [2:0] bc_bits_latch_3_channel; // @[Reg.scala 16:16]
  reg [2:0] bc_bits_latch_3_opcode; // @[Reg.scala 16:16]
  reg [2:0] bc_bits_latch_3_param; // @[Reg.scala 16:16]
  reg [2:0] bc_bits_latch_3_size; // @[Reg.scala 16:16]
  reg [2:0] bc_bits_latch_3_way; // @[Reg.scala 16:16]
  reg [5:0] bc_bits_latch_3_off; // @[Reg.scala 16:16]
  reg  bc_bits_latch_3_useBypass; // @[Reg.scala 16:16]
  reg [2:0] bc_bits_latch_3_bufIdx; // @[Reg.scala 16:16]
  reg  bc_bits_latch_3_denied; // @[Reg.scala 16:16]
  reg [3:0] bc_bits_latch_3_sinkId; // @[Reg.scala 16:16]
  reg  bc_bits_latch_3_bypassPut; // @[Reg.scala 16:16]
  reg  bc_bits_latch_3_dirty; // @[Reg.scala 16:16]
  reg  bc_valid_latch_3; // @[Slice.scala 484:37]
  reg [5:0] c_bits_latch_3_sourceId; // @[Reg.scala 16:16]
  reg [9:0] c_bits_latch_3_set; // @[Reg.scala 16:16]
  reg [2:0] c_bits_latch_3_channel; // @[Reg.scala 16:16]
  reg [2:0] c_bits_latch_3_opcode; // @[Reg.scala 16:16]
  reg [2:0] c_bits_latch_3_param; // @[Reg.scala 16:16]
  reg [2:0] c_bits_latch_3_size; // @[Reg.scala 16:16]
  reg [2:0] c_bits_latch_3_way; // @[Reg.scala 16:16]
  reg [5:0] c_bits_latch_3_off; // @[Reg.scala 16:16]
  reg  c_bits_latch_3_useBypass; // @[Reg.scala 16:16]
  reg [2:0] c_bits_latch_3_bufIdx; // @[Reg.scala 16:16]
  reg  c_bits_latch_3_denied; // @[Reg.scala 16:16]
  reg [3:0] c_bits_latch_3_sinkId; // @[Reg.scala 16:16]
  reg  c_bits_latch_3_bypassPut; // @[Reg.scala 16:16]
  reg  c_bits_latch_3_dirty; // @[Reg.scala 16:16]
  reg  c_valid_latch_3; // @[Slice.scala 486:36]
  wire  bc_real_valid_3 = bc_mshr_io_tasks_source_d_valid & bc_valid_latch_3; // @[Slice.scala 487:38]
  wire  c_real_valid_3 = c_mshr_io_tasks_source_d_valid & c_valid_latch_3; // @[Slice.scala 488:36]
  wire [5:0] _sourceD_io_task_bits_T_sourceId = bc_real_valid_3 ? bc_bits_latch_3_sourceId :
    sourceD_task_arb_io_out_bits_sourceId; // @[Slice.scala 490:56]
  wire [9:0] _sourceD_io_task_bits_T_set = bc_real_valid_3 ? bc_bits_latch_3_set : sourceD_task_arb_io_out_bits_set; // @[Slice.scala 490:56]
  wire [2:0] _sourceD_io_task_bits_T_channel = bc_real_valid_3 ? bc_bits_latch_3_channel :
    sourceD_task_arb_io_out_bits_channel; // @[Slice.scala 490:56]
  wire [2:0] _sourceD_io_task_bits_T_opcode = bc_real_valid_3 ? bc_bits_latch_3_opcode :
    sourceD_task_arb_io_out_bits_opcode; // @[Slice.scala 490:56]
  wire [2:0] _sourceD_io_task_bits_T_param = bc_real_valid_3 ? bc_bits_latch_3_param :
    sourceD_task_arb_io_out_bits_param; // @[Slice.scala 490:56]
  wire [2:0] _sourceD_io_task_bits_T_size = bc_real_valid_3 ? bc_bits_latch_3_size : sourceD_task_arb_io_out_bits_size; // @[Slice.scala 490:56]
  wire [2:0] _sourceD_io_task_bits_T_way = bc_real_valid_3 ? bc_bits_latch_3_way : sourceD_task_arb_io_out_bits_way; // @[Slice.scala 490:56]
  wire [5:0] _sourceD_io_task_bits_T_off = bc_real_valid_3 ? bc_bits_latch_3_off : sourceD_task_arb_io_out_bits_off; // @[Slice.scala 490:56]
  wire  _sourceD_io_task_bits_T_useBypass = bc_real_valid_3 ? bc_bits_latch_3_useBypass :
    sourceD_task_arb_io_out_bits_useBypass; // @[Slice.scala 490:56]
  wire [2:0] _sourceD_io_task_bits_T_bufIdx = bc_real_valid_3 ? bc_bits_latch_3_bufIdx :
    sourceD_task_arb_io_out_bits_bufIdx; // @[Slice.scala 490:56]
  wire  _sourceD_io_task_bits_T_denied = bc_real_valid_3 ? bc_bits_latch_3_denied : sourceD_task_arb_io_out_bits_denied; // @[Slice.scala 490:56]
  wire [3:0] _sourceD_io_task_bits_T_sinkId = bc_real_valid_3 ? bc_bits_latch_3_sinkId :
    sourceD_task_arb_io_out_bits_sinkId; // @[Slice.scala 490:56]
  wire  _sourceD_io_task_bits_T_bypassPut = bc_real_valid_3 ? bc_bits_latch_3_bypassPut :
    sourceD_task_arb_io_out_bits_bypassPut; // @[Slice.scala 490:56]
  wire  _sourceD_io_task_bits_T_dirty = bc_real_valid_3 ? bc_bits_latch_3_dirty : sourceD_task_arb_io_out_bits_dirty; // @[Slice.scala 490:56]
  wire  _ms_14_io_tasks_source_d_ready_T_1 = ~c_real_valid_3; // @[Slice.scala 492:52]
  reg [2:0] bc_bits_latch_4_sink; // @[Reg.scala 16:16]
  reg  bc_valid_latch_4; // @[Slice.scala 484:37]
  reg [2:0] c_bits_latch_4_sink; // @[Reg.scala 16:16]
  reg  c_valid_latch_4; // @[Slice.scala 486:36]
  wire  bc_real_valid_4 = bc_mshr_io_tasks_source_e_valid & bc_valid_latch_4; // @[Slice.scala 487:38]
  wire  c_real_valid_4 = c_mshr_io_tasks_source_e_valid & c_valid_latch_4; // @[Slice.scala 488:36]
  wire [2:0] _sourceE_io_task_bits_T_sink = bc_real_valid_4 ? bc_bits_latch_4_sink : sourceE_task_arb_io_out_bits_sink; // @[Slice.scala 490:56]
  wire  _ms_14_io_tasks_source_e_ready_T_1 = ~c_real_valid_4; // @[Slice.scala 492:52]
  reg [9:0] bc_bits_latch_6_set; // @[Reg.scala 16:16]
  reg [19:0] bc_bits_latch_6_tag; // @[Reg.scala 16:16]
  reg [2:0] bc_bits_latch_6_way; // @[Reg.scala 16:16]
  reg [2:0] bc_bits_latch_6_bufIdx; // @[Reg.scala 16:16]
  reg [2:0] bc_bits_latch_6_opcode; // @[Reg.scala 16:16]
  reg [3:0] bc_bits_latch_6_source; // @[Reg.scala 16:16]
  reg  bc_bits_latch_6_save; // @[Reg.scala 16:16]
  reg  bc_bits_latch_6_drop; // @[Reg.scala 16:16]
  reg  bc_bits_latch_6_release; // @[Reg.scala 16:16]
  reg  bc_valid_latch_6; // @[Slice.scala 484:37]
  reg [9:0] c_bits_latch_6_set; // @[Reg.scala 16:16]
  reg [19:0] c_bits_latch_6_tag; // @[Reg.scala 16:16]
  reg [2:0] c_bits_latch_6_way; // @[Reg.scala 16:16]
  reg [2:0] c_bits_latch_6_bufIdx; // @[Reg.scala 16:16]
  reg [2:0] c_bits_latch_6_opcode; // @[Reg.scala 16:16]
  reg [3:0] c_bits_latch_6_source; // @[Reg.scala 16:16]
  reg  c_bits_latch_6_save; // @[Reg.scala 16:16]
  reg  c_bits_latch_6_drop; // @[Reg.scala 16:16]
  reg  c_bits_latch_6_release; // @[Reg.scala 16:16]
  reg  c_valid_latch_6; // @[Slice.scala 486:36]
  wire  bc_real_valid_6 = bc_mshr_io_tasks_sink_c_valid & bc_valid_latch_6; // @[Slice.scala 487:38]
  wire  c_real_valid_6 = c_mshr_io_tasks_sink_c_valid & c_valid_latch_6; // @[Slice.scala 488:36]
  wire [9:0] _sinkC_io_task_bits_T_set = bc_real_valid_6 ? bc_bits_latch_6_set : sinkC_task_arb_io_out_bits_set; // @[Slice.scala 490:56]
  wire [19:0] _sinkC_io_task_bits_T_tag = bc_real_valid_6 ? bc_bits_latch_6_tag : sinkC_task_arb_io_out_bits_tag; // @[Slice.scala 490:56]
  wire [2:0] _sinkC_io_task_bits_T_way = bc_real_valid_6 ? bc_bits_latch_6_way : sinkC_task_arb_io_out_bits_way; // @[Slice.scala 490:56]
  wire [2:0] _sinkC_io_task_bits_T_bufIdx = bc_real_valid_6 ? bc_bits_latch_6_bufIdx : sinkC_task_arb_io_out_bits_bufIdx
    ; // @[Slice.scala 490:56]
  wire [2:0] _sinkC_io_task_bits_T_opcode = bc_real_valid_6 ? bc_bits_latch_6_opcode : sinkC_task_arb_io_out_bits_opcode
    ; // @[Slice.scala 490:56]
  wire [3:0] _sinkC_io_task_bits_T_source = bc_real_valid_6 ? bc_bits_latch_6_source : sinkC_task_arb_io_out_bits_source
    ; // @[Slice.scala 490:56]
  wire  _sinkC_io_task_bits_T_save = bc_real_valid_6 ? bc_bits_latch_6_save : sinkC_task_arb_io_out_bits_save; // @[Slice.scala 490:56]
  wire  _sinkC_io_task_bits_T_drop = bc_real_valid_6 ? bc_bits_latch_6_drop : sinkC_task_arb_io_out_bits_drop; // @[Slice.scala 490:56]
  wire  _sinkC_io_task_bits_T_release = bc_real_valid_6 ? bc_bits_latch_6_release : sinkC_task_arb_io_out_bits_release; // @[Slice.scala 490:56]
  wire  _ms_14_io_tasks_sink_c_ready_T_1 = ~c_real_valid_6; // @[Slice.scala 492:52]
  reg [9:0] bc_bits_latch_7_set; // @[Reg.scala 16:16]
  reg [2:0] bc_bits_latch_7_way; // @[Reg.scala 16:16]
  reg [19:0] bc_bits_latch_7_tag; // @[Reg.scala 16:16]
  reg  bc_valid_latch_7; // @[Slice.scala 484:37]
  reg [9:0] c_bits_latch_7_set; // @[Reg.scala 16:16]
  reg [2:0] c_bits_latch_7_way; // @[Reg.scala 16:16]
  reg [19:0] c_bits_latch_7_tag; // @[Reg.scala 16:16]
  reg  c_valid_latch_7; // @[Slice.scala 486:36]
  wire  bc_real_valid_7 = bc_mshr_io_tasks_tag_write_valid & bc_valid_latch_7; // @[Slice.scala 487:38]
  wire  c_real_valid_7 = c_mshr_io_tasks_tag_write_valid & c_valid_latch_7; // @[Slice.scala 488:36]
  wire [9:0] _pipeline_io_in_bits_T_set = bc_real_valid_7 ? bc_bits_latch_7_set : tagWrite_task_arb_io_out_bits_set; // @[Slice.scala 490:56]
  wire [2:0] _pipeline_io_in_bits_T_way = bc_real_valid_7 ? bc_bits_latch_7_way : tagWrite_task_arb_io_out_bits_way; // @[Slice.scala 490:56]
  wire [19:0] _pipeline_io_in_bits_T_tag = bc_real_valid_7 ? bc_bits_latch_7_tag : tagWrite_task_arb_io_out_bits_tag; // @[Slice.scala 490:56]
  wire  _ms_14_io_tasks_tag_write_ready_T_1 = ~c_real_valid_7; // @[Slice.scala 492:52]
  reg [6:0] bc_bits_latch_8_set; // @[Reg.scala 16:16]
  reg [3:0] bc_bits_latch_8_way; // @[Reg.scala 16:16]
  reg [22:0] bc_bits_latch_8_tag; // @[Reg.scala 16:16]
  reg  bc_valid_latch_8; // @[Slice.scala 484:37]
  reg [6:0] c_bits_latch_8_set; // @[Reg.scala 16:16]
  reg [3:0] c_bits_latch_8_way; // @[Reg.scala 16:16]
  reg [22:0] c_bits_latch_8_tag; // @[Reg.scala 16:16]
  reg  c_valid_latch_8; // @[Slice.scala 486:36]
  wire  bc_real_valid_8 = bc_mshr_io_tasks_client_tag_write_valid & bc_valid_latch_8; // @[Slice.scala 487:38]
  wire  c_real_valid_8 = c_mshr_io_tasks_client_tag_write_valid & c_valid_latch_8; // @[Slice.scala 488:36]
  wire [6:0] _pipeline_io_in_bits_T_2_set = bc_real_valid_8 ? bc_bits_latch_8_set : arbiter_2_io_out_bits_set; // @[Slice.scala 490:56]
  wire [3:0] _pipeline_io_in_bits_T_2_way = bc_real_valid_8 ? bc_bits_latch_8_way : arbiter_2_io_out_bits_way; // @[Slice.scala 490:56]
  wire [22:0] _pipeline_io_in_bits_T_2_tag = bc_real_valid_8 ? bc_bits_latch_8_tag : arbiter_2_io_out_bits_tag; // @[Slice.scala 490:56]
  wire  _ms_14_io_tasks_client_tag_write_ready_T_1 = ~c_real_valid_8; // @[Slice.scala 492:52]
  wire  is_ctrl_dir_res = directory_io_result_bits_idOH[1:0] == 2'h3; // @[Slice.scala 550:61]
  reg  ms_0_io_dirResult_valid_REG; // @[Slice.scala 556:41]
  reg  ms_1_io_dirResult_valid_REG; // @[Slice.scala 556:41]
  reg  ms_2_io_dirResult_valid_REG; // @[Slice.scala 556:41]
  reg  ms_3_io_dirResult_valid_REG; // @[Slice.scala 556:41]
  reg  ms_4_io_dirResult_valid_REG; // @[Slice.scala 556:41]
  reg  ms_5_io_dirResult_valid_REG; // @[Slice.scala 556:41]
  reg  ms_6_io_dirResult_valid_REG; // @[Slice.scala 556:41]
  reg  ms_7_io_dirResult_valid_REG; // @[Slice.scala 556:41]
  reg  ms_8_io_dirResult_valid_REG; // @[Slice.scala 556:41]
  reg  ms_9_io_dirResult_valid_REG; // @[Slice.scala 556:41]
  reg  ms_10_io_dirResult_valid_REG; // @[Slice.scala 556:41]
  reg  ms_11_io_dirResult_valid_REG; // @[Slice.scala 556:41]
  reg  ms_12_io_dirResult_valid_REG; // @[Slice.scala 556:41]
  reg  ms_13_io_dirResult_valid_REG; // @[Slice.scala 556:41]
  reg  ms_14_io_dirResult_valid_REG; // @[Slice.scala 556:41]
  reg  ms_15_io_dirResult_valid_REG; // @[Slice.scala 556:41]
  reg  probeHelperOpt_io_dirResult_valid_REG; // @[Slice.scala 560:36]
  wire  _sinkD_status_T = 4'h0 == sinkD_io_resp_bits_source; // @[Slice.scala 576:25]
  wire  _sinkD_status_T_1 = 4'h1 == sinkD_io_resp_bits_source; // @[Slice.scala 576:25]
  wire  _sinkD_status_T_2 = 4'h2 == sinkD_io_resp_bits_source; // @[Slice.scala 576:25]
  wire  _sinkD_status_T_3 = 4'h3 == sinkD_io_resp_bits_source; // @[Slice.scala 576:25]
  wire  _sinkD_status_T_4 = 4'h4 == sinkD_io_resp_bits_source; // @[Slice.scala 576:25]
  wire  _sinkD_status_T_5 = 4'h5 == sinkD_io_resp_bits_source; // @[Slice.scala 576:25]
  wire  _sinkD_status_T_6 = 4'h6 == sinkD_io_resp_bits_source; // @[Slice.scala 576:25]
  wire  _sinkD_status_T_7 = 4'h7 == sinkD_io_resp_bits_source; // @[Slice.scala 576:25]
  wire  _sinkD_status_T_8 = 4'h8 == sinkD_io_resp_bits_source; // @[Slice.scala 576:25]
  wire  _sinkD_status_T_9 = 4'h9 == sinkD_io_resp_bits_source; // @[Slice.scala 576:25]
  wire  _sinkD_status_T_10 = 4'ha == sinkD_io_resp_bits_source; // @[Slice.scala 576:25]
  wire  _sinkD_status_T_11 = 4'hb == sinkD_io_resp_bits_source; // @[Slice.scala 576:25]
  wire  _sinkD_status_T_12 = 4'hc == sinkD_io_resp_bits_source; // @[Slice.scala 576:25]
  wire  _sinkD_status_T_13 = 4'hd == sinkD_io_resp_bits_source; // @[Slice.scala 576:25]
  wire  _sinkD_status_T_14 = 4'he == sinkD_io_resp_bits_source; // @[Slice.scala 576:25]
  wire  _sinkD_status_T_15 = 4'hf == sinkD_io_resp_bits_source; // @[Slice.scala 576:25]
  wire  _sinkD_status_T_93 = _sinkD_status_T_15 & c_mshr_io_status_bits_will_save_data; // @[Mux.scala 27:73]
  wire  _sinkD_status_T_124 = _sinkD_status_T_15 & c_mshr_io_status_bits_will_grant_data; // @[Mux.scala 27:73]
  wire [2:0] _sinkD_status_T_295 = _sinkD_status_T ? abc_mshr_0_io_status_bits_way_reg : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _sinkD_status_T_296 = _sinkD_status_T_1 ? abc_mshr_1_io_status_bits_way_reg : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _sinkD_status_T_297 = _sinkD_status_T_2 ? abc_mshr_2_io_status_bits_way_reg : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _sinkD_status_T_298 = _sinkD_status_T_3 ? abc_mshr_3_io_status_bits_way_reg : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _sinkD_status_T_299 = _sinkD_status_T_4 ? abc_mshr_4_io_status_bits_way_reg : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _sinkD_status_T_300 = _sinkD_status_T_5 ? abc_mshr_5_io_status_bits_way_reg : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _sinkD_status_T_301 = _sinkD_status_T_6 ? abc_mshr_6_io_status_bits_way_reg : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _sinkD_status_T_302 = _sinkD_status_T_7 ? abc_mshr_7_io_status_bits_way_reg : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _sinkD_status_T_303 = _sinkD_status_T_8 ? abc_mshr_8_io_status_bits_way_reg : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _sinkD_status_T_304 = _sinkD_status_T_9 ? abc_mshr_9_io_status_bits_way_reg : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _sinkD_status_T_305 = _sinkD_status_T_10 ? abc_mshr_10_io_status_bits_way_reg : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _sinkD_status_T_306 = _sinkD_status_T_11 ? abc_mshr_11_io_status_bits_way_reg : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _sinkD_status_T_307 = _sinkD_status_T_12 ? abc_mshr_12_io_status_bits_way_reg : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _sinkD_status_T_308 = _sinkD_status_T_13 ? abc_mshr_13_io_status_bits_way_reg : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _sinkD_status_T_309 = _sinkD_status_T_14 ? bc_mshr_io_status_bits_way_reg : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _sinkD_status_T_310 = _sinkD_status_T_15 ? c_mshr_io_status_bits_way_reg : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _sinkD_status_T_311 = _sinkD_status_T_295 | _sinkD_status_T_296; // @[Mux.scala 27:73]
  wire [2:0] _sinkD_status_T_312 = _sinkD_status_T_311 | _sinkD_status_T_297; // @[Mux.scala 27:73]
  wire [2:0] _sinkD_status_T_313 = _sinkD_status_T_312 | _sinkD_status_T_298; // @[Mux.scala 27:73]
  wire [2:0] _sinkD_status_T_314 = _sinkD_status_T_313 | _sinkD_status_T_299; // @[Mux.scala 27:73]
  wire [2:0] _sinkD_status_T_315 = _sinkD_status_T_314 | _sinkD_status_T_300; // @[Mux.scala 27:73]
  wire [2:0] _sinkD_status_T_316 = _sinkD_status_T_315 | _sinkD_status_T_301; // @[Mux.scala 27:73]
  wire [2:0] _sinkD_status_T_317 = _sinkD_status_T_316 | _sinkD_status_T_302; // @[Mux.scala 27:73]
  wire [2:0] _sinkD_status_T_318 = _sinkD_status_T_317 | _sinkD_status_T_303; // @[Mux.scala 27:73]
  wire [2:0] _sinkD_status_T_319 = _sinkD_status_T_318 | _sinkD_status_T_304; // @[Mux.scala 27:73]
  wire [2:0] _sinkD_status_T_320 = _sinkD_status_T_319 | _sinkD_status_T_305; // @[Mux.scala 27:73]
  wire [2:0] _sinkD_status_T_321 = _sinkD_status_T_320 | _sinkD_status_T_306; // @[Mux.scala 27:73]
  wire [2:0] _sinkD_status_T_322 = _sinkD_status_T_321 | _sinkD_status_T_307; // @[Mux.scala 27:73]
  wire [2:0] _sinkD_status_T_323 = _sinkD_status_T_322 | _sinkD_status_T_308; // @[Mux.scala 27:73]
  wire [2:0] _sinkD_status_T_324 = _sinkD_status_T_323 | _sinkD_status_T_309; // @[Mux.scala 27:73]
  wire [9:0] _sinkD_status_T_388 = _sinkD_status_T ? abc_mshr_0_io_status_bits_set : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _sinkD_status_T_389 = _sinkD_status_T_1 ? abc_mshr_1_io_status_bits_set : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _sinkD_status_T_390 = _sinkD_status_T_2 ? abc_mshr_2_io_status_bits_set : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _sinkD_status_T_391 = _sinkD_status_T_3 ? abc_mshr_3_io_status_bits_set : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _sinkD_status_T_392 = _sinkD_status_T_4 ? abc_mshr_4_io_status_bits_set : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _sinkD_status_T_393 = _sinkD_status_T_5 ? abc_mshr_5_io_status_bits_set : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _sinkD_status_T_394 = _sinkD_status_T_6 ? abc_mshr_6_io_status_bits_set : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _sinkD_status_T_395 = _sinkD_status_T_7 ? abc_mshr_7_io_status_bits_set : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _sinkD_status_T_396 = _sinkD_status_T_8 ? abc_mshr_8_io_status_bits_set : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _sinkD_status_T_397 = _sinkD_status_T_9 ? abc_mshr_9_io_status_bits_set : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _sinkD_status_T_398 = _sinkD_status_T_10 ? abc_mshr_10_io_status_bits_set : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _sinkD_status_T_399 = _sinkD_status_T_11 ? abc_mshr_11_io_status_bits_set : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _sinkD_status_T_400 = _sinkD_status_T_12 ? abc_mshr_12_io_status_bits_set : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _sinkD_status_T_401 = _sinkD_status_T_13 ? abc_mshr_13_io_status_bits_set : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _sinkD_status_T_402 = _sinkD_status_T_14 ? bc_mshr_io_status_bits_set : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _sinkD_status_T_403 = _sinkD_status_T_15 ? c_mshr_io_status_bits_set : 10'h0; // @[Mux.scala 27:73]
  wire [9:0] _sinkD_status_T_404 = _sinkD_status_T_388 | _sinkD_status_T_389; // @[Mux.scala 27:73]
  wire [9:0] _sinkD_status_T_405 = _sinkD_status_T_404 | _sinkD_status_T_390; // @[Mux.scala 27:73]
  wire [9:0] _sinkD_status_T_406 = _sinkD_status_T_405 | _sinkD_status_T_391; // @[Mux.scala 27:73]
  wire [9:0] _sinkD_status_T_407 = _sinkD_status_T_406 | _sinkD_status_T_392; // @[Mux.scala 27:73]
  wire [9:0] _sinkD_status_T_408 = _sinkD_status_T_407 | _sinkD_status_T_393; // @[Mux.scala 27:73]
  wire [9:0] _sinkD_status_T_409 = _sinkD_status_T_408 | _sinkD_status_T_394; // @[Mux.scala 27:73]
  wire [9:0] _sinkD_status_T_410 = _sinkD_status_T_409 | _sinkD_status_T_395; // @[Mux.scala 27:73]
  wire [9:0] _sinkD_status_T_411 = _sinkD_status_T_410 | _sinkD_status_T_396; // @[Mux.scala 27:73]
  wire [9:0] _sinkD_status_T_412 = _sinkD_status_T_411 | _sinkD_status_T_397; // @[Mux.scala 27:73]
  wire [9:0] _sinkD_status_T_413 = _sinkD_status_T_412 | _sinkD_status_T_398; // @[Mux.scala 27:73]
  wire [9:0] _sinkD_status_T_414 = _sinkD_status_T_413 | _sinkD_status_T_399; // @[Mux.scala 27:73]
  wire [9:0] _sinkD_status_T_415 = _sinkD_status_T_414 | _sinkD_status_T_400; // @[Mux.scala 27:73]
  wire [9:0] _sinkD_status_T_416 = _sinkD_status_T_415 | _sinkD_status_T_401; // @[Mux.scala 27:73]
  wire [9:0] _sinkD_status_T_417 = _sinkD_status_T_416 | _sinkD_status_T_402; // @[Mux.scala 27:73]
  SinkA sinkA ( // @[Slice.scala 56:21]
    .clock(sinkA_clock),
    .reset(sinkA_reset),
    .io_a_ready(sinkA_io_a_ready),
    .io_a_valid(sinkA_io_a_valid),
    .io_a_bits_opcode(sinkA_io_a_bits_opcode),
    .io_a_bits_param(sinkA_io_a_bits_param),
    .io_a_bits_size(sinkA_io_a_bits_size),
    .io_a_bits_source(sinkA_io_a_bits_source),
    .io_a_bits_address(sinkA_io_a_bits_address),
    .io_a_bits_user_preferCache(sinkA_io_a_bits_user_preferCache),
    .io_a_bits_mask(sinkA_io_a_bits_mask),
    .io_a_bits_data(sinkA_io_a_bits_data),
    .io_alloc_ready(sinkA_io_alloc_ready),
    .io_alloc_valid(sinkA_io_alloc_valid),
    .io_alloc_bits_opcode(sinkA_io_alloc_bits_opcode),
    .io_alloc_bits_param(sinkA_io_alloc_bits_param),
    .io_alloc_bits_size(sinkA_io_alloc_bits_size),
    .io_alloc_bits_source(sinkA_io_alloc_bits_source),
    .io_alloc_bits_set(sinkA_io_alloc_bits_set),
    .io_alloc_bits_tag(sinkA_io_alloc_bits_tag),
    .io_alloc_bits_off(sinkA_io_alloc_bits_off),
    .io_alloc_bits_mask(sinkA_io_alloc_bits_mask),
    .io_alloc_bits_bufIdx(sinkA_io_alloc_bits_bufIdx),
    .io_alloc_bits_preferCache(sinkA_io_alloc_bits_preferCache),
    .io_d_pb_pop_ready(sinkA_io_d_pb_pop_ready),
    .io_d_pb_pop_valid(sinkA_io_d_pb_pop_valid),
    .io_d_pb_pop_bits_bufIdx(sinkA_io_d_pb_pop_bits_bufIdx),
    .io_d_pb_pop_bits_count(sinkA_io_d_pb_pop_bits_count),
    .io_d_pb_pop_bits_last(sinkA_io_d_pb_pop_bits_last),
    .io_d_pb_beat_data(sinkA_io_d_pb_beat_data),
    .io_d_pb_beat_mask(sinkA_io_d_pb_beat_mask),
    .io_a_pb_pop_ready(sinkA_io_a_pb_pop_ready),
    .io_a_pb_pop_valid(sinkA_io_a_pb_pop_valid),
    .io_a_pb_pop_bits_bufIdx(sinkA_io_a_pb_pop_bits_bufIdx),
    .io_a_pb_pop_bits_count(sinkA_io_a_pb_pop_bits_count),
    .io_a_pb_pop_bits_last(sinkA_io_a_pb_pop_bits_last),
    .io_a_pb_beat_data(sinkA_io_a_pb_beat_data),
    .io_a_pb_beat_mask(sinkA_io_a_pb_beat_mask)
  );
  SourceB sourceB ( // @[Slice.scala 57:23]
    .clock(sourceB_clock),
    .reset(sourceB_reset),
    .io_bready(sourceB_io_bready),
    .io_bvalid(sourceB_io_bvalid),
    .io_bparam(sourceB_io_bparam),
    .io_bsource(sourceB_io_bsource),
    .io_baddress(sourceB_io_baddress),
    .io_bdata(sourceB_io_bdata),
    .io_task_ready(sourceB_io_task_ready),
    .io_task_valid(sourceB_io_task_valid),
    .io_task_bits_set(sourceB_io_task_bits_set),
    .io_task_bits_tag(sourceB_io_task_bits_tag),
    .io_task_bits_param(sourceB_io_task_bits_param),
    .io_task_bits_clients(sourceB_io_task_bits_clients),
    .io_task_bits_needData(sourceB_io_task_bits_needData)
  );
  SinkC sinkC ( // @[Slice.scala 58:21]
    .clock(sinkC_clock),
    .reset(sinkC_reset),
    .io_c_ready(sinkC_io_c_ready),
    .io_c_valid(sinkC_io_c_valid),
    .io_c_bits_opcode(sinkC_io_c_bits_opcode),
    .io_c_bits_param(sinkC_io_c_bits_param),
    .io_c_bits_size(sinkC_io_c_bits_size),
    .io_c_bits_source(sinkC_io_c_bits_source),
    .io_c_bits_address(sinkC_io_c_bits_address),
    .io_c_bits_echo_blockisdirty(sinkC_io_c_bits_echo_blockisdirty),
    .io_c_bits_data(sinkC_io_c_bits_data),
    .io_alloc_ready(sinkC_io_alloc_ready),
    .io_alloc_valid(sinkC_io_alloc_valid),
    .io_alloc_bits_opcode(sinkC_io_alloc_bits_opcode),
    .io_alloc_bits_param(sinkC_io_alloc_bits_param),
    .io_alloc_bits_size(sinkC_io_alloc_bits_size),
    .io_alloc_bits_source(sinkC_io_alloc_bits_source),
    .io_alloc_bits_set(sinkC_io_alloc_bits_set),
    .io_alloc_bits_tag(sinkC_io_alloc_bits_tag),
    .io_alloc_bits_off(sinkC_io_alloc_bits_off),
    .io_alloc_bits_bufIdx(sinkC_io_alloc_bits_bufIdx),
    .io_alloc_bits_dirty(sinkC_io_alloc_bits_dirty),
    .io_resp_valid(sinkC_io_resp_valid),
    .io_resp_bits_hasData(sinkC_io_resp_bits_hasData),
    .io_resp_bits_param(sinkC_io_resp_bits_param),
    .io_resp_bits_source(sinkC_io_resp_bits_source),
    .io_resp_bits_last(sinkC_io_resp_bits_last),
    .io_resp_bits_set(sinkC_io_resp_bits_set),
    .io_resp_bits_bufIdx(sinkC_io_resp_bits_bufIdx),
    .io_task_ready(sinkC_io_task_ready),
    .io_task_valid(sinkC_io_task_valid),
    .io_task_bits_set(sinkC_io_task_bits_set),
    .io_task_bits_tag(sinkC_io_task_bits_tag),
    .io_task_bits_way(sinkC_io_task_bits_way),
    .io_task_bits_bufIdx(sinkC_io_task_bits_bufIdx),
    .io_task_bits_opcode(sinkC_io_task_bits_opcode),
    .io_task_bits_source(sinkC_io_task_bits_source),
    .io_task_bits_save(sinkC_io_task_bits_save),
    .io_task_bits_drop(sinkC_io_task_bits_drop),
    .io_task_bits_release(sinkC_io_task_bits_release),
    .io_bs_waddr_ready(sinkC_io_bs_waddr_ready),
    .io_bs_waddr_valid(sinkC_io_bs_waddr_valid),
    .io_bs_waddr_bits_way(sinkC_io_bs_waddr_bits_way),
    .io_bs_waddr_bits_set(sinkC_io_bs_waddr_bits_set),
    .io_bs_waddr_bits_beat(sinkC_io_bs_waddr_bits_beat),
    .io_bs_waddr_bits_noop(sinkC_io_bs_waddr_bits_noop),
    .io_bs_wdata_data(sinkC_io_bs_wdata_data),
    .io_sourceD_rhazard_valid(sinkC_io_sourceD_rhazard_valid),
    .io_sourceD_rhazard_bits_way(sinkC_io_sourceD_rhazard_bits_way),
    .io_sourceD_rhazard_bits_set(sinkC_io_sourceD_rhazard_bits_set),
    .io_release_ready(sinkC_io_release_ready),
    .io_release_valid(sinkC_io_release_valid),
    .io_release_bits_opcode(sinkC_io_release_bits_opcode),
    .io_release_bits_source(sinkC_io_release_bits_source),
    .io_release_bits_address(sinkC_io_release_bits_address),
    .io_release_bits_data(sinkC_io_release_bits_data)
  );
  SourceD sourceD ( // @[Slice.scala 59:23]
    .clock(sourceD_clock),
    .reset(sourceD_reset),
    .io_d_ready(sourceD_io_d_ready),
    .io_d_valid(sourceD_io_d_valid),
    .io_d_bits_opcode(sourceD_io_d_bits_opcode),
    .io_d_bits_param(sourceD_io_d_bits_param),
    .io_d_bits_size(sourceD_io_d_bits_size),
    .io_d_bits_source(sourceD_io_d_bits_source),
    .io_d_bits_sink(sourceD_io_d_bits_sink),
    .io_d_bits_denied(sourceD_io_d_bits_denied),
    .io_d_bits_echo_blockisdirty(sourceD_io_d_bits_echo_blockisdirty),
    .io_d_bits_data(sourceD_io_d_bits_data),
    .io_d_bits_corrupt(sourceD_io_d_bits_corrupt),
    .io_task_ready(sourceD_io_task_ready),
    .io_task_valid(sourceD_io_task_valid),
    .io_task_bits_sourceId(sourceD_io_task_bits_sourceId),
    .io_task_bits_set(sourceD_io_task_bits_set),
    .io_task_bits_channel(sourceD_io_task_bits_channel),
    .io_task_bits_opcode(sourceD_io_task_bits_opcode),
    .io_task_bits_param(sourceD_io_task_bits_param),
    .io_task_bits_size(sourceD_io_task_bits_size),
    .io_task_bits_way(sourceD_io_task_bits_way),
    .io_task_bits_off(sourceD_io_task_bits_off),
    .io_task_bits_useBypass(sourceD_io_task_bits_useBypass),
    .io_task_bits_bufIdx(sourceD_io_task_bits_bufIdx),
    .io_task_bits_denied(sourceD_io_task_bits_denied),
    .io_task_bits_sinkId(sourceD_io_task_bits_sinkId),
    .io_task_bits_bypassPut(sourceD_io_task_bits_bypassPut),
    .io_task_bits_dirty(sourceD_io_task_bits_dirty),
    .io_bs_raddr_ready(sourceD_io_bs_raddr_ready),
    .io_bs_raddr_valid(sourceD_io_bs_raddr_valid),
    .io_bs_raddr_bits_way(sourceD_io_bs_raddr_bits_way),
    .io_bs_raddr_bits_set(sourceD_io_bs_raddr_bits_set),
    .io_bs_raddr_bits_beat(sourceD_io_bs_raddr_bits_beat),
    .io_bs_rdata_data(sourceD_io_bs_rdata_data),
    .io_bypass_read_valid(sourceD_io_bypass_read_valid),
    .io_bypass_read_beat(sourceD_io_bypass_read_beat),
    .io_bypass_read_id(sourceD_io_bypass_read_id),
    .io_bypass_read_ready(sourceD_io_bypass_read_ready),
    .io_bypass_read_buffer_data_data(sourceD_io_bypass_read_buffer_data_data),
    .io_bypass_read_last(sourceD_io_bypass_read_last),
    .io_bs_waddr_ready(sourceD_io_bs_waddr_ready),
    .io_bs_waddr_valid(sourceD_io_bs_waddr_valid),
    .io_bs_waddr_bits_way(sourceD_io_bs_waddr_bits_way),
    .io_bs_waddr_bits_set(sourceD_io_bs_waddr_bits_set),
    .io_bs_waddr_bits_beat(sourceD_io_bs_waddr_bits_beat),
    .io_bs_wdata_data(sourceD_io_bs_wdata_data),
    .io_sourceD_rhazard_valid(sourceD_io_sourceD_rhazard_valid),
    .io_sourceD_rhazard_bits_way(sourceD_io_sourceD_rhazard_bits_way),
    .io_sourceD_rhazard_bits_set(sourceD_io_sourceD_rhazard_bits_set),
    .io_pb_pop_ready(sourceD_io_pb_pop_ready),
    .io_pb_pop_valid(sourceD_io_pb_pop_valid),
    .io_pb_pop_bits_bufIdx(sourceD_io_pb_pop_bits_bufIdx),
    .io_pb_pop_bits_count(sourceD_io_pb_pop_bits_count),
    .io_pb_pop_bits_last(sourceD_io_pb_pop_bits_last),
    .io_pb_beat_data(sourceD_io_pb_beat_data),
    .io_pb_beat_mask(sourceD_io_pb_beat_mask),
    .io_resp_valid(sourceD_io_resp_valid),
    .io_resp_bits_sink(sourceD_io_resp_bits_sink)
  );
  SinkE sinkE ( // @[Slice.scala 60:21]
    .io_e_ready(sinkE_io_e_ready),
    .io_e_valid(sinkE_io_e_valid),
    .io_e_bits_sink(sinkE_io_e_bits_sink),
    .io_resp_valid(sinkE_io_resp_valid),
    .io_resp_bits_sink(sinkE_io_resp_bits_sink)
  );
  SourceA sourceA ( // @[Slice.scala 70:23]
    .clock(sourceA_clock),
    .reset(sourceA_reset),
    .io_a_ready(sourceA_io_a_ready),
    .io_a_valid(sourceA_io_a_valid),
    .io_a_bits_opcode(sourceA_io_a_bits_opcode),
    .io_a_bits_param(sourceA_io_a_bits_param),
    .io_a_bits_size(sourceA_io_a_bits_size),
    .io_a_bits_source(sourceA_io_a_bits_source),
    .io_a_bits_address(sourceA_io_a_bits_address),
    .io_a_bits_mask(sourceA_io_a_bits_mask),
    .io_a_bits_data(sourceA_io_a_bits_data),
    .io_task_ready(sourceA_io_task_ready),
    .io_task_valid(sourceA_io_task_valid),
    .io_task_bits_tag(sourceA_io_task_bits_tag),
    .io_task_bits_set(sourceA_io_task_bits_set),
    .io_task_bits_off(sourceA_io_task_bits_off),
    .io_task_bits_opcode(sourceA_io_task_bits_opcode),
    .io_task_bits_param(sourceA_io_task_bits_param),
    .io_task_bits_source(sourceA_io_task_bits_source),
    .io_task_bits_bufIdx(sourceA_io_task_bits_bufIdx),
    .io_task_bits_size(sourceA_io_task_bits_size),
    .io_task_bits_putData(sourceA_io_task_bits_putData),
    .io_pb_pop_ready(sourceA_io_pb_pop_ready),
    .io_pb_pop_valid(sourceA_io_pb_pop_valid),
    .io_pb_pop_bits_bufIdx(sourceA_io_pb_pop_bits_bufIdx),
    .io_pb_pop_bits_count(sourceA_io_pb_pop_bits_count),
    .io_pb_pop_bits_last(sourceA_io_pb_pop_bits_last),
    .io_pb_beat_data(sourceA_io_pb_beat_data),
    .io_pb_beat_mask(sourceA_io_pb_beat_mask)
  );
  SinkB sinkB ( // @[Slice.scala 71:21]
    .io_bready(sinkB_io_bready),
    .io_bvalid(sinkB_io_bvalid),
    .io_bopcode(sinkB_io_bopcode),
    .io_bparam(sinkB_io_bparam),
    .io_bsize(sinkB_io_bsize),
    .io_bsource(sinkB_io_bsource),
    .io_baddress(sinkB_io_baddress),
    .io_bmask(sinkB_io_bmask),
    .io_bdata(sinkB_io_bdata),
    .io_alloc_ready(sinkB_io_alloc_ready),
    .io_alloc_valid(sinkB_io_alloc_valid),
    .io_alloc_bits_opcode(sinkB_io_alloc_bits_opcode),
    .io_alloc_bits_param(sinkB_io_alloc_bits_param),
    .io_alloc_bits_size(sinkB_io_alloc_bits_size),
    .io_alloc_bits_source(sinkB_io_alloc_bits_source),
    .io_alloc_bits_set(sinkB_io_alloc_bits_set),
    .io_alloc_bits_tag(sinkB_io_alloc_bits_tag),
    .io_alloc_bits_off(sinkB_io_alloc_bits_off),
    .io_alloc_bits_mask(sinkB_io_alloc_bits_mask),
    .io_alloc_bits_needProbeAckData(sinkB_io_alloc_bits_needProbeAckData)
  );
  SourceC sourceC ( // @[Slice.scala 72:23]
    .clock(sourceC_clock),
    .reset(sourceC_reset),
    .io_c_ready(sourceC_io_c_ready),
    .io_c_valid(sourceC_io_c_valid),
    .io_c_bits_opcode(sourceC_io_c_bits_opcode),
    .io_c_bits_size(sourceC_io_c_bits_size),
    .io_c_bits_source(sourceC_io_c_bits_source),
    .io_c_bits_address(sourceC_io_c_bits_address),
    .io_c_bits_data(sourceC_io_c_bits_data),
    .io_bs_raddr_ready(sourceC_io_bs_raddr_ready),
    .io_bs_raddr_valid(sourceC_io_bs_raddr_valid),
    .io_bs_raddr_bits_way(sourceC_io_bs_raddr_bits_way),
    .io_bs_raddr_bits_set(sourceC_io_bs_raddr_bits_set),
    .io_bs_raddr_bits_beat(sourceC_io_bs_raddr_bits_beat),
    .io_bs_rdata_data(sourceC_io_bs_rdata_data),
    .io_task_ready(sourceC_io_task_ready),
    .io_task_valid(sourceC_io_task_valid),
    .io_task_bits_opcode(sourceC_io_task_bits_opcode),
    .io_task_bits_tag(sourceC_io_task_bits_tag),
    .io_task_bits_set(sourceC_io_task_bits_set),
    .io_task_bits_source(sourceC_io_task_bits_source),
    .io_task_bits_way(sourceC_io_task_bits_way)
  );
  SinkD sinkD ( // @[Slice.scala 73:21]
    .clock(sinkD_clock),
    .reset(sinkD_reset),
    .io_d_ready(sinkD_io_d_ready),
    .io_d_valid(sinkD_io_d_valid),
    .io_d_bits_opcode(sinkD_io_d_bits_opcode),
    .io_d_bits_param(sinkD_io_d_bits_param),
    .io_d_bits_size(sinkD_io_d_bits_size),
    .io_d_bits_source(sinkD_io_d_bits_source),
    .io_d_bits_sink(sinkD_io_d_bits_sink),
    .io_d_bits_denied(sinkD_io_d_bits_denied),
    .io_d_bits_data(sinkD_io_d_bits_data),
    .io_bs_waddr_ready(sinkD_io_bs_waddr_ready),
    .io_bs_waddr_valid(sinkD_io_bs_waddr_valid),
    .io_bs_waddr_bits_way(sinkD_io_bs_waddr_bits_way),
    .io_bs_waddr_bits_set(sinkD_io_bs_waddr_bits_set),
    .io_bs_waddr_bits_beat(sinkD_io_bs_waddr_bits_beat),
    .io_bs_waddr_bits_noop(sinkD_io_bs_waddr_bits_noop),
    .io_bs_wdata_data(sinkD_io_bs_wdata_data),
    .io_bypass_write_valid(sinkD_io_bypass_write_valid),
    .io_bypass_write_beat(sinkD_io_bypass_write_beat),
    .io_bypass_write_data_data(sinkD_io_bypass_write_data_data),
    .io_bypass_write_ready(sinkD_io_bypass_write_ready),
    .io_bypass_write_id(sinkD_io_bypass_write_id),
    .io_way(sinkD_io_way),
    .io_set(sinkD_io_set),
    .io_inner_grant(sinkD_io_inner_grant),
    .io_save_data_in_bs(sinkD_io_save_data_in_bs),
    .io_resp_valid(sinkD_io_resp_valid),
    .io_resp_bits_opcode(sinkD_io_resp_bits_opcode),
    .io_resp_bits_param(sinkD_io_resp_bits_param),
    .io_resp_bits_source(sinkD_io_resp_bits_source),
    .io_resp_bits_sink(sinkD_io_resp_bits_sink),
    .io_resp_bits_last(sinkD_io_resp_bits_last),
    .io_resp_bits_denied(sinkD_io_resp_bits_denied),
    .io_resp_bits_bufIdx(sinkD_io_resp_bits_bufIdx),
    .io_sourceD_rhazard_valid(sinkD_io_sourceD_rhazard_valid),
    .io_sourceD_rhazard_bits_way(sinkD_io_sourceD_rhazard_bits_way),
    .io_sourceD_rhazard_bits_set(sinkD_io_sourceD_rhazard_bits_set)
  );
  SourceE sourceE ( // @[Slice.scala 74:23]
    .io_e_ready(sourceE_io_e_ready),
    .io_e_valid(sourceE_io_e_valid),
    .io_e_bits_sink(sourceE_io_e_bits_sink),
    .io_task_ready(sourceE_io_task_ready),
    .io_task_valid(sourceE_io_task_valid),
    .io_task_bits_sink(sourceE_io_task_bits_sink)
  );
  RefillBuffer refillBuffer ( // @[Slice.scala 76:28]
    .clock(refillBuffer_clock),
    .reset(refillBuffer_reset),
    .io_rvalid(refillBuffer_io_rvalid),
    .io_rbeat(refillBuffer_io_rbeat),
    .io_rid(refillBuffer_io_rid),
    .io_rready(refillBuffer_io_rready),
    .io_rbuffer_data_data(refillBuffer_io_rbuffer_data_data),
    .io_rlast(refillBuffer_io_rlast),
    .io_wvalid(refillBuffer_io_wvalid),
    .io_wbeat(refillBuffer_io_wbeat),
    .io_wdata_data(refillBuffer_io_wdata_data),
    .io_wready(refillBuffer_io_wready),
    .io_wid(refillBuffer_io_wid)
  );
  Queue_193 io_out_a_q ( // @[Decoupled.scala 361:21]
    .clock(io_out_a_q_clock),
    .reset(io_out_a_q_reset),
    .io_enq_ready(io_out_a_q_io_enq_ready),
    .io_enq_valid(io_out_a_q_io_enq_valid),
    .io_enq_bits_opcode(io_out_a_q_io_enq_bits_opcode),
    .io_enq_bits_param(io_out_a_q_io_enq_bits_param),
    .io_enq_bits_size(io_out_a_q_io_enq_bits_size),
    .io_enq_bits_source(io_out_a_q_io_enq_bits_source),
    .io_enq_bits_address(io_out_a_q_io_enq_bits_address),
    .io_enq_bits_mask(io_out_a_q_io_enq_bits_mask),
    .io_enq_bits_data(io_out_a_q_io_enq_bits_data),
    .io_deq_ready(io_out_a_q_io_deq_ready),
    .io_deq_valid(io_out_a_q_io_deq_valid),
    .io_deq_bits_opcode(io_out_a_q_io_deq_bits_opcode),
    .io_deq_bits_param(io_out_a_q_io_deq_bits_param),
    .io_deq_bits_size(io_out_a_q_io_deq_bits_size),
    .io_deq_bits_source(io_out_a_q_io_deq_bits_source),
    .io_deq_bits_address(io_out_a_q_io_deq_bits_address),
    .io_deq_bits_mask(io_out_a_q_io_deq_bits_mask),
    .io_deq_bits_data(io_out_a_q_io_deq_bits_data)
  );
  Queue_159 sinkB_io_bq ( // @[Decoupled.scala 361:21]
    .clock(sinkB_io_bq_clock),
    .reset(sinkB_io_bq_reset),
    .io_enq_ready(sinkB_io_bq_io_enq_ready),
    .io_enq_valid(sinkB_io_bq_io_enq_valid),
    .io_enq_bits_opcode(sinkB_io_bq_io_enq_bits_opcode),
    .io_enq_bits_param(sinkB_io_bq_io_enq_bits_param),
    .io_enq_bits_size(sinkB_io_bq_io_enq_bits_size),
    .io_enq_bits_source(sinkB_io_bq_io_enq_bits_source),
    .io_enq_bits_address(sinkB_io_bq_io_enq_bits_address),
    .io_enq_bits_mask(sinkB_io_bq_io_enq_bits_mask),
    .io_enq_bits_data(sinkB_io_bq_io_enq_bits_data),
    .io_deq_ready(sinkB_io_bq_io_deq_ready),
    .io_deq_valid(sinkB_io_bq_io_deq_valid),
    .io_deq_bits_opcode(sinkB_io_bq_io_deq_bits_opcode),
    .io_deq_bits_param(sinkB_io_bq_io_deq_bits_param),
    .io_deq_bits_size(sinkB_io_bq_io_deq_bits_size),
    .io_deq_bits_source(sinkB_io_bq_io_deq_bits_source),
    .io_deq_bits_address(sinkB_io_bq_io_deq_bits_address),
    .io_deq_bits_mask(sinkB_io_bq_io_deq_bits_mask),
    .io_deq_bits_data(sinkB_io_bq_io_deq_bits_data)
  );
  Queue_195 io_out_c_q ( // @[Decoupled.scala 361:21]
    .clock(io_out_c_q_clock),
    .reset(io_out_c_q_reset),
    .io_enq_ready(io_out_c_q_io_enq_ready),
    .io_enq_valid(io_out_c_q_io_enq_valid),
    .io_enq_bits_opcode(io_out_c_q_io_enq_bits_opcode),
    .io_enq_bits_size(io_out_c_q_io_enq_bits_size),
    .io_enq_bits_source(io_out_c_q_io_enq_bits_source),
    .io_enq_bits_address(io_out_c_q_io_enq_bits_address),
    .io_enq_bits_data(io_out_c_q_io_enq_bits_data),
    .io_deq_ready(io_out_c_q_io_deq_ready),
    .io_deq_valid(io_out_c_q_io_deq_valid),
    .io_deq_bits_opcode(io_out_c_q_io_deq_bits_opcode),
    .io_deq_bits_size(io_out_c_q_io_deq_bits_size),
    .io_deq_bits_source(io_out_c_q_io_deq_bits_source),
    .io_deq_bits_address(io_out_c_q_io_deq_bits_address),
    .io_deq_bits_data(io_out_c_q_io_deq_bits_data)
  );
  Queue_4 sinkD_io_d_q ( // @[Decoupled.scala 361:21]
    .clock(sinkD_io_d_q_clock),
    .reset(sinkD_io_d_q_reset),
    .io_enq_ready(sinkD_io_d_q_io_enq_ready),
    .io_enq_valid(sinkD_io_d_q_io_enq_valid),
    .io_enq_bits_opcode(sinkD_io_d_q_io_enq_bits_opcode),
    .io_enq_bits_param(sinkD_io_d_q_io_enq_bits_param),
    .io_enq_bits_size(sinkD_io_d_q_io_enq_bits_size),
    .io_enq_bits_source(sinkD_io_d_q_io_enq_bits_source),
    .io_enq_bits_sink(sinkD_io_d_q_io_enq_bits_sink),
    .io_enq_bits_denied(sinkD_io_d_q_io_enq_bits_denied),
    .io_enq_bits_data(sinkD_io_d_q_io_enq_bits_data),
    .io_deq_ready(sinkD_io_d_q_io_deq_ready),
    .io_deq_valid(sinkD_io_d_q_io_deq_valid),
    .io_deq_bits_opcode(sinkD_io_d_q_io_deq_bits_opcode),
    .io_deq_bits_param(sinkD_io_d_q_io_deq_bits_param),
    .io_deq_bits_size(sinkD_io_d_q_io_deq_bits_size),
    .io_deq_bits_source(sinkD_io_d_q_io_deq_bits_source),
    .io_deq_bits_sink(sinkD_io_d_q_io_deq_bits_sink),
    .io_deq_bits_denied(sinkD_io_d_q_io_deq_bits_denied),
    .io_deq_bits_data(sinkD_io_d_q_io_deq_bits_data)
  );
  Queue_197 io_out_e_q ( // @[Decoupled.scala 361:21]
    .clock(io_out_e_q_clock),
    .reset(io_out_e_q_reset),
    .io_enq_ready(io_out_e_q_io_enq_ready),
    .io_enq_valid(io_out_e_q_io_enq_valid),
    .io_enq_bits_sink(io_out_e_q_io_enq_bits_sink),
    .io_deq_valid(io_out_e_q_io_deq_valid),
    .io_deq_bits_sink(io_out_e_q_io_deq_bits_sink)
  );
  MSHR abc_mshr_0 ( // @[Slice.scala 94:16]
    .clock(abc_mshr_0_clock),
    .reset(abc_mshr_0_reset),
    .io_id(abc_mshr_0_io_id),
    .io_enable(abc_mshr_0_io_enable),
    .io_alloc_valid(abc_mshr_0_io_alloc_valid),
    .io_alloc_bits_channel(abc_mshr_0_io_alloc_bits_channel),
    .io_alloc_bits_opcode(abc_mshr_0_io_alloc_bits_opcode),
    .io_alloc_bits_param(abc_mshr_0_io_alloc_bits_param),
    .io_alloc_bits_size(abc_mshr_0_io_alloc_bits_size),
    .io_alloc_bits_source(abc_mshr_0_io_alloc_bits_source),
    .io_alloc_bits_set(abc_mshr_0_io_alloc_bits_set),
    .io_alloc_bits_tag(abc_mshr_0_io_alloc_bits_tag),
    .io_alloc_bits_off(abc_mshr_0_io_alloc_bits_off),
    .io_alloc_bits_mask(abc_mshr_0_io_alloc_bits_mask),
    .io_alloc_bits_bufIdx(abc_mshr_0_io_alloc_bits_bufIdx),
    .io_alloc_bits_preferCache(abc_mshr_0_io_alloc_bits_preferCache),
    .io_alloc_bits_dirty(abc_mshr_0_io_alloc_bits_dirty),
    .io_alloc_bits_fromProbeHelper(abc_mshr_0_io_alloc_bits_fromProbeHelper),
    .io_alloc_bits_fromCmoHelper(abc_mshr_0_io_alloc_bits_fromCmoHelper),
    .io_alloc_bits_needProbeAckData(abc_mshr_0_io_alloc_bits_needProbeAckData),
    .io_status_valid(abc_mshr_0_io_status_valid),
    .io_status_bits_set(abc_mshr_0_io_status_bits_set),
    .io_status_bits_tag(abc_mshr_0_io_status_bits_tag),
    .io_status_bits_way(abc_mshr_0_io_status_bits_way),
    .io_status_bits_way_reg(abc_mshr_0_io_status_bits_way_reg),
    .io_status_bits_nestB(abc_mshr_0_io_status_bits_nestB),
    .io_status_bits_nestC(abc_mshr_0_io_status_bits_nestC),
    .io_status_bits_will_grant_data(abc_mshr_0_io_status_bits_will_grant_data),
    .io_status_bits_will_save_data(abc_mshr_0_io_status_bits_will_save_data),
    .io_status_bits_will_free(abc_mshr_0_io_status_bits_will_free),
    .io_resps_sink_c_valid(abc_mshr_0_io_resps_sink_c_valid),
    .io_resps_sink_c_bits_hasData(abc_mshr_0_io_resps_sink_c_bits_hasData),
    .io_resps_sink_c_bits_param(abc_mshr_0_io_resps_sink_c_bits_param),
    .io_resps_sink_c_bits_source(abc_mshr_0_io_resps_sink_c_bits_source),
    .io_resps_sink_c_bits_last(abc_mshr_0_io_resps_sink_c_bits_last),
    .io_resps_sink_c_bits_bufIdx(abc_mshr_0_io_resps_sink_c_bits_bufIdx),
    .io_resps_sink_d_valid(abc_mshr_0_io_resps_sink_d_valid),
    .io_resps_sink_d_bits_opcode(abc_mshr_0_io_resps_sink_d_bits_opcode),
    .io_resps_sink_d_bits_param(abc_mshr_0_io_resps_sink_d_bits_param),
    .io_resps_sink_d_bits_sink(abc_mshr_0_io_resps_sink_d_bits_sink),
    .io_resps_sink_d_bits_last(abc_mshr_0_io_resps_sink_d_bits_last),
    .io_resps_sink_d_bits_denied(abc_mshr_0_io_resps_sink_d_bits_denied),
    .io_resps_sink_d_bits_bufIdx(abc_mshr_0_io_resps_sink_d_bits_bufIdx),
    .io_resps_sink_e_valid(abc_mshr_0_io_resps_sink_e_valid),
    .io_resps_source_d_valid(abc_mshr_0_io_resps_source_d_valid),
    .io_nestedwb_set(abc_mshr_0_io_nestedwb_set),
    .io_nestedwb_tag(abc_mshr_0_io_nestedwb_tag),
    .io_nestedwb_btoN(abc_mshr_0_io_nestedwb_btoN),
    .io_nestedwb_btoB(abc_mshr_0_io_nestedwb_btoB),
    .io_nestedwb_bclr_dirty(abc_mshr_0_io_nestedwb_bclr_dirty),
    .io_nestedwb_bset_dirty(abc_mshr_0_io_nestedwb_bset_dirty),
    .io_nestedwb_c_set_dirty(abc_mshr_0_io_nestedwb_c_set_dirty),
    .io_nestedwb_c_set_hit(abc_mshr_0_io_nestedwb_c_set_hit),
    .io_nestedwb_clients_0_isToN(abc_mshr_0_io_nestedwb_clients_0_isToN),
    .io_nestedwb_clients_1_isToN(abc_mshr_0_io_nestedwb_clients_1_isToN),
    .io_tasks_sink_a_ready(abc_mshr_0_io_tasks_sink_a_ready),
    .io_tasks_sink_a_valid(abc_mshr_0_io_tasks_sink_a_valid),
    .io_tasks_sink_a_bits_sourceId(abc_mshr_0_io_tasks_sink_a_bits_sourceId),
    .io_tasks_sink_a_bits_set(abc_mshr_0_io_tasks_sink_a_bits_set),
    .io_tasks_sink_a_bits_tag(abc_mshr_0_io_tasks_sink_a_bits_tag),
    .io_tasks_sink_a_bits_size(abc_mshr_0_io_tasks_sink_a_bits_size),
    .io_tasks_sink_a_bits_off(abc_mshr_0_io_tasks_sink_a_bits_off),
    .io_tasks_source_bready(abc_mshr_0_io_tasks_source_bready),
    .io_tasks_source_bvalid(abc_mshr_0_io_tasks_source_bvalid),
    .io_tasks_source_bset(abc_mshr_0_io_tasks_source_bset),
    .io_tasks_source_btag(abc_mshr_0_io_tasks_source_btag),
    .io_tasks_source_bparam(abc_mshr_0_io_tasks_source_bparam),
    .io_tasks_source_bclients(abc_mshr_0_io_tasks_source_bclients),
    .io_tasks_source_bneedData(abc_mshr_0_io_tasks_source_bneedData),
    .io_tasks_sink_c_ready(abc_mshr_0_io_tasks_sink_c_ready),
    .io_tasks_sink_c_valid(abc_mshr_0_io_tasks_sink_c_valid),
    .io_tasks_sink_c_bits_sourceId(abc_mshr_0_io_tasks_sink_c_bits_sourceId),
    .io_tasks_sink_c_bits_set(abc_mshr_0_io_tasks_sink_c_bits_set),
    .io_tasks_sink_c_bits_tag(abc_mshr_0_io_tasks_sink_c_bits_tag),
    .io_tasks_sink_c_bits_size(abc_mshr_0_io_tasks_sink_c_bits_size),
    .io_tasks_sink_c_bits_way(abc_mshr_0_io_tasks_sink_c_bits_way),
    .io_tasks_sink_c_bits_off(abc_mshr_0_io_tasks_sink_c_bits_off),
    .io_tasks_sink_c_bits_bufIdx(abc_mshr_0_io_tasks_sink_c_bits_bufIdx),
    .io_tasks_sink_c_bits_opcode(abc_mshr_0_io_tasks_sink_c_bits_opcode),
    .io_tasks_sink_c_bits_param(abc_mshr_0_io_tasks_sink_c_bits_param),
    .io_tasks_sink_c_bits_source(abc_mshr_0_io_tasks_sink_c_bits_source),
    .io_tasks_sink_c_bits_save(abc_mshr_0_io_tasks_sink_c_bits_save),
    .io_tasks_sink_c_bits_drop(abc_mshr_0_io_tasks_sink_c_bits_drop),
    .io_tasks_sink_c_bits_release(abc_mshr_0_io_tasks_sink_c_bits_release),
    .io_tasks_sink_c_bits_dirty(abc_mshr_0_io_tasks_sink_c_bits_dirty),
    .io_tasks_source_d_ready(abc_mshr_0_io_tasks_source_d_ready),
    .io_tasks_source_d_valid(abc_mshr_0_io_tasks_source_d_valid),
    .io_tasks_source_d_bits_sourceId(abc_mshr_0_io_tasks_source_d_bits_sourceId),
    .io_tasks_source_d_bits_set(abc_mshr_0_io_tasks_source_d_bits_set),
    .io_tasks_source_d_bits_tag(abc_mshr_0_io_tasks_source_d_bits_tag),
    .io_tasks_source_d_bits_channel(abc_mshr_0_io_tasks_source_d_bits_channel),
    .io_tasks_source_d_bits_opcode(abc_mshr_0_io_tasks_source_d_bits_opcode),
    .io_tasks_source_d_bits_param(abc_mshr_0_io_tasks_source_d_bits_param),
    .io_tasks_source_d_bits_size(abc_mshr_0_io_tasks_source_d_bits_size),
    .io_tasks_source_d_bits_way(abc_mshr_0_io_tasks_source_d_bits_way),
    .io_tasks_source_d_bits_off(abc_mshr_0_io_tasks_source_d_bits_off),
    .io_tasks_source_d_bits_useBypass(abc_mshr_0_io_tasks_source_d_bits_useBypass),
    .io_tasks_source_d_bits_bufIdx(abc_mshr_0_io_tasks_source_d_bits_bufIdx),
    .io_tasks_source_d_bits_denied(abc_mshr_0_io_tasks_source_d_bits_denied),
    .io_tasks_source_d_bits_sinkId(abc_mshr_0_io_tasks_source_d_bits_sinkId),
    .io_tasks_source_d_bits_bypassPut(abc_mshr_0_io_tasks_source_d_bits_bypassPut),
    .io_tasks_source_d_bits_dirty(abc_mshr_0_io_tasks_source_d_bits_dirty),
    .io_tasks_source_a_ready(abc_mshr_0_io_tasks_source_a_ready),
    .io_tasks_source_a_valid(abc_mshr_0_io_tasks_source_a_valid),
    .io_tasks_source_a_bits_tag(abc_mshr_0_io_tasks_source_a_bits_tag),
    .io_tasks_source_a_bits_set(abc_mshr_0_io_tasks_source_a_bits_set),
    .io_tasks_source_a_bits_off(abc_mshr_0_io_tasks_source_a_bits_off),
    .io_tasks_source_a_bits_mask(abc_mshr_0_io_tasks_source_a_bits_mask),
    .io_tasks_source_a_bits_opcode(abc_mshr_0_io_tasks_source_a_bits_opcode),
    .io_tasks_source_a_bits_param(abc_mshr_0_io_tasks_source_a_bits_param),
    .io_tasks_source_a_bits_source(abc_mshr_0_io_tasks_source_a_bits_source),
    .io_tasks_source_a_bits_bufIdx(abc_mshr_0_io_tasks_source_a_bits_bufIdx),
    .io_tasks_source_a_bits_size(abc_mshr_0_io_tasks_source_a_bits_size),
    .io_tasks_source_a_bits_needData(abc_mshr_0_io_tasks_source_a_bits_needData),
    .io_tasks_source_a_bits_putData(abc_mshr_0_io_tasks_source_a_bits_putData),
    .io_tasks_source_c_ready(abc_mshr_0_io_tasks_source_c_ready),
    .io_tasks_source_c_valid(abc_mshr_0_io_tasks_source_c_valid),
    .io_tasks_source_c_bits_opcode(abc_mshr_0_io_tasks_source_c_bits_opcode),
    .io_tasks_source_c_bits_tag(abc_mshr_0_io_tasks_source_c_bits_tag),
    .io_tasks_source_c_bits_set(abc_mshr_0_io_tasks_source_c_bits_set),
    .io_tasks_source_c_bits_param(abc_mshr_0_io_tasks_source_c_bits_param),
    .io_tasks_source_c_bits_source(abc_mshr_0_io_tasks_source_c_bits_source),
    .io_tasks_source_c_bits_way(abc_mshr_0_io_tasks_source_c_bits_way),
    .io_tasks_source_c_bits_dirty(abc_mshr_0_io_tasks_source_c_bits_dirty),
    .io_tasks_source_e_ready(abc_mshr_0_io_tasks_source_e_ready),
    .io_tasks_source_e_valid(abc_mshr_0_io_tasks_source_e_valid),
    .io_tasks_source_e_bits_sink(abc_mshr_0_io_tasks_source_e_bits_sink),
    .io_tasks_dir_write_ready(abc_mshr_0_io_tasks_dir_write_ready),
    .io_tasks_dir_write_valid(abc_mshr_0_io_tasks_dir_write_valid),
    .io_tasks_dir_write_bits_set(abc_mshr_0_io_tasks_dir_write_bits_set),
    .io_tasks_dir_write_bits_way(abc_mshr_0_io_tasks_dir_write_bits_way),
    .io_tasks_dir_write_bits_data_dirty(abc_mshr_0_io_tasks_dir_write_bits_data_dirty),
    .io_tasks_dir_write_bits_data_state(abc_mshr_0_io_tasks_dir_write_bits_data_state),
    .io_tasks_dir_write_bits_data_clientStates_0(abc_mshr_0_io_tasks_dir_write_bits_data_clientStates_0),
    .io_tasks_dir_write_bits_data_clientStates_1(abc_mshr_0_io_tasks_dir_write_bits_data_clientStates_1),
    .io_tasks_tag_write_ready(abc_mshr_0_io_tasks_tag_write_ready),
    .io_tasks_tag_write_valid(abc_mshr_0_io_tasks_tag_write_valid),
    .io_tasks_tag_write_bits_set(abc_mshr_0_io_tasks_tag_write_bits_set),
    .io_tasks_tag_write_bits_way(abc_mshr_0_io_tasks_tag_write_bits_way),
    .io_tasks_tag_write_bits_tag(abc_mshr_0_io_tasks_tag_write_bits_tag),
    .io_tasks_client_dir_write_ready(abc_mshr_0_io_tasks_client_dir_write_ready),
    .io_tasks_client_dir_write_valid(abc_mshr_0_io_tasks_client_dir_write_valid),
    .io_tasks_client_dir_write_bits_set(abc_mshr_0_io_tasks_client_dir_write_bits_set),
    .io_tasks_client_dir_write_bits_way(abc_mshr_0_io_tasks_client_dir_write_bits_way),
    .io_tasks_client_dir_write_bits_data_0_state(abc_mshr_0_io_tasks_client_dir_write_bits_data_0_state),
    .io_tasks_client_dir_write_bits_data_1_state(abc_mshr_0_io_tasks_client_dir_write_bits_data_1_state),
    .io_tasks_client_tag_write_ready(abc_mshr_0_io_tasks_client_tag_write_ready),
    .io_tasks_client_tag_write_valid(abc_mshr_0_io_tasks_client_tag_write_valid),
    .io_tasks_client_tag_write_bits_set(abc_mshr_0_io_tasks_client_tag_write_bits_set),
    .io_tasks_client_tag_write_bits_way(abc_mshr_0_io_tasks_client_tag_write_bits_way),
    .io_tasks_client_tag_write_bits_tag(abc_mshr_0_io_tasks_client_tag_write_bits_tag),
    .io_dirResult_valid(abc_mshr_0_io_dirResult_valid),
    .io_dirResult_bits_self_dirty(abc_mshr_0_io_dirResult_bits_self_dirty),
    .io_dirResult_bits_self_state(abc_mshr_0_io_dirResult_bits_self_state),
    .io_dirResult_bits_self_clientStates_0(abc_mshr_0_io_dirResult_bits_self_clientStates_0),
    .io_dirResult_bits_self_clientStates_1(abc_mshr_0_io_dirResult_bits_self_clientStates_1),
    .io_dirResult_bits_self_hit(abc_mshr_0_io_dirResult_bits_self_hit),
    .io_dirResult_bits_self_way(abc_mshr_0_io_dirResult_bits_self_way),
    .io_dirResult_bits_self_tag(abc_mshr_0_io_dirResult_bits_self_tag),
    .io_dirResult_bits_clients_states_0_state(abc_mshr_0_io_dirResult_bits_clients_states_0_state),
    .io_dirResult_bits_clients_states_0_hit(abc_mshr_0_io_dirResult_bits_clients_states_0_hit),
    .io_dirResult_bits_clients_states_1_state(abc_mshr_0_io_dirResult_bits_clients_states_1_state),
    .io_dirResult_bits_clients_states_1_hit(abc_mshr_0_io_dirResult_bits_clients_states_1_hit),
    .io_dirResult_bits_clients_tag(abc_mshr_0_io_dirResult_bits_clients_tag),
    .io_dirResult_bits_clients_way(abc_mshr_0_io_dirResult_bits_clients_way),
    .io_c_status_set(abc_mshr_0_io_c_status_set),
    .io_c_status_tag(abc_mshr_0_io_c_status_tag),
    .io_c_status_way(abc_mshr_0_io_c_status_way),
    .io_c_status_nestedReleaseData(abc_mshr_0_io_c_status_nestedReleaseData),
    .io_c_status_releaseThrough(abc_mshr_0_io_c_status_releaseThrough),
    .io_bstatus_set(abc_mshr_0_io_bstatus_set),
    .io_bstatus_tag(abc_mshr_0_io_bstatus_tag),
    .io_bstatus_way(abc_mshr_0_io_bstatus_way),
    .io_bstatus_nestedProbeAckData(abc_mshr_0_io_bstatus_nestedProbeAckData),
    .io_bstatus_probeHelperFinish(abc_mshr_0_io_bstatus_probeHelperFinish),
    .io_bstatus_probeAckDataThrough(abc_mshr_0_io_bstatus_probeAckDataThrough),
    .io_releaseThrough(abc_mshr_0_io_releaseThrough),
    .io_probeAckDataThrough(abc_mshr_0_io_probeAckDataThrough),
    .io_is_nestedReleaseData(abc_mshr_0_io_is_nestedReleaseData),
    .io_is_nestedProbeAckData(abc_mshr_0_io_is_nestedProbeAckData),
    .io_probeHelperFinish(abc_mshr_0_io_probeHelperFinish)
  );
  MSHR abc_mshr_1 ( // @[Slice.scala 94:16]
    .clock(abc_mshr_1_clock),
    .reset(abc_mshr_1_reset),
    .io_id(abc_mshr_1_io_id),
    .io_enable(abc_mshr_1_io_enable),
    .io_alloc_valid(abc_mshr_1_io_alloc_valid),
    .io_alloc_bits_channel(abc_mshr_1_io_alloc_bits_channel),
    .io_alloc_bits_opcode(abc_mshr_1_io_alloc_bits_opcode),
    .io_alloc_bits_param(abc_mshr_1_io_alloc_bits_param),
    .io_alloc_bits_size(abc_mshr_1_io_alloc_bits_size),
    .io_alloc_bits_source(abc_mshr_1_io_alloc_bits_source),
    .io_alloc_bits_set(abc_mshr_1_io_alloc_bits_set),
    .io_alloc_bits_tag(abc_mshr_1_io_alloc_bits_tag),
    .io_alloc_bits_off(abc_mshr_1_io_alloc_bits_off),
    .io_alloc_bits_mask(abc_mshr_1_io_alloc_bits_mask),
    .io_alloc_bits_bufIdx(abc_mshr_1_io_alloc_bits_bufIdx),
    .io_alloc_bits_preferCache(abc_mshr_1_io_alloc_bits_preferCache),
    .io_alloc_bits_dirty(abc_mshr_1_io_alloc_bits_dirty),
    .io_alloc_bits_fromProbeHelper(abc_mshr_1_io_alloc_bits_fromProbeHelper),
    .io_alloc_bits_fromCmoHelper(abc_mshr_1_io_alloc_bits_fromCmoHelper),
    .io_alloc_bits_needProbeAckData(abc_mshr_1_io_alloc_bits_needProbeAckData),
    .io_status_valid(abc_mshr_1_io_status_valid),
    .io_status_bits_set(abc_mshr_1_io_status_bits_set),
    .io_status_bits_tag(abc_mshr_1_io_status_bits_tag),
    .io_status_bits_way(abc_mshr_1_io_status_bits_way),
    .io_status_bits_way_reg(abc_mshr_1_io_status_bits_way_reg),
    .io_status_bits_nestB(abc_mshr_1_io_status_bits_nestB),
    .io_status_bits_nestC(abc_mshr_1_io_status_bits_nestC),
    .io_status_bits_will_grant_data(abc_mshr_1_io_status_bits_will_grant_data),
    .io_status_bits_will_save_data(abc_mshr_1_io_status_bits_will_save_data),
    .io_status_bits_will_free(abc_mshr_1_io_status_bits_will_free),
    .io_resps_sink_c_valid(abc_mshr_1_io_resps_sink_c_valid),
    .io_resps_sink_c_bits_hasData(abc_mshr_1_io_resps_sink_c_bits_hasData),
    .io_resps_sink_c_bits_param(abc_mshr_1_io_resps_sink_c_bits_param),
    .io_resps_sink_c_bits_source(abc_mshr_1_io_resps_sink_c_bits_source),
    .io_resps_sink_c_bits_last(abc_mshr_1_io_resps_sink_c_bits_last),
    .io_resps_sink_c_bits_bufIdx(abc_mshr_1_io_resps_sink_c_bits_bufIdx),
    .io_resps_sink_d_valid(abc_mshr_1_io_resps_sink_d_valid),
    .io_resps_sink_d_bits_opcode(abc_mshr_1_io_resps_sink_d_bits_opcode),
    .io_resps_sink_d_bits_param(abc_mshr_1_io_resps_sink_d_bits_param),
    .io_resps_sink_d_bits_sink(abc_mshr_1_io_resps_sink_d_bits_sink),
    .io_resps_sink_d_bits_last(abc_mshr_1_io_resps_sink_d_bits_last),
    .io_resps_sink_d_bits_denied(abc_mshr_1_io_resps_sink_d_bits_denied),
    .io_resps_sink_d_bits_bufIdx(abc_mshr_1_io_resps_sink_d_bits_bufIdx),
    .io_resps_sink_e_valid(abc_mshr_1_io_resps_sink_e_valid),
    .io_resps_source_d_valid(abc_mshr_1_io_resps_source_d_valid),
    .io_nestedwb_set(abc_mshr_1_io_nestedwb_set),
    .io_nestedwb_tag(abc_mshr_1_io_nestedwb_tag),
    .io_nestedwb_btoN(abc_mshr_1_io_nestedwb_btoN),
    .io_nestedwb_btoB(abc_mshr_1_io_nestedwb_btoB),
    .io_nestedwb_bclr_dirty(abc_mshr_1_io_nestedwb_bclr_dirty),
    .io_nestedwb_bset_dirty(abc_mshr_1_io_nestedwb_bset_dirty),
    .io_nestedwb_c_set_dirty(abc_mshr_1_io_nestedwb_c_set_dirty),
    .io_nestedwb_c_set_hit(abc_mshr_1_io_nestedwb_c_set_hit),
    .io_nestedwb_clients_0_isToN(abc_mshr_1_io_nestedwb_clients_0_isToN),
    .io_nestedwb_clients_1_isToN(abc_mshr_1_io_nestedwb_clients_1_isToN),
    .io_tasks_sink_a_ready(abc_mshr_1_io_tasks_sink_a_ready),
    .io_tasks_sink_a_valid(abc_mshr_1_io_tasks_sink_a_valid),
    .io_tasks_sink_a_bits_sourceId(abc_mshr_1_io_tasks_sink_a_bits_sourceId),
    .io_tasks_sink_a_bits_set(abc_mshr_1_io_tasks_sink_a_bits_set),
    .io_tasks_sink_a_bits_tag(abc_mshr_1_io_tasks_sink_a_bits_tag),
    .io_tasks_sink_a_bits_size(abc_mshr_1_io_tasks_sink_a_bits_size),
    .io_tasks_sink_a_bits_off(abc_mshr_1_io_tasks_sink_a_bits_off),
    .io_tasks_source_bready(abc_mshr_1_io_tasks_source_bready),
    .io_tasks_source_bvalid(abc_mshr_1_io_tasks_source_bvalid),
    .io_tasks_source_bset(abc_mshr_1_io_tasks_source_bset),
    .io_tasks_source_btag(abc_mshr_1_io_tasks_source_btag),
    .io_tasks_source_bparam(abc_mshr_1_io_tasks_source_bparam),
    .io_tasks_source_bclients(abc_mshr_1_io_tasks_source_bclients),
    .io_tasks_source_bneedData(abc_mshr_1_io_tasks_source_bneedData),
    .io_tasks_sink_c_ready(abc_mshr_1_io_tasks_sink_c_ready),
    .io_tasks_sink_c_valid(abc_mshr_1_io_tasks_sink_c_valid),
    .io_tasks_sink_c_bits_sourceId(abc_mshr_1_io_tasks_sink_c_bits_sourceId),
    .io_tasks_sink_c_bits_set(abc_mshr_1_io_tasks_sink_c_bits_set),
    .io_tasks_sink_c_bits_tag(abc_mshr_1_io_tasks_sink_c_bits_tag),
    .io_tasks_sink_c_bits_size(abc_mshr_1_io_tasks_sink_c_bits_size),
    .io_tasks_sink_c_bits_way(abc_mshr_1_io_tasks_sink_c_bits_way),
    .io_tasks_sink_c_bits_off(abc_mshr_1_io_tasks_sink_c_bits_off),
    .io_tasks_sink_c_bits_bufIdx(abc_mshr_1_io_tasks_sink_c_bits_bufIdx),
    .io_tasks_sink_c_bits_opcode(abc_mshr_1_io_tasks_sink_c_bits_opcode),
    .io_tasks_sink_c_bits_param(abc_mshr_1_io_tasks_sink_c_bits_param),
    .io_tasks_sink_c_bits_source(abc_mshr_1_io_tasks_sink_c_bits_source),
    .io_tasks_sink_c_bits_save(abc_mshr_1_io_tasks_sink_c_bits_save),
    .io_tasks_sink_c_bits_drop(abc_mshr_1_io_tasks_sink_c_bits_drop),
    .io_tasks_sink_c_bits_release(abc_mshr_1_io_tasks_sink_c_bits_release),
    .io_tasks_sink_c_bits_dirty(abc_mshr_1_io_tasks_sink_c_bits_dirty),
    .io_tasks_source_d_ready(abc_mshr_1_io_tasks_source_d_ready),
    .io_tasks_source_d_valid(abc_mshr_1_io_tasks_source_d_valid),
    .io_tasks_source_d_bits_sourceId(abc_mshr_1_io_tasks_source_d_bits_sourceId),
    .io_tasks_source_d_bits_set(abc_mshr_1_io_tasks_source_d_bits_set),
    .io_tasks_source_d_bits_tag(abc_mshr_1_io_tasks_source_d_bits_tag),
    .io_tasks_source_d_bits_channel(abc_mshr_1_io_tasks_source_d_bits_channel),
    .io_tasks_source_d_bits_opcode(abc_mshr_1_io_tasks_source_d_bits_opcode),
    .io_tasks_source_d_bits_param(abc_mshr_1_io_tasks_source_d_bits_param),
    .io_tasks_source_d_bits_size(abc_mshr_1_io_tasks_source_d_bits_size),
    .io_tasks_source_d_bits_way(abc_mshr_1_io_tasks_source_d_bits_way),
    .io_tasks_source_d_bits_off(abc_mshr_1_io_tasks_source_d_bits_off),
    .io_tasks_source_d_bits_useBypass(abc_mshr_1_io_tasks_source_d_bits_useBypass),
    .io_tasks_source_d_bits_bufIdx(abc_mshr_1_io_tasks_source_d_bits_bufIdx),
    .io_tasks_source_d_bits_denied(abc_mshr_1_io_tasks_source_d_bits_denied),
    .io_tasks_source_d_bits_sinkId(abc_mshr_1_io_tasks_source_d_bits_sinkId),
    .io_tasks_source_d_bits_bypassPut(abc_mshr_1_io_tasks_source_d_bits_bypassPut),
    .io_tasks_source_d_bits_dirty(abc_mshr_1_io_tasks_source_d_bits_dirty),
    .io_tasks_source_a_ready(abc_mshr_1_io_tasks_source_a_ready),
    .io_tasks_source_a_valid(abc_mshr_1_io_tasks_source_a_valid),
    .io_tasks_source_a_bits_tag(abc_mshr_1_io_tasks_source_a_bits_tag),
    .io_tasks_source_a_bits_set(abc_mshr_1_io_tasks_source_a_bits_set),
    .io_tasks_source_a_bits_off(abc_mshr_1_io_tasks_source_a_bits_off),
    .io_tasks_source_a_bits_mask(abc_mshr_1_io_tasks_source_a_bits_mask),
    .io_tasks_source_a_bits_opcode(abc_mshr_1_io_tasks_source_a_bits_opcode),
    .io_tasks_source_a_bits_param(abc_mshr_1_io_tasks_source_a_bits_param),
    .io_tasks_source_a_bits_source(abc_mshr_1_io_tasks_source_a_bits_source),
    .io_tasks_source_a_bits_bufIdx(abc_mshr_1_io_tasks_source_a_bits_bufIdx),
    .io_tasks_source_a_bits_size(abc_mshr_1_io_tasks_source_a_bits_size),
    .io_tasks_source_a_bits_needData(abc_mshr_1_io_tasks_source_a_bits_needData),
    .io_tasks_source_a_bits_putData(abc_mshr_1_io_tasks_source_a_bits_putData),
    .io_tasks_source_c_ready(abc_mshr_1_io_tasks_source_c_ready),
    .io_tasks_source_c_valid(abc_mshr_1_io_tasks_source_c_valid),
    .io_tasks_source_c_bits_opcode(abc_mshr_1_io_tasks_source_c_bits_opcode),
    .io_tasks_source_c_bits_tag(abc_mshr_1_io_tasks_source_c_bits_tag),
    .io_tasks_source_c_bits_set(abc_mshr_1_io_tasks_source_c_bits_set),
    .io_tasks_source_c_bits_param(abc_mshr_1_io_tasks_source_c_bits_param),
    .io_tasks_source_c_bits_source(abc_mshr_1_io_tasks_source_c_bits_source),
    .io_tasks_source_c_bits_way(abc_mshr_1_io_tasks_source_c_bits_way),
    .io_tasks_source_c_bits_dirty(abc_mshr_1_io_tasks_source_c_bits_dirty),
    .io_tasks_source_e_ready(abc_mshr_1_io_tasks_source_e_ready),
    .io_tasks_source_e_valid(abc_mshr_1_io_tasks_source_e_valid),
    .io_tasks_source_e_bits_sink(abc_mshr_1_io_tasks_source_e_bits_sink),
    .io_tasks_dir_write_ready(abc_mshr_1_io_tasks_dir_write_ready),
    .io_tasks_dir_write_valid(abc_mshr_1_io_tasks_dir_write_valid),
    .io_tasks_dir_write_bits_set(abc_mshr_1_io_tasks_dir_write_bits_set),
    .io_tasks_dir_write_bits_way(abc_mshr_1_io_tasks_dir_write_bits_way),
    .io_tasks_dir_write_bits_data_dirty(abc_mshr_1_io_tasks_dir_write_bits_data_dirty),
    .io_tasks_dir_write_bits_data_state(abc_mshr_1_io_tasks_dir_write_bits_data_state),
    .io_tasks_dir_write_bits_data_clientStates_0(abc_mshr_1_io_tasks_dir_write_bits_data_clientStates_0),
    .io_tasks_dir_write_bits_data_clientStates_1(abc_mshr_1_io_tasks_dir_write_bits_data_clientStates_1),
    .io_tasks_tag_write_ready(abc_mshr_1_io_tasks_tag_write_ready),
    .io_tasks_tag_write_valid(abc_mshr_1_io_tasks_tag_write_valid),
    .io_tasks_tag_write_bits_set(abc_mshr_1_io_tasks_tag_write_bits_set),
    .io_tasks_tag_write_bits_way(abc_mshr_1_io_tasks_tag_write_bits_way),
    .io_tasks_tag_write_bits_tag(abc_mshr_1_io_tasks_tag_write_bits_tag),
    .io_tasks_client_dir_write_ready(abc_mshr_1_io_tasks_client_dir_write_ready),
    .io_tasks_client_dir_write_valid(abc_mshr_1_io_tasks_client_dir_write_valid),
    .io_tasks_client_dir_write_bits_set(abc_mshr_1_io_tasks_client_dir_write_bits_set),
    .io_tasks_client_dir_write_bits_way(abc_mshr_1_io_tasks_client_dir_write_bits_way),
    .io_tasks_client_dir_write_bits_data_0_state(abc_mshr_1_io_tasks_client_dir_write_bits_data_0_state),
    .io_tasks_client_dir_write_bits_data_1_state(abc_mshr_1_io_tasks_client_dir_write_bits_data_1_state),
    .io_tasks_client_tag_write_ready(abc_mshr_1_io_tasks_client_tag_write_ready),
    .io_tasks_client_tag_write_valid(abc_mshr_1_io_tasks_client_tag_write_valid),
    .io_tasks_client_tag_write_bits_set(abc_mshr_1_io_tasks_client_tag_write_bits_set),
    .io_tasks_client_tag_write_bits_way(abc_mshr_1_io_tasks_client_tag_write_bits_way),
    .io_tasks_client_tag_write_bits_tag(abc_mshr_1_io_tasks_client_tag_write_bits_tag),
    .io_dirResult_valid(abc_mshr_1_io_dirResult_valid),
    .io_dirResult_bits_self_dirty(abc_mshr_1_io_dirResult_bits_self_dirty),
    .io_dirResult_bits_self_state(abc_mshr_1_io_dirResult_bits_self_state),
    .io_dirResult_bits_self_clientStates_0(abc_mshr_1_io_dirResult_bits_self_clientStates_0),
    .io_dirResult_bits_self_clientStates_1(abc_mshr_1_io_dirResult_bits_self_clientStates_1),
    .io_dirResult_bits_self_hit(abc_mshr_1_io_dirResult_bits_self_hit),
    .io_dirResult_bits_self_way(abc_mshr_1_io_dirResult_bits_self_way),
    .io_dirResult_bits_self_tag(abc_mshr_1_io_dirResult_bits_self_tag),
    .io_dirResult_bits_clients_states_0_state(abc_mshr_1_io_dirResult_bits_clients_states_0_state),
    .io_dirResult_bits_clients_states_0_hit(abc_mshr_1_io_dirResult_bits_clients_states_0_hit),
    .io_dirResult_bits_clients_states_1_state(abc_mshr_1_io_dirResult_bits_clients_states_1_state),
    .io_dirResult_bits_clients_states_1_hit(abc_mshr_1_io_dirResult_bits_clients_states_1_hit),
    .io_dirResult_bits_clients_tag(abc_mshr_1_io_dirResult_bits_clients_tag),
    .io_dirResult_bits_clients_way(abc_mshr_1_io_dirResult_bits_clients_way),
    .io_c_status_set(abc_mshr_1_io_c_status_set),
    .io_c_status_tag(abc_mshr_1_io_c_status_tag),
    .io_c_status_way(abc_mshr_1_io_c_status_way),
    .io_c_status_nestedReleaseData(abc_mshr_1_io_c_status_nestedReleaseData),
    .io_c_status_releaseThrough(abc_mshr_1_io_c_status_releaseThrough),
    .io_bstatus_set(abc_mshr_1_io_bstatus_set),
    .io_bstatus_tag(abc_mshr_1_io_bstatus_tag),
    .io_bstatus_way(abc_mshr_1_io_bstatus_way),
    .io_bstatus_nestedProbeAckData(abc_mshr_1_io_bstatus_nestedProbeAckData),
    .io_bstatus_probeHelperFinish(abc_mshr_1_io_bstatus_probeHelperFinish),
    .io_bstatus_probeAckDataThrough(abc_mshr_1_io_bstatus_probeAckDataThrough),
    .io_releaseThrough(abc_mshr_1_io_releaseThrough),
    .io_probeAckDataThrough(abc_mshr_1_io_probeAckDataThrough),
    .io_is_nestedReleaseData(abc_mshr_1_io_is_nestedReleaseData),
    .io_is_nestedProbeAckData(abc_mshr_1_io_is_nestedProbeAckData),
    .io_probeHelperFinish(abc_mshr_1_io_probeHelperFinish)
  );
  MSHR abc_mshr_2 ( // @[Slice.scala 94:16]
    .clock(abc_mshr_2_clock),
    .reset(abc_mshr_2_reset),
    .io_id(abc_mshr_2_io_id),
    .io_enable(abc_mshr_2_io_enable),
    .io_alloc_valid(abc_mshr_2_io_alloc_valid),
    .io_alloc_bits_channel(abc_mshr_2_io_alloc_bits_channel),
    .io_alloc_bits_opcode(abc_mshr_2_io_alloc_bits_opcode),
    .io_alloc_bits_param(abc_mshr_2_io_alloc_bits_param),
    .io_alloc_bits_size(abc_mshr_2_io_alloc_bits_size),
    .io_alloc_bits_source(abc_mshr_2_io_alloc_bits_source),
    .io_alloc_bits_set(abc_mshr_2_io_alloc_bits_set),
    .io_alloc_bits_tag(abc_mshr_2_io_alloc_bits_tag),
    .io_alloc_bits_off(abc_mshr_2_io_alloc_bits_off),
    .io_alloc_bits_mask(abc_mshr_2_io_alloc_bits_mask),
    .io_alloc_bits_bufIdx(abc_mshr_2_io_alloc_bits_bufIdx),
    .io_alloc_bits_preferCache(abc_mshr_2_io_alloc_bits_preferCache),
    .io_alloc_bits_dirty(abc_mshr_2_io_alloc_bits_dirty),
    .io_alloc_bits_fromProbeHelper(abc_mshr_2_io_alloc_bits_fromProbeHelper),
    .io_alloc_bits_fromCmoHelper(abc_mshr_2_io_alloc_bits_fromCmoHelper),
    .io_alloc_bits_needProbeAckData(abc_mshr_2_io_alloc_bits_needProbeAckData),
    .io_status_valid(abc_mshr_2_io_status_valid),
    .io_status_bits_set(abc_mshr_2_io_status_bits_set),
    .io_status_bits_tag(abc_mshr_2_io_status_bits_tag),
    .io_status_bits_way(abc_mshr_2_io_status_bits_way),
    .io_status_bits_way_reg(abc_mshr_2_io_status_bits_way_reg),
    .io_status_bits_nestB(abc_mshr_2_io_status_bits_nestB),
    .io_status_bits_nestC(abc_mshr_2_io_status_bits_nestC),
    .io_status_bits_will_grant_data(abc_mshr_2_io_status_bits_will_grant_data),
    .io_status_bits_will_save_data(abc_mshr_2_io_status_bits_will_save_data),
    .io_status_bits_will_free(abc_mshr_2_io_status_bits_will_free),
    .io_resps_sink_c_valid(abc_mshr_2_io_resps_sink_c_valid),
    .io_resps_sink_c_bits_hasData(abc_mshr_2_io_resps_sink_c_bits_hasData),
    .io_resps_sink_c_bits_param(abc_mshr_2_io_resps_sink_c_bits_param),
    .io_resps_sink_c_bits_source(abc_mshr_2_io_resps_sink_c_bits_source),
    .io_resps_sink_c_bits_last(abc_mshr_2_io_resps_sink_c_bits_last),
    .io_resps_sink_c_bits_bufIdx(abc_mshr_2_io_resps_sink_c_bits_bufIdx),
    .io_resps_sink_d_valid(abc_mshr_2_io_resps_sink_d_valid),
    .io_resps_sink_d_bits_opcode(abc_mshr_2_io_resps_sink_d_bits_opcode),
    .io_resps_sink_d_bits_param(abc_mshr_2_io_resps_sink_d_bits_param),
    .io_resps_sink_d_bits_sink(abc_mshr_2_io_resps_sink_d_bits_sink),
    .io_resps_sink_d_bits_last(abc_mshr_2_io_resps_sink_d_bits_last),
    .io_resps_sink_d_bits_denied(abc_mshr_2_io_resps_sink_d_bits_denied),
    .io_resps_sink_d_bits_bufIdx(abc_mshr_2_io_resps_sink_d_bits_bufIdx),
    .io_resps_sink_e_valid(abc_mshr_2_io_resps_sink_e_valid),
    .io_resps_source_d_valid(abc_mshr_2_io_resps_source_d_valid),
    .io_nestedwb_set(abc_mshr_2_io_nestedwb_set),
    .io_nestedwb_tag(abc_mshr_2_io_nestedwb_tag),
    .io_nestedwb_btoN(abc_mshr_2_io_nestedwb_btoN),
    .io_nestedwb_btoB(abc_mshr_2_io_nestedwb_btoB),
    .io_nestedwb_bclr_dirty(abc_mshr_2_io_nestedwb_bclr_dirty),
    .io_nestedwb_bset_dirty(abc_mshr_2_io_nestedwb_bset_dirty),
    .io_nestedwb_c_set_dirty(abc_mshr_2_io_nestedwb_c_set_dirty),
    .io_nestedwb_c_set_hit(abc_mshr_2_io_nestedwb_c_set_hit),
    .io_nestedwb_clients_0_isToN(abc_mshr_2_io_nestedwb_clients_0_isToN),
    .io_nestedwb_clients_1_isToN(abc_mshr_2_io_nestedwb_clients_1_isToN),
    .io_tasks_sink_a_ready(abc_mshr_2_io_tasks_sink_a_ready),
    .io_tasks_sink_a_valid(abc_mshr_2_io_tasks_sink_a_valid),
    .io_tasks_sink_a_bits_sourceId(abc_mshr_2_io_tasks_sink_a_bits_sourceId),
    .io_tasks_sink_a_bits_set(abc_mshr_2_io_tasks_sink_a_bits_set),
    .io_tasks_sink_a_bits_tag(abc_mshr_2_io_tasks_sink_a_bits_tag),
    .io_tasks_sink_a_bits_size(abc_mshr_2_io_tasks_sink_a_bits_size),
    .io_tasks_sink_a_bits_off(abc_mshr_2_io_tasks_sink_a_bits_off),
    .io_tasks_source_bready(abc_mshr_2_io_tasks_source_bready),
    .io_tasks_source_bvalid(abc_mshr_2_io_tasks_source_bvalid),
    .io_tasks_source_bset(abc_mshr_2_io_tasks_source_bset),
    .io_tasks_source_btag(abc_mshr_2_io_tasks_source_btag),
    .io_tasks_source_bparam(abc_mshr_2_io_tasks_source_bparam),
    .io_tasks_source_bclients(abc_mshr_2_io_tasks_source_bclients),
    .io_tasks_source_bneedData(abc_mshr_2_io_tasks_source_bneedData),
    .io_tasks_sink_c_ready(abc_mshr_2_io_tasks_sink_c_ready),
    .io_tasks_sink_c_valid(abc_mshr_2_io_tasks_sink_c_valid),
    .io_tasks_sink_c_bits_sourceId(abc_mshr_2_io_tasks_sink_c_bits_sourceId),
    .io_tasks_sink_c_bits_set(abc_mshr_2_io_tasks_sink_c_bits_set),
    .io_tasks_sink_c_bits_tag(abc_mshr_2_io_tasks_sink_c_bits_tag),
    .io_tasks_sink_c_bits_size(abc_mshr_2_io_tasks_sink_c_bits_size),
    .io_tasks_sink_c_bits_way(abc_mshr_2_io_tasks_sink_c_bits_way),
    .io_tasks_sink_c_bits_off(abc_mshr_2_io_tasks_sink_c_bits_off),
    .io_tasks_sink_c_bits_bufIdx(abc_mshr_2_io_tasks_sink_c_bits_bufIdx),
    .io_tasks_sink_c_bits_opcode(abc_mshr_2_io_tasks_sink_c_bits_opcode),
    .io_tasks_sink_c_bits_param(abc_mshr_2_io_tasks_sink_c_bits_param),
    .io_tasks_sink_c_bits_source(abc_mshr_2_io_tasks_sink_c_bits_source),
    .io_tasks_sink_c_bits_save(abc_mshr_2_io_tasks_sink_c_bits_save),
    .io_tasks_sink_c_bits_drop(abc_mshr_2_io_tasks_sink_c_bits_drop),
    .io_tasks_sink_c_bits_release(abc_mshr_2_io_tasks_sink_c_bits_release),
    .io_tasks_sink_c_bits_dirty(abc_mshr_2_io_tasks_sink_c_bits_dirty),
    .io_tasks_source_d_ready(abc_mshr_2_io_tasks_source_d_ready),
    .io_tasks_source_d_valid(abc_mshr_2_io_tasks_source_d_valid),
    .io_tasks_source_d_bits_sourceId(abc_mshr_2_io_tasks_source_d_bits_sourceId),
    .io_tasks_source_d_bits_set(abc_mshr_2_io_tasks_source_d_bits_set),
    .io_tasks_source_d_bits_tag(abc_mshr_2_io_tasks_source_d_bits_tag),
    .io_tasks_source_d_bits_channel(abc_mshr_2_io_tasks_source_d_bits_channel),
    .io_tasks_source_d_bits_opcode(abc_mshr_2_io_tasks_source_d_bits_opcode),
    .io_tasks_source_d_bits_param(abc_mshr_2_io_tasks_source_d_bits_param),
    .io_tasks_source_d_bits_size(abc_mshr_2_io_tasks_source_d_bits_size),
    .io_tasks_source_d_bits_way(abc_mshr_2_io_tasks_source_d_bits_way),
    .io_tasks_source_d_bits_off(abc_mshr_2_io_tasks_source_d_bits_off),
    .io_tasks_source_d_bits_useBypass(abc_mshr_2_io_tasks_source_d_bits_useBypass),
    .io_tasks_source_d_bits_bufIdx(abc_mshr_2_io_tasks_source_d_bits_bufIdx),
    .io_tasks_source_d_bits_denied(abc_mshr_2_io_tasks_source_d_bits_denied),
    .io_tasks_source_d_bits_sinkId(abc_mshr_2_io_tasks_source_d_bits_sinkId),
    .io_tasks_source_d_bits_bypassPut(abc_mshr_2_io_tasks_source_d_bits_bypassPut),
    .io_tasks_source_d_bits_dirty(abc_mshr_2_io_tasks_source_d_bits_dirty),
    .io_tasks_source_a_ready(abc_mshr_2_io_tasks_source_a_ready),
    .io_tasks_source_a_valid(abc_mshr_2_io_tasks_source_a_valid),
    .io_tasks_source_a_bits_tag(abc_mshr_2_io_tasks_source_a_bits_tag),
    .io_tasks_source_a_bits_set(abc_mshr_2_io_tasks_source_a_bits_set),
    .io_tasks_source_a_bits_off(abc_mshr_2_io_tasks_source_a_bits_off),
    .io_tasks_source_a_bits_mask(abc_mshr_2_io_tasks_source_a_bits_mask),
    .io_tasks_source_a_bits_opcode(abc_mshr_2_io_tasks_source_a_bits_opcode),
    .io_tasks_source_a_bits_param(abc_mshr_2_io_tasks_source_a_bits_param),
    .io_tasks_source_a_bits_source(abc_mshr_2_io_tasks_source_a_bits_source),
    .io_tasks_source_a_bits_bufIdx(abc_mshr_2_io_tasks_source_a_bits_bufIdx),
    .io_tasks_source_a_bits_size(abc_mshr_2_io_tasks_source_a_bits_size),
    .io_tasks_source_a_bits_needData(abc_mshr_2_io_tasks_source_a_bits_needData),
    .io_tasks_source_a_bits_putData(abc_mshr_2_io_tasks_source_a_bits_putData),
    .io_tasks_source_c_ready(abc_mshr_2_io_tasks_source_c_ready),
    .io_tasks_source_c_valid(abc_mshr_2_io_tasks_source_c_valid),
    .io_tasks_source_c_bits_opcode(abc_mshr_2_io_tasks_source_c_bits_opcode),
    .io_tasks_source_c_bits_tag(abc_mshr_2_io_tasks_source_c_bits_tag),
    .io_tasks_source_c_bits_set(abc_mshr_2_io_tasks_source_c_bits_set),
    .io_tasks_source_c_bits_param(abc_mshr_2_io_tasks_source_c_bits_param),
    .io_tasks_source_c_bits_source(abc_mshr_2_io_tasks_source_c_bits_source),
    .io_tasks_source_c_bits_way(abc_mshr_2_io_tasks_source_c_bits_way),
    .io_tasks_source_c_bits_dirty(abc_mshr_2_io_tasks_source_c_bits_dirty),
    .io_tasks_source_e_ready(abc_mshr_2_io_tasks_source_e_ready),
    .io_tasks_source_e_valid(abc_mshr_2_io_tasks_source_e_valid),
    .io_tasks_source_e_bits_sink(abc_mshr_2_io_tasks_source_e_bits_sink),
    .io_tasks_dir_write_ready(abc_mshr_2_io_tasks_dir_write_ready),
    .io_tasks_dir_write_valid(abc_mshr_2_io_tasks_dir_write_valid),
    .io_tasks_dir_write_bits_set(abc_mshr_2_io_tasks_dir_write_bits_set),
    .io_tasks_dir_write_bits_way(abc_mshr_2_io_tasks_dir_write_bits_way),
    .io_tasks_dir_write_bits_data_dirty(abc_mshr_2_io_tasks_dir_write_bits_data_dirty),
    .io_tasks_dir_write_bits_data_state(abc_mshr_2_io_tasks_dir_write_bits_data_state),
    .io_tasks_dir_write_bits_data_clientStates_0(abc_mshr_2_io_tasks_dir_write_bits_data_clientStates_0),
    .io_tasks_dir_write_bits_data_clientStates_1(abc_mshr_2_io_tasks_dir_write_bits_data_clientStates_1),
    .io_tasks_tag_write_ready(abc_mshr_2_io_tasks_tag_write_ready),
    .io_tasks_tag_write_valid(abc_mshr_2_io_tasks_tag_write_valid),
    .io_tasks_tag_write_bits_set(abc_mshr_2_io_tasks_tag_write_bits_set),
    .io_tasks_tag_write_bits_way(abc_mshr_2_io_tasks_tag_write_bits_way),
    .io_tasks_tag_write_bits_tag(abc_mshr_2_io_tasks_tag_write_bits_tag),
    .io_tasks_client_dir_write_ready(abc_mshr_2_io_tasks_client_dir_write_ready),
    .io_tasks_client_dir_write_valid(abc_mshr_2_io_tasks_client_dir_write_valid),
    .io_tasks_client_dir_write_bits_set(abc_mshr_2_io_tasks_client_dir_write_bits_set),
    .io_tasks_client_dir_write_bits_way(abc_mshr_2_io_tasks_client_dir_write_bits_way),
    .io_tasks_client_dir_write_bits_data_0_state(abc_mshr_2_io_tasks_client_dir_write_bits_data_0_state),
    .io_tasks_client_dir_write_bits_data_1_state(abc_mshr_2_io_tasks_client_dir_write_bits_data_1_state),
    .io_tasks_client_tag_write_ready(abc_mshr_2_io_tasks_client_tag_write_ready),
    .io_tasks_client_tag_write_valid(abc_mshr_2_io_tasks_client_tag_write_valid),
    .io_tasks_client_tag_write_bits_set(abc_mshr_2_io_tasks_client_tag_write_bits_set),
    .io_tasks_client_tag_write_bits_way(abc_mshr_2_io_tasks_client_tag_write_bits_way),
    .io_tasks_client_tag_write_bits_tag(abc_mshr_2_io_tasks_client_tag_write_bits_tag),
    .io_dirResult_valid(abc_mshr_2_io_dirResult_valid),
    .io_dirResult_bits_self_dirty(abc_mshr_2_io_dirResult_bits_self_dirty),
    .io_dirResult_bits_self_state(abc_mshr_2_io_dirResult_bits_self_state),
    .io_dirResult_bits_self_clientStates_0(abc_mshr_2_io_dirResult_bits_self_clientStates_0),
    .io_dirResult_bits_self_clientStates_1(abc_mshr_2_io_dirResult_bits_self_clientStates_1),
    .io_dirResult_bits_self_hit(abc_mshr_2_io_dirResult_bits_self_hit),
    .io_dirResult_bits_self_way(abc_mshr_2_io_dirResult_bits_self_way),
    .io_dirResult_bits_self_tag(abc_mshr_2_io_dirResult_bits_self_tag),
    .io_dirResult_bits_clients_states_0_state(abc_mshr_2_io_dirResult_bits_clients_states_0_state),
    .io_dirResult_bits_clients_states_0_hit(abc_mshr_2_io_dirResult_bits_clients_states_0_hit),
    .io_dirResult_bits_clients_states_1_state(abc_mshr_2_io_dirResult_bits_clients_states_1_state),
    .io_dirResult_bits_clients_states_1_hit(abc_mshr_2_io_dirResult_bits_clients_states_1_hit),
    .io_dirResult_bits_clients_tag(abc_mshr_2_io_dirResult_bits_clients_tag),
    .io_dirResult_bits_clients_way(abc_mshr_2_io_dirResult_bits_clients_way),
    .io_c_status_set(abc_mshr_2_io_c_status_set),
    .io_c_status_tag(abc_mshr_2_io_c_status_tag),
    .io_c_status_way(abc_mshr_2_io_c_status_way),
    .io_c_status_nestedReleaseData(abc_mshr_2_io_c_status_nestedReleaseData),
    .io_c_status_releaseThrough(abc_mshr_2_io_c_status_releaseThrough),
    .io_bstatus_set(abc_mshr_2_io_bstatus_set),
    .io_bstatus_tag(abc_mshr_2_io_bstatus_tag),
    .io_bstatus_way(abc_mshr_2_io_bstatus_way),
    .io_bstatus_nestedProbeAckData(abc_mshr_2_io_bstatus_nestedProbeAckData),
    .io_bstatus_probeHelperFinish(abc_mshr_2_io_bstatus_probeHelperFinish),
    .io_bstatus_probeAckDataThrough(abc_mshr_2_io_bstatus_probeAckDataThrough),
    .io_releaseThrough(abc_mshr_2_io_releaseThrough),
    .io_probeAckDataThrough(abc_mshr_2_io_probeAckDataThrough),
    .io_is_nestedReleaseData(abc_mshr_2_io_is_nestedReleaseData),
    .io_is_nestedProbeAckData(abc_mshr_2_io_is_nestedProbeAckData),
    .io_probeHelperFinish(abc_mshr_2_io_probeHelperFinish)
  );
  MSHR abc_mshr_3 ( // @[Slice.scala 94:16]
    .clock(abc_mshr_3_clock),
    .reset(abc_mshr_3_reset),
    .io_id(abc_mshr_3_io_id),
    .io_enable(abc_mshr_3_io_enable),
    .io_alloc_valid(abc_mshr_3_io_alloc_valid),
    .io_alloc_bits_channel(abc_mshr_3_io_alloc_bits_channel),
    .io_alloc_bits_opcode(abc_mshr_3_io_alloc_bits_opcode),
    .io_alloc_bits_param(abc_mshr_3_io_alloc_bits_param),
    .io_alloc_bits_size(abc_mshr_3_io_alloc_bits_size),
    .io_alloc_bits_source(abc_mshr_3_io_alloc_bits_source),
    .io_alloc_bits_set(abc_mshr_3_io_alloc_bits_set),
    .io_alloc_bits_tag(abc_mshr_3_io_alloc_bits_tag),
    .io_alloc_bits_off(abc_mshr_3_io_alloc_bits_off),
    .io_alloc_bits_mask(abc_mshr_3_io_alloc_bits_mask),
    .io_alloc_bits_bufIdx(abc_mshr_3_io_alloc_bits_bufIdx),
    .io_alloc_bits_preferCache(abc_mshr_3_io_alloc_bits_preferCache),
    .io_alloc_bits_dirty(abc_mshr_3_io_alloc_bits_dirty),
    .io_alloc_bits_fromProbeHelper(abc_mshr_3_io_alloc_bits_fromProbeHelper),
    .io_alloc_bits_fromCmoHelper(abc_mshr_3_io_alloc_bits_fromCmoHelper),
    .io_alloc_bits_needProbeAckData(abc_mshr_3_io_alloc_bits_needProbeAckData),
    .io_status_valid(abc_mshr_3_io_status_valid),
    .io_status_bits_set(abc_mshr_3_io_status_bits_set),
    .io_status_bits_tag(abc_mshr_3_io_status_bits_tag),
    .io_status_bits_way(abc_mshr_3_io_status_bits_way),
    .io_status_bits_way_reg(abc_mshr_3_io_status_bits_way_reg),
    .io_status_bits_nestB(abc_mshr_3_io_status_bits_nestB),
    .io_status_bits_nestC(abc_mshr_3_io_status_bits_nestC),
    .io_status_bits_will_grant_data(abc_mshr_3_io_status_bits_will_grant_data),
    .io_status_bits_will_save_data(abc_mshr_3_io_status_bits_will_save_data),
    .io_status_bits_will_free(abc_mshr_3_io_status_bits_will_free),
    .io_resps_sink_c_valid(abc_mshr_3_io_resps_sink_c_valid),
    .io_resps_sink_c_bits_hasData(abc_mshr_3_io_resps_sink_c_bits_hasData),
    .io_resps_sink_c_bits_param(abc_mshr_3_io_resps_sink_c_bits_param),
    .io_resps_sink_c_bits_source(abc_mshr_3_io_resps_sink_c_bits_source),
    .io_resps_sink_c_bits_last(abc_mshr_3_io_resps_sink_c_bits_last),
    .io_resps_sink_c_bits_bufIdx(abc_mshr_3_io_resps_sink_c_bits_bufIdx),
    .io_resps_sink_d_valid(abc_mshr_3_io_resps_sink_d_valid),
    .io_resps_sink_d_bits_opcode(abc_mshr_3_io_resps_sink_d_bits_opcode),
    .io_resps_sink_d_bits_param(abc_mshr_3_io_resps_sink_d_bits_param),
    .io_resps_sink_d_bits_sink(abc_mshr_3_io_resps_sink_d_bits_sink),
    .io_resps_sink_d_bits_last(abc_mshr_3_io_resps_sink_d_bits_last),
    .io_resps_sink_d_bits_denied(abc_mshr_3_io_resps_sink_d_bits_denied),
    .io_resps_sink_d_bits_bufIdx(abc_mshr_3_io_resps_sink_d_bits_bufIdx),
    .io_resps_sink_e_valid(abc_mshr_3_io_resps_sink_e_valid),
    .io_resps_source_d_valid(abc_mshr_3_io_resps_source_d_valid),
    .io_nestedwb_set(abc_mshr_3_io_nestedwb_set),
    .io_nestedwb_tag(abc_mshr_3_io_nestedwb_tag),
    .io_nestedwb_btoN(abc_mshr_3_io_nestedwb_btoN),
    .io_nestedwb_btoB(abc_mshr_3_io_nestedwb_btoB),
    .io_nestedwb_bclr_dirty(abc_mshr_3_io_nestedwb_bclr_dirty),
    .io_nestedwb_bset_dirty(abc_mshr_3_io_nestedwb_bset_dirty),
    .io_nestedwb_c_set_dirty(abc_mshr_3_io_nestedwb_c_set_dirty),
    .io_nestedwb_c_set_hit(abc_mshr_3_io_nestedwb_c_set_hit),
    .io_nestedwb_clients_0_isToN(abc_mshr_3_io_nestedwb_clients_0_isToN),
    .io_nestedwb_clients_1_isToN(abc_mshr_3_io_nestedwb_clients_1_isToN),
    .io_tasks_sink_a_ready(abc_mshr_3_io_tasks_sink_a_ready),
    .io_tasks_sink_a_valid(abc_mshr_3_io_tasks_sink_a_valid),
    .io_tasks_sink_a_bits_sourceId(abc_mshr_3_io_tasks_sink_a_bits_sourceId),
    .io_tasks_sink_a_bits_set(abc_mshr_3_io_tasks_sink_a_bits_set),
    .io_tasks_sink_a_bits_tag(abc_mshr_3_io_tasks_sink_a_bits_tag),
    .io_tasks_sink_a_bits_size(abc_mshr_3_io_tasks_sink_a_bits_size),
    .io_tasks_sink_a_bits_off(abc_mshr_3_io_tasks_sink_a_bits_off),
    .io_tasks_source_bready(abc_mshr_3_io_tasks_source_bready),
    .io_tasks_source_bvalid(abc_mshr_3_io_tasks_source_bvalid),
    .io_tasks_source_bset(abc_mshr_3_io_tasks_source_bset),
    .io_tasks_source_btag(abc_mshr_3_io_tasks_source_btag),
    .io_tasks_source_bparam(abc_mshr_3_io_tasks_source_bparam),
    .io_tasks_source_bclients(abc_mshr_3_io_tasks_source_bclients),
    .io_tasks_source_bneedData(abc_mshr_3_io_tasks_source_bneedData),
    .io_tasks_sink_c_ready(abc_mshr_3_io_tasks_sink_c_ready),
    .io_tasks_sink_c_valid(abc_mshr_3_io_tasks_sink_c_valid),
    .io_tasks_sink_c_bits_sourceId(abc_mshr_3_io_tasks_sink_c_bits_sourceId),
    .io_tasks_sink_c_bits_set(abc_mshr_3_io_tasks_sink_c_bits_set),
    .io_tasks_sink_c_bits_tag(abc_mshr_3_io_tasks_sink_c_bits_tag),
    .io_tasks_sink_c_bits_size(abc_mshr_3_io_tasks_sink_c_bits_size),
    .io_tasks_sink_c_bits_way(abc_mshr_3_io_tasks_sink_c_bits_way),
    .io_tasks_sink_c_bits_off(abc_mshr_3_io_tasks_sink_c_bits_off),
    .io_tasks_sink_c_bits_bufIdx(abc_mshr_3_io_tasks_sink_c_bits_bufIdx),
    .io_tasks_sink_c_bits_opcode(abc_mshr_3_io_tasks_sink_c_bits_opcode),
    .io_tasks_sink_c_bits_param(abc_mshr_3_io_tasks_sink_c_bits_param),
    .io_tasks_sink_c_bits_source(abc_mshr_3_io_tasks_sink_c_bits_source),
    .io_tasks_sink_c_bits_save(abc_mshr_3_io_tasks_sink_c_bits_save),
    .io_tasks_sink_c_bits_drop(abc_mshr_3_io_tasks_sink_c_bits_drop),
    .io_tasks_sink_c_bits_release(abc_mshr_3_io_tasks_sink_c_bits_release),
    .io_tasks_sink_c_bits_dirty(abc_mshr_3_io_tasks_sink_c_bits_dirty),
    .io_tasks_source_d_ready(abc_mshr_3_io_tasks_source_d_ready),
    .io_tasks_source_d_valid(abc_mshr_3_io_tasks_source_d_valid),
    .io_tasks_source_d_bits_sourceId(abc_mshr_3_io_tasks_source_d_bits_sourceId),
    .io_tasks_source_d_bits_set(abc_mshr_3_io_tasks_source_d_bits_set),
    .io_tasks_source_d_bits_tag(abc_mshr_3_io_tasks_source_d_bits_tag),
    .io_tasks_source_d_bits_channel(abc_mshr_3_io_tasks_source_d_bits_channel),
    .io_tasks_source_d_bits_opcode(abc_mshr_3_io_tasks_source_d_bits_opcode),
    .io_tasks_source_d_bits_param(abc_mshr_3_io_tasks_source_d_bits_param),
    .io_tasks_source_d_bits_size(abc_mshr_3_io_tasks_source_d_bits_size),
    .io_tasks_source_d_bits_way(abc_mshr_3_io_tasks_source_d_bits_way),
    .io_tasks_source_d_bits_off(abc_mshr_3_io_tasks_source_d_bits_off),
    .io_tasks_source_d_bits_useBypass(abc_mshr_3_io_tasks_source_d_bits_useBypass),
    .io_tasks_source_d_bits_bufIdx(abc_mshr_3_io_tasks_source_d_bits_bufIdx),
    .io_tasks_source_d_bits_denied(abc_mshr_3_io_tasks_source_d_bits_denied),
    .io_tasks_source_d_bits_sinkId(abc_mshr_3_io_tasks_source_d_bits_sinkId),
    .io_tasks_source_d_bits_bypassPut(abc_mshr_3_io_tasks_source_d_bits_bypassPut),
    .io_tasks_source_d_bits_dirty(abc_mshr_3_io_tasks_source_d_bits_dirty),
    .io_tasks_source_a_ready(abc_mshr_3_io_tasks_source_a_ready),
    .io_tasks_source_a_valid(abc_mshr_3_io_tasks_source_a_valid),
    .io_tasks_source_a_bits_tag(abc_mshr_3_io_tasks_source_a_bits_tag),
    .io_tasks_source_a_bits_set(abc_mshr_3_io_tasks_source_a_bits_set),
    .io_tasks_source_a_bits_off(abc_mshr_3_io_tasks_source_a_bits_off),
    .io_tasks_source_a_bits_mask(abc_mshr_3_io_tasks_source_a_bits_mask),
    .io_tasks_source_a_bits_opcode(abc_mshr_3_io_tasks_source_a_bits_opcode),
    .io_tasks_source_a_bits_param(abc_mshr_3_io_tasks_source_a_bits_param),
    .io_tasks_source_a_bits_source(abc_mshr_3_io_tasks_source_a_bits_source),
    .io_tasks_source_a_bits_bufIdx(abc_mshr_3_io_tasks_source_a_bits_bufIdx),
    .io_tasks_source_a_bits_size(abc_mshr_3_io_tasks_source_a_bits_size),
    .io_tasks_source_a_bits_needData(abc_mshr_3_io_tasks_source_a_bits_needData),
    .io_tasks_source_a_bits_putData(abc_mshr_3_io_tasks_source_a_bits_putData),
    .io_tasks_source_c_ready(abc_mshr_3_io_tasks_source_c_ready),
    .io_tasks_source_c_valid(abc_mshr_3_io_tasks_source_c_valid),
    .io_tasks_source_c_bits_opcode(abc_mshr_3_io_tasks_source_c_bits_opcode),
    .io_tasks_source_c_bits_tag(abc_mshr_3_io_tasks_source_c_bits_tag),
    .io_tasks_source_c_bits_set(abc_mshr_3_io_tasks_source_c_bits_set),
    .io_tasks_source_c_bits_param(abc_mshr_3_io_tasks_source_c_bits_param),
    .io_tasks_source_c_bits_source(abc_mshr_3_io_tasks_source_c_bits_source),
    .io_tasks_source_c_bits_way(abc_mshr_3_io_tasks_source_c_bits_way),
    .io_tasks_source_c_bits_dirty(abc_mshr_3_io_tasks_source_c_bits_dirty),
    .io_tasks_source_e_ready(abc_mshr_3_io_tasks_source_e_ready),
    .io_tasks_source_e_valid(abc_mshr_3_io_tasks_source_e_valid),
    .io_tasks_source_e_bits_sink(abc_mshr_3_io_tasks_source_e_bits_sink),
    .io_tasks_dir_write_ready(abc_mshr_3_io_tasks_dir_write_ready),
    .io_tasks_dir_write_valid(abc_mshr_3_io_tasks_dir_write_valid),
    .io_tasks_dir_write_bits_set(abc_mshr_3_io_tasks_dir_write_bits_set),
    .io_tasks_dir_write_bits_way(abc_mshr_3_io_tasks_dir_write_bits_way),
    .io_tasks_dir_write_bits_data_dirty(abc_mshr_3_io_tasks_dir_write_bits_data_dirty),
    .io_tasks_dir_write_bits_data_state(abc_mshr_3_io_tasks_dir_write_bits_data_state),
    .io_tasks_dir_write_bits_data_clientStates_0(abc_mshr_3_io_tasks_dir_write_bits_data_clientStates_0),
    .io_tasks_dir_write_bits_data_clientStates_1(abc_mshr_3_io_tasks_dir_write_bits_data_clientStates_1),
    .io_tasks_tag_write_ready(abc_mshr_3_io_tasks_tag_write_ready),
    .io_tasks_tag_write_valid(abc_mshr_3_io_tasks_tag_write_valid),
    .io_tasks_tag_write_bits_set(abc_mshr_3_io_tasks_tag_write_bits_set),
    .io_tasks_tag_write_bits_way(abc_mshr_3_io_tasks_tag_write_bits_way),
    .io_tasks_tag_write_bits_tag(abc_mshr_3_io_tasks_tag_write_bits_tag),
    .io_tasks_client_dir_write_ready(abc_mshr_3_io_tasks_client_dir_write_ready),
    .io_tasks_client_dir_write_valid(abc_mshr_3_io_tasks_client_dir_write_valid),
    .io_tasks_client_dir_write_bits_set(abc_mshr_3_io_tasks_client_dir_write_bits_set),
    .io_tasks_client_dir_write_bits_way(abc_mshr_3_io_tasks_client_dir_write_bits_way),
    .io_tasks_client_dir_write_bits_data_0_state(abc_mshr_3_io_tasks_client_dir_write_bits_data_0_state),
    .io_tasks_client_dir_write_bits_data_1_state(abc_mshr_3_io_tasks_client_dir_write_bits_data_1_state),
    .io_tasks_client_tag_write_ready(abc_mshr_3_io_tasks_client_tag_write_ready),
    .io_tasks_client_tag_write_valid(abc_mshr_3_io_tasks_client_tag_write_valid),
    .io_tasks_client_tag_write_bits_set(abc_mshr_3_io_tasks_client_tag_write_bits_set),
    .io_tasks_client_tag_write_bits_way(abc_mshr_3_io_tasks_client_tag_write_bits_way),
    .io_tasks_client_tag_write_bits_tag(abc_mshr_3_io_tasks_client_tag_write_bits_tag),
    .io_dirResult_valid(abc_mshr_3_io_dirResult_valid),
    .io_dirResult_bits_self_dirty(abc_mshr_3_io_dirResult_bits_self_dirty),
    .io_dirResult_bits_self_state(abc_mshr_3_io_dirResult_bits_self_state),
    .io_dirResult_bits_self_clientStates_0(abc_mshr_3_io_dirResult_bits_self_clientStates_0),
    .io_dirResult_bits_self_clientStates_1(abc_mshr_3_io_dirResult_bits_self_clientStates_1),
    .io_dirResult_bits_self_hit(abc_mshr_3_io_dirResult_bits_self_hit),
    .io_dirResult_bits_self_way(abc_mshr_3_io_dirResult_bits_self_way),
    .io_dirResult_bits_self_tag(abc_mshr_3_io_dirResult_bits_self_tag),
    .io_dirResult_bits_clients_states_0_state(abc_mshr_3_io_dirResult_bits_clients_states_0_state),
    .io_dirResult_bits_clients_states_0_hit(abc_mshr_3_io_dirResult_bits_clients_states_0_hit),
    .io_dirResult_bits_clients_states_1_state(abc_mshr_3_io_dirResult_bits_clients_states_1_state),
    .io_dirResult_bits_clients_states_1_hit(abc_mshr_3_io_dirResult_bits_clients_states_1_hit),
    .io_dirResult_bits_clients_tag(abc_mshr_3_io_dirResult_bits_clients_tag),
    .io_dirResult_bits_clients_way(abc_mshr_3_io_dirResult_bits_clients_way),
    .io_c_status_set(abc_mshr_3_io_c_status_set),
    .io_c_status_tag(abc_mshr_3_io_c_status_tag),
    .io_c_status_way(abc_mshr_3_io_c_status_way),
    .io_c_status_nestedReleaseData(abc_mshr_3_io_c_status_nestedReleaseData),
    .io_c_status_releaseThrough(abc_mshr_3_io_c_status_releaseThrough),
    .io_bstatus_set(abc_mshr_3_io_bstatus_set),
    .io_bstatus_tag(abc_mshr_3_io_bstatus_tag),
    .io_bstatus_way(abc_mshr_3_io_bstatus_way),
    .io_bstatus_nestedProbeAckData(abc_mshr_3_io_bstatus_nestedProbeAckData),
    .io_bstatus_probeHelperFinish(abc_mshr_3_io_bstatus_probeHelperFinish),
    .io_bstatus_probeAckDataThrough(abc_mshr_3_io_bstatus_probeAckDataThrough),
    .io_releaseThrough(abc_mshr_3_io_releaseThrough),
    .io_probeAckDataThrough(abc_mshr_3_io_probeAckDataThrough),
    .io_is_nestedReleaseData(abc_mshr_3_io_is_nestedReleaseData),
    .io_is_nestedProbeAckData(abc_mshr_3_io_is_nestedProbeAckData),
    .io_probeHelperFinish(abc_mshr_3_io_probeHelperFinish)
  );
  MSHR abc_mshr_4 ( // @[Slice.scala 94:16]
    .clock(abc_mshr_4_clock),
    .reset(abc_mshr_4_reset),
    .io_id(abc_mshr_4_io_id),
    .io_enable(abc_mshr_4_io_enable),
    .io_alloc_valid(abc_mshr_4_io_alloc_valid),
    .io_alloc_bits_channel(abc_mshr_4_io_alloc_bits_channel),
    .io_alloc_bits_opcode(abc_mshr_4_io_alloc_bits_opcode),
    .io_alloc_bits_param(abc_mshr_4_io_alloc_bits_param),
    .io_alloc_bits_size(abc_mshr_4_io_alloc_bits_size),
    .io_alloc_bits_source(abc_mshr_4_io_alloc_bits_source),
    .io_alloc_bits_set(abc_mshr_4_io_alloc_bits_set),
    .io_alloc_bits_tag(abc_mshr_4_io_alloc_bits_tag),
    .io_alloc_bits_off(abc_mshr_4_io_alloc_bits_off),
    .io_alloc_bits_mask(abc_mshr_4_io_alloc_bits_mask),
    .io_alloc_bits_bufIdx(abc_mshr_4_io_alloc_bits_bufIdx),
    .io_alloc_bits_preferCache(abc_mshr_4_io_alloc_bits_preferCache),
    .io_alloc_bits_dirty(abc_mshr_4_io_alloc_bits_dirty),
    .io_alloc_bits_fromProbeHelper(abc_mshr_4_io_alloc_bits_fromProbeHelper),
    .io_alloc_bits_fromCmoHelper(abc_mshr_4_io_alloc_bits_fromCmoHelper),
    .io_alloc_bits_needProbeAckData(abc_mshr_4_io_alloc_bits_needProbeAckData),
    .io_status_valid(abc_mshr_4_io_status_valid),
    .io_status_bits_set(abc_mshr_4_io_status_bits_set),
    .io_status_bits_tag(abc_mshr_4_io_status_bits_tag),
    .io_status_bits_way(abc_mshr_4_io_status_bits_way),
    .io_status_bits_way_reg(abc_mshr_4_io_status_bits_way_reg),
    .io_status_bits_nestB(abc_mshr_4_io_status_bits_nestB),
    .io_status_bits_nestC(abc_mshr_4_io_status_bits_nestC),
    .io_status_bits_will_grant_data(abc_mshr_4_io_status_bits_will_grant_data),
    .io_status_bits_will_save_data(abc_mshr_4_io_status_bits_will_save_data),
    .io_status_bits_will_free(abc_mshr_4_io_status_bits_will_free),
    .io_resps_sink_c_valid(abc_mshr_4_io_resps_sink_c_valid),
    .io_resps_sink_c_bits_hasData(abc_mshr_4_io_resps_sink_c_bits_hasData),
    .io_resps_sink_c_bits_param(abc_mshr_4_io_resps_sink_c_bits_param),
    .io_resps_sink_c_bits_source(abc_mshr_4_io_resps_sink_c_bits_source),
    .io_resps_sink_c_bits_last(abc_mshr_4_io_resps_sink_c_bits_last),
    .io_resps_sink_c_bits_bufIdx(abc_mshr_4_io_resps_sink_c_bits_bufIdx),
    .io_resps_sink_d_valid(abc_mshr_4_io_resps_sink_d_valid),
    .io_resps_sink_d_bits_opcode(abc_mshr_4_io_resps_sink_d_bits_opcode),
    .io_resps_sink_d_bits_param(abc_mshr_4_io_resps_sink_d_bits_param),
    .io_resps_sink_d_bits_sink(abc_mshr_4_io_resps_sink_d_bits_sink),
    .io_resps_sink_d_bits_last(abc_mshr_4_io_resps_sink_d_bits_last),
    .io_resps_sink_d_bits_denied(abc_mshr_4_io_resps_sink_d_bits_denied),
    .io_resps_sink_d_bits_bufIdx(abc_mshr_4_io_resps_sink_d_bits_bufIdx),
    .io_resps_sink_e_valid(abc_mshr_4_io_resps_sink_e_valid),
    .io_resps_source_d_valid(abc_mshr_4_io_resps_source_d_valid),
    .io_nestedwb_set(abc_mshr_4_io_nestedwb_set),
    .io_nestedwb_tag(abc_mshr_4_io_nestedwb_tag),
    .io_nestedwb_btoN(abc_mshr_4_io_nestedwb_btoN),
    .io_nestedwb_btoB(abc_mshr_4_io_nestedwb_btoB),
    .io_nestedwb_bclr_dirty(abc_mshr_4_io_nestedwb_bclr_dirty),
    .io_nestedwb_bset_dirty(abc_mshr_4_io_nestedwb_bset_dirty),
    .io_nestedwb_c_set_dirty(abc_mshr_4_io_nestedwb_c_set_dirty),
    .io_nestedwb_c_set_hit(abc_mshr_4_io_nestedwb_c_set_hit),
    .io_nestedwb_clients_0_isToN(abc_mshr_4_io_nestedwb_clients_0_isToN),
    .io_nestedwb_clients_1_isToN(abc_mshr_4_io_nestedwb_clients_1_isToN),
    .io_tasks_sink_a_ready(abc_mshr_4_io_tasks_sink_a_ready),
    .io_tasks_sink_a_valid(abc_mshr_4_io_tasks_sink_a_valid),
    .io_tasks_sink_a_bits_sourceId(abc_mshr_4_io_tasks_sink_a_bits_sourceId),
    .io_tasks_sink_a_bits_set(abc_mshr_4_io_tasks_sink_a_bits_set),
    .io_tasks_sink_a_bits_tag(abc_mshr_4_io_tasks_sink_a_bits_tag),
    .io_tasks_sink_a_bits_size(abc_mshr_4_io_tasks_sink_a_bits_size),
    .io_tasks_sink_a_bits_off(abc_mshr_4_io_tasks_sink_a_bits_off),
    .io_tasks_source_bready(abc_mshr_4_io_tasks_source_bready),
    .io_tasks_source_bvalid(abc_mshr_4_io_tasks_source_bvalid),
    .io_tasks_source_bset(abc_mshr_4_io_tasks_source_bset),
    .io_tasks_source_btag(abc_mshr_4_io_tasks_source_btag),
    .io_tasks_source_bparam(abc_mshr_4_io_tasks_source_bparam),
    .io_tasks_source_bclients(abc_mshr_4_io_tasks_source_bclients),
    .io_tasks_source_bneedData(abc_mshr_4_io_tasks_source_bneedData),
    .io_tasks_sink_c_ready(abc_mshr_4_io_tasks_sink_c_ready),
    .io_tasks_sink_c_valid(abc_mshr_4_io_tasks_sink_c_valid),
    .io_tasks_sink_c_bits_sourceId(abc_mshr_4_io_tasks_sink_c_bits_sourceId),
    .io_tasks_sink_c_bits_set(abc_mshr_4_io_tasks_sink_c_bits_set),
    .io_tasks_sink_c_bits_tag(abc_mshr_4_io_tasks_sink_c_bits_tag),
    .io_tasks_sink_c_bits_size(abc_mshr_4_io_tasks_sink_c_bits_size),
    .io_tasks_sink_c_bits_way(abc_mshr_4_io_tasks_sink_c_bits_way),
    .io_tasks_sink_c_bits_off(abc_mshr_4_io_tasks_sink_c_bits_off),
    .io_tasks_sink_c_bits_bufIdx(abc_mshr_4_io_tasks_sink_c_bits_bufIdx),
    .io_tasks_sink_c_bits_opcode(abc_mshr_4_io_tasks_sink_c_bits_opcode),
    .io_tasks_sink_c_bits_param(abc_mshr_4_io_tasks_sink_c_bits_param),
    .io_tasks_sink_c_bits_source(abc_mshr_4_io_tasks_sink_c_bits_source),
    .io_tasks_sink_c_bits_save(abc_mshr_4_io_tasks_sink_c_bits_save),
    .io_tasks_sink_c_bits_drop(abc_mshr_4_io_tasks_sink_c_bits_drop),
    .io_tasks_sink_c_bits_release(abc_mshr_4_io_tasks_sink_c_bits_release),
    .io_tasks_sink_c_bits_dirty(abc_mshr_4_io_tasks_sink_c_bits_dirty),
    .io_tasks_source_d_ready(abc_mshr_4_io_tasks_source_d_ready),
    .io_tasks_source_d_valid(abc_mshr_4_io_tasks_source_d_valid),
    .io_tasks_source_d_bits_sourceId(abc_mshr_4_io_tasks_source_d_bits_sourceId),
    .io_tasks_source_d_bits_set(abc_mshr_4_io_tasks_source_d_bits_set),
    .io_tasks_source_d_bits_tag(abc_mshr_4_io_tasks_source_d_bits_tag),
    .io_tasks_source_d_bits_channel(abc_mshr_4_io_tasks_source_d_bits_channel),
    .io_tasks_source_d_bits_opcode(abc_mshr_4_io_tasks_source_d_bits_opcode),
    .io_tasks_source_d_bits_param(abc_mshr_4_io_tasks_source_d_bits_param),
    .io_tasks_source_d_bits_size(abc_mshr_4_io_tasks_source_d_bits_size),
    .io_tasks_source_d_bits_way(abc_mshr_4_io_tasks_source_d_bits_way),
    .io_tasks_source_d_bits_off(abc_mshr_4_io_tasks_source_d_bits_off),
    .io_tasks_source_d_bits_useBypass(abc_mshr_4_io_tasks_source_d_bits_useBypass),
    .io_tasks_source_d_bits_bufIdx(abc_mshr_4_io_tasks_source_d_bits_bufIdx),
    .io_tasks_source_d_bits_denied(abc_mshr_4_io_tasks_source_d_bits_denied),
    .io_tasks_source_d_bits_sinkId(abc_mshr_4_io_tasks_source_d_bits_sinkId),
    .io_tasks_source_d_bits_bypassPut(abc_mshr_4_io_tasks_source_d_bits_bypassPut),
    .io_tasks_source_d_bits_dirty(abc_mshr_4_io_tasks_source_d_bits_dirty),
    .io_tasks_source_a_ready(abc_mshr_4_io_tasks_source_a_ready),
    .io_tasks_source_a_valid(abc_mshr_4_io_tasks_source_a_valid),
    .io_tasks_source_a_bits_tag(abc_mshr_4_io_tasks_source_a_bits_tag),
    .io_tasks_source_a_bits_set(abc_mshr_4_io_tasks_source_a_bits_set),
    .io_tasks_source_a_bits_off(abc_mshr_4_io_tasks_source_a_bits_off),
    .io_tasks_source_a_bits_mask(abc_mshr_4_io_tasks_source_a_bits_mask),
    .io_tasks_source_a_bits_opcode(abc_mshr_4_io_tasks_source_a_bits_opcode),
    .io_tasks_source_a_bits_param(abc_mshr_4_io_tasks_source_a_bits_param),
    .io_tasks_source_a_bits_source(abc_mshr_4_io_tasks_source_a_bits_source),
    .io_tasks_source_a_bits_bufIdx(abc_mshr_4_io_tasks_source_a_bits_bufIdx),
    .io_tasks_source_a_bits_size(abc_mshr_4_io_tasks_source_a_bits_size),
    .io_tasks_source_a_bits_needData(abc_mshr_4_io_tasks_source_a_bits_needData),
    .io_tasks_source_a_bits_putData(abc_mshr_4_io_tasks_source_a_bits_putData),
    .io_tasks_source_c_ready(abc_mshr_4_io_tasks_source_c_ready),
    .io_tasks_source_c_valid(abc_mshr_4_io_tasks_source_c_valid),
    .io_tasks_source_c_bits_opcode(abc_mshr_4_io_tasks_source_c_bits_opcode),
    .io_tasks_source_c_bits_tag(abc_mshr_4_io_tasks_source_c_bits_tag),
    .io_tasks_source_c_bits_set(abc_mshr_4_io_tasks_source_c_bits_set),
    .io_tasks_source_c_bits_param(abc_mshr_4_io_tasks_source_c_bits_param),
    .io_tasks_source_c_bits_source(abc_mshr_4_io_tasks_source_c_bits_source),
    .io_tasks_source_c_bits_way(abc_mshr_4_io_tasks_source_c_bits_way),
    .io_tasks_source_c_bits_dirty(abc_mshr_4_io_tasks_source_c_bits_dirty),
    .io_tasks_source_e_ready(abc_mshr_4_io_tasks_source_e_ready),
    .io_tasks_source_e_valid(abc_mshr_4_io_tasks_source_e_valid),
    .io_tasks_source_e_bits_sink(abc_mshr_4_io_tasks_source_e_bits_sink),
    .io_tasks_dir_write_ready(abc_mshr_4_io_tasks_dir_write_ready),
    .io_tasks_dir_write_valid(abc_mshr_4_io_tasks_dir_write_valid),
    .io_tasks_dir_write_bits_set(abc_mshr_4_io_tasks_dir_write_bits_set),
    .io_tasks_dir_write_bits_way(abc_mshr_4_io_tasks_dir_write_bits_way),
    .io_tasks_dir_write_bits_data_dirty(abc_mshr_4_io_tasks_dir_write_bits_data_dirty),
    .io_tasks_dir_write_bits_data_state(abc_mshr_4_io_tasks_dir_write_bits_data_state),
    .io_tasks_dir_write_bits_data_clientStates_0(abc_mshr_4_io_tasks_dir_write_bits_data_clientStates_0),
    .io_tasks_dir_write_bits_data_clientStates_1(abc_mshr_4_io_tasks_dir_write_bits_data_clientStates_1),
    .io_tasks_tag_write_ready(abc_mshr_4_io_tasks_tag_write_ready),
    .io_tasks_tag_write_valid(abc_mshr_4_io_tasks_tag_write_valid),
    .io_tasks_tag_write_bits_set(abc_mshr_4_io_tasks_tag_write_bits_set),
    .io_tasks_tag_write_bits_way(abc_mshr_4_io_tasks_tag_write_bits_way),
    .io_tasks_tag_write_bits_tag(abc_mshr_4_io_tasks_tag_write_bits_tag),
    .io_tasks_client_dir_write_ready(abc_mshr_4_io_tasks_client_dir_write_ready),
    .io_tasks_client_dir_write_valid(abc_mshr_4_io_tasks_client_dir_write_valid),
    .io_tasks_client_dir_write_bits_set(abc_mshr_4_io_tasks_client_dir_write_bits_set),
    .io_tasks_client_dir_write_bits_way(abc_mshr_4_io_tasks_client_dir_write_bits_way),
    .io_tasks_client_dir_write_bits_data_0_state(abc_mshr_4_io_tasks_client_dir_write_bits_data_0_state),
    .io_tasks_client_dir_write_bits_data_1_state(abc_mshr_4_io_tasks_client_dir_write_bits_data_1_state),
    .io_tasks_client_tag_write_ready(abc_mshr_4_io_tasks_client_tag_write_ready),
    .io_tasks_client_tag_write_valid(abc_mshr_4_io_tasks_client_tag_write_valid),
    .io_tasks_client_tag_write_bits_set(abc_mshr_4_io_tasks_client_tag_write_bits_set),
    .io_tasks_client_tag_write_bits_way(abc_mshr_4_io_tasks_client_tag_write_bits_way),
    .io_tasks_client_tag_write_bits_tag(abc_mshr_4_io_tasks_client_tag_write_bits_tag),
    .io_dirResult_valid(abc_mshr_4_io_dirResult_valid),
    .io_dirResult_bits_self_dirty(abc_mshr_4_io_dirResult_bits_self_dirty),
    .io_dirResult_bits_self_state(abc_mshr_4_io_dirResult_bits_self_state),
    .io_dirResult_bits_self_clientStates_0(abc_mshr_4_io_dirResult_bits_self_clientStates_0),
    .io_dirResult_bits_self_clientStates_1(abc_mshr_4_io_dirResult_bits_self_clientStates_1),
    .io_dirResult_bits_self_hit(abc_mshr_4_io_dirResult_bits_self_hit),
    .io_dirResult_bits_self_way(abc_mshr_4_io_dirResult_bits_self_way),
    .io_dirResult_bits_self_tag(abc_mshr_4_io_dirResult_bits_self_tag),
    .io_dirResult_bits_clients_states_0_state(abc_mshr_4_io_dirResult_bits_clients_states_0_state),
    .io_dirResult_bits_clients_states_0_hit(abc_mshr_4_io_dirResult_bits_clients_states_0_hit),
    .io_dirResult_bits_clients_states_1_state(abc_mshr_4_io_dirResult_bits_clients_states_1_state),
    .io_dirResult_bits_clients_states_1_hit(abc_mshr_4_io_dirResult_bits_clients_states_1_hit),
    .io_dirResult_bits_clients_tag(abc_mshr_4_io_dirResult_bits_clients_tag),
    .io_dirResult_bits_clients_way(abc_mshr_4_io_dirResult_bits_clients_way),
    .io_c_status_set(abc_mshr_4_io_c_status_set),
    .io_c_status_tag(abc_mshr_4_io_c_status_tag),
    .io_c_status_way(abc_mshr_4_io_c_status_way),
    .io_c_status_nestedReleaseData(abc_mshr_4_io_c_status_nestedReleaseData),
    .io_c_status_releaseThrough(abc_mshr_4_io_c_status_releaseThrough),
    .io_bstatus_set(abc_mshr_4_io_bstatus_set),
    .io_bstatus_tag(abc_mshr_4_io_bstatus_tag),
    .io_bstatus_way(abc_mshr_4_io_bstatus_way),
    .io_bstatus_nestedProbeAckData(abc_mshr_4_io_bstatus_nestedProbeAckData),
    .io_bstatus_probeHelperFinish(abc_mshr_4_io_bstatus_probeHelperFinish),
    .io_bstatus_probeAckDataThrough(abc_mshr_4_io_bstatus_probeAckDataThrough),
    .io_releaseThrough(abc_mshr_4_io_releaseThrough),
    .io_probeAckDataThrough(abc_mshr_4_io_probeAckDataThrough),
    .io_is_nestedReleaseData(abc_mshr_4_io_is_nestedReleaseData),
    .io_is_nestedProbeAckData(abc_mshr_4_io_is_nestedProbeAckData),
    .io_probeHelperFinish(abc_mshr_4_io_probeHelperFinish)
  );
  MSHR abc_mshr_5 ( // @[Slice.scala 94:16]
    .clock(abc_mshr_5_clock),
    .reset(abc_mshr_5_reset),
    .io_id(abc_mshr_5_io_id),
    .io_enable(abc_mshr_5_io_enable),
    .io_alloc_valid(abc_mshr_5_io_alloc_valid),
    .io_alloc_bits_channel(abc_mshr_5_io_alloc_bits_channel),
    .io_alloc_bits_opcode(abc_mshr_5_io_alloc_bits_opcode),
    .io_alloc_bits_param(abc_mshr_5_io_alloc_bits_param),
    .io_alloc_bits_size(abc_mshr_5_io_alloc_bits_size),
    .io_alloc_bits_source(abc_mshr_5_io_alloc_bits_source),
    .io_alloc_bits_set(abc_mshr_5_io_alloc_bits_set),
    .io_alloc_bits_tag(abc_mshr_5_io_alloc_bits_tag),
    .io_alloc_bits_off(abc_mshr_5_io_alloc_bits_off),
    .io_alloc_bits_mask(abc_mshr_5_io_alloc_bits_mask),
    .io_alloc_bits_bufIdx(abc_mshr_5_io_alloc_bits_bufIdx),
    .io_alloc_bits_preferCache(abc_mshr_5_io_alloc_bits_preferCache),
    .io_alloc_bits_dirty(abc_mshr_5_io_alloc_bits_dirty),
    .io_alloc_bits_fromProbeHelper(abc_mshr_5_io_alloc_bits_fromProbeHelper),
    .io_alloc_bits_fromCmoHelper(abc_mshr_5_io_alloc_bits_fromCmoHelper),
    .io_alloc_bits_needProbeAckData(abc_mshr_5_io_alloc_bits_needProbeAckData),
    .io_status_valid(abc_mshr_5_io_status_valid),
    .io_status_bits_set(abc_mshr_5_io_status_bits_set),
    .io_status_bits_tag(abc_mshr_5_io_status_bits_tag),
    .io_status_bits_way(abc_mshr_5_io_status_bits_way),
    .io_status_bits_way_reg(abc_mshr_5_io_status_bits_way_reg),
    .io_status_bits_nestB(abc_mshr_5_io_status_bits_nestB),
    .io_status_bits_nestC(abc_mshr_5_io_status_bits_nestC),
    .io_status_bits_will_grant_data(abc_mshr_5_io_status_bits_will_grant_data),
    .io_status_bits_will_save_data(abc_mshr_5_io_status_bits_will_save_data),
    .io_status_bits_will_free(abc_mshr_5_io_status_bits_will_free),
    .io_resps_sink_c_valid(abc_mshr_5_io_resps_sink_c_valid),
    .io_resps_sink_c_bits_hasData(abc_mshr_5_io_resps_sink_c_bits_hasData),
    .io_resps_sink_c_bits_param(abc_mshr_5_io_resps_sink_c_bits_param),
    .io_resps_sink_c_bits_source(abc_mshr_5_io_resps_sink_c_bits_source),
    .io_resps_sink_c_bits_last(abc_mshr_5_io_resps_sink_c_bits_last),
    .io_resps_sink_c_bits_bufIdx(abc_mshr_5_io_resps_sink_c_bits_bufIdx),
    .io_resps_sink_d_valid(abc_mshr_5_io_resps_sink_d_valid),
    .io_resps_sink_d_bits_opcode(abc_mshr_5_io_resps_sink_d_bits_opcode),
    .io_resps_sink_d_bits_param(abc_mshr_5_io_resps_sink_d_bits_param),
    .io_resps_sink_d_bits_sink(abc_mshr_5_io_resps_sink_d_bits_sink),
    .io_resps_sink_d_bits_last(abc_mshr_5_io_resps_sink_d_bits_last),
    .io_resps_sink_d_bits_denied(abc_mshr_5_io_resps_sink_d_bits_denied),
    .io_resps_sink_d_bits_bufIdx(abc_mshr_5_io_resps_sink_d_bits_bufIdx),
    .io_resps_sink_e_valid(abc_mshr_5_io_resps_sink_e_valid),
    .io_resps_source_d_valid(abc_mshr_5_io_resps_source_d_valid),
    .io_nestedwb_set(abc_mshr_5_io_nestedwb_set),
    .io_nestedwb_tag(abc_mshr_5_io_nestedwb_tag),
    .io_nestedwb_btoN(abc_mshr_5_io_nestedwb_btoN),
    .io_nestedwb_btoB(abc_mshr_5_io_nestedwb_btoB),
    .io_nestedwb_bclr_dirty(abc_mshr_5_io_nestedwb_bclr_dirty),
    .io_nestedwb_bset_dirty(abc_mshr_5_io_nestedwb_bset_dirty),
    .io_nestedwb_c_set_dirty(abc_mshr_5_io_nestedwb_c_set_dirty),
    .io_nestedwb_c_set_hit(abc_mshr_5_io_nestedwb_c_set_hit),
    .io_nestedwb_clients_0_isToN(abc_mshr_5_io_nestedwb_clients_0_isToN),
    .io_nestedwb_clients_1_isToN(abc_mshr_5_io_nestedwb_clients_1_isToN),
    .io_tasks_sink_a_ready(abc_mshr_5_io_tasks_sink_a_ready),
    .io_tasks_sink_a_valid(abc_mshr_5_io_tasks_sink_a_valid),
    .io_tasks_sink_a_bits_sourceId(abc_mshr_5_io_tasks_sink_a_bits_sourceId),
    .io_tasks_sink_a_bits_set(abc_mshr_5_io_tasks_sink_a_bits_set),
    .io_tasks_sink_a_bits_tag(abc_mshr_5_io_tasks_sink_a_bits_tag),
    .io_tasks_sink_a_bits_size(abc_mshr_5_io_tasks_sink_a_bits_size),
    .io_tasks_sink_a_bits_off(abc_mshr_5_io_tasks_sink_a_bits_off),
    .io_tasks_source_bready(abc_mshr_5_io_tasks_source_bready),
    .io_tasks_source_bvalid(abc_mshr_5_io_tasks_source_bvalid),
    .io_tasks_source_bset(abc_mshr_5_io_tasks_source_bset),
    .io_tasks_source_btag(abc_mshr_5_io_tasks_source_btag),
    .io_tasks_source_bparam(abc_mshr_5_io_tasks_source_bparam),
    .io_tasks_source_bclients(abc_mshr_5_io_tasks_source_bclients),
    .io_tasks_source_bneedData(abc_mshr_5_io_tasks_source_bneedData),
    .io_tasks_sink_c_ready(abc_mshr_5_io_tasks_sink_c_ready),
    .io_tasks_sink_c_valid(abc_mshr_5_io_tasks_sink_c_valid),
    .io_tasks_sink_c_bits_sourceId(abc_mshr_5_io_tasks_sink_c_bits_sourceId),
    .io_tasks_sink_c_bits_set(abc_mshr_5_io_tasks_sink_c_bits_set),
    .io_tasks_sink_c_bits_tag(abc_mshr_5_io_tasks_sink_c_bits_tag),
    .io_tasks_sink_c_bits_size(abc_mshr_5_io_tasks_sink_c_bits_size),
    .io_tasks_sink_c_bits_way(abc_mshr_5_io_tasks_sink_c_bits_way),
    .io_tasks_sink_c_bits_off(abc_mshr_5_io_tasks_sink_c_bits_off),
    .io_tasks_sink_c_bits_bufIdx(abc_mshr_5_io_tasks_sink_c_bits_bufIdx),
    .io_tasks_sink_c_bits_opcode(abc_mshr_5_io_tasks_sink_c_bits_opcode),
    .io_tasks_sink_c_bits_param(abc_mshr_5_io_tasks_sink_c_bits_param),
    .io_tasks_sink_c_bits_source(abc_mshr_5_io_tasks_sink_c_bits_source),
    .io_tasks_sink_c_bits_save(abc_mshr_5_io_tasks_sink_c_bits_save),
    .io_tasks_sink_c_bits_drop(abc_mshr_5_io_tasks_sink_c_bits_drop),
    .io_tasks_sink_c_bits_release(abc_mshr_5_io_tasks_sink_c_bits_release),
    .io_tasks_sink_c_bits_dirty(abc_mshr_5_io_tasks_sink_c_bits_dirty),
    .io_tasks_source_d_ready(abc_mshr_5_io_tasks_source_d_ready),
    .io_tasks_source_d_valid(abc_mshr_5_io_tasks_source_d_valid),
    .io_tasks_source_d_bits_sourceId(abc_mshr_5_io_tasks_source_d_bits_sourceId),
    .io_tasks_source_d_bits_set(abc_mshr_5_io_tasks_source_d_bits_set),
    .io_tasks_source_d_bits_tag(abc_mshr_5_io_tasks_source_d_bits_tag),
    .io_tasks_source_d_bits_channel(abc_mshr_5_io_tasks_source_d_bits_channel),
    .io_tasks_source_d_bits_opcode(abc_mshr_5_io_tasks_source_d_bits_opcode),
    .io_tasks_source_d_bits_param(abc_mshr_5_io_tasks_source_d_bits_param),
    .io_tasks_source_d_bits_size(abc_mshr_5_io_tasks_source_d_bits_size),
    .io_tasks_source_d_bits_way(abc_mshr_5_io_tasks_source_d_bits_way),
    .io_tasks_source_d_bits_off(abc_mshr_5_io_tasks_source_d_bits_off),
    .io_tasks_source_d_bits_useBypass(abc_mshr_5_io_tasks_source_d_bits_useBypass),
    .io_tasks_source_d_bits_bufIdx(abc_mshr_5_io_tasks_source_d_bits_bufIdx),
    .io_tasks_source_d_bits_denied(abc_mshr_5_io_tasks_source_d_bits_denied),
    .io_tasks_source_d_bits_sinkId(abc_mshr_5_io_tasks_source_d_bits_sinkId),
    .io_tasks_source_d_bits_bypassPut(abc_mshr_5_io_tasks_source_d_bits_bypassPut),
    .io_tasks_source_d_bits_dirty(abc_mshr_5_io_tasks_source_d_bits_dirty),
    .io_tasks_source_a_ready(abc_mshr_5_io_tasks_source_a_ready),
    .io_tasks_source_a_valid(abc_mshr_5_io_tasks_source_a_valid),
    .io_tasks_source_a_bits_tag(abc_mshr_5_io_tasks_source_a_bits_tag),
    .io_tasks_source_a_bits_set(abc_mshr_5_io_tasks_source_a_bits_set),
    .io_tasks_source_a_bits_off(abc_mshr_5_io_tasks_source_a_bits_off),
    .io_tasks_source_a_bits_mask(abc_mshr_5_io_tasks_source_a_bits_mask),
    .io_tasks_source_a_bits_opcode(abc_mshr_5_io_tasks_source_a_bits_opcode),
    .io_tasks_source_a_bits_param(abc_mshr_5_io_tasks_source_a_bits_param),
    .io_tasks_source_a_bits_source(abc_mshr_5_io_tasks_source_a_bits_source),
    .io_tasks_source_a_bits_bufIdx(abc_mshr_5_io_tasks_source_a_bits_bufIdx),
    .io_tasks_source_a_bits_size(abc_mshr_5_io_tasks_source_a_bits_size),
    .io_tasks_source_a_bits_needData(abc_mshr_5_io_tasks_source_a_bits_needData),
    .io_tasks_source_a_bits_putData(abc_mshr_5_io_tasks_source_a_bits_putData),
    .io_tasks_source_c_ready(abc_mshr_5_io_tasks_source_c_ready),
    .io_tasks_source_c_valid(abc_mshr_5_io_tasks_source_c_valid),
    .io_tasks_source_c_bits_opcode(abc_mshr_5_io_tasks_source_c_bits_opcode),
    .io_tasks_source_c_bits_tag(abc_mshr_5_io_tasks_source_c_bits_tag),
    .io_tasks_source_c_bits_set(abc_mshr_5_io_tasks_source_c_bits_set),
    .io_tasks_source_c_bits_param(abc_mshr_5_io_tasks_source_c_bits_param),
    .io_tasks_source_c_bits_source(abc_mshr_5_io_tasks_source_c_bits_source),
    .io_tasks_source_c_bits_way(abc_mshr_5_io_tasks_source_c_bits_way),
    .io_tasks_source_c_bits_dirty(abc_mshr_5_io_tasks_source_c_bits_dirty),
    .io_tasks_source_e_ready(abc_mshr_5_io_tasks_source_e_ready),
    .io_tasks_source_e_valid(abc_mshr_5_io_tasks_source_e_valid),
    .io_tasks_source_e_bits_sink(abc_mshr_5_io_tasks_source_e_bits_sink),
    .io_tasks_dir_write_ready(abc_mshr_5_io_tasks_dir_write_ready),
    .io_tasks_dir_write_valid(abc_mshr_5_io_tasks_dir_write_valid),
    .io_tasks_dir_write_bits_set(abc_mshr_5_io_tasks_dir_write_bits_set),
    .io_tasks_dir_write_bits_way(abc_mshr_5_io_tasks_dir_write_bits_way),
    .io_tasks_dir_write_bits_data_dirty(abc_mshr_5_io_tasks_dir_write_bits_data_dirty),
    .io_tasks_dir_write_bits_data_state(abc_mshr_5_io_tasks_dir_write_bits_data_state),
    .io_tasks_dir_write_bits_data_clientStates_0(abc_mshr_5_io_tasks_dir_write_bits_data_clientStates_0),
    .io_tasks_dir_write_bits_data_clientStates_1(abc_mshr_5_io_tasks_dir_write_bits_data_clientStates_1),
    .io_tasks_tag_write_ready(abc_mshr_5_io_tasks_tag_write_ready),
    .io_tasks_tag_write_valid(abc_mshr_5_io_tasks_tag_write_valid),
    .io_tasks_tag_write_bits_set(abc_mshr_5_io_tasks_tag_write_bits_set),
    .io_tasks_tag_write_bits_way(abc_mshr_5_io_tasks_tag_write_bits_way),
    .io_tasks_tag_write_bits_tag(abc_mshr_5_io_tasks_tag_write_bits_tag),
    .io_tasks_client_dir_write_ready(abc_mshr_5_io_tasks_client_dir_write_ready),
    .io_tasks_client_dir_write_valid(abc_mshr_5_io_tasks_client_dir_write_valid),
    .io_tasks_client_dir_write_bits_set(abc_mshr_5_io_tasks_client_dir_write_bits_set),
    .io_tasks_client_dir_write_bits_way(abc_mshr_5_io_tasks_client_dir_write_bits_way),
    .io_tasks_client_dir_write_bits_data_0_state(abc_mshr_5_io_tasks_client_dir_write_bits_data_0_state),
    .io_tasks_client_dir_write_bits_data_1_state(abc_mshr_5_io_tasks_client_dir_write_bits_data_1_state),
    .io_tasks_client_tag_write_ready(abc_mshr_5_io_tasks_client_tag_write_ready),
    .io_tasks_client_tag_write_valid(abc_mshr_5_io_tasks_client_tag_write_valid),
    .io_tasks_client_tag_write_bits_set(abc_mshr_5_io_tasks_client_tag_write_bits_set),
    .io_tasks_client_tag_write_bits_way(abc_mshr_5_io_tasks_client_tag_write_bits_way),
    .io_tasks_client_tag_write_bits_tag(abc_mshr_5_io_tasks_client_tag_write_bits_tag),
    .io_dirResult_valid(abc_mshr_5_io_dirResult_valid),
    .io_dirResult_bits_self_dirty(abc_mshr_5_io_dirResult_bits_self_dirty),
    .io_dirResult_bits_self_state(abc_mshr_5_io_dirResult_bits_self_state),
    .io_dirResult_bits_self_clientStates_0(abc_mshr_5_io_dirResult_bits_self_clientStates_0),
    .io_dirResult_bits_self_clientStates_1(abc_mshr_5_io_dirResult_bits_self_clientStates_1),
    .io_dirResult_bits_self_hit(abc_mshr_5_io_dirResult_bits_self_hit),
    .io_dirResult_bits_self_way(abc_mshr_5_io_dirResult_bits_self_way),
    .io_dirResult_bits_self_tag(abc_mshr_5_io_dirResult_bits_self_tag),
    .io_dirResult_bits_clients_states_0_state(abc_mshr_5_io_dirResult_bits_clients_states_0_state),
    .io_dirResult_bits_clients_states_0_hit(abc_mshr_5_io_dirResult_bits_clients_states_0_hit),
    .io_dirResult_bits_clients_states_1_state(abc_mshr_5_io_dirResult_bits_clients_states_1_state),
    .io_dirResult_bits_clients_states_1_hit(abc_mshr_5_io_dirResult_bits_clients_states_1_hit),
    .io_dirResult_bits_clients_tag(abc_mshr_5_io_dirResult_bits_clients_tag),
    .io_dirResult_bits_clients_way(abc_mshr_5_io_dirResult_bits_clients_way),
    .io_c_status_set(abc_mshr_5_io_c_status_set),
    .io_c_status_tag(abc_mshr_5_io_c_status_tag),
    .io_c_status_way(abc_mshr_5_io_c_status_way),
    .io_c_status_nestedReleaseData(abc_mshr_5_io_c_status_nestedReleaseData),
    .io_c_status_releaseThrough(abc_mshr_5_io_c_status_releaseThrough),
    .io_bstatus_set(abc_mshr_5_io_bstatus_set),
    .io_bstatus_tag(abc_mshr_5_io_bstatus_tag),
    .io_bstatus_way(abc_mshr_5_io_bstatus_way),
    .io_bstatus_nestedProbeAckData(abc_mshr_5_io_bstatus_nestedProbeAckData),
    .io_bstatus_probeHelperFinish(abc_mshr_5_io_bstatus_probeHelperFinish),
    .io_bstatus_probeAckDataThrough(abc_mshr_5_io_bstatus_probeAckDataThrough),
    .io_releaseThrough(abc_mshr_5_io_releaseThrough),
    .io_probeAckDataThrough(abc_mshr_5_io_probeAckDataThrough),
    .io_is_nestedReleaseData(abc_mshr_5_io_is_nestedReleaseData),
    .io_is_nestedProbeAckData(abc_mshr_5_io_is_nestedProbeAckData),
    .io_probeHelperFinish(abc_mshr_5_io_probeHelperFinish)
  );
  MSHR abc_mshr_6 ( // @[Slice.scala 94:16]
    .clock(abc_mshr_6_clock),
    .reset(abc_mshr_6_reset),
    .io_id(abc_mshr_6_io_id),
    .io_enable(abc_mshr_6_io_enable),
    .io_alloc_valid(abc_mshr_6_io_alloc_valid),
    .io_alloc_bits_channel(abc_mshr_6_io_alloc_bits_channel),
    .io_alloc_bits_opcode(abc_mshr_6_io_alloc_bits_opcode),
    .io_alloc_bits_param(abc_mshr_6_io_alloc_bits_param),
    .io_alloc_bits_size(abc_mshr_6_io_alloc_bits_size),
    .io_alloc_bits_source(abc_mshr_6_io_alloc_bits_source),
    .io_alloc_bits_set(abc_mshr_6_io_alloc_bits_set),
    .io_alloc_bits_tag(abc_mshr_6_io_alloc_bits_tag),
    .io_alloc_bits_off(abc_mshr_6_io_alloc_bits_off),
    .io_alloc_bits_mask(abc_mshr_6_io_alloc_bits_mask),
    .io_alloc_bits_bufIdx(abc_mshr_6_io_alloc_bits_bufIdx),
    .io_alloc_bits_preferCache(abc_mshr_6_io_alloc_bits_preferCache),
    .io_alloc_bits_dirty(abc_mshr_6_io_alloc_bits_dirty),
    .io_alloc_bits_fromProbeHelper(abc_mshr_6_io_alloc_bits_fromProbeHelper),
    .io_alloc_bits_fromCmoHelper(abc_mshr_6_io_alloc_bits_fromCmoHelper),
    .io_alloc_bits_needProbeAckData(abc_mshr_6_io_alloc_bits_needProbeAckData),
    .io_status_valid(abc_mshr_6_io_status_valid),
    .io_status_bits_set(abc_mshr_6_io_status_bits_set),
    .io_status_bits_tag(abc_mshr_6_io_status_bits_tag),
    .io_status_bits_way(abc_mshr_6_io_status_bits_way),
    .io_status_bits_way_reg(abc_mshr_6_io_status_bits_way_reg),
    .io_status_bits_nestB(abc_mshr_6_io_status_bits_nestB),
    .io_status_bits_nestC(abc_mshr_6_io_status_bits_nestC),
    .io_status_bits_will_grant_data(abc_mshr_6_io_status_bits_will_grant_data),
    .io_status_bits_will_save_data(abc_mshr_6_io_status_bits_will_save_data),
    .io_status_bits_will_free(abc_mshr_6_io_status_bits_will_free),
    .io_resps_sink_c_valid(abc_mshr_6_io_resps_sink_c_valid),
    .io_resps_sink_c_bits_hasData(abc_mshr_6_io_resps_sink_c_bits_hasData),
    .io_resps_sink_c_bits_param(abc_mshr_6_io_resps_sink_c_bits_param),
    .io_resps_sink_c_bits_source(abc_mshr_6_io_resps_sink_c_bits_source),
    .io_resps_sink_c_bits_last(abc_mshr_6_io_resps_sink_c_bits_last),
    .io_resps_sink_c_bits_bufIdx(abc_mshr_6_io_resps_sink_c_bits_bufIdx),
    .io_resps_sink_d_valid(abc_mshr_6_io_resps_sink_d_valid),
    .io_resps_sink_d_bits_opcode(abc_mshr_6_io_resps_sink_d_bits_opcode),
    .io_resps_sink_d_bits_param(abc_mshr_6_io_resps_sink_d_bits_param),
    .io_resps_sink_d_bits_sink(abc_mshr_6_io_resps_sink_d_bits_sink),
    .io_resps_sink_d_bits_last(abc_mshr_6_io_resps_sink_d_bits_last),
    .io_resps_sink_d_bits_denied(abc_mshr_6_io_resps_sink_d_bits_denied),
    .io_resps_sink_d_bits_bufIdx(abc_mshr_6_io_resps_sink_d_bits_bufIdx),
    .io_resps_sink_e_valid(abc_mshr_6_io_resps_sink_e_valid),
    .io_resps_source_d_valid(abc_mshr_6_io_resps_source_d_valid),
    .io_nestedwb_set(abc_mshr_6_io_nestedwb_set),
    .io_nestedwb_tag(abc_mshr_6_io_nestedwb_tag),
    .io_nestedwb_btoN(abc_mshr_6_io_nestedwb_btoN),
    .io_nestedwb_btoB(abc_mshr_6_io_nestedwb_btoB),
    .io_nestedwb_bclr_dirty(abc_mshr_6_io_nestedwb_bclr_dirty),
    .io_nestedwb_bset_dirty(abc_mshr_6_io_nestedwb_bset_dirty),
    .io_nestedwb_c_set_dirty(abc_mshr_6_io_nestedwb_c_set_dirty),
    .io_nestedwb_c_set_hit(abc_mshr_6_io_nestedwb_c_set_hit),
    .io_nestedwb_clients_0_isToN(abc_mshr_6_io_nestedwb_clients_0_isToN),
    .io_nestedwb_clients_1_isToN(abc_mshr_6_io_nestedwb_clients_1_isToN),
    .io_tasks_sink_a_ready(abc_mshr_6_io_tasks_sink_a_ready),
    .io_tasks_sink_a_valid(abc_mshr_6_io_tasks_sink_a_valid),
    .io_tasks_sink_a_bits_sourceId(abc_mshr_6_io_tasks_sink_a_bits_sourceId),
    .io_tasks_sink_a_bits_set(abc_mshr_6_io_tasks_sink_a_bits_set),
    .io_tasks_sink_a_bits_tag(abc_mshr_6_io_tasks_sink_a_bits_tag),
    .io_tasks_sink_a_bits_size(abc_mshr_6_io_tasks_sink_a_bits_size),
    .io_tasks_sink_a_bits_off(abc_mshr_6_io_tasks_sink_a_bits_off),
    .io_tasks_source_bready(abc_mshr_6_io_tasks_source_bready),
    .io_tasks_source_bvalid(abc_mshr_6_io_tasks_source_bvalid),
    .io_tasks_source_bset(abc_mshr_6_io_tasks_source_bset),
    .io_tasks_source_btag(abc_mshr_6_io_tasks_source_btag),
    .io_tasks_source_bparam(abc_mshr_6_io_tasks_source_bparam),
    .io_tasks_source_bclients(abc_mshr_6_io_tasks_source_bclients),
    .io_tasks_source_bneedData(abc_mshr_6_io_tasks_source_bneedData),
    .io_tasks_sink_c_ready(abc_mshr_6_io_tasks_sink_c_ready),
    .io_tasks_sink_c_valid(abc_mshr_6_io_tasks_sink_c_valid),
    .io_tasks_sink_c_bits_sourceId(abc_mshr_6_io_tasks_sink_c_bits_sourceId),
    .io_tasks_sink_c_bits_set(abc_mshr_6_io_tasks_sink_c_bits_set),
    .io_tasks_sink_c_bits_tag(abc_mshr_6_io_tasks_sink_c_bits_tag),
    .io_tasks_sink_c_bits_size(abc_mshr_6_io_tasks_sink_c_bits_size),
    .io_tasks_sink_c_bits_way(abc_mshr_6_io_tasks_sink_c_bits_way),
    .io_tasks_sink_c_bits_off(abc_mshr_6_io_tasks_sink_c_bits_off),
    .io_tasks_sink_c_bits_bufIdx(abc_mshr_6_io_tasks_sink_c_bits_bufIdx),
    .io_tasks_sink_c_bits_opcode(abc_mshr_6_io_tasks_sink_c_bits_opcode),
    .io_tasks_sink_c_bits_param(abc_mshr_6_io_tasks_sink_c_bits_param),
    .io_tasks_sink_c_bits_source(abc_mshr_6_io_tasks_sink_c_bits_source),
    .io_tasks_sink_c_bits_save(abc_mshr_6_io_tasks_sink_c_bits_save),
    .io_tasks_sink_c_bits_drop(abc_mshr_6_io_tasks_sink_c_bits_drop),
    .io_tasks_sink_c_bits_release(abc_mshr_6_io_tasks_sink_c_bits_release),
    .io_tasks_sink_c_bits_dirty(abc_mshr_6_io_tasks_sink_c_bits_dirty),
    .io_tasks_source_d_ready(abc_mshr_6_io_tasks_source_d_ready),
    .io_tasks_source_d_valid(abc_mshr_6_io_tasks_source_d_valid),
    .io_tasks_source_d_bits_sourceId(abc_mshr_6_io_tasks_source_d_bits_sourceId),
    .io_tasks_source_d_bits_set(abc_mshr_6_io_tasks_source_d_bits_set),
    .io_tasks_source_d_bits_tag(abc_mshr_6_io_tasks_source_d_bits_tag),
    .io_tasks_source_d_bits_channel(abc_mshr_6_io_tasks_source_d_bits_channel),
    .io_tasks_source_d_bits_opcode(abc_mshr_6_io_tasks_source_d_bits_opcode),
    .io_tasks_source_d_bits_param(abc_mshr_6_io_tasks_source_d_bits_param),
    .io_tasks_source_d_bits_size(abc_mshr_6_io_tasks_source_d_bits_size),
    .io_tasks_source_d_bits_way(abc_mshr_6_io_tasks_source_d_bits_way),
    .io_tasks_source_d_bits_off(abc_mshr_6_io_tasks_source_d_bits_off),
    .io_tasks_source_d_bits_useBypass(abc_mshr_6_io_tasks_source_d_bits_useBypass),
    .io_tasks_source_d_bits_bufIdx(abc_mshr_6_io_tasks_source_d_bits_bufIdx),
    .io_tasks_source_d_bits_denied(abc_mshr_6_io_tasks_source_d_bits_denied),
    .io_tasks_source_d_bits_sinkId(abc_mshr_6_io_tasks_source_d_bits_sinkId),
    .io_tasks_source_d_bits_bypassPut(abc_mshr_6_io_tasks_source_d_bits_bypassPut),
    .io_tasks_source_d_bits_dirty(abc_mshr_6_io_tasks_source_d_bits_dirty),
    .io_tasks_source_a_ready(abc_mshr_6_io_tasks_source_a_ready),
    .io_tasks_source_a_valid(abc_mshr_6_io_tasks_source_a_valid),
    .io_tasks_source_a_bits_tag(abc_mshr_6_io_tasks_source_a_bits_tag),
    .io_tasks_source_a_bits_set(abc_mshr_6_io_tasks_source_a_bits_set),
    .io_tasks_source_a_bits_off(abc_mshr_6_io_tasks_source_a_bits_off),
    .io_tasks_source_a_bits_mask(abc_mshr_6_io_tasks_source_a_bits_mask),
    .io_tasks_source_a_bits_opcode(abc_mshr_6_io_tasks_source_a_bits_opcode),
    .io_tasks_source_a_bits_param(abc_mshr_6_io_tasks_source_a_bits_param),
    .io_tasks_source_a_bits_source(abc_mshr_6_io_tasks_source_a_bits_source),
    .io_tasks_source_a_bits_bufIdx(abc_mshr_6_io_tasks_source_a_bits_bufIdx),
    .io_tasks_source_a_bits_size(abc_mshr_6_io_tasks_source_a_bits_size),
    .io_tasks_source_a_bits_needData(abc_mshr_6_io_tasks_source_a_bits_needData),
    .io_tasks_source_a_bits_putData(abc_mshr_6_io_tasks_source_a_bits_putData),
    .io_tasks_source_c_ready(abc_mshr_6_io_tasks_source_c_ready),
    .io_tasks_source_c_valid(abc_mshr_6_io_tasks_source_c_valid),
    .io_tasks_source_c_bits_opcode(abc_mshr_6_io_tasks_source_c_bits_opcode),
    .io_tasks_source_c_bits_tag(abc_mshr_6_io_tasks_source_c_bits_tag),
    .io_tasks_source_c_bits_set(abc_mshr_6_io_tasks_source_c_bits_set),
    .io_tasks_source_c_bits_param(abc_mshr_6_io_tasks_source_c_bits_param),
    .io_tasks_source_c_bits_source(abc_mshr_6_io_tasks_source_c_bits_source),
    .io_tasks_source_c_bits_way(abc_mshr_6_io_tasks_source_c_bits_way),
    .io_tasks_source_c_bits_dirty(abc_mshr_6_io_tasks_source_c_bits_dirty),
    .io_tasks_source_e_ready(abc_mshr_6_io_tasks_source_e_ready),
    .io_tasks_source_e_valid(abc_mshr_6_io_tasks_source_e_valid),
    .io_tasks_source_e_bits_sink(abc_mshr_6_io_tasks_source_e_bits_sink),
    .io_tasks_dir_write_ready(abc_mshr_6_io_tasks_dir_write_ready),
    .io_tasks_dir_write_valid(abc_mshr_6_io_tasks_dir_write_valid),
    .io_tasks_dir_write_bits_set(abc_mshr_6_io_tasks_dir_write_bits_set),
    .io_tasks_dir_write_bits_way(abc_mshr_6_io_tasks_dir_write_bits_way),
    .io_tasks_dir_write_bits_data_dirty(abc_mshr_6_io_tasks_dir_write_bits_data_dirty),
    .io_tasks_dir_write_bits_data_state(abc_mshr_6_io_tasks_dir_write_bits_data_state),
    .io_tasks_dir_write_bits_data_clientStates_0(abc_mshr_6_io_tasks_dir_write_bits_data_clientStates_0),
    .io_tasks_dir_write_bits_data_clientStates_1(abc_mshr_6_io_tasks_dir_write_bits_data_clientStates_1),
    .io_tasks_tag_write_ready(abc_mshr_6_io_tasks_tag_write_ready),
    .io_tasks_tag_write_valid(abc_mshr_6_io_tasks_tag_write_valid),
    .io_tasks_tag_write_bits_set(abc_mshr_6_io_tasks_tag_write_bits_set),
    .io_tasks_tag_write_bits_way(abc_mshr_6_io_tasks_tag_write_bits_way),
    .io_tasks_tag_write_bits_tag(abc_mshr_6_io_tasks_tag_write_bits_tag),
    .io_tasks_client_dir_write_ready(abc_mshr_6_io_tasks_client_dir_write_ready),
    .io_tasks_client_dir_write_valid(abc_mshr_6_io_tasks_client_dir_write_valid),
    .io_tasks_client_dir_write_bits_set(abc_mshr_6_io_tasks_client_dir_write_bits_set),
    .io_tasks_client_dir_write_bits_way(abc_mshr_6_io_tasks_client_dir_write_bits_way),
    .io_tasks_client_dir_write_bits_data_0_state(abc_mshr_6_io_tasks_client_dir_write_bits_data_0_state),
    .io_tasks_client_dir_write_bits_data_1_state(abc_mshr_6_io_tasks_client_dir_write_bits_data_1_state),
    .io_tasks_client_tag_write_ready(abc_mshr_6_io_tasks_client_tag_write_ready),
    .io_tasks_client_tag_write_valid(abc_mshr_6_io_tasks_client_tag_write_valid),
    .io_tasks_client_tag_write_bits_set(abc_mshr_6_io_tasks_client_tag_write_bits_set),
    .io_tasks_client_tag_write_bits_way(abc_mshr_6_io_tasks_client_tag_write_bits_way),
    .io_tasks_client_tag_write_bits_tag(abc_mshr_6_io_tasks_client_tag_write_bits_tag),
    .io_dirResult_valid(abc_mshr_6_io_dirResult_valid),
    .io_dirResult_bits_self_dirty(abc_mshr_6_io_dirResult_bits_self_dirty),
    .io_dirResult_bits_self_state(abc_mshr_6_io_dirResult_bits_self_state),
    .io_dirResult_bits_self_clientStates_0(abc_mshr_6_io_dirResult_bits_self_clientStates_0),
    .io_dirResult_bits_self_clientStates_1(abc_mshr_6_io_dirResult_bits_self_clientStates_1),
    .io_dirResult_bits_self_hit(abc_mshr_6_io_dirResult_bits_self_hit),
    .io_dirResult_bits_self_way(abc_mshr_6_io_dirResult_bits_self_way),
    .io_dirResult_bits_self_tag(abc_mshr_6_io_dirResult_bits_self_tag),
    .io_dirResult_bits_clients_states_0_state(abc_mshr_6_io_dirResult_bits_clients_states_0_state),
    .io_dirResult_bits_clients_states_0_hit(abc_mshr_6_io_dirResult_bits_clients_states_0_hit),
    .io_dirResult_bits_clients_states_1_state(abc_mshr_6_io_dirResult_bits_clients_states_1_state),
    .io_dirResult_bits_clients_states_1_hit(abc_mshr_6_io_dirResult_bits_clients_states_1_hit),
    .io_dirResult_bits_clients_tag(abc_mshr_6_io_dirResult_bits_clients_tag),
    .io_dirResult_bits_clients_way(abc_mshr_6_io_dirResult_bits_clients_way),
    .io_c_status_set(abc_mshr_6_io_c_status_set),
    .io_c_status_tag(abc_mshr_6_io_c_status_tag),
    .io_c_status_way(abc_mshr_6_io_c_status_way),
    .io_c_status_nestedReleaseData(abc_mshr_6_io_c_status_nestedReleaseData),
    .io_c_status_releaseThrough(abc_mshr_6_io_c_status_releaseThrough),
    .io_bstatus_set(abc_mshr_6_io_bstatus_set),
    .io_bstatus_tag(abc_mshr_6_io_bstatus_tag),
    .io_bstatus_way(abc_mshr_6_io_bstatus_way),
    .io_bstatus_nestedProbeAckData(abc_mshr_6_io_bstatus_nestedProbeAckData),
    .io_bstatus_probeHelperFinish(abc_mshr_6_io_bstatus_probeHelperFinish),
    .io_bstatus_probeAckDataThrough(abc_mshr_6_io_bstatus_probeAckDataThrough),
    .io_releaseThrough(abc_mshr_6_io_releaseThrough),
    .io_probeAckDataThrough(abc_mshr_6_io_probeAckDataThrough),
    .io_is_nestedReleaseData(abc_mshr_6_io_is_nestedReleaseData),
    .io_is_nestedProbeAckData(abc_mshr_6_io_is_nestedProbeAckData),
    .io_probeHelperFinish(abc_mshr_6_io_probeHelperFinish)
  );
  MSHR abc_mshr_7 ( // @[Slice.scala 94:16]
    .clock(abc_mshr_7_clock),
    .reset(abc_mshr_7_reset),
    .io_id(abc_mshr_7_io_id),
    .io_enable(abc_mshr_7_io_enable),
    .io_alloc_valid(abc_mshr_7_io_alloc_valid),
    .io_alloc_bits_channel(abc_mshr_7_io_alloc_bits_channel),
    .io_alloc_bits_opcode(abc_mshr_7_io_alloc_bits_opcode),
    .io_alloc_bits_param(abc_mshr_7_io_alloc_bits_param),
    .io_alloc_bits_size(abc_mshr_7_io_alloc_bits_size),
    .io_alloc_bits_source(abc_mshr_7_io_alloc_bits_source),
    .io_alloc_bits_set(abc_mshr_7_io_alloc_bits_set),
    .io_alloc_bits_tag(abc_mshr_7_io_alloc_bits_tag),
    .io_alloc_bits_off(abc_mshr_7_io_alloc_bits_off),
    .io_alloc_bits_mask(abc_mshr_7_io_alloc_bits_mask),
    .io_alloc_bits_bufIdx(abc_mshr_7_io_alloc_bits_bufIdx),
    .io_alloc_bits_preferCache(abc_mshr_7_io_alloc_bits_preferCache),
    .io_alloc_bits_dirty(abc_mshr_7_io_alloc_bits_dirty),
    .io_alloc_bits_fromProbeHelper(abc_mshr_7_io_alloc_bits_fromProbeHelper),
    .io_alloc_bits_fromCmoHelper(abc_mshr_7_io_alloc_bits_fromCmoHelper),
    .io_alloc_bits_needProbeAckData(abc_mshr_7_io_alloc_bits_needProbeAckData),
    .io_status_valid(abc_mshr_7_io_status_valid),
    .io_status_bits_set(abc_mshr_7_io_status_bits_set),
    .io_status_bits_tag(abc_mshr_7_io_status_bits_tag),
    .io_status_bits_way(abc_mshr_7_io_status_bits_way),
    .io_status_bits_way_reg(abc_mshr_7_io_status_bits_way_reg),
    .io_status_bits_nestB(abc_mshr_7_io_status_bits_nestB),
    .io_status_bits_nestC(abc_mshr_7_io_status_bits_nestC),
    .io_status_bits_will_grant_data(abc_mshr_7_io_status_bits_will_grant_data),
    .io_status_bits_will_save_data(abc_mshr_7_io_status_bits_will_save_data),
    .io_status_bits_will_free(abc_mshr_7_io_status_bits_will_free),
    .io_resps_sink_c_valid(abc_mshr_7_io_resps_sink_c_valid),
    .io_resps_sink_c_bits_hasData(abc_mshr_7_io_resps_sink_c_bits_hasData),
    .io_resps_sink_c_bits_param(abc_mshr_7_io_resps_sink_c_bits_param),
    .io_resps_sink_c_bits_source(abc_mshr_7_io_resps_sink_c_bits_source),
    .io_resps_sink_c_bits_last(abc_mshr_7_io_resps_sink_c_bits_last),
    .io_resps_sink_c_bits_bufIdx(abc_mshr_7_io_resps_sink_c_bits_bufIdx),
    .io_resps_sink_d_valid(abc_mshr_7_io_resps_sink_d_valid),
    .io_resps_sink_d_bits_opcode(abc_mshr_7_io_resps_sink_d_bits_opcode),
    .io_resps_sink_d_bits_param(abc_mshr_7_io_resps_sink_d_bits_param),
    .io_resps_sink_d_bits_sink(abc_mshr_7_io_resps_sink_d_bits_sink),
    .io_resps_sink_d_bits_last(abc_mshr_7_io_resps_sink_d_bits_last),
    .io_resps_sink_d_bits_denied(abc_mshr_7_io_resps_sink_d_bits_denied),
    .io_resps_sink_d_bits_bufIdx(abc_mshr_7_io_resps_sink_d_bits_bufIdx),
    .io_resps_sink_e_valid(abc_mshr_7_io_resps_sink_e_valid),
    .io_resps_source_d_valid(abc_mshr_7_io_resps_source_d_valid),
    .io_nestedwb_set(abc_mshr_7_io_nestedwb_set),
    .io_nestedwb_tag(abc_mshr_7_io_nestedwb_tag),
    .io_nestedwb_btoN(abc_mshr_7_io_nestedwb_btoN),
    .io_nestedwb_btoB(abc_mshr_7_io_nestedwb_btoB),
    .io_nestedwb_bclr_dirty(abc_mshr_7_io_nestedwb_bclr_dirty),
    .io_nestedwb_bset_dirty(abc_mshr_7_io_nestedwb_bset_dirty),
    .io_nestedwb_c_set_dirty(abc_mshr_7_io_nestedwb_c_set_dirty),
    .io_nestedwb_c_set_hit(abc_mshr_7_io_nestedwb_c_set_hit),
    .io_nestedwb_clients_0_isToN(abc_mshr_7_io_nestedwb_clients_0_isToN),
    .io_nestedwb_clients_1_isToN(abc_mshr_7_io_nestedwb_clients_1_isToN),
    .io_tasks_sink_a_ready(abc_mshr_7_io_tasks_sink_a_ready),
    .io_tasks_sink_a_valid(abc_mshr_7_io_tasks_sink_a_valid),
    .io_tasks_sink_a_bits_sourceId(abc_mshr_7_io_tasks_sink_a_bits_sourceId),
    .io_tasks_sink_a_bits_set(abc_mshr_7_io_tasks_sink_a_bits_set),
    .io_tasks_sink_a_bits_tag(abc_mshr_7_io_tasks_sink_a_bits_tag),
    .io_tasks_sink_a_bits_size(abc_mshr_7_io_tasks_sink_a_bits_size),
    .io_tasks_sink_a_bits_off(abc_mshr_7_io_tasks_sink_a_bits_off),
    .io_tasks_source_bready(abc_mshr_7_io_tasks_source_bready),
    .io_tasks_source_bvalid(abc_mshr_7_io_tasks_source_bvalid),
    .io_tasks_source_bset(abc_mshr_7_io_tasks_source_bset),
    .io_tasks_source_btag(abc_mshr_7_io_tasks_source_btag),
    .io_tasks_source_bparam(abc_mshr_7_io_tasks_source_bparam),
    .io_tasks_source_bclients(abc_mshr_7_io_tasks_source_bclients),
    .io_tasks_source_bneedData(abc_mshr_7_io_tasks_source_bneedData),
    .io_tasks_sink_c_ready(abc_mshr_7_io_tasks_sink_c_ready),
    .io_tasks_sink_c_valid(abc_mshr_7_io_tasks_sink_c_valid),
    .io_tasks_sink_c_bits_sourceId(abc_mshr_7_io_tasks_sink_c_bits_sourceId),
    .io_tasks_sink_c_bits_set(abc_mshr_7_io_tasks_sink_c_bits_set),
    .io_tasks_sink_c_bits_tag(abc_mshr_7_io_tasks_sink_c_bits_tag),
    .io_tasks_sink_c_bits_size(abc_mshr_7_io_tasks_sink_c_bits_size),
    .io_tasks_sink_c_bits_way(abc_mshr_7_io_tasks_sink_c_bits_way),
    .io_tasks_sink_c_bits_off(abc_mshr_7_io_tasks_sink_c_bits_off),
    .io_tasks_sink_c_bits_bufIdx(abc_mshr_7_io_tasks_sink_c_bits_bufIdx),
    .io_tasks_sink_c_bits_opcode(abc_mshr_7_io_tasks_sink_c_bits_opcode),
    .io_tasks_sink_c_bits_param(abc_mshr_7_io_tasks_sink_c_bits_param),
    .io_tasks_sink_c_bits_source(abc_mshr_7_io_tasks_sink_c_bits_source),
    .io_tasks_sink_c_bits_save(abc_mshr_7_io_tasks_sink_c_bits_save),
    .io_tasks_sink_c_bits_drop(abc_mshr_7_io_tasks_sink_c_bits_drop),
    .io_tasks_sink_c_bits_release(abc_mshr_7_io_tasks_sink_c_bits_release),
    .io_tasks_sink_c_bits_dirty(abc_mshr_7_io_tasks_sink_c_bits_dirty),
    .io_tasks_source_d_ready(abc_mshr_7_io_tasks_source_d_ready),
    .io_tasks_source_d_valid(abc_mshr_7_io_tasks_source_d_valid),
    .io_tasks_source_d_bits_sourceId(abc_mshr_7_io_tasks_source_d_bits_sourceId),
    .io_tasks_source_d_bits_set(abc_mshr_7_io_tasks_source_d_bits_set),
    .io_tasks_source_d_bits_tag(abc_mshr_7_io_tasks_source_d_bits_tag),
    .io_tasks_source_d_bits_channel(abc_mshr_7_io_tasks_source_d_bits_channel),
    .io_tasks_source_d_bits_opcode(abc_mshr_7_io_tasks_source_d_bits_opcode),
    .io_tasks_source_d_bits_param(abc_mshr_7_io_tasks_source_d_bits_param),
    .io_tasks_source_d_bits_size(abc_mshr_7_io_tasks_source_d_bits_size),
    .io_tasks_source_d_bits_way(abc_mshr_7_io_tasks_source_d_bits_way),
    .io_tasks_source_d_bits_off(abc_mshr_7_io_tasks_source_d_bits_off),
    .io_tasks_source_d_bits_useBypass(abc_mshr_7_io_tasks_source_d_bits_useBypass),
    .io_tasks_source_d_bits_bufIdx(abc_mshr_7_io_tasks_source_d_bits_bufIdx),
    .io_tasks_source_d_bits_denied(abc_mshr_7_io_tasks_source_d_bits_denied),
    .io_tasks_source_d_bits_sinkId(abc_mshr_7_io_tasks_source_d_bits_sinkId),
    .io_tasks_source_d_bits_bypassPut(abc_mshr_7_io_tasks_source_d_bits_bypassPut),
    .io_tasks_source_d_bits_dirty(abc_mshr_7_io_tasks_source_d_bits_dirty),
    .io_tasks_source_a_ready(abc_mshr_7_io_tasks_source_a_ready),
    .io_tasks_source_a_valid(abc_mshr_7_io_tasks_source_a_valid),
    .io_tasks_source_a_bits_tag(abc_mshr_7_io_tasks_source_a_bits_tag),
    .io_tasks_source_a_bits_set(abc_mshr_7_io_tasks_source_a_bits_set),
    .io_tasks_source_a_bits_off(abc_mshr_7_io_tasks_source_a_bits_off),
    .io_tasks_source_a_bits_mask(abc_mshr_7_io_tasks_source_a_bits_mask),
    .io_tasks_source_a_bits_opcode(abc_mshr_7_io_tasks_source_a_bits_opcode),
    .io_tasks_source_a_bits_param(abc_mshr_7_io_tasks_source_a_bits_param),
    .io_tasks_source_a_bits_source(abc_mshr_7_io_tasks_source_a_bits_source),
    .io_tasks_source_a_bits_bufIdx(abc_mshr_7_io_tasks_source_a_bits_bufIdx),
    .io_tasks_source_a_bits_size(abc_mshr_7_io_tasks_source_a_bits_size),
    .io_tasks_source_a_bits_needData(abc_mshr_7_io_tasks_source_a_bits_needData),
    .io_tasks_source_a_bits_putData(abc_mshr_7_io_tasks_source_a_bits_putData),
    .io_tasks_source_c_ready(abc_mshr_7_io_tasks_source_c_ready),
    .io_tasks_source_c_valid(abc_mshr_7_io_tasks_source_c_valid),
    .io_tasks_source_c_bits_opcode(abc_mshr_7_io_tasks_source_c_bits_opcode),
    .io_tasks_source_c_bits_tag(abc_mshr_7_io_tasks_source_c_bits_tag),
    .io_tasks_source_c_bits_set(abc_mshr_7_io_tasks_source_c_bits_set),
    .io_tasks_source_c_bits_param(abc_mshr_7_io_tasks_source_c_bits_param),
    .io_tasks_source_c_bits_source(abc_mshr_7_io_tasks_source_c_bits_source),
    .io_tasks_source_c_bits_way(abc_mshr_7_io_tasks_source_c_bits_way),
    .io_tasks_source_c_bits_dirty(abc_mshr_7_io_tasks_source_c_bits_dirty),
    .io_tasks_source_e_ready(abc_mshr_7_io_tasks_source_e_ready),
    .io_tasks_source_e_valid(abc_mshr_7_io_tasks_source_e_valid),
    .io_tasks_source_e_bits_sink(abc_mshr_7_io_tasks_source_e_bits_sink),
    .io_tasks_dir_write_ready(abc_mshr_7_io_tasks_dir_write_ready),
    .io_tasks_dir_write_valid(abc_mshr_7_io_tasks_dir_write_valid),
    .io_tasks_dir_write_bits_set(abc_mshr_7_io_tasks_dir_write_bits_set),
    .io_tasks_dir_write_bits_way(abc_mshr_7_io_tasks_dir_write_bits_way),
    .io_tasks_dir_write_bits_data_dirty(abc_mshr_7_io_tasks_dir_write_bits_data_dirty),
    .io_tasks_dir_write_bits_data_state(abc_mshr_7_io_tasks_dir_write_bits_data_state),
    .io_tasks_dir_write_bits_data_clientStates_0(abc_mshr_7_io_tasks_dir_write_bits_data_clientStates_0),
    .io_tasks_dir_write_bits_data_clientStates_1(abc_mshr_7_io_tasks_dir_write_bits_data_clientStates_1),
    .io_tasks_tag_write_ready(abc_mshr_7_io_tasks_tag_write_ready),
    .io_tasks_tag_write_valid(abc_mshr_7_io_tasks_tag_write_valid),
    .io_tasks_tag_write_bits_set(abc_mshr_7_io_tasks_tag_write_bits_set),
    .io_tasks_tag_write_bits_way(abc_mshr_7_io_tasks_tag_write_bits_way),
    .io_tasks_tag_write_bits_tag(abc_mshr_7_io_tasks_tag_write_bits_tag),
    .io_tasks_client_dir_write_ready(abc_mshr_7_io_tasks_client_dir_write_ready),
    .io_tasks_client_dir_write_valid(abc_mshr_7_io_tasks_client_dir_write_valid),
    .io_tasks_client_dir_write_bits_set(abc_mshr_7_io_tasks_client_dir_write_bits_set),
    .io_tasks_client_dir_write_bits_way(abc_mshr_7_io_tasks_client_dir_write_bits_way),
    .io_tasks_client_dir_write_bits_data_0_state(abc_mshr_7_io_tasks_client_dir_write_bits_data_0_state),
    .io_tasks_client_dir_write_bits_data_1_state(abc_mshr_7_io_tasks_client_dir_write_bits_data_1_state),
    .io_tasks_client_tag_write_ready(abc_mshr_7_io_tasks_client_tag_write_ready),
    .io_tasks_client_tag_write_valid(abc_mshr_7_io_tasks_client_tag_write_valid),
    .io_tasks_client_tag_write_bits_set(abc_mshr_7_io_tasks_client_tag_write_bits_set),
    .io_tasks_client_tag_write_bits_way(abc_mshr_7_io_tasks_client_tag_write_bits_way),
    .io_tasks_client_tag_write_bits_tag(abc_mshr_7_io_tasks_client_tag_write_bits_tag),
    .io_dirResult_valid(abc_mshr_7_io_dirResult_valid),
    .io_dirResult_bits_self_dirty(abc_mshr_7_io_dirResult_bits_self_dirty),
    .io_dirResult_bits_self_state(abc_mshr_7_io_dirResult_bits_self_state),
    .io_dirResult_bits_self_clientStates_0(abc_mshr_7_io_dirResult_bits_self_clientStates_0),
    .io_dirResult_bits_self_clientStates_1(abc_mshr_7_io_dirResult_bits_self_clientStates_1),
    .io_dirResult_bits_self_hit(abc_mshr_7_io_dirResult_bits_self_hit),
    .io_dirResult_bits_self_way(abc_mshr_7_io_dirResult_bits_self_way),
    .io_dirResult_bits_self_tag(abc_mshr_7_io_dirResult_bits_self_tag),
    .io_dirResult_bits_clients_states_0_state(abc_mshr_7_io_dirResult_bits_clients_states_0_state),
    .io_dirResult_bits_clients_states_0_hit(abc_mshr_7_io_dirResult_bits_clients_states_0_hit),
    .io_dirResult_bits_clients_states_1_state(abc_mshr_7_io_dirResult_bits_clients_states_1_state),
    .io_dirResult_bits_clients_states_1_hit(abc_mshr_7_io_dirResult_bits_clients_states_1_hit),
    .io_dirResult_bits_clients_tag(abc_mshr_7_io_dirResult_bits_clients_tag),
    .io_dirResult_bits_clients_way(abc_mshr_7_io_dirResult_bits_clients_way),
    .io_c_status_set(abc_mshr_7_io_c_status_set),
    .io_c_status_tag(abc_mshr_7_io_c_status_tag),
    .io_c_status_way(abc_mshr_7_io_c_status_way),
    .io_c_status_nestedReleaseData(abc_mshr_7_io_c_status_nestedReleaseData),
    .io_c_status_releaseThrough(abc_mshr_7_io_c_status_releaseThrough),
    .io_bstatus_set(abc_mshr_7_io_bstatus_set),
    .io_bstatus_tag(abc_mshr_7_io_bstatus_tag),
    .io_bstatus_way(abc_mshr_7_io_bstatus_way),
    .io_bstatus_nestedProbeAckData(abc_mshr_7_io_bstatus_nestedProbeAckData),
    .io_bstatus_probeHelperFinish(abc_mshr_7_io_bstatus_probeHelperFinish),
    .io_bstatus_probeAckDataThrough(abc_mshr_7_io_bstatus_probeAckDataThrough),
    .io_releaseThrough(abc_mshr_7_io_releaseThrough),
    .io_probeAckDataThrough(abc_mshr_7_io_probeAckDataThrough),
    .io_is_nestedReleaseData(abc_mshr_7_io_is_nestedReleaseData),
    .io_is_nestedProbeAckData(abc_mshr_7_io_is_nestedProbeAckData),
    .io_probeHelperFinish(abc_mshr_7_io_probeHelperFinish)
  );
  MSHR abc_mshr_8 ( // @[Slice.scala 94:16]
    .clock(abc_mshr_8_clock),
    .reset(abc_mshr_8_reset),
    .io_id(abc_mshr_8_io_id),
    .io_enable(abc_mshr_8_io_enable),
    .io_alloc_valid(abc_mshr_8_io_alloc_valid),
    .io_alloc_bits_channel(abc_mshr_8_io_alloc_bits_channel),
    .io_alloc_bits_opcode(abc_mshr_8_io_alloc_bits_opcode),
    .io_alloc_bits_param(abc_mshr_8_io_alloc_bits_param),
    .io_alloc_bits_size(abc_mshr_8_io_alloc_bits_size),
    .io_alloc_bits_source(abc_mshr_8_io_alloc_bits_source),
    .io_alloc_bits_set(abc_mshr_8_io_alloc_bits_set),
    .io_alloc_bits_tag(abc_mshr_8_io_alloc_bits_tag),
    .io_alloc_bits_off(abc_mshr_8_io_alloc_bits_off),
    .io_alloc_bits_mask(abc_mshr_8_io_alloc_bits_mask),
    .io_alloc_bits_bufIdx(abc_mshr_8_io_alloc_bits_bufIdx),
    .io_alloc_bits_preferCache(abc_mshr_8_io_alloc_bits_preferCache),
    .io_alloc_bits_dirty(abc_mshr_8_io_alloc_bits_dirty),
    .io_alloc_bits_fromProbeHelper(abc_mshr_8_io_alloc_bits_fromProbeHelper),
    .io_alloc_bits_fromCmoHelper(abc_mshr_8_io_alloc_bits_fromCmoHelper),
    .io_alloc_bits_needProbeAckData(abc_mshr_8_io_alloc_bits_needProbeAckData),
    .io_status_valid(abc_mshr_8_io_status_valid),
    .io_status_bits_set(abc_mshr_8_io_status_bits_set),
    .io_status_bits_tag(abc_mshr_8_io_status_bits_tag),
    .io_status_bits_way(abc_mshr_8_io_status_bits_way),
    .io_status_bits_way_reg(abc_mshr_8_io_status_bits_way_reg),
    .io_status_bits_nestB(abc_mshr_8_io_status_bits_nestB),
    .io_status_bits_nestC(abc_mshr_8_io_status_bits_nestC),
    .io_status_bits_will_grant_data(abc_mshr_8_io_status_bits_will_grant_data),
    .io_status_bits_will_save_data(abc_mshr_8_io_status_bits_will_save_data),
    .io_status_bits_will_free(abc_mshr_8_io_status_bits_will_free),
    .io_resps_sink_c_valid(abc_mshr_8_io_resps_sink_c_valid),
    .io_resps_sink_c_bits_hasData(abc_mshr_8_io_resps_sink_c_bits_hasData),
    .io_resps_sink_c_bits_param(abc_mshr_8_io_resps_sink_c_bits_param),
    .io_resps_sink_c_bits_source(abc_mshr_8_io_resps_sink_c_bits_source),
    .io_resps_sink_c_bits_last(abc_mshr_8_io_resps_sink_c_bits_last),
    .io_resps_sink_c_bits_bufIdx(abc_mshr_8_io_resps_sink_c_bits_bufIdx),
    .io_resps_sink_d_valid(abc_mshr_8_io_resps_sink_d_valid),
    .io_resps_sink_d_bits_opcode(abc_mshr_8_io_resps_sink_d_bits_opcode),
    .io_resps_sink_d_bits_param(abc_mshr_8_io_resps_sink_d_bits_param),
    .io_resps_sink_d_bits_sink(abc_mshr_8_io_resps_sink_d_bits_sink),
    .io_resps_sink_d_bits_last(abc_mshr_8_io_resps_sink_d_bits_last),
    .io_resps_sink_d_bits_denied(abc_mshr_8_io_resps_sink_d_bits_denied),
    .io_resps_sink_d_bits_bufIdx(abc_mshr_8_io_resps_sink_d_bits_bufIdx),
    .io_resps_sink_e_valid(abc_mshr_8_io_resps_sink_e_valid),
    .io_resps_source_d_valid(abc_mshr_8_io_resps_source_d_valid),
    .io_nestedwb_set(abc_mshr_8_io_nestedwb_set),
    .io_nestedwb_tag(abc_mshr_8_io_nestedwb_tag),
    .io_nestedwb_btoN(abc_mshr_8_io_nestedwb_btoN),
    .io_nestedwb_btoB(abc_mshr_8_io_nestedwb_btoB),
    .io_nestedwb_bclr_dirty(abc_mshr_8_io_nestedwb_bclr_dirty),
    .io_nestedwb_bset_dirty(abc_mshr_8_io_nestedwb_bset_dirty),
    .io_nestedwb_c_set_dirty(abc_mshr_8_io_nestedwb_c_set_dirty),
    .io_nestedwb_c_set_hit(abc_mshr_8_io_nestedwb_c_set_hit),
    .io_nestedwb_clients_0_isToN(abc_mshr_8_io_nestedwb_clients_0_isToN),
    .io_nestedwb_clients_1_isToN(abc_mshr_8_io_nestedwb_clients_1_isToN),
    .io_tasks_sink_a_ready(abc_mshr_8_io_tasks_sink_a_ready),
    .io_tasks_sink_a_valid(abc_mshr_8_io_tasks_sink_a_valid),
    .io_tasks_sink_a_bits_sourceId(abc_mshr_8_io_tasks_sink_a_bits_sourceId),
    .io_tasks_sink_a_bits_set(abc_mshr_8_io_tasks_sink_a_bits_set),
    .io_tasks_sink_a_bits_tag(abc_mshr_8_io_tasks_sink_a_bits_tag),
    .io_tasks_sink_a_bits_size(abc_mshr_8_io_tasks_sink_a_bits_size),
    .io_tasks_sink_a_bits_off(abc_mshr_8_io_tasks_sink_a_bits_off),
    .io_tasks_source_bready(abc_mshr_8_io_tasks_source_bready),
    .io_tasks_source_bvalid(abc_mshr_8_io_tasks_source_bvalid),
    .io_tasks_source_bset(abc_mshr_8_io_tasks_source_bset),
    .io_tasks_source_btag(abc_mshr_8_io_tasks_source_btag),
    .io_tasks_source_bparam(abc_mshr_8_io_tasks_source_bparam),
    .io_tasks_source_bclients(abc_mshr_8_io_tasks_source_bclients),
    .io_tasks_source_bneedData(abc_mshr_8_io_tasks_source_bneedData),
    .io_tasks_sink_c_ready(abc_mshr_8_io_tasks_sink_c_ready),
    .io_tasks_sink_c_valid(abc_mshr_8_io_tasks_sink_c_valid),
    .io_tasks_sink_c_bits_sourceId(abc_mshr_8_io_tasks_sink_c_bits_sourceId),
    .io_tasks_sink_c_bits_set(abc_mshr_8_io_tasks_sink_c_bits_set),
    .io_tasks_sink_c_bits_tag(abc_mshr_8_io_tasks_sink_c_bits_tag),
    .io_tasks_sink_c_bits_size(abc_mshr_8_io_tasks_sink_c_bits_size),
    .io_tasks_sink_c_bits_way(abc_mshr_8_io_tasks_sink_c_bits_way),
    .io_tasks_sink_c_bits_off(abc_mshr_8_io_tasks_sink_c_bits_off),
    .io_tasks_sink_c_bits_bufIdx(abc_mshr_8_io_tasks_sink_c_bits_bufIdx),
    .io_tasks_sink_c_bits_opcode(abc_mshr_8_io_tasks_sink_c_bits_opcode),
    .io_tasks_sink_c_bits_param(abc_mshr_8_io_tasks_sink_c_bits_param),
    .io_tasks_sink_c_bits_source(abc_mshr_8_io_tasks_sink_c_bits_source),
    .io_tasks_sink_c_bits_save(abc_mshr_8_io_tasks_sink_c_bits_save),
    .io_tasks_sink_c_bits_drop(abc_mshr_8_io_tasks_sink_c_bits_drop),
    .io_tasks_sink_c_bits_release(abc_mshr_8_io_tasks_sink_c_bits_release),
    .io_tasks_sink_c_bits_dirty(abc_mshr_8_io_tasks_sink_c_bits_dirty),
    .io_tasks_source_d_ready(abc_mshr_8_io_tasks_source_d_ready),
    .io_tasks_source_d_valid(abc_mshr_8_io_tasks_source_d_valid),
    .io_tasks_source_d_bits_sourceId(abc_mshr_8_io_tasks_source_d_bits_sourceId),
    .io_tasks_source_d_bits_set(abc_mshr_8_io_tasks_source_d_bits_set),
    .io_tasks_source_d_bits_tag(abc_mshr_8_io_tasks_source_d_bits_tag),
    .io_tasks_source_d_bits_channel(abc_mshr_8_io_tasks_source_d_bits_channel),
    .io_tasks_source_d_bits_opcode(abc_mshr_8_io_tasks_source_d_bits_opcode),
    .io_tasks_source_d_bits_param(abc_mshr_8_io_tasks_source_d_bits_param),
    .io_tasks_source_d_bits_size(abc_mshr_8_io_tasks_source_d_bits_size),
    .io_tasks_source_d_bits_way(abc_mshr_8_io_tasks_source_d_bits_way),
    .io_tasks_source_d_bits_off(abc_mshr_8_io_tasks_source_d_bits_off),
    .io_tasks_source_d_bits_useBypass(abc_mshr_8_io_tasks_source_d_bits_useBypass),
    .io_tasks_source_d_bits_bufIdx(abc_mshr_8_io_tasks_source_d_bits_bufIdx),
    .io_tasks_source_d_bits_denied(abc_mshr_8_io_tasks_source_d_bits_denied),
    .io_tasks_source_d_bits_sinkId(abc_mshr_8_io_tasks_source_d_bits_sinkId),
    .io_tasks_source_d_bits_bypassPut(abc_mshr_8_io_tasks_source_d_bits_bypassPut),
    .io_tasks_source_d_bits_dirty(abc_mshr_8_io_tasks_source_d_bits_dirty),
    .io_tasks_source_a_ready(abc_mshr_8_io_tasks_source_a_ready),
    .io_tasks_source_a_valid(abc_mshr_8_io_tasks_source_a_valid),
    .io_tasks_source_a_bits_tag(abc_mshr_8_io_tasks_source_a_bits_tag),
    .io_tasks_source_a_bits_set(abc_mshr_8_io_tasks_source_a_bits_set),
    .io_tasks_source_a_bits_off(abc_mshr_8_io_tasks_source_a_bits_off),
    .io_tasks_source_a_bits_mask(abc_mshr_8_io_tasks_source_a_bits_mask),
    .io_tasks_source_a_bits_opcode(abc_mshr_8_io_tasks_source_a_bits_opcode),
    .io_tasks_source_a_bits_param(abc_mshr_8_io_tasks_source_a_bits_param),
    .io_tasks_source_a_bits_source(abc_mshr_8_io_tasks_source_a_bits_source),
    .io_tasks_source_a_bits_bufIdx(abc_mshr_8_io_tasks_source_a_bits_bufIdx),
    .io_tasks_source_a_bits_size(abc_mshr_8_io_tasks_source_a_bits_size),
    .io_tasks_source_a_bits_needData(abc_mshr_8_io_tasks_source_a_bits_needData),
    .io_tasks_source_a_bits_putData(abc_mshr_8_io_tasks_source_a_bits_putData),
    .io_tasks_source_c_ready(abc_mshr_8_io_tasks_source_c_ready),
    .io_tasks_source_c_valid(abc_mshr_8_io_tasks_source_c_valid),
    .io_tasks_source_c_bits_opcode(abc_mshr_8_io_tasks_source_c_bits_opcode),
    .io_tasks_source_c_bits_tag(abc_mshr_8_io_tasks_source_c_bits_tag),
    .io_tasks_source_c_bits_set(abc_mshr_8_io_tasks_source_c_bits_set),
    .io_tasks_source_c_bits_param(abc_mshr_8_io_tasks_source_c_bits_param),
    .io_tasks_source_c_bits_source(abc_mshr_8_io_tasks_source_c_bits_source),
    .io_tasks_source_c_bits_way(abc_mshr_8_io_tasks_source_c_bits_way),
    .io_tasks_source_c_bits_dirty(abc_mshr_8_io_tasks_source_c_bits_dirty),
    .io_tasks_source_e_ready(abc_mshr_8_io_tasks_source_e_ready),
    .io_tasks_source_e_valid(abc_mshr_8_io_tasks_source_e_valid),
    .io_tasks_source_e_bits_sink(abc_mshr_8_io_tasks_source_e_bits_sink),
    .io_tasks_dir_write_ready(abc_mshr_8_io_tasks_dir_write_ready),
    .io_tasks_dir_write_valid(abc_mshr_8_io_tasks_dir_write_valid),
    .io_tasks_dir_write_bits_set(abc_mshr_8_io_tasks_dir_write_bits_set),
    .io_tasks_dir_write_bits_way(abc_mshr_8_io_tasks_dir_write_bits_way),
    .io_tasks_dir_write_bits_data_dirty(abc_mshr_8_io_tasks_dir_write_bits_data_dirty),
    .io_tasks_dir_write_bits_data_state(abc_mshr_8_io_tasks_dir_write_bits_data_state),
    .io_tasks_dir_write_bits_data_clientStates_0(abc_mshr_8_io_tasks_dir_write_bits_data_clientStates_0),
    .io_tasks_dir_write_bits_data_clientStates_1(abc_mshr_8_io_tasks_dir_write_bits_data_clientStates_1),
    .io_tasks_tag_write_ready(abc_mshr_8_io_tasks_tag_write_ready),
    .io_tasks_tag_write_valid(abc_mshr_8_io_tasks_tag_write_valid),
    .io_tasks_tag_write_bits_set(abc_mshr_8_io_tasks_tag_write_bits_set),
    .io_tasks_tag_write_bits_way(abc_mshr_8_io_tasks_tag_write_bits_way),
    .io_tasks_tag_write_bits_tag(abc_mshr_8_io_tasks_tag_write_bits_tag),
    .io_tasks_client_dir_write_ready(abc_mshr_8_io_tasks_client_dir_write_ready),
    .io_tasks_client_dir_write_valid(abc_mshr_8_io_tasks_client_dir_write_valid),
    .io_tasks_client_dir_write_bits_set(abc_mshr_8_io_tasks_client_dir_write_bits_set),
    .io_tasks_client_dir_write_bits_way(abc_mshr_8_io_tasks_client_dir_write_bits_way),
    .io_tasks_client_dir_write_bits_data_0_state(abc_mshr_8_io_tasks_client_dir_write_bits_data_0_state),
    .io_tasks_client_dir_write_bits_data_1_state(abc_mshr_8_io_tasks_client_dir_write_bits_data_1_state),
    .io_tasks_client_tag_write_ready(abc_mshr_8_io_tasks_client_tag_write_ready),
    .io_tasks_client_tag_write_valid(abc_mshr_8_io_tasks_client_tag_write_valid),
    .io_tasks_client_tag_write_bits_set(abc_mshr_8_io_tasks_client_tag_write_bits_set),
    .io_tasks_client_tag_write_bits_way(abc_mshr_8_io_tasks_client_tag_write_bits_way),
    .io_tasks_client_tag_write_bits_tag(abc_mshr_8_io_tasks_client_tag_write_bits_tag),
    .io_dirResult_valid(abc_mshr_8_io_dirResult_valid),
    .io_dirResult_bits_self_dirty(abc_mshr_8_io_dirResult_bits_self_dirty),
    .io_dirResult_bits_self_state(abc_mshr_8_io_dirResult_bits_self_state),
    .io_dirResult_bits_self_clientStates_0(abc_mshr_8_io_dirResult_bits_self_clientStates_0),
    .io_dirResult_bits_self_clientStates_1(abc_mshr_8_io_dirResult_bits_self_clientStates_1),
    .io_dirResult_bits_self_hit(abc_mshr_8_io_dirResult_bits_self_hit),
    .io_dirResult_bits_self_way(abc_mshr_8_io_dirResult_bits_self_way),
    .io_dirResult_bits_self_tag(abc_mshr_8_io_dirResult_bits_self_tag),
    .io_dirResult_bits_clients_states_0_state(abc_mshr_8_io_dirResult_bits_clients_states_0_state),
    .io_dirResult_bits_clients_states_0_hit(abc_mshr_8_io_dirResult_bits_clients_states_0_hit),
    .io_dirResult_bits_clients_states_1_state(abc_mshr_8_io_dirResult_bits_clients_states_1_state),
    .io_dirResult_bits_clients_states_1_hit(abc_mshr_8_io_dirResult_bits_clients_states_1_hit),
    .io_dirResult_bits_clients_tag(abc_mshr_8_io_dirResult_bits_clients_tag),
    .io_dirResult_bits_clients_way(abc_mshr_8_io_dirResult_bits_clients_way),
    .io_c_status_set(abc_mshr_8_io_c_status_set),
    .io_c_status_tag(abc_mshr_8_io_c_status_tag),
    .io_c_status_way(abc_mshr_8_io_c_status_way),
    .io_c_status_nestedReleaseData(abc_mshr_8_io_c_status_nestedReleaseData),
    .io_c_status_releaseThrough(abc_mshr_8_io_c_status_releaseThrough),
    .io_bstatus_set(abc_mshr_8_io_bstatus_set),
    .io_bstatus_tag(abc_mshr_8_io_bstatus_tag),
    .io_bstatus_way(abc_mshr_8_io_bstatus_way),
    .io_bstatus_nestedProbeAckData(abc_mshr_8_io_bstatus_nestedProbeAckData),
    .io_bstatus_probeHelperFinish(abc_mshr_8_io_bstatus_probeHelperFinish),
    .io_bstatus_probeAckDataThrough(abc_mshr_8_io_bstatus_probeAckDataThrough),
    .io_releaseThrough(abc_mshr_8_io_releaseThrough),
    .io_probeAckDataThrough(abc_mshr_8_io_probeAckDataThrough),
    .io_is_nestedReleaseData(abc_mshr_8_io_is_nestedReleaseData),
    .io_is_nestedProbeAckData(abc_mshr_8_io_is_nestedProbeAckData),
    .io_probeHelperFinish(abc_mshr_8_io_probeHelperFinish)
  );
  MSHR abc_mshr_9 ( // @[Slice.scala 94:16]
    .clock(abc_mshr_9_clock),
    .reset(abc_mshr_9_reset),
    .io_id(abc_mshr_9_io_id),
    .io_enable(abc_mshr_9_io_enable),
    .io_alloc_valid(abc_mshr_9_io_alloc_valid),
    .io_alloc_bits_channel(abc_mshr_9_io_alloc_bits_channel),
    .io_alloc_bits_opcode(abc_mshr_9_io_alloc_bits_opcode),
    .io_alloc_bits_param(abc_mshr_9_io_alloc_bits_param),
    .io_alloc_bits_size(abc_mshr_9_io_alloc_bits_size),
    .io_alloc_bits_source(abc_mshr_9_io_alloc_bits_source),
    .io_alloc_bits_set(abc_mshr_9_io_alloc_bits_set),
    .io_alloc_bits_tag(abc_mshr_9_io_alloc_bits_tag),
    .io_alloc_bits_off(abc_mshr_9_io_alloc_bits_off),
    .io_alloc_bits_mask(abc_mshr_9_io_alloc_bits_mask),
    .io_alloc_bits_bufIdx(abc_mshr_9_io_alloc_bits_bufIdx),
    .io_alloc_bits_preferCache(abc_mshr_9_io_alloc_bits_preferCache),
    .io_alloc_bits_dirty(abc_mshr_9_io_alloc_bits_dirty),
    .io_alloc_bits_fromProbeHelper(abc_mshr_9_io_alloc_bits_fromProbeHelper),
    .io_alloc_bits_fromCmoHelper(abc_mshr_9_io_alloc_bits_fromCmoHelper),
    .io_alloc_bits_needProbeAckData(abc_mshr_9_io_alloc_bits_needProbeAckData),
    .io_status_valid(abc_mshr_9_io_status_valid),
    .io_status_bits_set(abc_mshr_9_io_status_bits_set),
    .io_status_bits_tag(abc_mshr_9_io_status_bits_tag),
    .io_status_bits_way(abc_mshr_9_io_status_bits_way),
    .io_status_bits_way_reg(abc_mshr_9_io_status_bits_way_reg),
    .io_status_bits_nestB(abc_mshr_9_io_status_bits_nestB),
    .io_status_bits_nestC(abc_mshr_9_io_status_bits_nestC),
    .io_status_bits_will_grant_data(abc_mshr_9_io_status_bits_will_grant_data),
    .io_status_bits_will_save_data(abc_mshr_9_io_status_bits_will_save_data),
    .io_status_bits_will_free(abc_mshr_9_io_status_bits_will_free),
    .io_resps_sink_c_valid(abc_mshr_9_io_resps_sink_c_valid),
    .io_resps_sink_c_bits_hasData(abc_mshr_9_io_resps_sink_c_bits_hasData),
    .io_resps_sink_c_bits_param(abc_mshr_9_io_resps_sink_c_bits_param),
    .io_resps_sink_c_bits_source(abc_mshr_9_io_resps_sink_c_bits_source),
    .io_resps_sink_c_bits_last(abc_mshr_9_io_resps_sink_c_bits_last),
    .io_resps_sink_c_bits_bufIdx(abc_mshr_9_io_resps_sink_c_bits_bufIdx),
    .io_resps_sink_d_valid(abc_mshr_9_io_resps_sink_d_valid),
    .io_resps_sink_d_bits_opcode(abc_mshr_9_io_resps_sink_d_bits_opcode),
    .io_resps_sink_d_bits_param(abc_mshr_9_io_resps_sink_d_bits_param),
    .io_resps_sink_d_bits_sink(abc_mshr_9_io_resps_sink_d_bits_sink),
    .io_resps_sink_d_bits_last(abc_mshr_9_io_resps_sink_d_bits_last),
    .io_resps_sink_d_bits_denied(abc_mshr_9_io_resps_sink_d_bits_denied),
    .io_resps_sink_d_bits_bufIdx(abc_mshr_9_io_resps_sink_d_bits_bufIdx),
    .io_resps_sink_e_valid(abc_mshr_9_io_resps_sink_e_valid),
    .io_resps_source_d_valid(abc_mshr_9_io_resps_source_d_valid),
    .io_nestedwb_set(abc_mshr_9_io_nestedwb_set),
    .io_nestedwb_tag(abc_mshr_9_io_nestedwb_tag),
    .io_nestedwb_btoN(abc_mshr_9_io_nestedwb_btoN),
    .io_nestedwb_btoB(abc_mshr_9_io_nestedwb_btoB),
    .io_nestedwb_bclr_dirty(abc_mshr_9_io_nestedwb_bclr_dirty),
    .io_nestedwb_bset_dirty(abc_mshr_9_io_nestedwb_bset_dirty),
    .io_nestedwb_c_set_dirty(abc_mshr_9_io_nestedwb_c_set_dirty),
    .io_nestedwb_c_set_hit(abc_mshr_9_io_nestedwb_c_set_hit),
    .io_nestedwb_clients_0_isToN(abc_mshr_9_io_nestedwb_clients_0_isToN),
    .io_nestedwb_clients_1_isToN(abc_mshr_9_io_nestedwb_clients_1_isToN),
    .io_tasks_sink_a_ready(abc_mshr_9_io_tasks_sink_a_ready),
    .io_tasks_sink_a_valid(abc_mshr_9_io_tasks_sink_a_valid),
    .io_tasks_sink_a_bits_sourceId(abc_mshr_9_io_tasks_sink_a_bits_sourceId),
    .io_tasks_sink_a_bits_set(abc_mshr_9_io_tasks_sink_a_bits_set),
    .io_tasks_sink_a_bits_tag(abc_mshr_9_io_tasks_sink_a_bits_tag),
    .io_tasks_sink_a_bits_size(abc_mshr_9_io_tasks_sink_a_bits_size),
    .io_tasks_sink_a_bits_off(abc_mshr_9_io_tasks_sink_a_bits_off),
    .io_tasks_source_bready(abc_mshr_9_io_tasks_source_bready),
    .io_tasks_source_bvalid(abc_mshr_9_io_tasks_source_bvalid),
    .io_tasks_source_bset(abc_mshr_9_io_tasks_source_bset),
    .io_tasks_source_btag(abc_mshr_9_io_tasks_source_btag),
    .io_tasks_source_bparam(abc_mshr_9_io_tasks_source_bparam),
    .io_tasks_source_bclients(abc_mshr_9_io_tasks_source_bclients),
    .io_tasks_source_bneedData(abc_mshr_9_io_tasks_source_bneedData),
    .io_tasks_sink_c_ready(abc_mshr_9_io_tasks_sink_c_ready),
    .io_tasks_sink_c_valid(abc_mshr_9_io_tasks_sink_c_valid),
    .io_tasks_sink_c_bits_sourceId(abc_mshr_9_io_tasks_sink_c_bits_sourceId),
    .io_tasks_sink_c_bits_set(abc_mshr_9_io_tasks_sink_c_bits_set),
    .io_tasks_sink_c_bits_tag(abc_mshr_9_io_tasks_sink_c_bits_tag),
    .io_tasks_sink_c_bits_size(abc_mshr_9_io_tasks_sink_c_bits_size),
    .io_tasks_sink_c_bits_way(abc_mshr_9_io_tasks_sink_c_bits_way),
    .io_tasks_sink_c_bits_off(abc_mshr_9_io_tasks_sink_c_bits_off),
    .io_tasks_sink_c_bits_bufIdx(abc_mshr_9_io_tasks_sink_c_bits_bufIdx),
    .io_tasks_sink_c_bits_opcode(abc_mshr_9_io_tasks_sink_c_bits_opcode),
    .io_tasks_sink_c_bits_param(abc_mshr_9_io_tasks_sink_c_bits_param),
    .io_tasks_sink_c_bits_source(abc_mshr_9_io_tasks_sink_c_bits_source),
    .io_tasks_sink_c_bits_save(abc_mshr_9_io_tasks_sink_c_bits_save),
    .io_tasks_sink_c_bits_drop(abc_mshr_9_io_tasks_sink_c_bits_drop),
    .io_tasks_sink_c_bits_release(abc_mshr_9_io_tasks_sink_c_bits_release),
    .io_tasks_sink_c_bits_dirty(abc_mshr_9_io_tasks_sink_c_bits_dirty),
    .io_tasks_source_d_ready(abc_mshr_9_io_tasks_source_d_ready),
    .io_tasks_source_d_valid(abc_mshr_9_io_tasks_source_d_valid),
    .io_tasks_source_d_bits_sourceId(abc_mshr_9_io_tasks_source_d_bits_sourceId),
    .io_tasks_source_d_bits_set(abc_mshr_9_io_tasks_source_d_bits_set),
    .io_tasks_source_d_bits_tag(abc_mshr_9_io_tasks_source_d_bits_tag),
    .io_tasks_source_d_bits_channel(abc_mshr_9_io_tasks_source_d_bits_channel),
    .io_tasks_source_d_bits_opcode(abc_mshr_9_io_tasks_source_d_bits_opcode),
    .io_tasks_source_d_bits_param(abc_mshr_9_io_tasks_source_d_bits_param),
    .io_tasks_source_d_bits_size(abc_mshr_9_io_tasks_source_d_bits_size),
    .io_tasks_source_d_bits_way(abc_mshr_9_io_tasks_source_d_bits_way),
    .io_tasks_source_d_bits_off(abc_mshr_9_io_tasks_source_d_bits_off),
    .io_tasks_source_d_bits_useBypass(abc_mshr_9_io_tasks_source_d_bits_useBypass),
    .io_tasks_source_d_bits_bufIdx(abc_mshr_9_io_tasks_source_d_bits_bufIdx),
    .io_tasks_source_d_bits_denied(abc_mshr_9_io_tasks_source_d_bits_denied),
    .io_tasks_source_d_bits_sinkId(abc_mshr_9_io_tasks_source_d_bits_sinkId),
    .io_tasks_source_d_bits_bypassPut(abc_mshr_9_io_tasks_source_d_bits_bypassPut),
    .io_tasks_source_d_bits_dirty(abc_mshr_9_io_tasks_source_d_bits_dirty),
    .io_tasks_source_a_ready(abc_mshr_9_io_tasks_source_a_ready),
    .io_tasks_source_a_valid(abc_mshr_9_io_tasks_source_a_valid),
    .io_tasks_source_a_bits_tag(abc_mshr_9_io_tasks_source_a_bits_tag),
    .io_tasks_source_a_bits_set(abc_mshr_9_io_tasks_source_a_bits_set),
    .io_tasks_source_a_bits_off(abc_mshr_9_io_tasks_source_a_bits_off),
    .io_tasks_source_a_bits_mask(abc_mshr_9_io_tasks_source_a_bits_mask),
    .io_tasks_source_a_bits_opcode(abc_mshr_9_io_tasks_source_a_bits_opcode),
    .io_tasks_source_a_bits_param(abc_mshr_9_io_tasks_source_a_bits_param),
    .io_tasks_source_a_bits_source(abc_mshr_9_io_tasks_source_a_bits_source),
    .io_tasks_source_a_bits_bufIdx(abc_mshr_9_io_tasks_source_a_bits_bufIdx),
    .io_tasks_source_a_bits_size(abc_mshr_9_io_tasks_source_a_bits_size),
    .io_tasks_source_a_bits_needData(abc_mshr_9_io_tasks_source_a_bits_needData),
    .io_tasks_source_a_bits_putData(abc_mshr_9_io_tasks_source_a_bits_putData),
    .io_tasks_source_c_ready(abc_mshr_9_io_tasks_source_c_ready),
    .io_tasks_source_c_valid(abc_mshr_9_io_tasks_source_c_valid),
    .io_tasks_source_c_bits_opcode(abc_mshr_9_io_tasks_source_c_bits_opcode),
    .io_tasks_source_c_bits_tag(abc_mshr_9_io_tasks_source_c_bits_tag),
    .io_tasks_source_c_bits_set(abc_mshr_9_io_tasks_source_c_bits_set),
    .io_tasks_source_c_bits_param(abc_mshr_9_io_tasks_source_c_bits_param),
    .io_tasks_source_c_bits_source(abc_mshr_9_io_tasks_source_c_bits_source),
    .io_tasks_source_c_bits_way(abc_mshr_9_io_tasks_source_c_bits_way),
    .io_tasks_source_c_bits_dirty(abc_mshr_9_io_tasks_source_c_bits_dirty),
    .io_tasks_source_e_ready(abc_mshr_9_io_tasks_source_e_ready),
    .io_tasks_source_e_valid(abc_mshr_9_io_tasks_source_e_valid),
    .io_tasks_source_e_bits_sink(abc_mshr_9_io_tasks_source_e_bits_sink),
    .io_tasks_dir_write_ready(abc_mshr_9_io_tasks_dir_write_ready),
    .io_tasks_dir_write_valid(abc_mshr_9_io_tasks_dir_write_valid),
    .io_tasks_dir_write_bits_set(abc_mshr_9_io_tasks_dir_write_bits_set),
    .io_tasks_dir_write_bits_way(abc_mshr_9_io_tasks_dir_write_bits_way),
    .io_tasks_dir_write_bits_data_dirty(abc_mshr_9_io_tasks_dir_write_bits_data_dirty),
    .io_tasks_dir_write_bits_data_state(abc_mshr_9_io_tasks_dir_write_bits_data_state),
    .io_tasks_dir_write_bits_data_clientStates_0(abc_mshr_9_io_tasks_dir_write_bits_data_clientStates_0),
    .io_tasks_dir_write_bits_data_clientStates_1(abc_mshr_9_io_tasks_dir_write_bits_data_clientStates_1),
    .io_tasks_tag_write_ready(abc_mshr_9_io_tasks_tag_write_ready),
    .io_tasks_tag_write_valid(abc_mshr_9_io_tasks_tag_write_valid),
    .io_tasks_tag_write_bits_set(abc_mshr_9_io_tasks_tag_write_bits_set),
    .io_tasks_tag_write_bits_way(abc_mshr_9_io_tasks_tag_write_bits_way),
    .io_tasks_tag_write_bits_tag(abc_mshr_9_io_tasks_tag_write_bits_tag),
    .io_tasks_client_dir_write_ready(abc_mshr_9_io_tasks_client_dir_write_ready),
    .io_tasks_client_dir_write_valid(abc_mshr_9_io_tasks_client_dir_write_valid),
    .io_tasks_client_dir_write_bits_set(abc_mshr_9_io_tasks_client_dir_write_bits_set),
    .io_tasks_client_dir_write_bits_way(abc_mshr_9_io_tasks_client_dir_write_bits_way),
    .io_tasks_client_dir_write_bits_data_0_state(abc_mshr_9_io_tasks_client_dir_write_bits_data_0_state),
    .io_tasks_client_dir_write_bits_data_1_state(abc_mshr_9_io_tasks_client_dir_write_bits_data_1_state),
    .io_tasks_client_tag_write_ready(abc_mshr_9_io_tasks_client_tag_write_ready),
    .io_tasks_client_tag_write_valid(abc_mshr_9_io_tasks_client_tag_write_valid),
    .io_tasks_client_tag_write_bits_set(abc_mshr_9_io_tasks_client_tag_write_bits_set),
    .io_tasks_client_tag_write_bits_way(abc_mshr_9_io_tasks_client_tag_write_bits_way),
    .io_tasks_client_tag_write_bits_tag(abc_mshr_9_io_tasks_client_tag_write_bits_tag),
    .io_dirResult_valid(abc_mshr_9_io_dirResult_valid),
    .io_dirResult_bits_self_dirty(abc_mshr_9_io_dirResult_bits_self_dirty),
    .io_dirResult_bits_self_state(abc_mshr_9_io_dirResult_bits_self_state),
    .io_dirResult_bits_self_clientStates_0(abc_mshr_9_io_dirResult_bits_self_clientStates_0),
    .io_dirResult_bits_self_clientStates_1(abc_mshr_9_io_dirResult_bits_self_clientStates_1),
    .io_dirResult_bits_self_hit(abc_mshr_9_io_dirResult_bits_self_hit),
    .io_dirResult_bits_self_way(abc_mshr_9_io_dirResult_bits_self_way),
    .io_dirResult_bits_self_tag(abc_mshr_9_io_dirResult_bits_self_tag),
    .io_dirResult_bits_clients_states_0_state(abc_mshr_9_io_dirResult_bits_clients_states_0_state),
    .io_dirResult_bits_clients_states_0_hit(abc_mshr_9_io_dirResult_bits_clients_states_0_hit),
    .io_dirResult_bits_clients_states_1_state(abc_mshr_9_io_dirResult_bits_clients_states_1_state),
    .io_dirResult_bits_clients_states_1_hit(abc_mshr_9_io_dirResult_bits_clients_states_1_hit),
    .io_dirResult_bits_clients_tag(abc_mshr_9_io_dirResult_bits_clients_tag),
    .io_dirResult_bits_clients_way(abc_mshr_9_io_dirResult_bits_clients_way),
    .io_c_status_set(abc_mshr_9_io_c_status_set),
    .io_c_status_tag(abc_mshr_9_io_c_status_tag),
    .io_c_status_way(abc_mshr_9_io_c_status_way),
    .io_c_status_nestedReleaseData(abc_mshr_9_io_c_status_nestedReleaseData),
    .io_c_status_releaseThrough(abc_mshr_9_io_c_status_releaseThrough),
    .io_bstatus_set(abc_mshr_9_io_bstatus_set),
    .io_bstatus_tag(abc_mshr_9_io_bstatus_tag),
    .io_bstatus_way(abc_mshr_9_io_bstatus_way),
    .io_bstatus_nestedProbeAckData(abc_mshr_9_io_bstatus_nestedProbeAckData),
    .io_bstatus_probeHelperFinish(abc_mshr_9_io_bstatus_probeHelperFinish),
    .io_bstatus_probeAckDataThrough(abc_mshr_9_io_bstatus_probeAckDataThrough),
    .io_releaseThrough(abc_mshr_9_io_releaseThrough),
    .io_probeAckDataThrough(abc_mshr_9_io_probeAckDataThrough),
    .io_is_nestedReleaseData(abc_mshr_9_io_is_nestedReleaseData),
    .io_is_nestedProbeAckData(abc_mshr_9_io_is_nestedProbeAckData),
    .io_probeHelperFinish(abc_mshr_9_io_probeHelperFinish)
  );
  MSHR abc_mshr_10 ( // @[Slice.scala 94:16]
    .clock(abc_mshr_10_clock),
    .reset(abc_mshr_10_reset),
    .io_id(abc_mshr_10_io_id),
    .io_enable(abc_mshr_10_io_enable),
    .io_alloc_valid(abc_mshr_10_io_alloc_valid),
    .io_alloc_bits_channel(abc_mshr_10_io_alloc_bits_channel),
    .io_alloc_bits_opcode(abc_mshr_10_io_alloc_bits_opcode),
    .io_alloc_bits_param(abc_mshr_10_io_alloc_bits_param),
    .io_alloc_bits_size(abc_mshr_10_io_alloc_bits_size),
    .io_alloc_bits_source(abc_mshr_10_io_alloc_bits_source),
    .io_alloc_bits_set(abc_mshr_10_io_alloc_bits_set),
    .io_alloc_bits_tag(abc_mshr_10_io_alloc_bits_tag),
    .io_alloc_bits_off(abc_mshr_10_io_alloc_bits_off),
    .io_alloc_bits_mask(abc_mshr_10_io_alloc_bits_mask),
    .io_alloc_bits_bufIdx(abc_mshr_10_io_alloc_bits_bufIdx),
    .io_alloc_bits_preferCache(abc_mshr_10_io_alloc_bits_preferCache),
    .io_alloc_bits_dirty(abc_mshr_10_io_alloc_bits_dirty),
    .io_alloc_bits_fromProbeHelper(abc_mshr_10_io_alloc_bits_fromProbeHelper),
    .io_alloc_bits_fromCmoHelper(abc_mshr_10_io_alloc_bits_fromCmoHelper),
    .io_alloc_bits_needProbeAckData(abc_mshr_10_io_alloc_bits_needProbeAckData),
    .io_status_valid(abc_mshr_10_io_status_valid),
    .io_status_bits_set(abc_mshr_10_io_status_bits_set),
    .io_status_bits_tag(abc_mshr_10_io_status_bits_tag),
    .io_status_bits_way(abc_mshr_10_io_status_bits_way),
    .io_status_bits_way_reg(abc_mshr_10_io_status_bits_way_reg),
    .io_status_bits_nestB(abc_mshr_10_io_status_bits_nestB),
    .io_status_bits_nestC(abc_mshr_10_io_status_bits_nestC),
    .io_status_bits_will_grant_data(abc_mshr_10_io_status_bits_will_grant_data),
    .io_status_bits_will_save_data(abc_mshr_10_io_status_bits_will_save_data),
    .io_status_bits_will_free(abc_mshr_10_io_status_bits_will_free),
    .io_resps_sink_c_valid(abc_mshr_10_io_resps_sink_c_valid),
    .io_resps_sink_c_bits_hasData(abc_mshr_10_io_resps_sink_c_bits_hasData),
    .io_resps_sink_c_bits_param(abc_mshr_10_io_resps_sink_c_bits_param),
    .io_resps_sink_c_bits_source(abc_mshr_10_io_resps_sink_c_bits_source),
    .io_resps_sink_c_bits_last(abc_mshr_10_io_resps_sink_c_bits_last),
    .io_resps_sink_c_bits_bufIdx(abc_mshr_10_io_resps_sink_c_bits_bufIdx),
    .io_resps_sink_d_valid(abc_mshr_10_io_resps_sink_d_valid),
    .io_resps_sink_d_bits_opcode(abc_mshr_10_io_resps_sink_d_bits_opcode),
    .io_resps_sink_d_bits_param(abc_mshr_10_io_resps_sink_d_bits_param),
    .io_resps_sink_d_bits_sink(abc_mshr_10_io_resps_sink_d_bits_sink),
    .io_resps_sink_d_bits_last(abc_mshr_10_io_resps_sink_d_bits_last),
    .io_resps_sink_d_bits_denied(abc_mshr_10_io_resps_sink_d_bits_denied),
    .io_resps_sink_d_bits_bufIdx(abc_mshr_10_io_resps_sink_d_bits_bufIdx),
    .io_resps_sink_e_valid(abc_mshr_10_io_resps_sink_e_valid),
    .io_resps_source_d_valid(abc_mshr_10_io_resps_source_d_valid),
    .io_nestedwb_set(abc_mshr_10_io_nestedwb_set),
    .io_nestedwb_tag(abc_mshr_10_io_nestedwb_tag),
    .io_nestedwb_btoN(abc_mshr_10_io_nestedwb_btoN),
    .io_nestedwb_btoB(abc_mshr_10_io_nestedwb_btoB),
    .io_nestedwb_bclr_dirty(abc_mshr_10_io_nestedwb_bclr_dirty),
    .io_nestedwb_bset_dirty(abc_mshr_10_io_nestedwb_bset_dirty),
    .io_nestedwb_c_set_dirty(abc_mshr_10_io_nestedwb_c_set_dirty),
    .io_nestedwb_c_set_hit(abc_mshr_10_io_nestedwb_c_set_hit),
    .io_nestedwb_clients_0_isToN(abc_mshr_10_io_nestedwb_clients_0_isToN),
    .io_nestedwb_clients_1_isToN(abc_mshr_10_io_nestedwb_clients_1_isToN),
    .io_tasks_sink_a_ready(abc_mshr_10_io_tasks_sink_a_ready),
    .io_tasks_sink_a_valid(abc_mshr_10_io_tasks_sink_a_valid),
    .io_tasks_sink_a_bits_sourceId(abc_mshr_10_io_tasks_sink_a_bits_sourceId),
    .io_tasks_sink_a_bits_set(abc_mshr_10_io_tasks_sink_a_bits_set),
    .io_tasks_sink_a_bits_tag(abc_mshr_10_io_tasks_sink_a_bits_tag),
    .io_tasks_sink_a_bits_size(abc_mshr_10_io_tasks_sink_a_bits_size),
    .io_tasks_sink_a_bits_off(abc_mshr_10_io_tasks_sink_a_bits_off),
    .io_tasks_source_bready(abc_mshr_10_io_tasks_source_bready),
    .io_tasks_source_bvalid(abc_mshr_10_io_tasks_source_bvalid),
    .io_tasks_source_bset(abc_mshr_10_io_tasks_source_bset),
    .io_tasks_source_btag(abc_mshr_10_io_tasks_source_btag),
    .io_tasks_source_bparam(abc_mshr_10_io_tasks_source_bparam),
    .io_tasks_source_bclients(abc_mshr_10_io_tasks_source_bclients),
    .io_tasks_source_bneedData(abc_mshr_10_io_tasks_source_bneedData),
    .io_tasks_sink_c_ready(abc_mshr_10_io_tasks_sink_c_ready),
    .io_tasks_sink_c_valid(abc_mshr_10_io_tasks_sink_c_valid),
    .io_tasks_sink_c_bits_sourceId(abc_mshr_10_io_tasks_sink_c_bits_sourceId),
    .io_tasks_sink_c_bits_set(abc_mshr_10_io_tasks_sink_c_bits_set),
    .io_tasks_sink_c_bits_tag(abc_mshr_10_io_tasks_sink_c_bits_tag),
    .io_tasks_sink_c_bits_size(abc_mshr_10_io_tasks_sink_c_bits_size),
    .io_tasks_sink_c_bits_way(abc_mshr_10_io_tasks_sink_c_bits_way),
    .io_tasks_sink_c_bits_off(abc_mshr_10_io_tasks_sink_c_bits_off),
    .io_tasks_sink_c_bits_bufIdx(abc_mshr_10_io_tasks_sink_c_bits_bufIdx),
    .io_tasks_sink_c_bits_opcode(abc_mshr_10_io_tasks_sink_c_bits_opcode),
    .io_tasks_sink_c_bits_param(abc_mshr_10_io_tasks_sink_c_bits_param),
    .io_tasks_sink_c_bits_source(abc_mshr_10_io_tasks_sink_c_bits_source),
    .io_tasks_sink_c_bits_save(abc_mshr_10_io_tasks_sink_c_bits_save),
    .io_tasks_sink_c_bits_drop(abc_mshr_10_io_tasks_sink_c_bits_drop),
    .io_tasks_sink_c_bits_release(abc_mshr_10_io_tasks_sink_c_bits_release),
    .io_tasks_sink_c_bits_dirty(abc_mshr_10_io_tasks_sink_c_bits_dirty),
    .io_tasks_source_d_ready(abc_mshr_10_io_tasks_source_d_ready),
    .io_tasks_source_d_valid(abc_mshr_10_io_tasks_source_d_valid),
    .io_tasks_source_d_bits_sourceId(abc_mshr_10_io_tasks_source_d_bits_sourceId),
    .io_tasks_source_d_bits_set(abc_mshr_10_io_tasks_source_d_bits_set),
    .io_tasks_source_d_bits_tag(abc_mshr_10_io_tasks_source_d_bits_tag),
    .io_tasks_source_d_bits_channel(abc_mshr_10_io_tasks_source_d_bits_channel),
    .io_tasks_source_d_bits_opcode(abc_mshr_10_io_tasks_source_d_bits_opcode),
    .io_tasks_source_d_bits_param(abc_mshr_10_io_tasks_source_d_bits_param),
    .io_tasks_source_d_bits_size(abc_mshr_10_io_tasks_source_d_bits_size),
    .io_tasks_source_d_bits_way(abc_mshr_10_io_tasks_source_d_bits_way),
    .io_tasks_source_d_bits_off(abc_mshr_10_io_tasks_source_d_bits_off),
    .io_tasks_source_d_bits_useBypass(abc_mshr_10_io_tasks_source_d_bits_useBypass),
    .io_tasks_source_d_bits_bufIdx(abc_mshr_10_io_tasks_source_d_bits_bufIdx),
    .io_tasks_source_d_bits_denied(abc_mshr_10_io_tasks_source_d_bits_denied),
    .io_tasks_source_d_bits_sinkId(abc_mshr_10_io_tasks_source_d_bits_sinkId),
    .io_tasks_source_d_bits_bypassPut(abc_mshr_10_io_tasks_source_d_bits_bypassPut),
    .io_tasks_source_d_bits_dirty(abc_mshr_10_io_tasks_source_d_bits_dirty),
    .io_tasks_source_a_ready(abc_mshr_10_io_tasks_source_a_ready),
    .io_tasks_source_a_valid(abc_mshr_10_io_tasks_source_a_valid),
    .io_tasks_source_a_bits_tag(abc_mshr_10_io_tasks_source_a_bits_tag),
    .io_tasks_source_a_bits_set(abc_mshr_10_io_tasks_source_a_bits_set),
    .io_tasks_source_a_bits_off(abc_mshr_10_io_tasks_source_a_bits_off),
    .io_tasks_source_a_bits_mask(abc_mshr_10_io_tasks_source_a_bits_mask),
    .io_tasks_source_a_bits_opcode(abc_mshr_10_io_tasks_source_a_bits_opcode),
    .io_tasks_source_a_bits_param(abc_mshr_10_io_tasks_source_a_bits_param),
    .io_tasks_source_a_bits_source(abc_mshr_10_io_tasks_source_a_bits_source),
    .io_tasks_source_a_bits_bufIdx(abc_mshr_10_io_tasks_source_a_bits_bufIdx),
    .io_tasks_source_a_bits_size(abc_mshr_10_io_tasks_source_a_bits_size),
    .io_tasks_source_a_bits_needData(abc_mshr_10_io_tasks_source_a_bits_needData),
    .io_tasks_source_a_bits_putData(abc_mshr_10_io_tasks_source_a_bits_putData),
    .io_tasks_source_c_ready(abc_mshr_10_io_tasks_source_c_ready),
    .io_tasks_source_c_valid(abc_mshr_10_io_tasks_source_c_valid),
    .io_tasks_source_c_bits_opcode(abc_mshr_10_io_tasks_source_c_bits_opcode),
    .io_tasks_source_c_bits_tag(abc_mshr_10_io_tasks_source_c_bits_tag),
    .io_tasks_source_c_bits_set(abc_mshr_10_io_tasks_source_c_bits_set),
    .io_tasks_source_c_bits_param(abc_mshr_10_io_tasks_source_c_bits_param),
    .io_tasks_source_c_bits_source(abc_mshr_10_io_tasks_source_c_bits_source),
    .io_tasks_source_c_bits_way(abc_mshr_10_io_tasks_source_c_bits_way),
    .io_tasks_source_c_bits_dirty(abc_mshr_10_io_tasks_source_c_bits_dirty),
    .io_tasks_source_e_ready(abc_mshr_10_io_tasks_source_e_ready),
    .io_tasks_source_e_valid(abc_mshr_10_io_tasks_source_e_valid),
    .io_tasks_source_e_bits_sink(abc_mshr_10_io_tasks_source_e_bits_sink),
    .io_tasks_dir_write_ready(abc_mshr_10_io_tasks_dir_write_ready),
    .io_tasks_dir_write_valid(abc_mshr_10_io_tasks_dir_write_valid),
    .io_tasks_dir_write_bits_set(abc_mshr_10_io_tasks_dir_write_bits_set),
    .io_tasks_dir_write_bits_way(abc_mshr_10_io_tasks_dir_write_bits_way),
    .io_tasks_dir_write_bits_data_dirty(abc_mshr_10_io_tasks_dir_write_bits_data_dirty),
    .io_tasks_dir_write_bits_data_state(abc_mshr_10_io_tasks_dir_write_bits_data_state),
    .io_tasks_dir_write_bits_data_clientStates_0(abc_mshr_10_io_tasks_dir_write_bits_data_clientStates_0),
    .io_tasks_dir_write_bits_data_clientStates_1(abc_mshr_10_io_tasks_dir_write_bits_data_clientStates_1),
    .io_tasks_tag_write_ready(abc_mshr_10_io_tasks_tag_write_ready),
    .io_tasks_tag_write_valid(abc_mshr_10_io_tasks_tag_write_valid),
    .io_tasks_tag_write_bits_set(abc_mshr_10_io_tasks_tag_write_bits_set),
    .io_tasks_tag_write_bits_way(abc_mshr_10_io_tasks_tag_write_bits_way),
    .io_tasks_tag_write_bits_tag(abc_mshr_10_io_tasks_tag_write_bits_tag),
    .io_tasks_client_dir_write_ready(abc_mshr_10_io_tasks_client_dir_write_ready),
    .io_tasks_client_dir_write_valid(abc_mshr_10_io_tasks_client_dir_write_valid),
    .io_tasks_client_dir_write_bits_set(abc_mshr_10_io_tasks_client_dir_write_bits_set),
    .io_tasks_client_dir_write_bits_way(abc_mshr_10_io_tasks_client_dir_write_bits_way),
    .io_tasks_client_dir_write_bits_data_0_state(abc_mshr_10_io_tasks_client_dir_write_bits_data_0_state),
    .io_tasks_client_dir_write_bits_data_1_state(abc_mshr_10_io_tasks_client_dir_write_bits_data_1_state),
    .io_tasks_client_tag_write_ready(abc_mshr_10_io_tasks_client_tag_write_ready),
    .io_tasks_client_tag_write_valid(abc_mshr_10_io_tasks_client_tag_write_valid),
    .io_tasks_client_tag_write_bits_set(abc_mshr_10_io_tasks_client_tag_write_bits_set),
    .io_tasks_client_tag_write_bits_way(abc_mshr_10_io_tasks_client_tag_write_bits_way),
    .io_tasks_client_tag_write_bits_tag(abc_mshr_10_io_tasks_client_tag_write_bits_tag),
    .io_dirResult_valid(abc_mshr_10_io_dirResult_valid),
    .io_dirResult_bits_self_dirty(abc_mshr_10_io_dirResult_bits_self_dirty),
    .io_dirResult_bits_self_state(abc_mshr_10_io_dirResult_bits_self_state),
    .io_dirResult_bits_self_clientStates_0(abc_mshr_10_io_dirResult_bits_self_clientStates_0),
    .io_dirResult_bits_self_clientStates_1(abc_mshr_10_io_dirResult_bits_self_clientStates_1),
    .io_dirResult_bits_self_hit(abc_mshr_10_io_dirResult_bits_self_hit),
    .io_dirResult_bits_self_way(abc_mshr_10_io_dirResult_bits_self_way),
    .io_dirResult_bits_self_tag(abc_mshr_10_io_dirResult_bits_self_tag),
    .io_dirResult_bits_clients_states_0_state(abc_mshr_10_io_dirResult_bits_clients_states_0_state),
    .io_dirResult_bits_clients_states_0_hit(abc_mshr_10_io_dirResult_bits_clients_states_0_hit),
    .io_dirResult_bits_clients_states_1_state(abc_mshr_10_io_dirResult_bits_clients_states_1_state),
    .io_dirResult_bits_clients_states_1_hit(abc_mshr_10_io_dirResult_bits_clients_states_1_hit),
    .io_dirResult_bits_clients_tag(abc_mshr_10_io_dirResult_bits_clients_tag),
    .io_dirResult_bits_clients_way(abc_mshr_10_io_dirResult_bits_clients_way),
    .io_c_status_set(abc_mshr_10_io_c_status_set),
    .io_c_status_tag(abc_mshr_10_io_c_status_tag),
    .io_c_status_way(abc_mshr_10_io_c_status_way),
    .io_c_status_nestedReleaseData(abc_mshr_10_io_c_status_nestedReleaseData),
    .io_c_status_releaseThrough(abc_mshr_10_io_c_status_releaseThrough),
    .io_bstatus_set(abc_mshr_10_io_bstatus_set),
    .io_bstatus_tag(abc_mshr_10_io_bstatus_tag),
    .io_bstatus_way(abc_mshr_10_io_bstatus_way),
    .io_bstatus_nestedProbeAckData(abc_mshr_10_io_bstatus_nestedProbeAckData),
    .io_bstatus_probeHelperFinish(abc_mshr_10_io_bstatus_probeHelperFinish),
    .io_bstatus_probeAckDataThrough(abc_mshr_10_io_bstatus_probeAckDataThrough),
    .io_releaseThrough(abc_mshr_10_io_releaseThrough),
    .io_probeAckDataThrough(abc_mshr_10_io_probeAckDataThrough),
    .io_is_nestedReleaseData(abc_mshr_10_io_is_nestedReleaseData),
    .io_is_nestedProbeAckData(abc_mshr_10_io_is_nestedProbeAckData),
    .io_probeHelperFinish(abc_mshr_10_io_probeHelperFinish)
  );
  MSHR abc_mshr_11 ( // @[Slice.scala 94:16]
    .clock(abc_mshr_11_clock),
    .reset(abc_mshr_11_reset),
    .io_id(abc_mshr_11_io_id),
    .io_enable(abc_mshr_11_io_enable),
    .io_alloc_valid(abc_mshr_11_io_alloc_valid),
    .io_alloc_bits_channel(abc_mshr_11_io_alloc_bits_channel),
    .io_alloc_bits_opcode(abc_mshr_11_io_alloc_bits_opcode),
    .io_alloc_bits_param(abc_mshr_11_io_alloc_bits_param),
    .io_alloc_bits_size(abc_mshr_11_io_alloc_bits_size),
    .io_alloc_bits_source(abc_mshr_11_io_alloc_bits_source),
    .io_alloc_bits_set(abc_mshr_11_io_alloc_bits_set),
    .io_alloc_bits_tag(abc_mshr_11_io_alloc_bits_tag),
    .io_alloc_bits_off(abc_mshr_11_io_alloc_bits_off),
    .io_alloc_bits_mask(abc_mshr_11_io_alloc_bits_mask),
    .io_alloc_bits_bufIdx(abc_mshr_11_io_alloc_bits_bufIdx),
    .io_alloc_bits_preferCache(abc_mshr_11_io_alloc_bits_preferCache),
    .io_alloc_bits_dirty(abc_mshr_11_io_alloc_bits_dirty),
    .io_alloc_bits_fromProbeHelper(abc_mshr_11_io_alloc_bits_fromProbeHelper),
    .io_alloc_bits_fromCmoHelper(abc_mshr_11_io_alloc_bits_fromCmoHelper),
    .io_alloc_bits_needProbeAckData(abc_mshr_11_io_alloc_bits_needProbeAckData),
    .io_status_valid(abc_mshr_11_io_status_valid),
    .io_status_bits_set(abc_mshr_11_io_status_bits_set),
    .io_status_bits_tag(abc_mshr_11_io_status_bits_tag),
    .io_status_bits_way(abc_mshr_11_io_status_bits_way),
    .io_status_bits_way_reg(abc_mshr_11_io_status_bits_way_reg),
    .io_status_bits_nestB(abc_mshr_11_io_status_bits_nestB),
    .io_status_bits_nestC(abc_mshr_11_io_status_bits_nestC),
    .io_status_bits_will_grant_data(abc_mshr_11_io_status_bits_will_grant_data),
    .io_status_bits_will_save_data(abc_mshr_11_io_status_bits_will_save_data),
    .io_status_bits_will_free(abc_mshr_11_io_status_bits_will_free),
    .io_resps_sink_c_valid(abc_mshr_11_io_resps_sink_c_valid),
    .io_resps_sink_c_bits_hasData(abc_mshr_11_io_resps_sink_c_bits_hasData),
    .io_resps_sink_c_bits_param(abc_mshr_11_io_resps_sink_c_bits_param),
    .io_resps_sink_c_bits_source(abc_mshr_11_io_resps_sink_c_bits_source),
    .io_resps_sink_c_bits_last(abc_mshr_11_io_resps_sink_c_bits_last),
    .io_resps_sink_c_bits_bufIdx(abc_mshr_11_io_resps_sink_c_bits_bufIdx),
    .io_resps_sink_d_valid(abc_mshr_11_io_resps_sink_d_valid),
    .io_resps_sink_d_bits_opcode(abc_mshr_11_io_resps_sink_d_bits_opcode),
    .io_resps_sink_d_bits_param(abc_mshr_11_io_resps_sink_d_bits_param),
    .io_resps_sink_d_bits_sink(abc_mshr_11_io_resps_sink_d_bits_sink),
    .io_resps_sink_d_bits_last(abc_mshr_11_io_resps_sink_d_bits_last),
    .io_resps_sink_d_bits_denied(abc_mshr_11_io_resps_sink_d_bits_denied),
    .io_resps_sink_d_bits_bufIdx(abc_mshr_11_io_resps_sink_d_bits_bufIdx),
    .io_resps_sink_e_valid(abc_mshr_11_io_resps_sink_e_valid),
    .io_resps_source_d_valid(abc_mshr_11_io_resps_source_d_valid),
    .io_nestedwb_set(abc_mshr_11_io_nestedwb_set),
    .io_nestedwb_tag(abc_mshr_11_io_nestedwb_tag),
    .io_nestedwb_btoN(abc_mshr_11_io_nestedwb_btoN),
    .io_nestedwb_btoB(abc_mshr_11_io_nestedwb_btoB),
    .io_nestedwb_bclr_dirty(abc_mshr_11_io_nestedwb_bclr_dirty),
    .io_nestedwb_bset_dirty(abc_mshr_11_io_nestedwb_bset_dirty),
    .io_nestedwb_c_set_dirty(abc_mshr_11_io_nestedwb_c_set_dirty),
    .io_nestedwb_c_set_hit(abc_mshr_11_io_nestedwb_c_set_hit),
    .io_nestedwb_clients_0_isToN(abc_mshr_11_io_nestedwb_clients_0_isToN),
    .io_nestedwb_clients_1_isToN(abc_mshr_11_io_nestedwb_clients_1_isToN),
    .io_tasks_sink_a_ready(abc_mshr_11_io_tasks_sink_a_ready),
    .io_tasks_sink_a_valid(abc_mshr_11_io_tasks_sink_a_valid),
    .io_tasks_sink_a_bits_sourceId(abc_mshr_11_io_tasks_sink_a_bits_sourceId),
    .io_tasks_sink_a_bits_set(abc_mshr_11_io_tasks_sink_a_bits_set),
    .io_tasks_sink_a_bits_tag(abc_mshr_11_io_tasks_sink_a_bits_tag),
    .io_tasks_sink_a_bits_size(abc_mshr_11_io_tasks_sink_a_bits_size),
    .io_tasks_sink_a_bits_off(abc_mshr_11_io_tasks_sink_a_bits_off),
    .io_tasks_source_bready(abc_mshr_11_io_tasks_source_bready),
    .io_tasks_source_bvalid(abc_mshr_11_io_tasks_source_bvalid),
    .io_tasks_source_bset(abc_mshr_11_io_tasks_source_bset),
    .io_tasks_source_btag(abc_mshr_11_io_tasks_source_btag),
    .io_tasks_source_bparam(abc_mshr_11_io_tasks_source_bparam),
    .io_tasks_source_bclients(abc_mshr_11_io_tasks_source_bclients),
    .io_tasks_source_bneedData(abc_mshr_11_io_tasks_source_bneedData),
    .io_tasks_sink_c_ready(abc_mshr_11_io_tasks_sink_c_ready),
    .io_tasks_sink_c_valid(abc_mshr_11_io_tasks_sink_c_valid),
    .io_tasks_sink_c_bits_sourceId(abc_mshr_11_io_tasks_sink_c_bits_sourceId),
    .io_tasks_sink_c_bits_set(abc_mshr_11_io_tasks_sink_c_bits_set),
    .io_tasks_sink_c_bits_tag(abc_mshr_11_io_tasks_sink_c_bits_tag),
    .io_tasks_sink_c_bits_size(abc_mshr_11_io_tasks_sink_c_bits_size),
    .io_tasks_sink_c_bits_way(abc_mshr_11_io_tasks_sink_c_bits_way),
    .io_tasks_sink_c_bits_off(abc_mshr_11_io_tasks_sink_c_bits_off),
    .io_tasks_sink_c_bits_bufIdx(abc_mshr_11_io_tasks_sink_c_bits_bufIdx),
    .io_tasks_sink_c_bits_opcode(abc_mshr_11_io_tasks_sink_c_bits_opcode),
    .io_tasks_sink_c_bits_param(abc_mshr_11_io_tasks_sink_c_bits_param),
    .io_tasks_sink_c_bits_source(abc_mshr_11_io_tasks_sink_c_bits_source),
    .io_tasks_sink_c_bits_save(abc_mshr_11_io_tasks_sink_c_bits_save),
    .io_tasks_sink_c_bits_drop(abc_mshr_11_io_tasks_sink_c_bits_drop),
    .io_tasks_sink_c_bits_release(abc_mshr_11_io_tasks_sink_c_bits_release),
    .io_tasks_sink_c_bits_dirty(abc_mshr_11_io_tasks_sink_c_bits_dirty),
    .io_tasks_source_d_ready(abc_mshr_11_io_tasks_source_d_ready),
    .io_tasks_source_d_valid(abc_mshr_11_io_tasks_source_d_valid),
    .io_tasks_source_d_bits_sourceId(abc_mshr_11_io_tasks_source_d_bits_sourceId),
    .io_tasks_source_d_bits_set(abc_mshr_11_io_tasks_source_d_bits_set),
    .io_tasks_source_d_bits_tag(abc_mshr_11_io_tasks_source_d_bits_tag),
    .io_tasks_source_d_bits_channel(abc_mshr_11_io_tasks_source_d_bits_channel),
    .io_tasks_source_d_bits_opcode(abc_mshr_11_io_tasks_source_d_bits_opcode),
    .io_tasks_source_d_bits_param(abc_mshr_11_io_tasks_source_d_bits_param),
    .io_tasks_source_d_bits_size(abc_mshr_11_io_tasks_source_d_bits_size),
    .io_tasks_source_d_bits_way(abc_mshr_11_io_tasks_source_d_bits_way),
    .io_tasks_source_d_bits_off(abc_mshr_11_io_tasks_source_d_bits_off),
    .io_tasks_source_d_bits_useBypass(abc_mshr_11_io_tasks_source_d_bits_useBypass),
    .io_tasks_source_d_bits_bufIdx(abc_mshr_11_io_tasks_source_d_bits_bufIdx),
    .io_tasks_source_d_bits_denied(abc_mshr_11_io_tasks_source_d_bits_denied),
    .io_tasks_source_d_bits_sinkId(abc_mshr_11_io_tasks_source_d_bits_sinkId),
    .io_tasks_source_d_bits_bypassPut(abc_mshr_11_io_tasks_source_d_bits_bypassPut),
    .io_tasks_source_d_bits_dirty(abc_mshr_11_io_tasks_source_d_bits_dirty),
    .io_tasks_source_a_ready(abc_mshr_11_io_tasks_source_a_ready),
    .io_tasks_source_a_valid(abc_mshr_11_io_tasks_source_a_valid),
    .io_tasks_source_a_bits_tag(abc_mshr_11_io_tasks_source_a_bits_tag),
    .io_tasks_source_a_bits_set(abc_mshr_11_io_tasks_source_a_bits_set),
    .io_tasks_source_a_bits_off(abc_mshr_11_io_tasks_source_a_bits_off),
    .io_tasks_source_a_bits_mask(abc_mshr_11_io_tasks_source_a_bits_mask),
    .io_tasks_source_a_bits_opcode(abc_mshr_11_io_tasks_source_a_bits_opcode),
    .io_tasks_source_a_bits_param(abc_mshr_11_io_tasks_source_a_bits_param),
    .io_tasks_source_a_bits_source(abc_mshr_11_io_tasks_source_a_bits_source),
    .io_tasks_source_a_bits_bufIdx(abc_mshr_11_io_tasks_source_a_bits_bufIdx),
    .io_tasks_source_a_bits_size(abc_mshr_11_io_tasks_source_a_bits_size),
    .io_tasks_source_a_bits_needData(abc_mshr_11_io_tasks_source_a_bits_needData),
    .io_tasks_source_a_bits_putData(abc_mshr_11_io_tasks_source_a_bits_putData),
    .io_tasks_source_c_ready(abc_mshr_11_io_tasks_source_c_ready),
    .io_tasks_source_c_valid(abc_mshr_11_io_tasks_source_c_valid),
    .io_tasks_source_c_bits_opcode(abc_mshr_11_io_tasks_source_c_bits_opcode),
    .io_tasks_source_c_bits_tag(abc_mshr_11_io_tasks_source_c_bits_tag),
    .io_tasks_source_c_bits_set(abc_mshr_11_io_tasks_source_c_bits_set),
    .io_tasks_source_c_bits_param(abc_mshr_11_io_tasks_source_c_bits_param),
    .io_tasks_source_c_bits_source(abc_mshr_11_io_tasks_source_c_bits_source),
    .io_tasks_source_c_bits_way(abc_mshr_11_io_tasks_source_c_bits_way),
    .io_tasks_source_c_bits_dirty(abc_mshr_11_io_tasks_source_c_bits_dirty),
    .io_tasks_source_e_ready(abc_mshr_11_io_tasks_source_e_ready),
    .io_tasks_source_e_valid(abc_mshr_11_io_tasks_source_e_valid),
    .io_tasks_source_e_bits_sink(abc_mshr_11_io_tasks_source_e_bits_sink),
    .io_tasks_dir_write_ready(abc_mshr_11_io_tasks_dir_write_ready),
    .io_tasks_dir_write_valid(abc_mshr_11_io_tasks_dir_write_valid),
    .io_tasks_dir_write_bits_set(abc_mshr_11_io_tasks_dir_write_bits_set),
    .io_tasks_dir_write_bits_way(abc_mshr_11_io_tasks_dir_write_bits_way),
    .io_tasks_dir_write_bits_data_dirty(abc_mshr_11_io_tasks_dir_write_bits_data_dirty),
    .io_tasks_dir_write_bits_data_state(abc_mshr_11_io_tasks_dir_write_bits_data_state),
    .io_tasks_dir_write_bits_data_clientStates_0(abc_mshr_11_io_tasks_dir_write_bits_data_clientStates_0),
    .io_tasks_dir_write_bits_data_clientStates_1(abc_mshr_11_io_tasks_dir_write_bits_data_clientStates_1),
    .io_tasks_tag_write_ready(abc_mshr_11_io_tasks_tag_write_ready),
    .io_tasks_tag_write_valid(abc_mshr_11_io_tasks_tag_write_valid),
    .io_tasks_tag_write_bits_set(abc_mshr_11_io_tasks_tag_write_bits_set),
    .io_tasks_tag_write_bits_way(abc_mshr_11_io_tasks_tag_write_bits_way),
    .io_tasks_tag_write_bits_tag(abc_mshr_11_io_tasks_tag_write_bits_tag),
    .io_tasks_client_dir_write_ready(abc_mshr_11_io_tasks_client_dir_write_ready),
    .io_tasks_client_dir_write_valid(abc_mshr_11_io_tasks_client_dir_write_valid),
    .io_tasks_client_dir_write_bits_set(abc_mshr_11_io_tasks_client_dir_write_bits_set),
    .io_tasks_client_dir_write_bits_way(abc_mshr_11_io_tasks_client_dir_write_bits_way),
    .io_tasks_client_dir_write_bits_data_0_state(abc_mshr_11_io_tasks_client_dir_write_bits_data_0_state),
    .io_tasks_client_dir_write_bits_data_1_state(abc_mshr_11_io_tasks_client_dir_write_bits_data_1_state),
    .io_tasks_client_tag_write_ready(abc_mshr_11_io_tasks_client_tag_write_ready),
    .io_tasks_client_tag_write_valid(abc_mshr_11_io_tasks_client_tag_write_valid),
    .io_tasks_client_tag_write_bits_set(abc_mshr_11_io_tasks_client_tag_write_bits_set),
    .io_tasks_client_tag_write_bits_way(abc_mshr_11_io_tasks_client_tag_write_bits_way),
    .io_tasks_client_tag_write_bits_tag(abc_mshr_11_io_tasks_client_tag_write_bits_tag),
    .io_dirResult_valid(abc_mshr_11_io_dirResult_valid),
    .io_dirResult_bits_self_dirty(abc_mshr_11_io_dirResult_bits_self_dirty),
    .io_dirResult_bits_self_state(abc_mshr_11_io_dirResult_bits_self_state),
    .io_dirResult_bits_self_clientStates_0(abc_mshr_11_io_dirResult_bits_self_clientStates_0),
    .io_dirResult_bits_self_clientStates_1(abc_mshr_11_io_dirResult_bits_self_clientStates_1),
    .io_dirResult_bits_self_hit(abc_mshr_11_io_dirResult_bits_self_hit),
    .io_dirResult_bits_self_way(abc_mshr_11_io_dirResult_bits_self_way),
    .io_dirResult_bits_self_tag(abc_mshr_11_io_dirResult_bits_self_tag),
    .io_dirResult_bits_clients_states_0_state(abc_mshr_11_io_dirResult_bits_clients_states_0_state),
    .io_dirResult_bits_clients_states_0_hit(abc_mshr_11_io_dirResult_bits_clients_states_0_hit),
    .io_dirResult_bits_clients_states_1_state(abc_mshr_11_io_dirResult_bits_clients_states_1_state),
    .io_dirResult_bits_clients_states_1_hit(abc_mshr_11_io_dirResult_bits_clients_states_1_hit),
    .io_dirResult_bits_clients_tag(abc_mshr_11_io_dirResult_bits_clients_tag),
    .io_dirResult_bits_clients_way(abc_mshr_11_io_dirResult_bits_clients_way),
    .io_c_status_set(abc_mshr_11_io_c_status_set),
    .io_c_status_tag(abc_mshr_11_io_c_status_tag),
    .io_c_status_way(abc_mshr_11_io_c_status_way),
    .io_c_status_nestedReleaseData(abc_mshr_11_io_c_status_nestedReleaseData),
    .io_c_status_releaseThrough(abc_mshr_11_io_c_status_releaseThrough),
    .io_bstatus_set(abc_mshr_11_io_bstatus_set),
    .io_bstatus_tag(abc_mshr_11_io_bstatus_tag),
    .io_bstatus_way(abc_mshr_11_io_bstatus_way),
    .io_bstatus_nestedProbeAckData(abc_mshr_11_io_bstatus_nestedProbeAckData),
    .io_bstatus_probeHelperFinish(abc_mshr_11_io_bstatus_probeHelperFinish),
    .io_bstatus_probeAckDataThrough(abc_mshr_11_io_bstatus_probeAckDataThrough),
    .io_releaseThrough(abc_mshr_11_io_releaseThrough),
    .io_probeAckDataThrough(abc_mshr_11_io_probeAckDataThrough),
    .io_is_nestedReleaseData(abc_mshr_11_io_is_nestedReleaseData),
    .io_is_nestedProbeAckData(abc_mshr_11_io_is_nestedProbeAckData),
    .io_probeHelperFinish(abc_mshr_11_io_probeHelperFinish)
  );
  MSHR abc_mshr_12 ( // @[Slice.scala 94:16]
    .clock(abc_mshr_12_clock),
    .reset(abc_mshr_12_reset),
    .io_id(abc_mshr_12_io_id),
    .io_enable(abc_mshr_12_io_enable),
    .io_alloc_valid(abc_mshr_12_io_alloc_valid),
    .io_alloc_bits_channel(abc_mshr_12_io_alloc_bits_channel),
    .io_alloc_bits_opcode(abc_mshr_12_io_alloc_bits_opcode),
    .io_alloc_bits_param(abc_mshr_12_io_alloc_bits_param),
    .io_alloc_bits_size(abc_mshr_12_io_alloc_bits_size),
    .io_alloc_bits_source(abc_mshr_12_io_alloc_bits_source),
    .io_alloc_bits_set(abc_mshr_12_io_alloc_bits_set),
    .io_alloc_bits_tag(abc_mshr_12_io_alloc_bits_tag),
    .io_alloc_bits_off(abc_mshr_12_io_alloc_bits_off),
    .io_alloc_bits_mask(abc_mshr_12_io_alloc_bits_mask),
    .io_alloc_bits_bufIdx(abc_mshr_12_io_alloc_bits_bufIdx),
    .io_alloc_bits_preferCache(abc_mshr_12_io_alloc_bits_preferCache),
    .io_alloc_bits_dirty(abc_mshr_12_io_alloc_bits_dirty),
    .io_alloc_bits_fromProbeHelper(abc_mshr_12_io_alloc_bits_fromProbeHelper),
    .io_alloc_bits_fromCmoHelper(abc_mshr_12_io_alloc_bits_fromCmoHelper),
    .io_alloc_bits_needProbeAckData(abc_mshr_12_io_alloc_bits_needProbeAckData),
    .io_status_valid(abc_mshr_12_io_status_valid),
    .io_status_bits_set(abc_mshr_12_io_status_bits_set),
    .io_status_bits_tag(abc_mshr_12_io_status_bits_tag),
    .io_status_bits_way(abc_mshr_12_io_status_bits_way),
    .io_status_bits_way_reg(abc_mshr_12_io_status_bits_way_reg),
    .io_status_bits_nestB(abc_mshr_12_io_status_bits_nestB),
    .io_status_bits_nestC(abc_mshr_12_io_status_bits_nestC),
    .io_status_bits_will_grant_data(abc_mshr_12_io_status_bits_will_grant_data),
    .io_status_bits_will_save_data(abc_mshr_12_io_status_bits_will_save_data),
    .io_status_bits_will_free(abc_mshr_12_io_status_bits_will_free),
    .io_resps_sink_c_valid(abc_mshr_12_io_resps_sink_c_valid),
    .io_resps_sink_c_bits_hasData(abc_mshr_12_io_resps_sink_c_bits_hasData),
    .io_resps_sink_c_bits_param(abc_mshr_12_io_resps_sink_c_bits_param),
    .io_resps_sink_c_bits_source(abc_mshr_12_io_resps_sink_c_bits_source),
    .io_resps_sink_c_bits_last(abc_mshr_12_io_resps_sink_c_bits_last),
    .io_resps_sink_c_bits_bufIdx(abc_mshr_12_io_resps_sink_c_bits_bufIdx),
    .io_resps_sink_d_valid(abc_mshr_12_io_resps_sink_d_valid),
    .io_resps_sink_d_bits_opcode(abc_mshr_12_io_resps_sink_d_bits_opcode),
    .io_resps_sink_d_bits_param(abc_mshr_12_io_resps_sink_d_bits_param),
    .io_resps_sink_d_bits_sink(abc_mshr_12_io_resps_sink_d_bits_sink),
    .io_resps_sink_d_bits_last(abc_mshr_12_io_resps_sink_d_bits_last),
    .io_resps_sink_d_bits_denied(abc_mshr_12_io_resps_sink_d_bits_denied),
    .io_resps_sink_d_bits_bufIdx(abc_mshr_12_io_resps_sink_d_bits_bufIdx),
    .io_resps_sink_e_valid(abc_mshr_12_io_resps_sink_e_valid),
    .io_resps_source_d_valid(abc_mshr_12_io_resps_source_d_valid),
    .io_nestedwb_set(abc_mshr_12_io_nestedwb_set),
    .io_nestedwb_tag(abc_mshr_12_io_nestedwb_tag),
    .io_nestedwb_btoN(abc_mshr_12_io_nestedwb_btoN),
    .io_nestedwb_btoB(abc_mshr_12_io_nestedwb_btoB),
    .io_nestedwb_bclr_dirty(abc_mshr_12_io_nestedwb_bclr_dirty),
    .io_nestedwb_bset_dirty(abc_mshr_12_io_nestedwb_bset_dirty),
    .io_nestedwb_c_set_dirty(abc_mshr_12_io_nestedwb_c_set_dirty),
    .io_nestedwb_c_set_hit(abc_mshr_12_io_nestedwb_c_set_hit),
    .io_nestedwb_clients_0_isToN(abc_mshr_12_io_nestedwb_clients_0_isToN),
    .io_nestedwb_clients_1_isToN(abc_mshr_12_io_nestedwb_clients_1_isToN),
    .io_tasks_sink_a_ready(abc_mshr_12_io_tasks_sink_a_ready),
    .io_tasks_sink_a_valid(abc_mshr_12_io_tasks_sink_a_valid),
    .io_tasks_sink_a_bits_sourceId(abc_mshr_12_io_tasks_sink_a_bits_sourceId),
    .io_tasks_sink_a_bits_set(abc_mshr_12_io_tasks_sink_a_bits_set),
    .io_tasks_sink_a_bits_tag(abc_mshr_12_io_tasks_sink_a_bits_tag),
    .io_tasks_sink_a_bits_size(abc_mshr_12_io_tasks_sink_a_bits_size),
    .io_tasks_sink_a_bits_off(abc_mshr_12_io_tasks_sink_a_bits_off),
    .io_tasks_source_bready(abc_mshr_12_io_tasks_source_bready),
    .io_tasks_source_bvalid(abc_mshr_12_io_tasks_source_bvalid),
    .io_tasks_source_bset(abc_mshr_12_io_tasks_source_bset),
    .io_tasks_source_btag(abc_mshr_12_io_tasks_source_btag),
    .io_tasks_source_bparam(abc_mshr_12_io_tasks_source_bparam),
    .io_tasks_source_bclients(abc_mshr_12_io_tasks_source_bclients),
    .io_tasks_source_bneedData(abc_mshr_12_io_tasks_source_bneedData),
    .io_tasks_sink_c_ready(abc_mshr_12_io_tasks_sink_c_ready),
    .io_tasks_sink_c_valid(abc_mshr_12_io_tasks_sink_c_valid),
    .io_tasks_sink_c_bits_sourceId(abc_mshr_12_io_tasks_sink_c_bits_sourceId),
    .io_tasks_sink_c_bits_set(abc_mshr_12_io_tasks_sink_c_bits_set),
    .io_tasks_sink_c_bits_tag(abc_mshr_12_io_tasks_sink_c_bits_tag),
    .io_tasks_sink_c_bits_size(abc_mshr_12_io_tasks_sink_c_bits_size),
    .io_tasks_sink_c_bits_way(abc_mshr_12_io_tasks_sink_c_bits_way),
    .io_tasks_sink_c_bits_off(abc_mshr_12_io_tasks_sink_c_bits_off),
    .io_tasks_sink_c_bits_bufIdx(abc_mshr_12_io_tasks_sink_c_bits_bufIdx),
    .io_tasks_sink_c_bits_opcode(abc_mshr_12_io_tasks_sink_c_bits_opcode),
    .io_tasks_sink_c_bits_param(abc_mshr_12_io_tasks_sink_c_bits_param),
    .io_tasks_sink_c_bits_source(abc_mshr_12_io_tasks_sink_c_bits_source),
    .io_tasks_sink_c_bits_save(abc_mshr_12_io_tasks_sink_c_bits_save),
    .io_tasks_sink_c_bits_drop(abc_mshr_12_io_tasks_sink_c_bits_drop),
    .io_tasks_sink_c_bits_release(abc_mshr_12_io_tasks_sink_c_bits_release),
    .io_tasks_sink_c_bits_dirty(abc_mshr_12_io_tasks_sink_c_bits_dirty),
    .io_tasks_source_d_ready(abc_mshr_12_io_tasks_source_d_ready),
    .io_tasks_source_d_valid(abc_mshr_12_io_tasks_source_d_valid),
    .io_tasks_source_d_bits_sourceId(abc_mshr_12_io_tasks_source_d_bits_sourceId),
    .io_tasks_source_d_bits_set(abc_mshr_12_io_tasks_source_d_bits_set),
    .io_tasks_source_d_bits_tag(abc_mshr_12_io_tasks_source_d_bits_tag),
    .io_tasks_source_d_bits_channel(abc_mshr_12_io_tasks_source_d_bits_channel),
    .io_tasks_source_d_bits_opcode(abc_mshr_12_io_tasks_source_d_bits_opcode),
    .io_tasks_source_d_bits_param(abc_mshr_12_io_tasks_source_d_bits_param),
    .io_tasks_source_d_bits_size(abc_mshr_12_io_tasks_source_d_bits_size),
    .io_tasks_source_d_bits_way(abc_mshr_12_io_tasks_source_d_bits_way),
    .io_tasks_source_d_bits_off(abc_mshr_12_io_tasks_source_d_bits_off),
    .io_tasks_source_d_bits_useBypass(abc_mshr_12_io_tasks_source_d_bits_useBypass),
    .io_tasks_source_d_bits_bufIdx(abc_mshr_12_io_tasks_source_d_bits_bufIdx),
    .io_tasks_source_d_bits_denied(abc_mshr_12_io_tasks_source_d_bits_denied),
    .io_tasks_source_d_bits_sinkId(abc_mshr_12_io_tasks_source_d_bits_sinkId),
    .io_tasks_source_d_bits_bypassPut(abc_mshr_12_io_tasks_source_d_bits_bypassPut),
    .io_tasks_source_d_bits_dirty(abc_mshr_12_io_tasks_source_d_bits_dirty),
    .io_tasks_source_a_ready(abc_mshr_12_io_tasks_source_a_ready),
    .io_tasks_source_a_valid(abc_mshr_12_io_tasks_source_a_valid),
    .io_tasks_source_a_bits_tag(abc_mshr_12_io_tasks_source_a_bits_tag),
    .io_tasks_source_a_bits_set(abc_mshr_12_io_tasks_source_a_bits_set),
    .io_tasks_source_a_bits_off(abc_mshr_12_io_tasks_source_a_bits_off),
    .io_tasks_source_a_bits_mask(abc_mshr_12_io_tasks_source_a_bits_mask),
    .io_tasks_source_a_bits_opcode(abc_mshr_12_io_tasks_source_a_bits_opcode),
    .io_tasks_source_a_bits_param(abc_mshr_12_io_tasks_source_a_bits_param),
    .io_tasks_source_a_bits_source(abc_mshr_12_io_tasks_source_a_bits_source),
    .io_tasks_source_a_bits_bufIdx(abc_mshr_12_io_tasks_source_a_bits_bufIdx),
    .io_tasks_source_a_bits_size(abc_mshr_12_io_tasks_source_a_bits_size),
    .io_tasks_source_a_bits_needData(abc_mshr_12_io_tasks_source_a_bits_needData),
    .io_tasks_source_a_bits_putData(abc_mshr_12_io_tasks_source_a_bits_putData),
    .io_tasks_source_c_ready(abc_mshr_12_io_tasks_source_c_ready),
    .io_tasks_source_c_valid(abc_mshr_12_io_tasks_source_c_valid),
    .io_tasks_source_c_bits_opcode(abc_mshr_12_io_tasks_source_c_bits_opcode),
    .io_tasks_source_c_bits_tag(abc_mshr_12_io_tasks_source_c_bits_tag),
    .io_tasks_source_c_bits_set(abc_mshr_12_io_tasks_source_c_bits_set),
    .io_tasks_source_c_bits_param(abc_mshr_12_io_tasks_source_c_bits_param),
    .io_tasks_source_c_bits_source(abc_mshr_12_io_tasks_source_c_bits_source),
    .io_tasks_source_c_bits_way(abc_mshr_12_io_tasks_source_c_bits_way),
    .io_tasks_source_c_bits_dirty(abc_mshr_12_io_tasks_source_c_bits_dirty),
    .io_tasks_source_e_ready(abc_mshr_12_io_tasks_source_e_ready),
    .io_tasks_source_e_valid(abc_mshr_12_io_tasks_source_e_valid),
    .io_tasks_source_e_bits_sink(abc_mshr_12_io_tasks_source_e_bits_sink),
    .io_tasks_dir_write_ready(abc_mshr_12_io_tasks_dir_write_ready),
    .io_tasks_dir_write_valid(abc_mshr_12_io_tasks_dir_write_valid),
    .io_tasks_dir_write_bits_set(abc_mshr_12_io_tasks_dir_write_bits_set),
    .io_tasks_dir_write_bits_way(abc_mshr_12_io_tasks_dir_write_bits_way),
    .io_tasks_dir_write_bits_data_dirty(abc_mshr_12_io_tasks_dir_write_bits_data_dirty),
    .io_tasks_dir_write_bits_data_state(abc_mshr_12_io_tasks_dir_write_bits_data_state),
    .io_tasks_dir_write_bits_data_clientStates_0(abc_mshr_12_io_tasks_dir_write_bits_data_clientStates_0),
    .io_tasks_dir_write_bits_data_clientStates_1(abc_mshr_12_io_tasks_dir_write_bits_data_clientStates_1),
    .io_tasks_tag_write_ready(abc_mshr_12_io_tasks_tag_write_ready),
    .io_tasks_tag_write_valid(abc_mshr_12_io_tasks_tag_write_valid),
    .io_tasks_tag_write_bits_set(abc_mshr_12_io_tasks_tag_write_bits_set),
    .io_tasks_tag_write_bits_way(abc_mshr_12_io_tasks_tag_write_bits_way),
    .io_tasks_tag_write_bits_tag(abc_mshr_12_io_tasks_tag_write_bits_tag),
    .io_tasks_client_dir_write_ready(abc_mshr_12_io_tasks_client_dir_write_ready),
    .io_tasks_client_dir_write_valid(abc_mshr_12_io_tasks_client_dir_write_valid),
    .io_tasks_client_dir_write_bits_set(abc_mshr_12_io_tasks_client_dir_write_bits_set),
    .io_tasks_client_dir_write_bits_way(abc_mshr_12_io_tasks_client_dir_write_bits_way),
    .io_tasks_client_dir_write_bits_data_0_state(abc_mshr_12_io_tasks_client_dir_write_bits_data_0_state),
    .io_tasks_client_dir_write_bits_data_1_state(abc_mshr_12_io_tasks_client_dir_write_bits_data_1_state),
    .io_tasks_client_tag_write_ready(abc_mshr_12_io_tasks_client_tag_write_ready),
    .io_tasks_client_tag_write_valid(abc_mshr_12_io_tasks_client_tag_write_valid),
    .io_tasks_client_tag_write_bits_set(abc_mshr_12_io_tasks_client_tag_write_bits_set),
    .io_tasks_client_tag_write_bits_way(abc_mshr_12_io_tasks_client_tag_write_bits_way),
    .io_tasks_client_tag_write_bits_tag(abc_mshr_12_io_tasks_client_tag_write_bits_tag),
    .io_dirResult_valid(abc_mshr_12_io_dirResult_valid),
    .io_dirResult_bits_self_dirty(abc_mshr_12_io_dirResult_bits_self_dirty),
    .io_dirResult_bits_self_state(abc_mshr_12_io_dirResult_bits_self_state),
    .io_dirResult_bits_self_clientStates_0(abc_mshr_12_io_dirResult_bits_self_clientStates_0),
    .io_dirResult_bits_self_clientStates_1(abc_mshr_12_io_dirResult_bits_self_clientStates_1),
    .io_dirResult_bits_self_hit(abc_mshr_12_io_dirResult_bits_self_hit),
    .io_dirResult_bits_self_way(abc_mshr_12_io_dirResult_bits_self_way),
    .io_dirResult_bits_self_tag(abc_mshr_12_io_dirResult_bits_self_tag),
    .io_dirResult_bits_clients_states_0_state(abc_mshr_12_io_dirResult_bits_clients_states_0_state),
    .io_dirResult_bits_clients_states_0_hit(abc_mshr_12_io_dirResult_bits_clients_states_0_hit),
    .io_dirResult_bits_clients_states_1_state(abc_mshr_12_io_dirResult_bits_clients_states_1_state),
    .io_dirResult_bits_clients_states_1_hit(abc_mshr_12_io_dirResult_bits_clients_states_1_hit),
    .io_dirResult_bits_clients_tag(abc_mshr_12_io_dirResult_bits_clients_tag),
    .io_dirResult_bits_clients_way(abc_mshr_12_io_dirResult_bits_clients_way),
    .io_c_status_set(abc_mshr_12_io_c_status_set),
    .io_c_status_tag(abc_mshr_12_io_c_status_tag),
    .io_c_status_way(abc_mshr_12_io_c_status_way),
    .io_c_status_nestedReleaseData(abc_mshr_12_io_c_status_nestedReleaseData),
    .io_c_status_releaseThrough(abc_mshr_12_io_c_status_releaseThrough),
    .io_bstatus_set(abc_mshr_12_io_bstatus_set),
    .io_bstatus_tag(abc_mshr_12_io_bstatus_tag),
    .io_bstatus_way(abc_mshr_12_io_bstatus_way),
    .io_bstatus_nestedProbeAckData(abc_mshr_12_io_bstatus_nestedProbeAckData),
    .io_bstatus_probeHelperFinish(abc_mshr_12_io_bstatus_probeHelperFinish),
    .io_bstatus_probeAckDataThrough(abc_mshr_12_io_bstatus_probeAckDataThrough),
    .io_releaseThrough(abc_mshr_12_io_releaseThrough),
    .io_probeAckDataThrough(abc_mshr_12_io_probeAckDataThrough),
    .io_is_nestedReleaseData(abc_mshr_12_io_is_nestedReleaseData),
    .io_is_nestedProbeAckData(abc_mshr_12_io_is_nestedProbeAckData),
    .io_probeHelperFinish(abc_mshr_12_io_probeHelperFinish)
  );
  MSHR abc_mshr_13 ( // @[Slice.scala 94:16]
    .clock(abc_mshr_13_clock),
    .reset(abc_mshr_13_reset),
    .io_id(abc_mshr_13_io_id),
    .io_enable(abc_mshr_13_io_enable),
    .io_alloc_valid(abc_mshr_13_io_alloc_valid),
    .io_alloc_bits_channel(abc_mshr_13_io_alloc_bits_channel),
    .io_alloc_bits_opcode(abc_mshr_13_io_alloc_bits_opcode),
    .io_alloc_bits_param(abc_mshr_13_io_alloc_bits_param),
    .io_alloc_bits_size(abc_mshr_13_io_alloc_bits_size),
    .io_alloc_bits_source(abc_mshr_13_io_alloc_bits_source),
    .io_alloc_bits_set(abc_mshr_13_io_alloc_bits_set),
    .io_alloc_bits_tag(abc_mshr_13_io_alloc_bits_tag),
    .io_alloc_bits_off(abc_mshr_13_io_alloc_bits_off),
    .io_alloc_bits_mask(abc_mshr_13_io_alloc_bits_mask),
    .io_alloc_bits_bufIdx(abc_mshr_13_io_alloc_bits_bufIdx),
    .io_alloc_bits_preferCache(abc_mshr_13_io_alloc_bits_preferCache),
    .io_alloc_bits_dirty(abc_mshr_13_io_alloc_bits_dirty),
    .io_alloc_bits_fromProbeHelper(abc_mshr_13_io_alloc_bits_fromProbeHelper),
    .io_alloc_bits_fromCmoHelper(abc_mshr_13_io_alloc_bits_fromCmoHelper),
    .io_alloc_bits_needProbeAckData(abc_mshr_13_io_alloc_bits_needProbeAckData),
    .io_status_valid(abc_mshr_13_io_status_valid),
    .io_status_bits_set(abc_mshr_13_io_status_bits_set),
    .io_status_bits_tag(abc_mshr_13_io_status_bits_tag),
    .io_status_bits_way(abc_mshr_13_io_status_bits_way),
    .io_status_bits_way_reg(abc_mshr_13_io_status_bits_way_reg),
    .io_status_bits_nestB(abc_mshr_13_io_status_bits_nestB),
    .io_status_bits_nestC(abc_mshr_13_io_status_bits_nestC),
    .io_status_bits_will_grant_data(abc_mshr_13_io_status_bits_will_grant_data),
    .io_status_bits_will_save_data(abc_mshr_13_io_status_bits_will_save_data),
    .io_status_bits_will_free(abc_mshr_13_io_status_bits_will_free),
    .io_resps_sink_c_valid(abc_mshr_13_io_resps_sink_c_valid),
    .io_resps_sink_c_bits_hasData(abc_mshr_13_io_resps_sink_c_bits_hasData),
    .io_resps_sink_c_bits_param(abc_mshr_13_io_resps_sink_c_bits_param),
    .io_resps_sink_c_bits_source(abc_mshr_13_io_resps_sink_c_bits_source),
    .io_resps_sink_c_bits_last(abc_mshr_13_io_resps_sink_c_bits_last),
    .io_resps_sink_c_bits_bufIdx(abc_mshr_13_io_resps_sink_c_bits_bufIdx),
    .io_resps_sink_d_valid(abc_mshr_13_io_resps_sink_d_valid),
    .io_resps_sink_d_bits_opcode(abc_mshr_13_io_resps_sink_d_bits_opcode),
    .io_resps_sink_d_bits_param(abc_mshr_13_io_resps_sink_d_bits_param),
    .io_resps_sink_d_bits_sink(abc_mshr_13_io_resps_sink_d_bits_sink),
    .io_resps_sink_d_bits_last(abc_mshr_13_io_resps_sink_d_bits_last),
    .io_resps_sink_d_bits_denied(abc_mshr_13_io_resps_sink_d_bits_denied),
    .io_resps_sink_d_bits_bufIdx(abc_mshr_13_io_resps_sink_d_bits_bufIdx),
    .io_resps_sink_e_valid(abc_mshr_13_io_resps_sink_e_valid),
    .io_resps_source_d_valid(abc_mshr_13_io_resps_source_d_valid),
    .io_nestedwb_set(abc_mshr_13_io_nestedwb_set),
    .io_nestedwb_tag(abc_mshr_13_io_nestedwb_tag),
    .io_nestedwb_btoN(abc_mshr_13_io_nestedwb_btoN),
    .io_nestedwb_btoB(abc_mshr_13_io_nestedwb_btoB),
    .io_nestedwb_bclr_dirty(abc_mshr_13_io_nestedwb_bclr_dirty),
    .io_nestedwb_bset_dirty(abc_mshr_13_io_nestedwb_bset_dirty),
    .io_nestedwb_c_set_dirty(abc_mshr_13_io_nestedwb_c_set_dirty),
    .io_nestedwb_c_set_hit(abc_mshr_13_io_nestedwb_c_set_hit),
    .io_nestedwb_clients_0_isToN(abc_mshr_13_io_nestedwb_clients_0_isToN),
    .io_nestedwb_clients_1_isToN(abc_mshr_13_io_nestedwb_clients_1_isToN),
    .io_tasks_sink_a_ready(abc_mshr_13_io_tasks_sink_a_ready),
    .io_tasks_sink_a_valid(abc_mshr_13_io_tasks_sink_a_valid),
    .io_tasks_sink_a_bits_sourceId(abc_mshr_13_io_tasks_sink_a_bits_sourceId),
    .io_tasks_sink_a_bits_set(abc_mshr_13_io_tasks_sink_a_bits_set),
    .io_tasks_sink_a_bits_tag(abc_mshr_13_io_tasks_sink_a_bits_tag),
    .io_tasks_sink_a_bits_size(abc_mshr_13_io_tasks_sink_a_bits_size),
    .io_tasks_sink_a_bits_off(abc_mshr_13_io_tasks_sink_a_bits_off),
    .io_tasks_source_bready(abc_mshr_13_io_tasks_source_bready),
    .io_tasks_source_bvalid(abc_mshr_13_io_tasks_source_bvalid),
    .io_tasks_source_bset(abc_mshr_13_io_tasks_source_bset),
    .io_tasks_source_btag(abc_mshr_13_io_tasks_source_btag),
    .io_tasks_source_bparam(abc_mshr_13_io_tasks_source_bparam),
    .io_tasks_source_bclients(abc_mshr_13_io_tasks_source_bclients),
    .io_tasks_source_bneedData(abc_mshr_13_io_tasks_source_bneedData),
    .io_tasks_sink_c_ready(abc_mshr_13_io_tasks_sink_c_ready),
    .io_tasks_sink_c_valid(abc_mshr_13_io_tasks_sink_c_valid),
    .io_tasks_sink_c_bits_sourceId(abc_mshr_13_io_tasks_sink_c_bits_sourceId),
    .io_tasks_sink_c_bits_set(abc_mshr_13_io_tasks_sink_c_bits_set),
    .io_tasks_sink_c_bits_tag(abc_mshr_13_io_tasks_sink_c_bits_tag),
    .io_tasks_sink_c_bits_size(abc_mshr_13_io_tasks_sink_c_bits_size),
    .io_tasks_sink_c_bits_way(abc_mshr_13_io_tasks_sink_c_bits_way),
    .io_tasks_sink_c_bits_off(abc_mshr_13_io_tasks_sink_c_bits_off),
    .io_tasks_sink_c_bits_bufIdx(abc_mshr_13_io_tasks_sink_c_bits_bufIdx),
    .io_tasks_sink_c_bits_opcode(abc_mshr_13_io_tasks_sink_c_bits_opcode),
    .io_tasks_sink_c_bits_param(abc_mshr_13_io_tasks_sink_c_bits_param),
    .io_tasks_sink_c_bits_source(abc_mshr_13_io_tasks_sink_c_bits_source),
    .io_tasks_sink_c_bits_save(abc_mshr_13_io_tasks_sink_c_bits_save),
    .io_tasks_sink_c_bits_drop(abc_mshr_13_io_tasks_sink_c_bits_drop),
    .io_tasks_sink_c_bits_release(abc_mshr_13_io_tasks_sink_c_bits_release),
    .io_tasks_sink_c_bits_dirty(abc_mshr_13_io_tasks_sink_c_bits_dirty),
    .io_tasks_source_d_ready(abc_mshr_13_io_tasks_source_d_ready),
    .io_tasks_source_d_valid(abc_mshr_13_io_tasks_source_d_valid),
    .io_tasks_source_d_bits_sourceId(abc_mshr_13_io_tasks_source_d_bits_sourceId),
    .io_tasks_source_d_bits_set(abc_mshr_13_io_tasks_source_d_bits_set),
    .io_tasks_source_d_bits_tag(abc_mshr_13_io_tasks_source_d_bits_tag),
    .io_tasks_source_d_bits_channel(abc_mshr_13_io_tasks_source_d_bits_channel),
    .io_tasks_source_d_bits_opcode(abc_mshr_13_io_tasks_source_d_bits_opcode),
    .io_tasks_source_d_bits_param(abc_mshr_13_io_tasks_source_d_bits_param),
    .io_tasks_source_d_bits_size(abc_mshr_13_io_tasks_source_d_bits_size),
    .io_tasks_source_d_bits_way(abc_mshr_13_io_tasks_source_d_bits_way),
    .io_tasks_source_d_bits_off(abc_mshr_13_io_tasks_source_d_bits_off),
    .io_tasks_source_d_bits_useBypass(abc_mshr_13_io_tasks_source_d_bits_useBypass),
    .io_tasks_source_d_bits_bufIdx(abc_mshr_13_io_tasks_source_d_bits_bufIdx),
    .io_tasks_source_d_bits_denied(abc_mshr_13_io_tasks_source_d_bits_denied),
    .io_tasks_source_d_bits_sinkId(abc_mshr_13_io_tasks_source_d_bits_sinkId),
    .io_tasks_source_d_bits_bypassPut(abc_mshr_13_io_tasks_source_d_bits_bypassPut),
    .io_tasks_source_d_bits_dirty(abc_mshr_13_io_tasks_source_d_bits_dirty),
    .io_tasks_source_a_ready(abc_mshr_13_io_tasks_source_a_ready),
    .io_tasks_source_a_valid(abc_mshr_13_io_tasks_source_a_valid),
    .io_tasks_source_a_bits_tag(abc_mshr_13_io_tasks_source_a_bits_tag),
    .io_tasks_source_a_bits_set(abc_mshr_13_io_tasks_source_a_bits_set),
    .io_tasks_source_a_bits_off(abc_mshr_13_io_tasks_source_a_bits_off),
    .io_tasks_source_a_bits_mask(abc_mshr_13_io_tasks_source_a_bits_mask),
    .io_tasks_source_a_bits_opcode(abc_mshr_13_io_tasks_source_a_bits_opcode),
    .io_tasks_source_a_bits_param(abc_mshr_13_io_tasks_source_a_bits_param),
    .io_tasks_source_a_bits_source(abc_mshr_13_io_tasks_source_a_bits_source),
    .io_tasks_source_a_bits_bufIdx(abc_mshr_13_io_tasks_source_a_bits_bufIdx),
    .io_tasks_source_a_bits_size(abc_mshr_13_io_tasks_source_a_bits_size),
    .io_tasks_source_a_bits_needData(abc_mshr_13_io_tasks_source_a_bits_needData),
    .io_tasks_source_a_bits_putData(abc_mshr_13_io_tasks_source_a_bits_putData),
    .io_tasks_source_c_ready(abc_mshr_13_io_tasks_source_c_ready),
    .io_tasks_source_c_valid(abc_mshr_13_io_tasks_source_c_valid),
    .io_tasks_source_c_bits_opcode(abc_mshr_13_io_tasks_source_c_bits_opcode),
    .io_tasks_source_c_bits_tag(abc_mshr_13_io_tasks_source_c_bits_tag),
    .io_tasks_source_c_bits_set(abc_mshr_13_io_tasks_source_c_bits_set),
    .io_tasks_source_c_bits_param(abc_mshr_13_io_tasks_source_c_bits_param),
    .io_tasks_source_c_bits_source(abc_mshr_13_io_tasks_source_c_bits_source),
    .io_tasks_source_c_bits_way(abc_mshr_13_io_tasks_source_c_bits_way),
    .io_tasks_source_c_bits_dirty(abc_mshr_13_io_tasks_source_c_bits_dirty),
    .io_tasks_source_e_ready(abc_mshr_13_io_tasks_source_e_ready),
    .io_tasks_source_e_valid(abc_mshr_13_io_tasks_source_e_valid),
    .io_tasks_source_e_bits_sink(abc_mshr_13_io_tasks_source_e_bits_sink),
    .io_tasks_dir_write_ready(abc_mshr_13_io_tasks_dir_write_ready),
    .io_tasks_dir_write_valid(abc_mshr_13_io_tasks_dir_write_valid),
    .io_tasks_dir_write_bits_set(abc_mshr_13_io_tasks_dir_write_bits_set),
    .io_tasks_dir_write_bits_way(abc_mshr_13_io_tasks_dir_write_bits_way),
    .io_tasks_dir_write_bits_data_dirty(abc_mshr_13_io_tasks_dir_write_bits_data_dirty),
    .io_tasks_dir_write_bits_data_state(abc_mshr_13_io_tasks_dir_write_bits_data_state),
    .io_tasks_dir_write_bits_data_clientStates_0(abc_mshr_13_io_tasks_dir_write_bits_data_clientStates_0),
    .io_tasks_dir_write_bits_data_clientStates_1(abc_mshr_13_io_tasks_dir_write_bits_data_clientStates_1),
    .io_tasks_tag_write_ready(abc_mshr_13_io_tasks_tag_write_ready),
    .io_tasks_tag_write_valid(abc_mshr_13_io_tasks_tag_write_valid),
    .io_tasks_tag_write_bits_set(abc_mshr_13_io_tasks_tag_write_bits_set),
    .io_tasks_tag_write_bits_way(abc_mshr_13_io_tasks_tag_write_bits_way),
    .io_tasks_tag_write_bits_tag(abc_mshr_13_io_tasks_tag_write_bits_tag),
    .io_tasks_client_dir_write_ready(abc_mshr_13_io_tasks_client_dir_write_ready),
    .io_tasks_client_dir_write_valid(abc_mshr_13_io_tasks_client_dir_write_valid),
    .io_tasks_client_dir_write_bits_set(abc_mshr_13_io_tasks_client_dir_write_bits_set),
    .io_tasks_client_dir_write_bits_way(abc_mshr_13_io_tasks_client_dir_write_bits_way),
    .io_tasks_client_dir_write_bits_data_0_state(abc_mshr_13_io_tasks_client_dir_write_bits_data_0_state),
    .io_tasks_client_dir_write_bits_data_1_state(abc_mshr_13_io_tasks_client_dir_write_bits_data_1_state),
    .io_tasks_client_tag_write_ready(abc_mshr_13_io_tasks_client_tag_write_ready),
    .io_tasks_client_tag_write_valid(abc_mshr_13_io_tasks_client_tag_write_valid),
    .io_tasks_client_tag_write_bits_set(abc_mshr_13_io_tasks_client_tag_write_bits_set),
    .io_tasks_client_tag_write_bits_way(abc_mshr_13_io_tasks_client_tag_write_bits_way),
    .io_tasks_client_tag_write_bits_tag(abc_mshr_13_io_tasks_client_tag_write_bits_tag),
    .io_dirResult_valid(abc_mshr_13_io_dirResult_valid),
    .io_dirResult_bits_self_dirty(abc_mshr_13_io_dirResult_bits_self_dirty),
    .io_dirResult_bits_self_state(abc_mshr_13_io_dirResult_bits_self_state),
    .io_dirResult_bits_self_clientStates_0(abc_mshr_13_io_dirResult_bits_self_clientStates_0),
    .io_dirResult_bits_self_clientStates_1(abc_mshr_13_io_dirResult_bits_self_clientStates_1),
    .io_dirResult_bits_self_hit(abc_mshr_13_io_dirResult_bits_self_hit),
    .io_dirResult_bits_self_way(abc_mshr_13_io_dirResult_bits_self_way),
    .io_dirResult_bits_self_tag(abc_mshr_13_io_dirResult_bits_self_tag),
    .io_dirResult_bits_clients_states_0_state(abc_mshr_13_io_dirResult_bits_clients_states_0_state),
    .io_dirResult_bits_clients_states_0_hit(abc_mshr_13_io_dirResult_bits_clients_states_0_hit),
    .io_dirResult_bits_clients_states_1_state(abc_mshr_13_io_dirResult_bits_clients_states_1_state),
    .io_dirResult_bits_clients_states_1_hit(abc_mshr_13_io_dirResult_bits_clients_states_1_hit),
    .io_dirResult_bits_clients_tag(abc_mshr_13_io_dirResult_bits_clients_tag),
    .io_dirResult_bits_clients_way(abc_mshr_13_io_dirResult_bits_clients_way),
    .io_c_status_set(abc_mshr_13_io_c_status_set),
    .io_c_status_tag(abc_mshr_13_io_c_status_tag),
    .io_c_status_way(abc_mshr_13_io_c_status_way),
    .io_c_status_nestedReleaseData(abc_mshr_13_io_c_status_nestedReleaseData),
    .io_c_status_releaseThrough(abc_mshr_13_io_c_status_releaseThrough),
    .io_bstatus_set(abc_mshr_13_io_bstatus_set),
    .io_bstatus_tag(abc_mshr_13_io_bstatus_tag),
    .io_bstatus_way(abc_mshr_13_io_bstatus_way),
    .io_bstatus_nestedProbeAckData(abc_mshr_13_io_bstatus_nestedProbeAckData),
    .io_bstatus_probeHelperFinish(abc_mshr_13_io_bstatus_probeHelperFinish),
    .io_bstatus_probeAckDataThrough(abc_mshr_13_io_bstatus_probeAckDataThrough),
    .io_releaseThrough(abc_mshr_13_io_releaseThrough),
    .io_probeAckDataThrough(abc_mshr_13_io_probeAckDataThrough),
    .io_is_nestedReleaseData(abc_mshr_13_io_is_nestedReleaseData),
    .io_is_nestedProbeAckData(abc_mshr_13_io_is_nestedProbeAckData),
    .io_probeHelperFinish(abc_mshr_13_io_probeHelperFinish)
  );
  MSHR bc_mshr ( // @[Slice.scala 94:16]
    .clock(bc_mshr_clock),
    .reset(bc_mshr_reset),
    .io_id(bc_mshr_io_id),
    .io_enable(bc_mshr_io_enable),
    .io_alloc_valid(bc_mshr_io_alloc_valid),
    .io_alloc_bits_channel(bc_mshr_io_alloc_bits_channel),
    .io_alloc_bits_opcode(bc_mshr_io_alloc_bits_opcode),
    .io_alloc_bits_param(bc_mshr_io_alloc_bits_param),
    .io_alloc_bits_size(bc_mshr_io_alloc_bits_size),
    .io_alloc_bits_source(bc_mshr_io_alloc_bits_source),
    .io_alloc_bits_set(bc_mshr_io_alloc_bits_set),
    .io_alloc_bits_tag(bc_mshr_io_alloc_bits_tag),
    .io_alloc_bits_off(bc_mshr_io_alloc_bits_off),
    .io_alloc_bits_mask(bc_mshr_io_alloc_bits_mask),
    .io_alloc_bits_bufIdx(bc_mshr_io_alloc_bits_bufIdx),
    .io_alloc_bits_preferCache(bc_mshr_io_alloc_bits_preferCache),
    .io_alloc_bits_dirty(bc_mshr_io_alloc_bits_dirty),
    .io_alloc_bits_fromProbeHelper(bc_mshr_io_alloc_bits_fromProbeHelper),
    .io_alloc_bits_fromCmoHelper(bc_mshr_io_alloc_bits_fromCmoHelper),
    .io_alloc_bits_needProbeAckData(bc_mshr_io_alloc_bits_needProbeAckData),
    .io_status_valid(bc_mshr_io_status_valid),
    .io_status_bits_set(bc_mshr_io_status_bits_set),
    .io_status_bits_tag(bc_mshr_io_status_bits_tag),
    .io_status_bits_way(bc_mshr_io_status_bits_way),
    .io_status_bits_way_reg(bc_mshr_io_status_bits_way_reg),
    .io_status_bits_nestB(bc_mshr_io_status_bits_nestB),
    .io_status_bits_nestC(bc_mshr_io_status_bits_nestC),
    .io_status_bits_will_grant_data(bc_mshr_io_status_bits_will_grant_data),
    .io_status_bits_will_save_data(bc_mshr_io_status_bits_will_save_data),
    .io_status_bits_will_free(bc_mshr_io_status_bits_will_free),
    .io_resps_sink_c_valid(bc_mshr_io_resps_sink_c_valid),
    .io_resps_sink_c_bits_hasData(bc_mshr_io_resps_sink_c_bits_hasData),
    .io_resps_sink_c_bits_param(bc_mshr_io_resps_sink_c_bits_param),
    .io_resps_sink_c_bits_source(bc_mshr_io_resps_sink_c_bits_source),
    .io_resps_sink_c_bits_last(bc_mshr_io_resps_sink_c_bits_last),
    .io_resps_sink_c_bits_bufIdx(bc_mshr_io_resps_sink_c_bits_bufIdx),
    .io_resps_sink_d_valid(bc_mshr_io_resps_sink_d_valid),
    .io_resps_sink_d_bits_opcode(bc_mshr_io_resps_sink_d_bits_opcode),
    .io_resps_sink_d_bits_param(bc_mshr_io_resps_sink_d_bits_param),
    .io_resps_sink_d_bits_sink(bc_mshr_io_resps_sink_d_bits_sink),
    .io_resps_sink_d_bits_last(bc_mshr_io_resps_sink_d_bits_last),
    .io_resps_sink_d_bits_denied(bc_mshr_io_resps_sink_d_bits_denied),
    .io_resps_sink_d_bits_bufIdx(bc_mshr_io_resps_sink_d_bits_bufIdx),
    .io_resps_sink_e_valid(bc_mshr_io_resps_sink_e_valid),
    .io_resps_source_d_valid(bc_mshr_io_resps_source_d_valid),
    .io_nestedwb_set(bc_mshr_io_nestedwb_set),
    .io_nestedwb_tag(bc_mshr_io_nestedwb_tag),
    .io_nestedwb_btoN(bc_mshr_io_nestedwb_btoN),
    .io_nestedwb_btoB(bc_mshr_io_nestedwb_btoB),
    .io_nestedwb_bclr_dirty(bc_mshr_io_nestedwb_bclr_dirty),
    .io_nestedwb_bset_dirty(bc_mshr_io_nestedwb_bset_dirty),
    .io_nestedwb_c_set_dirty(bc_mshr_io_nestedwb_c_set_dirty),
    .io_nestedwb_c_set_hit(bc_mshr_io_nestedwb_c_set_hit),
    .io_nestedwb_clients_0_isToN(bc_mshr_io_nestedwb_clients_0_isToN),
    .io_nestedwb_clients_1_isToN(bc_mshr_io_nestedwb_clients_1_isToN),
    .io_tasks_sink_a_ready(bc_mshr_io_tasks_sink_a_ready),
    .io_tasks_sink_a_valid(bc_mshr_io_tasks_sink_a_valid),
    .io_tasks_sink_a_bits_sourceId(bc_mshr_io_tasks_sink_a_bits_sourceId),
    .io_tasks_sink_a_bits_set(bc_mshr_io_tasks_sink_a_bits_set),
    .io_tasks_sink_a_bits_tag(bc_mshr_io_tasks_sink_a_bits_tag),
    .io_tasks_sink_a_bits_size(bc_mshr_io_tasks_sink_a_bits_size),
    .io_tasks_sink_a_bits_off(bc_mshr_io_tasks_sink_a_bits_off),
    .io_tasks_source_bready(bc_mshr_io_tasks_source_bready),
    .io_tasks_source_bvalid(bc_mshr_io_tasks_source_bvalid),
    .io_tasks_source_bset(bc_mshr_io_tasks_source_bset),
    .io_tasks_source_btag(bc_mshr_io_tasks_source_btag),
    .io_tasks_source_bparam(bc_mshr_io_tasks_source_bparam),
    .io_tasks_source_bclients(bc_mshr_io_tasks_source_bclients),
    .io_tasks_source_bneedData(bc_mshr_io_tasks_source_bneedData),
    .io_tasks_sink_c_ready(bc_mshr_io_tasks_sink_c_ready),
    .io_tasks_sink_c_valid(bc_mshr_io_tasks_sink_c_valid),
    .io_tasks_sink_c_bits_sourceId(bc_mshr_io_tasks_sink_c_bits_sourceId),
    .io_tasks_sink_c_bits_set(bc_mshr_io_tasks_sink_c_bits_set),
    .io_tasks_sink_c_bits_tag(bc_mshr_io_tasks_sink_c_bits_tag),
    .io_tasks_sink_c_bits_size(bc_mshr_io_tasks_sink_c_bits_size),
    .io_tasks_sink_c_bits_way(bc_mshr_io_tasks_sink_c_bits_way),
    .io_tasks_sink_c_bits_off(bc_mshr_io_tasks_sink_c_bits_off),
    .io_tasks_sink_c_bits_bufIdx(bc_mshr_io_tasks_sink_c_bits_bufIdx),
    .io_tasks_sink_c_bits_opcode(bc_mshr_io_tasks_sink_c_bits_opcode),
    .io_tasks_sink_c_bits_param(bc_mshr_io_tasks_sink_c_bits_param),
    .io_tasks_sink_c_bits_source(bc_mshr_io_tasks_sink_c_bits_source),
    .io_tasks_sink_c_bits_save(bc_mshr_io_tasks_sink_c_bits_save),
    .io_tasks_sink_c_bits_drop(bc_mshr_io_tasks_sink_c_bits_drop),
    .io_tasks_sink_c_bits_release(bc_mshr_io_tasks_sink_c_bits_release),
    .io_tasks_sink_c_bits_dirty(bc_mshr_io_tasks_sink_c_bits_dirty),
    .io_tasks_source_d_ready(bc_mshr_io_tasks_source_d_ready),
    .io_tasks_source_d_valid(bc_mshr_io_tasks_source_d_valid),
    .io_tasks_source_d_bits_sourceId(bc_mshr_io_tasks_source_d_bits_sourceId),
    .io_tasks_source_d_bits_set(bc_mshr_io_tasks_source_d_bits_set),
    .io_tasks_source_d_bits_tag(bc_mshr_io_tasks_source_d_bits_tag),
    .io_tasks_source_d_bits_channel(bc_mshr_io_tasks_source_d_bits_channel),
    .io_tasks_source_d_bits_opcode(bc_mshr_io_tasks_source_d_bits_opcode),
    .io_tasks_source_d_bits_param(bc_mshr_io_tasks_source_d_bits_param),
    .io_tasks_source_d_bits_size(bc_mshr_io_tasks_source_d_bits_size),
    .io_tasks_source_d_bits_way(bc_mshr_io_tasks_source_d_bits_way),
    .io_tasks_source_d_bits_off(bc_mshr_io_tasks_source_d_bits_off),
    .io_tasks_source_d_bits_useBypass(bc_mshr_io_tasks_source_d_bits_useBypass),
    .io_tasks_source_d_bits_bufIdx(bc_mshr_io_tasks_source_d_bits_bufIdx),
    .io_tasks_source_d_bits_denied(bc_mshr_io_tasks_source_d_bits_denied),
    .io_tasks_source_d_bits_sinkId(bc_mshr_io_tasks_source_d_bits_sinkId),
    .io_tasks_source_d_bits_bypassPut(bc_mshr_io_tasks_source_d_bits_bypassPut),
    .io_tasks_source_d_bits_dirty(bc_mshr_io_tasks_source_d_bits_dirty),
    .io_tasks_source_a_ready(bc_mshr_io_tasks_source_a_ready),
    .io_tasks_source_a_valid(bc_mshr_io_tasks_source_a_valid),
    .io_tasks_source_a_bits_tag(bc_mshr_io_tasks_source_a_bits_tag),
    .io_tasks_source_a_bits_set(bc_mshr_io_tasks_source_a_bits_set),
    .io_tasks_source_a_bits_off(bc_mshr_io_tasks_source_a_bits_off),
    .io_tasks_source_a_bits_mask(bc_mshr_io_tasks_source_a_bits_mask),
    .io_tasks_source_a_bits_opcode(bc_mshr_io_tasks_source_a_bits_opcode),
    .io_tasks_source_a_bits_param(bc_mshr_io_tasks_source_a_bits_param),
    .io_tasks_source_a_bits_source(bc_mshr_io_tasks_source_a_bits_source),
    .io_tasks_source_a_bits_bufIdx(bc_mshr_io_tasks_source_a_bits_bufIdx),
    .io_tasks_source_a_bits_size(bc_mshr_io_tasks_source_a_bits_size),
    .io_tasks_source_a_bits_needData(bc_mshr_io_tasks_source_a_bits_needData),
    .io_tasks_source_a_bits_putData(bc_mshr_io_tasks_source_a_bits_putData),
    .io_tasks_source_c_ready(bc_mshr_io_tasks_source_c_ready),
    .io_tasks_source_c_valid(bc_mshr_io_tasks_source_c_valid),
    .io_tasks_source_c_bits_opcode(bc_mshr_io_tasks_source_c_bits_opcode),
    .io_tasks_source_c_bits_tag(bc_mshr_io_tasks_source_c_bits_tag),
    .io_tasks_source_c_bits_set(bc_mshr_io_tasks_source_c_bits_set),
    .io_tasks_source_c_bits_param(bc_mshr_io_tasks_source_c_bits_param),
    .io_tasks_source_c_bits_source(bc_mshr_io_tasks_source_c_bits_source),
    .io_tasks_source_c_bits_way(bc_mshr_io_tasks_source_c_bits_way),
    .io_tasks_source_c_bits_dirty(bc_mshr_io_tasks_source_c_bits_dirty),
    .io_tasks_source_e_ready(bc_mshr_io_tasks_source_e_ready),
    .io_tasks_source_e_valid(bc_mshr_io_tasks_source_e_valid),
    .io_tasks_source_e_bits_sink(bc_mshr_io_tasks_source_e_bits_sink),
    .io_tasks_dir_write_ready(bc_mshr_io_tasks_dir_write_ready),
    .io_tasks_dir_write_valid(bc_mshr_io_tasks_dir_write_valid),
    .io_tasks_dir_write_bits_set(bc_mshr_io_tasks_dir_write_bits_set),
    .io_tasks_dir_write_bits_way(bc_mshr_io_tasks_dir_write_bits_way),
    .io_tasks_dir_write_bits_data_dirty(bc_mshr_io_tasks_dir_write_bits_data_dirty),
    .io_tasks_dir_write_bits_data_state(bc_mshr_io_tasks_dir_write_bits_data_state),
    .io_tasks_dir_write_bits_data_clientStates_0(bc_mshr_io_tasks_dir_write_bits_data_clientStates_0),
    .io_tasks_dir_write_bits_data_clientStates_1(bc_mshr_io_tasks_dir_write_bits_data_clientStates_1),
    .io_tasks_tag_write_ready(bc_mshr_io_tasks_tag_write_ready),
    .io_tasks_tag_write_valid(bc_mshr_io_tasks_tag_write_valid),
    .io_tasks_tag_write_bits_set(bc_mshr_io_tasks_tag_write_bits_set),
    .io_tasks_tag_write_bits_way(bc_mshr_io_tasks_tag_write_bits_way),
    .io_tasks_tag_write_bits_tag(bc_mshr_io_tasks_tag_write_bits_tag),
    .io_tasks_client_dir_write_ready(bc_mshr_io_tasks_client_dir_write_ready),
    .io_tasks_client_dir_write_valid(bc_mshr_io_tasks_client_dir_write_valid),
    .io_tasks_client_dir_write_bits_set(bc_mshr_io_tasks_client_dir_write_bits_set),
    .io_tasks_client_dir_write_bits_way(bc_mshr_io_tasks_client_dir_write_bits_way),
    .io_tasks_client_dir_write_bits_data_0_state(bc_mshr_io_tasks_client_dir_write_bits_data_0_state),
    .io_tasks_client_dir_write_bits_data_1_state(bc_mshr_io_tasks_client_dir_write_bits_data_1_state),
    .io_tasks_client_tag_write_ready(bc_mshr_io_tasks_client_tag_write_ready),
    .io_tasks_client_tag_write_valid(bc_mshr_io_tasks_client_tag_write_valid),
    .io_tasks_client_tag_write_bits_set(bc_mshr_io_tasks_client_tag_write_bits_set),
    .io_tasks_client_tag_write_bits_way(bc_mshr_io_tasks_client_tag_write_bits_way),
    .io_tasks_client_tag_write_bits_tag(bc_mshr_io_tasks_client_tag_write_bits_tag),
    .io_dirResult_valid(bc_mshr_io_dirResult_valid),
    .io_dirResult_bits_self_dirty(bc_mshr_io_dirResult_bits_self_dirty),
    .io_dirResult_bits_self_state(bc_mshr_io_dirResult_bits_self_state),
    .io_dirResult_bits_self_clientStates_0(bc_mshr_io_dirResult_bits_self_clientStates_0),
    .io_dirResult_bits_self_clientStates_1(bc_mshr_io_dirResult_bits_self_clientStates_1),
    .io_dirResult_bits_self_hit(bc_mshr_io_dirResult_bits_self_hit),
    .io_dirResult_bits_self_way(bc_mshr_io_dirResult_bits_self_way),
    .io_dirResult_bits_self_tag(bc_mshr_io_dirResult_bits_self_tag),
    .io_dirResult_bits_clients_states_0_state(bc_mshr_io_dirResult_bits_clients_states_0_state),
    .io_dirResult_bits_clients_states_0_hit(bc_mshr_io_dirResult_bits_clients_states_0_hit),
    .io_dirResult_bits_clients_states_1_state(bc_mshr_io_dirResult_bits_clients_states_1_state),
    .io_dirResult_bits_clients_states_1_hit(bc_mshr_io_dirResult_bits_clients_states_1_hit),
    .io_dirResult_bits_clients_tag(bc_mshr_io_dirResult_bits_clients_tag),
    .io_dirResult_bits_clients_way(bc_mshr_io_dirResult_bits_clients_way),
    .io_c_status_set(bc_mshr_io_c_status_set),
    .io_c_status_tag(bc_mshr_io_c_status_tag),
    .io_c_status_way(bc_mshr_io_c_status_way),
    .io_c_status_nestedReleaseData(bc_mshr_io_c_status_nestedReleaseData),
    .io_c_status_releaseThrough(bc_mshr_io_c_status_releaseThrough),
    .io_bstatus_set(bc_mshr_io_bstatus_set),
    .io_bstatus_tag(bc_mshr_io_bstatus_tag),
    .io_bstatus_way(bc_mshr_io_bstatus_way),
    .io_bstatus_nestedProbeAckData(bc_mshr_io_bstatus_nestedProbeAckData),
    .io_bstatus_probeHelperFinish(bc_mshr_io_bstatus_probeHelperFinish),
    .io_bstatus_probeAckDataThrough(bc_mshr_io_bstatus_probeAckDataThrough),
    .io_releaseThrough(bc_mshr_io_releaseThrough),
    .io_probeAckDataThrough(bc_mshr_io_probeAckDataThrough),
    .io_is_nestedReleaseData(bc_mshr_io_is_nestedReleaseData),
    .io_is_nestedProbeAckData(bc_mshr_io_is_nestedProbeAckData),
    .io_probeHelperFinish(bc_mshr_io_probeHelperFinish)
  );
  MSHR c_mshr ( // @[Slice.scala 94:16]
    .clock(c_mshr_clock),
    .reset(c_mshr_reset),
    .io_id(c_mshr_io_id),
    .io_enable(c_mshr_io_enable),
    .io_alloc_valid(c_mshr_io_alloc_valid),
    .io_alloc_bits_channel(c_mshr_io_alloc_bits_channel),
    .io_alloc_bits_opcode(c_mshr_io_alloc_bits_opcode),
    .io_alloc_bits_param(c_mshr_io_alloc_bits_param),
    .io_alloc_bits_size(c_mshr_io_alloc_bits_size),
    .io_alloc_bits_source(c_mshr_io_alloc_bits_source),
    .io_alloc_bits_set(c_mshr_io_alloc_bits_set),
    .io_alloc_bits_tag(c_mshr_io_alloc_bits_tag),
    .io_alloc_bits_off(c_mshr_io_alloc_bits_off),
    .io_alloc_bits_mask(c_mshr_io_alloc_bits_mask),
    .io_alloc_bits_bufIdx(c_mshr_io_alloc_bits_bufIdx),
    .io_alloc_bits_preferCache(c_mshr_io_alloc_bits_preferCache),
    .io_alloc_bits_dirty(c_mshr_io_alloc_bits_dirty),
    .io_alloc_bits_fromProbeHelper(c_mshr_io_alloc_bits_fromProbeHelper),
    .io_alloc_bits_fromCmoHelper(c_mshr_io_alloc_bits_fromCmoHelper),
    .io_alloc_bits_needProbeAckData(c_mshr_io_alloc_bits_needProbeAckData),
    .io_status_valid(c_mshr_io_status_valid),
    .io_status_bits_set(c_mshr_io_status_bits_set),
    .io_status_bits_tag(c_mshr_io_status_bits_tag),
    .io_status_bits_way(c_mshr_io_status_bits_way),
    .io_status_bits_way_reg(c_mshr_io_status_bits_way_reg),
    .io_status_bits_nestB(c_mshr_io_status_bits_nestB),
    .io_status_bits_nestC(c_mshr_io_status_bits_nestC),
    .io_status_bits_will_grant_data(c_mshr_io_status_bits_will_grant_data),
    .io_status_bits_will_save_data(c_mshr_io_status_bits_will_save_data),
    .io_status_bits_will_free(c_mshr_io_status_bits_will_free),
    .io_resps_sink_c_valid(c_mshr_io_resps_sink_c_valid),
    .io_resps_sink_c_bits_hasData(c_mshr_io_resps_sink_c_bits_hasData),
    .io_resps_sink_c_bits_param(c_mshr_io_resps_sink_c_bits_param),
    .io_resps_sink_c_bits_source(c_mshr_io_resps_sink_c_bits_source),
    .io_resps_sink_c_bits_last(c_mshr_io_resps_sink_c_bits_last),
    .io_resps_sink_c_bits_bufIdx(c_mshr_io_resps_sink_c_bits_bufIdx),
    .io_resps_sink_d_valid(c_mshr_io_resps_sink_d_valid),
    .io_resps_sink_d_bits_opcode(c_mshr_io_resps_sink_d_bits_opcode),
    .io_resps_sink_d_bits_param(c_mshr_io_resps_sink_d_bits_param),
    .io_resps_sink_d_bits_sink(c_mshr_io_resps_sink_d_bits_sink),
    .io_resps_sink_d_bits_last(c_mshr_io_resps_sink_d_bits_last),
    .io_resps_sink_d_bits_denied(c_mshr_io_resps_sink_d_bits_denied),
    .io_resps_sink_d_bits_bufIdx(c_mshr_io_resps_sink_d_bits_bufIdx),
    .io_resps_sink_e_valid(c_mshr_io_resps_sink_e_valid),
    .io_resps_source_d_valid(c_mshr_io_resps_source_d_valid),
    .io_nestedwb_set(c_mshr_io_nestedwb_set),
    .io_nestedwb_tag(c_mshr_io_nestedwb_tag),
    .io_nestedwb_btoN(c_mshr_io_nestedwb_btoN),
    .io_nestedwb_btoB(c_mshr_io_nestedwb_btoB),
    .io_nestedwb_bclr_dirty(c_mshr_io_nestedwb_bclr_dirty),
    .io_nestedwb_bset_dirty(c_mshr_io_nestedwb_bset_dirty),
    .io_nestedwb_c_set_dirty(c_mshr_io_nestedwb_c_set_dirty),
    .io_nestedwb_c_set_hit(c_mshr_io_nestedwb_c_set_hit),
    .io_nestedwb_clients_0_isToN(c_mshr_io_nestedwb_clients_0_isToN),
    .io_nestedwb_clients_1_isToN(c_mshr_io_nestedwb_clients_1_isToN),
    .io_tasks_sink_a_ready(c_mshr_io_tasks_sink_a_ready),
    .io_tasks_sink_a_valid(c_mshr_io_tasks_sink_a_valid),
    .io_tasks_sink_a_bits_sourceId(c_mshr_io_tasks_sink_a_bits_sourceId),
    .io_tasks_sink_a_bits_set(c_mshr_io_tasks_sink_a_bits_set),
    .io_tasks_sink_a_bits_tag(c_mshr_io_tasks_sink_a_bits_tag),
    .io_tasks_sink_a_bits_size(c_mshr_io_tasks_sink_a_bits_size),
    .io_tasks_sink_a_bits_off(c_mshr_io_tasks_sink_a_bits_off),
    .io_tasks_source_bready(c_mshr_io_tasks_source_bready),
    .io_tasks_source_bvalid(c_mshr_io_tasks_source_bvalid),
    .io_tasks_source_bset(c_mshr_io_tasks_source_bset),
    .io_tasks_source_btag(c_mshr_io_tasks_source_btag),
    .io_tasks_source_bparam(c_mshr_io_tasks_source_bparam),
    .io_tasks_source_bclients(c_mshr_io_tasks_source_bclients),
    .io_tasks_source_bneedData(c_mshr_io_tasks_source_bneedData),
    .io_tasks_sink_c_ready(c_mshr_io_tasks_sink_c_ready),
    .io_tasks_sink_c_valid(c_mshr_io_tasks_sink_c_valid),
    .io_tasks_sink_c_bits_sourceId(c_mshr_io_tasks_sink_c_bits_sourceId),
    .io_tasks_sink_c_bits_set(c_mshr_io_tasks_sink_c_bits_set),
    .io_tasks_sink_c_bits_tag(c_mshr_io_tasks_sink_c_bits_tag),
    .io_tasks_sink_c_bits_size(c_mshr_io_tasks_sink_c_bits_size),
    .io_tasks_sink_c_bits_way(c_mshr_io_tasks_sink_c_bits_way),
    .io_tasks_sink_c_bits_off(c_mshr_io_tasks_sink_c_bits_off),
    .io_tasks_sink_c_bits_bufIdx(c_mshr_io_tasks_sink_c_bits_bufIdx),
    .io_tasks_sink_c_bits_opcode(c_mshr_io_tasks_sink_c_bits_opcode),
    .io_tasks_sink_c_bits_param(c_mshr_io_tasks_sink_c_bits_param),
    .io_tasks_sink_c_bits_source(c_mshr_io_tasks_sink_c_bits_source),
    .io_tasks_sink_c_bits_save(c_mshr_io_tasks_sink_c_bits_save),
    .io_tasks_sink_c_bits_drop(c_mshr_io_tasks_sink_c_bits_drop),
    .io_tasks_sink_c_bits_release(c_mshr_io_tasks_sink_c_bits_release),
    .io_tasks_sink_c_bits_dirty(c_mshr_io_tasks_sink_c_bits_dirty),
    .io_tasks_source_d_ready(c_mshr_io_tasks_source_d_ready),
    .io_tasks_source_d_valid(c_mshr_io_tasks_source_d_valid),
    .io_tasks_source_d_bits_sourceId(c_mshr_io_tasks_source_d_bits_sourceId),
    .io_tasks_source_d_bits_set(c_mshr_io_tasks_source_d_bits_set),
    .io_tasks_source_d_bits_tag(c_mshr_io_tasks_source_d_bits_tag),
    .io_tasks_source_d_bits_channel(c_mshr_io_tasks_source_d_bits_channel),
    .io_tasks_source_d_bits_opcode(c_mshr_io_tasks_source_d_bits_opcode),
    .io_tasks_source_d_bits_param(c_mshr_io_tasks_source_d_bits_param),
    .io_tasks_source_d_bits_size(c_mshr_io_tasks_source_d_bits_size),
    .io_tasks_source_d_bits_way(c_mshr_io_tasks_source_d_bits_way),
    .io_tasks_source_d_bits_off(c_mshr_io_tasks_source_d_bits_off),
    .io_tasks_source_d_bits_useBypass(c_mshr_io_tasks_source_d_bits_useBypass),
    .io_tasks_source_d_bits_bufIdx(c_mshr_io_tasks_source_d_bits_bufIdx),
    .io_tasks_source_d_bits_denied(c_mshr_io_tasks_source_d_bits_denied),
    .io_tasks_source_d_bits_sinkId(c_mshr_io_tasks_source_d_bits_sinkId),
    .io_tasks_source_d_bits_bypassPut(c_mshr_io_tasks_source_d_bits_bypassPut),
    .io_tasks_source_d_bits_dirty(c_mshr_io_tasks_source_d_bits_dirty),
    .io_tasks_source_a_ready(c_mshr_io_tasks_source_a_ready),
    .io_tasks_source_a_valid(c_mshr_io_tasks_source_a_valid),
    .io_tasks_source_a_bits_tag(c_mshr_io_tasks_source_a_bits_tag),
    .io_tasks_source_a_bits_set(c_mshr_io_tasks_source_a_bits_set),
    .io_tasks_source_a_bits_off(c_mshr_io_tasks_source_a_bits_off),
    .io_tasks_source_a_bits_mask(c_mshr_io_tasks_source_a_bits_mask),
    .io_tasks_source_a_bits_opcode(c_mshr_io_tasks_source_a_bits_opcode),
    .io_tasks_source_a_bits_param(c_mshr_io_tasks_source_a_bits_param),
    .io_tasks_source_a_bits_source(c_mshr_io_tasks_source_a_bits_source),
    .io_tasks_source_a_bits_bufIdx(c_mshr_io_tasks_source_a_bits_bufIdx),
    .io_tasks_source_a_bits_size(c_mshr_io_tasks_source_a_bits_size),
    .io_tasks_source_a_bits_needData(c_mshr_io_tasks_source_a_bits_needData),
    .io_tasks_source_a_bits_putData(c_mshr_io_tasks_source_a_bits_putData),
    .io_tasks_source_c_ready(c_mshr_io_tasks_source_c_ready),
    .io_tasks_source_c_valid(c_mshr_io_tasks_source_c_valid),
    .io_tasks_source_c_bits_opcode(c_mshr_io_tasks_source_c_bits_opcode),
    .io_tasks_source_c_bits_tag(c_mshr_io_tasks_source_c_bits_tag),
    .io_tasks_source_c_bits_set(c_mshr_io_tasks_source_c_bits_set),
    .io_tasks_source_c_bits_param(c_mshr_io_tasks_source_c_bits_param),
    .io_tasks_source_c_bits_source(c_mshr_io_tasks_source_c_bits_source),
    .io_tasks_source_c_bits_way(c_mshr_io_tasks_source_c_bits_way),
    .io_tasks_source_c_bits_dirty(c_mshr_io_tasks_source_c_bits_dirty),
    .io_tasks_source_e_ready(c_mshr_io_tasks_source_e_ready),
    .io_tasks_source_e_valid(c_mshr_io_tasks_source_e_valid),
    .io_tasks_source_e_bits_sink(c_mshr_io_tasks_source_e_bits_sink),
    .io_tasks_dir_write_ready(c_mshr_io_tasks_dir_write_ready),
    .io_tasks_dir_write_valid(c_mshr_io_tasks_dir_write_valid),
    .io_tasks_dir_write_bits_set(c_mshr_io_tasks_dir_write_bits_set),
    .io_tasks_dir_write_bits_way(c_mshr_io_tasks_dir_write_bits_way),
    .io_tasks_dir_write_bits_data_dirty(c_mshr_io_tasks_dir_write_bits_data_dirty),
    .io_tasks_dir_write_bits_data_state(c_mshr_io_tasks_dir_write_bits_data_state),
    .io_tasks_dir_write_bits_data_clientStates_0(c_mshr_io_tasks_dir_write_bits_data_clientStates_0),
    .io_tasks_dir_write_bits_data_clientStates_1(c_mshr_io_tasks_dir_write_bits_data_clientStates_1),
    .io_tasks_tag_write_ready(c_mshr_io_tasks_tag_write_ready),
    .io_tasks_tag_write_valid(c_mshr_io_tasks_tag_write_valid),
    .io_tasks_tag_write_bits_set(c_mshr_io_tasks_tag_write_bits_set),
    .io_tasks_tag_write_bits_way(c_mshr_io_tasks_tag_write_bits_way),
    .io_tasks_tag_write_bits_tag(c_mshr_io_tasks_tag_write_bits_tag),
    .io_tasks_client_dir_write_ready(c_mshr_io_tasks_client_dir_write_ready),
    .io_tasks_client_dir_write_valid(c_mshr_io_tasks_client_dir_write_valid),
    .io_tasks_client_dir_write_bits_set(c_mshr_io_tasks_client_dir_write_bits_set),
    .io_tasks_client_dir_write_bits_way(c_mshr_io_tasks_client_dir_write_bits_way),
    .io_tasks_client_dir_write_bits_data_0_state(c_mshr_io_tasks_client_dir_write_bits_data_0_state),
    .io_tasks_client_dir_write_bits_data_1_state(c_mshr_io_tasks_client_dir_write_bits_data_1_state),
    .io_tasks_client_tag_write_ready(c_mshr_io_tasks_client_tag_write_ready),
    .io_tasks_client_tag_write_valid(c_mshr_io_tasks_client_tag_write_valid),
    .io_tasks_client_tag_write_bits_set(c_mshr_io_tasks_client_tag_write_bits_set),
    .io_tasks_client_tag_write_bits_way(c_mshr_io_tasks_client_tag_write_bits_way),
    .io_tasks_client_tag_write_bits_tag(c_mshr_io_tasks_client_tag_write_bits_tag),
    .io_dirResult_valid(c_mshr_io_dirResult_valid),
    .io_dirResult_bits_self_dirty(c_mshr_io_dirResult_bits_self_dirty),
    .io_dirResult_bits_self_state(c_mshr_io_dirResult_bits_self_state),
    .io_dirResult_bits_self_clientStates_0(c_mshr_io_dirResult_bits_self_clientStates_0),
    .io_dirResult_bits_self_clientStates_1(c_mshr_io_dirResult_bits_self_clientStates_1),
    .io_dirResult_bits_self_hit(c_mshr_io_dirResult_bits_self_hit),
    .io_dirResult_bits_self_way(c_mshr_io_dirResult_bits_self_way),
    .io_dirResult_bits_self_tag(c_mshr_io_dirResult_bits_self_tag),
    .io_dirResult_bits_clients_states_0_state(c_mshr_io_dirResult_bits_clients_states_0_state),
    .io_dirResult_bits_clients_states_0_hit(c_mshr_io_dirResult_bits_clients_states_0_hit),
    .io_dirResult_bits_clients_states_1_state(c_mshr_io_dirResult_bits_clients_states_1_state),
    .io_dirResult_bits_clients_states_1_hit(c_mshr_io_dirResult_bits_clients_states_1_hit),
    .io_dirResult_bits_clients_tag(c_mshr_io_dirResult_bits_clients_tag),
    .io_dirResult_bits_clients_way(c_mshr_io_dirResult_bits_clients_way),
    .io_c_status_set(c_mshr_io_c_status_set),
    .io_c_status_tag(c_mshr_io_c_status_tag),
    .io_c_status_way(c_mshr_io_c_status_way),
    .io_c_status_nestedReleaseData(c_mshr_io_c_status_nestedReleaseData),
    .io_c_status_releaseThrough(c_mshr_io_c_status_releaseThrough),
    .io_bstatus_set(c_mshr_io_bstatus_set),
    .io_bstatus_tag(c_mshr_io_bstatus_tag),
    .io_bstatus_way(c_mshr_io_bstatus_way),
    .io_bstatus_nestedProbeAckData(c_mshr_io_bstatus_nestedProbeAckData),
    .io_bstatus_probeHelperFinish(c_mshr_io_bstatus_probeHelperFinish),
    .io_bstatus_probeAckDataThrough(c_mshr_io_bstatus_probeAckDataThrough),
    .io_releaseThrough(c_mshr_io_releaseThrough),
    .io_probeAckDataThrough(c_mshr_io_probeAckDataThrough),
    .io_is_nestedReleaseData(c_mshr_io_is_nestedReleaseData),
    .io_is_nestedProbeAckData(c_mshr_io_is_nestedProbeAckData),
    .io_probeHelperFinish(c_mshr_io_probeHelperFinish)
  );
  DataStorage dataStorage ( // @[Slice.scala 101:27]
    .clock(dataStorage_clock),
    .reset(dataStorage_reset),
    .io_sourceC_raddr_ready(dataStorage_io_sourceC_raddr_ready),
    .io_sourceC_raddr_valid(dataStorage_io_sourceC_raddr_valid),
    .io_sourceC_raddr_bits_way(dataStorage_io_sourceC_raddr_bits_way),
    .io_sourceC_raddr_bits_set(dataStorage_io_sourceC_raddr_bits_set),
    .io_sourceC_raddr_bits_beat(dataStorage_io_sourceC_raddr_bits_beat),
    .io_sourceC_rdata_data(dataStorage_io_sourceC_rdata_data),
    .io_sinkD_waddr_ready(dataStorage_io_sinkD_waddr_ready),
    .io_sinkD_waddr_valid(dataStorage_io_sinkD_waddr_valid),
    .io_sinkD_waddr_bits_way(dataStorage_io_sinkD_waddr_bits_way),
    .io_sinkD_waddr_bits_set(dataStorage_io_sinkD_waddr_bits_set),
    .io_sinkD_waddr_bits_beat(dataStorage_io_sinkD_waddr_bits_beat),
    .io_sinkD_waddr_bits_noop(dataStorage_io_sinkD_waddr_bits_noop),
    .io_sinkD_wdata_data(dataStorage_io_sinkD_wdata_data),
    .io_sourceD_raddr_ready(dataStorage_io_sourceD_raddr_ready),
    .io_sourceD_raddr_valid(dataStorage_io_sourceD_raddr_valid),
    .io_sourceD_raddr_bits_way(dataStorage_io_sourceD_raddr_bits_way),
    .io_sourceD_raddr_bits_set(dataStorage_io_sourceD_raddr_bits_set),
    .io_sourceD_raddr_bits_beat(dataStorage_io_sourceD_raddr_bits_beat),
    .io_sourceD_rdata_data(dataStorage_io_sourceD_rdata_data),
    .io_sourceD_waddr_ready(dataStorage_io_sourceD_waddr_ready),
    .io_sourceD_waddr_valid(dataStorage_io_sourceD_waddr_valid),
    .io_sourceD_waddr_bits_way(dataStorage_io_sourceD_waddr_bits_way),
    .io_sourceD_waddr_bits_set(dataStorage_io_sourceD_waddr_bits_set),
    .io_sourceD_waddr_bits_beat(dataStorage_io_sourceD_waddr_bits_beat),
    .io_sourceD_wdata_data(dataStorage_io_sourceD_wdata_data),
    .io_sinkC_waddr_ready(dataStorage_io_sinkC_waddr_ready),
    .io_sinkC_waddr_valid(dataStorage_io_sinkC_waddr_valid),
    .io_sinkC_waddr_bits_way(dataStorage_io_sinkC_waddr_bits_way),
    .io_sinkC_waddr_bits_set(dataStorage_io_sinkC_waddr_bits_set),
    .io_sinkC_waddr_bits_beat(dataStorage_io_sinkC_waddr_bits_beat),
    .io_sinkC_waddr_bits_noop(dataStorage_io_sinkC_waddr_bits_noop),
    .io_sinkC_wdata_data(dataStorage_io_sinkC_wdata_data)
  );
  MSHRAlloc mshrAlloc ( // @[Slice.scala 123:25]
    .io_a_req_ready(mshrAlloc_io_a_req_ready),
    .io_a_req_valid(mshrAlloc_io_a_req_valid),
    .io_a_req_bits_channel(mshrAlloc_io_a_req_bits_channel),
    .io_a_req_bits_opcode(mshrAlloc_io_a_req_bits_opcode),
    .io_a_req_bits_param(mshrAlloc_io_a_req_bits_param),
    .io_a_req_bits_size(mshrAlloc_io_a_req_bits_size),
    .io_a_req_bits_source(mshrAlloc_io_a_req_bits_source),
    .io_a_req_bits_set(mshrAlloc_io_a_req_bits_set),
    .io_a_req_bits_tag(mshrAlloc_io_a_req_bits_tag),
    .io_a_req_bits_off(mshrAlloc_io_a_req_bits_off),
    .io_a_req_bits_mask(mshrAlloc_io_a_req_bits_mask),
    .io_a_req_bits_bufIdx(mshrAlloc_io_a_req_bits_bufIdx),
    .io_a_req_bits_preferCache(mshrAlloc_io_a_req_bits_preferCache),
    .io_a_req_bits_dirty(mshrAlloc_io_a_req_bits_dirty),
    .io_a_req_bits_fromProbeHelper(mshrAlloc_io_a_req_bits_fromProbeHelper),
    .io_a_req_bits_fromCmoHelper(mshrAlloc_io_a_req_bits_fromCmoHelper),
    .io_a_req_bits_needProbeAckData(mshrAlloc_io_a_req_bits_needProbeAckData),
    .io_breq_ready(mshrAlloc_io_breq_ready),
    .io_breq_valid(mshrAlloc_io_breq_valid),
    .io_breq_bits_channel(mshrAlloc_io_breq_bits_channel),
    .io_breq_bits_opcode(mshrAlloc_io_breq_bits_opcode),
    .io_breq_bits_param(mshrAlloc_io_breq_bits_param),
    .io_breq_bits_size(mshrAlloc_io_breq_bits_size),
    .io_breq_bits_source(mshrAlloc_io_breq_bits_source),
    .io_breq_bits_set(mshrAlloc_io_breq_bits_set),
    .io_breq_bits_tag(mshrAlloc_io_breq_bits_tag),
    .io_breq_bits_off(mshrAlloc_io_breq_bits_off),
    .io_breq_bits_mask(mshrAlloc_io_breq_bits_mask),
    .io_breq_bits_bufIdx(mshrAlloc_io_breq_bits_bufIdx),
    .io_breq_bits_preferCache(mshrAlloc_io_breq_bits_preferCache),
    .io_breq_bits_dirty(mshrAlloc_io_breq_bits_dirty),
    .io_breq_bits_fromProbeHelper(mshrAlloc_io_breq_bits_fromProbeHelper),
    .io_breq_bits_fromCmoHelper(mshrAlloc_io_breq_bits_fromCmoHelper),
    .io_breq_bits_needProbeAckData(mshrAlloc_io_breq_bits_needProbeAckData),
    .io_c_req_ready(mshrAlloc_io_c_req_ready),
    .io_c_req_valid(mshrAlloc_io_c_req_valid),
    .io_c_req_bits_opcode(mshrAlloc_io_c_req_bits_opcode),
    .io_c_req_bits_param(mshrAlloc_io_c_req_bits_param),
    .io_c_req_bits_size(mshrAlloc_io_c_req_bits_size),
    .io_c_req_bits_source(mshrAlloc_io_c_req_bits_source),
    .io_c_req_bits_set(mshrAlloc_io_c_req_bits_set),
    .io_c_req_bits_tag(mshrAlloc_io_c_req_bits_tag),
    .io_c_req_bits_off(mshrAlloc_io_c_req_bits_off),
    .io_c_req_bits_bufIdx(mshrAlloc_io_c_req_bits_bufIdx),
    .io_c_req_bits_dirty(mshrAlloc_io_c_req_bits_dirty),
    .io_status_0_valid(mshrAlloc_io_status_0_valid),
    .io_status_0_bits_set(mshrAlloc_io_status_0_bits_set),
    .io_status_0_bits_nestB(mshrAlloc_io_status_0_bits_nestB),
    .io_status_0_bits_nestC(mshrAlloc_io_status_0_bits_nestC),
    .io_status_1_valid(mshrAlloc_io_status_1_valid),
    .io_status_1_bits_set(mshrAlloc_io_status_1_bits_set),
    .io_status_1_bits_nestB(mshrAlloc_io_status_1_bits_nestB),
    .io_status_1_bits_nestC(mshrAlloc_io_status_1_bits_nestC),
    .io_status_2_valid(mshrAlloc_io_status_2_valid),
    .io_status_2_bits_set(mshrAlloc_io_status_2_bits_set),
    .io_status_2_bits_nestB(mshrAlloc_io_status_2_bits_nestB),
    .io_status_2_bits_nestC(mshrAlloc_io_status_2_bits_nestC),
    .io_status_3_valid(mshrAlloc_io_status_3_valid),
    .io_status_3_bits_set(mshrAlloc_io_status_3_bits_set),
    .io_status_3_bits_nestB(mshrAlloc_io_status_3_bits_nestB),
    .io_status_3_bits_nestC(mshrAlloc_io_status_3_bits_nestC),
    .io_status_4_valid(mshrAlloc_io_status_4_valid),
    .io_status_4_bits_set(mshrAlloc_io_status_4_bits_set),
    .io_status_4_bits_nestB(mshrAlloc_io_status_4_bits_nestB),
    .io_status_4_bits_nestC(mshrAlloc_io_status_4_bits_nestC),
    .io_status_5_valid(mshrAlloc_io_status_5_valid),
    .io_status_5_bits_set(mshrAlloc_io_status_5_bits_set),
    .io_status_5_bits_nestB(mshrAlloc_io_status_5_bits_nestB),
    .io_status_5_bits_nestC(mshrAlloc_io_status_5_bits_nestC),
    .io_status_6_valid(mshrAlloc_io_status_6_valid),
    .io_status_6_bits_set(mshrAlloc_io_status_6_bits_set),
    .io_status_6_bits_nestB(mshrAlloc_io_status_6_bits_nestB),
    .io_status_6_bits_nestC(mshrAlloc_io_status_6_bits_nestC),
    .io_status_7_valid(mshrAlloc_io_status_7_valid),
    .io_status_7_bits_set(mshrAlloc_io_status_7_bits_set),
    .io_status_7_bits_nestB(mshrAlloc_io_status_7_bits_nestB),
    .io_status_7_bits_nestC(mshrAlloc_io_status_7_bits_nestC),
    .io_status_8_valid(mshrAlloc_io_status_8_valid),
    .io_status_8_bits_set(mshrAlloc_io_status_8_bits_set),
    .io_status_8_bits_nestB(mshrAlloc_io_status_8_bits_nestB),
    .io_status_8_bits_nestC(mshrAlloc_io_status_8_bits_nestC),
    .io_status_9_valid(mshrAlloc_io_status_9_valid),
    .io_status_9_bits_set(mshrAlloc_io_status_9_bits_set),
    .io_status_9_bits_nestB(mshrAlloc_io_status_9_bits_nestB),
    .io_status_9_bits_nestC(mshrAlloc_io_status_9_bits_nestC),
    .io_status_10_valid(mshrAlloc_io_status_10_valid),
    .io_status_10_bits_set(mshrAlloc_io_status_10_bits_set),
    .io_status_10_bits_nestB(mshrAlloc_io_status_10_bits_nestB),
    .io_status_10_bits_nestC(mshrAlloc_io_status_10_bits_nestC),
    .io_status_11_valid(mshrAlloc_io_status_11_valid),
    .io_status_11_bits_set(mshrAlloc_io_status_11_bits_set),
    .io_status_11_bits_nestB(mshrAlloc_io_status_11_bits_nestB),
    .io_status_11_bits_nestC(mshrAlloc_io_status_11_bits_nestC),
    .io_status_12_valid(mshrAlloc_io_status_12_valid),
    .io_status_12_bits_set(mshrAlloc_io_status_12_bits_set),
    .io_status_12_bits_nestB(mshrAlloc_io_status_12_bits_nestB),
    .io_status_12_bits_nestC(mshrAlloc_io_status_12_bits_nestC),
    .io_status_13_valid(mshrAlloc_io_status_13_valid),
    .io_status_13_bits_set(mshrAlloc_io_status_13_bits_set),
    .io_status_13_bits_nestB(mshrAlloc_io_status_13_bits_nestB),
    .io_status_13_bits_nestC(mshrAlloc_io_status_13_bits_nestC),
    .io_status_14_valid(mshrAlloc_io_status_14_valid),
    .io_status_14_bits_set(mshrAlloc_io_status_14_bits_set),
    .io_status_14_bits_nestC(mshrAlloc_io_status_14_bits_nestC),
    .io_status_15_valid(mshrAlloc_io_status_15_valid),
    .io_status_15_bits_set(mshrAlloc_io_status_15_bits_set),
    .io_alloc_0_valid(mshrAlloc_io_alloc_0_valid),
    .io_alloc_0_bits_channel(mshrAlloc_io_alloc_0_bits_channel),
    .io_alloc_0_bits_opcode(mshrAlloc_io_alloc_0_bits_opcode),
    .io_alloc_0_bits_param(mshrAlloc_io_alloc_0_bits_param),
    .io_alloc_0_bits_size(mshrAlloc_io_alloc_0_bits_size),
    .io_alloc_0_bits_source(mshrAlloc_io_alloc_0_bits_source),
    .io_alloc_0_bits_set(mshrAlloc_io_alloc_0_bits_set),
    .io_alloc_0_bits_tag(mshrAlloc_io_alloc_0_bits_tag),
    .io_alloc_0_bits_off(mshrAlloc_io_alloc_0_bits_off),
    .io_alloc_0_bits_mask(mshrAlloc_io_alloc_0_bits_mask),
    .io_alloc_0_bits_bufIdx(mshrAlloc_io_alloc_0_bits_bufIdx),
    .io_alloc_0_bits_preferCache(mshrAlloc_io_alloc_0_bits_preferCache),
    .io_alloc_0_bits_dirty(mshrAlloc_io_alloc_0_bits_dirty),
    .io_alloc_0_bits_fromProbeHelper(mshrAlloc_io_alloc_0_bits_fromProbeHelper),
    .io_alloc_0_bits_fromCmoHelper(mshrAlloc_io_alloc_0_bits_fromCmoHelper),
    .io_alloc_0_bits_needProbeAckData(mshrAlloc_io_alloc_0_bits_needProbeAckData),
    .io_alloc_1_valid(mshrAlloc_io_alloc_1_valid),
    .io_alloc_1_bits_channel(mshrAlloc_io_alloc_1_bits_channel),
    .io_alloc_1_bits_opcode(mshrAlloc_io_alloc_1_bits_opcode),
    .io_alloc_1_bits_param(mshrAlloc_io_alloc_1_bits_param),
    .io_alloc_1_bits_size(mshrAlloc_io_alloc_1_bits_size),
    .io_alloc_1_bits_source(mshrAlloc_io_alloc_1_bits_source),
    .io_alloc_1_bits_set(mshrAlloc_io_alloc_1_bits_set),
    .io_alloc_1_bits_tag(mshrAlloc_io_alloc_1_bits_tag),
    .io_alloc_1_bits_off(mshrAlloc_io_alloc_1_bits_off),
    .io_alloc_1_bits_mask(mshrAlloc_io_alloc_1_bits_mask),
    .io_alloc_1_bits_bufIdx(mshrAlloc_io_alloc_1_bits_bufIdx),
    .io_alloc_1_bits_preferCache(mshrAlloc_io_alloc_1_bits_preferCache),
    .io_alloc_1_bits_dirty(mshrAlloc_io_alloc_1_bits_dirty),
    .io_alloc_1_bits_fromProbeHelper(mshrAlloc_io_alloc_1_bits_fromProbeHelper),
    .io_alloc_1_bits_fromCmoHelper(mshrAlloc_io_alloc_1_bits_fromCmoHelper),
    .io_alloc_1_bits_needProbeAckData(mshrAlloc_io_alloc_1_bits_needProbeAckData),
    .io_alloc_2_valid(mshrAlloc_io_alloc_2_valid),
    .io_alloc_2_bits_channel(mshrAlloc_io_alloc_2_bits_channel),
    .io_alloc_2_bits_opcode(mshrAlloc_io_alloc_2_bits_opcode),
    .io_alloc_2_bits_param(mshrAlloc_io_alloc_2_bits_param),
    .io_alloc_2_bits_size(mshrAlloc_io_alloc_2_bits_size),
    .io_alloc_2_bits_source(mshrAlloc_io_alloc_2_bits_source),
    .io_alloc_2_bits_set(mshrAlloc_io_alloc_2_bits_set),
    .io_alloc_2_bits_tag(mshrAlloc_io_alloc_2_bits_tag),
    .io_alloc_2_bits_off(mshrAlloc_io_alloc_2_bits_off),
    .io_alloc_2_bits_mask(mshrAlloc_io_alloc_2_bits_mask),
    .io_alloc_2_bits_bufIdx(mshrAlloc_io_alloc_2_bits_bufIdx),
    .io_alloc_2_bits_preferCache(mshrAlloc_io_alloc_2_bits_preferCache),
    .io_alloc_2_bits_dirty(mshrAlloc_io_alloc_2_bits_dirty),
    .io_alloc_2_bits_fromProbeHelper(mshrAlloc_io_alloc_2_bits_fromProbeHelper),
    .io_alloc_2_bits_fromCmoHelper(mshrAlloc_io_alloc_2_bits_fromCmoHelper),
    .io_alloc_2_bits_needProbeAckData(mshrAlloc_io_alloc_2_bits_needProbeAckData),
    .io_alloc_3_valid(mshrAlloc_io_alloc_3_valid),
    .io_alloc_3_bits_channel(mshrAlloc_io_alloc_3_bits_channel),
    .io_alloc_3_bits_opcode(mshrAlloc_io_alloc_3_bits_opcode),
    .io_alloc_3_bits_param(mshrAlloc_io_alloc_3_bits_param),
    .io_alloc_3_bits_size(mshrAlloc_io_alloc_3_bits_size),
    .io_alloc_3_bits_source(mshrAlloc_io_alloc_3_bits_source),
    .io_alloc_3_bits_set(mshrAlloc_io_alloc_3_bits_set),
    .io_alloc_3_bits_tag(mshrAlloc_io_alloc_3_bits_tag),
    .io_alloc_3_bits_off(mshrAlloc_io_alloc_3_bits_off),
    .io_alloc_3_bits_mask(mshrAlloc_io_alloc_3_bits_mask),
    .io_alloc_3_bits_bufIdx(mshrAlloc_io_alloc_3_bits_bufIdx),
    .io_alloc_3_bits_preferCache(mshrAlloc_io_alloc_3_bits_preferCache),
    .io_alloc_3_bits_dirty(mshrAlloc_io_alloc_3_bits_dirty),
    .io_alloc_3_bits_fromProbeHelper(mshrAlloc_io_alloc_3_bits_fromProbeHelper),
    .io_alloc_3_bits_fromCmoHelper(mshrAlloc_io_alloc_3_bits_fromCmoHelper),
    .io_alloc_3_bits_needProbeAckData(mshrAlloc_io_alloc_3_bits_needProbeAckData),
    .io_alloc_4_valid(mshrAlloc_io_alloc_4_valid),
    .io_alloc_4_bits_channel(mshrAlloc_io_alloc_4_bits_channel),
    .io_alloc_4_bits_opcode(mshrAlloc_io_alloc_4_bits_opcode),
    .io_alloc_4_bits_param(mshrAlloc_io_alloc_4_bits_param),
    .io_alloc_4_bits_size(mshrAlloc_io_alloc_4_bits_size),
    .io_alloc_4_bits_source(mshrAlloc_io_alloc_4_bits_source),
    .io_alloc_4_bits_set(mshrAlloc_io_alloc_4_bits_set),
    .io_alloc_4_bits_tag(mshrAlloc_io_alloc_4_bits_tag),
    .io_alloc_4_bits_off(mshrAlloc_io_alloc_4_bits_off),
    .io_alloc_4_bits_mask(mshrAlloc_io_alloc_4_bits_mask),
    .io_alloc_4_bits_bufIdx(mshrAlloc_io_alloc_4_bits_bufIdx),
    .io_alloc_4_bits_preferCache(mshrAlloc_io_alloc_4_bits_preferCache),
    .io_alloc_4_bits_dirty(mshrAlloc_io_alloc_4_bits_dirty),
    .io_alloc_4_bits_fromProbeHelper(mshrAlloc_io_alloc_4_bits_fromProbeHelper),
    .io_alloc_4_bits_fromCmoHelper(mshrAlloc_io_alloc_4_bits_fromCmoHelper),
    .io_alloc_4_bits_needProbeAckData(mshrAlloc_io_alloc_4_bits_needProbeAckData),
    .io_alloc_5_valid(mshrAlloc_io_alloc_5_valid),
    .io_alloc_5_bits_channel(mshrAlloc_io_alloc_5_bits_channel),
    .io_alloc_5_bits_opcode(mshrAlloc_io_alloc_5_bits_opcode),
    .io_alloc_5_bits_param(mshrAlloc_io_alloc_5_bits_param),
    .io_alloc_5_bits_size(mshrAlloc_io_alloc_5_bits_size),
    .io_alloc_5_bits_source(mshrAlloc_io_alloc_5_bits_source),
    .io_alloc_5_bits_set(mshrAlloc_io_alloc_5_bits_set),
    .io_alloc_5_bits_tag(mshrAlloc_io_alloc_5_bits_tag),
    .io_alloc_5_bits_off(mshrAlloc_io_alloc_5_bits_off),
    .io_alloc_5_bits_mask(mshrAlloc_io_alloc_5_bits_mask),
    .io_alloc_5_bits_bufIdx(mshrAlloc_io_alloc_5_bits_bufIdx),
    .io_alloc_5_bits_preferCache(mshrAlloc_io_alloc_5_bits_preferCache),
    .io_alloc_5_bits_dirty(mshrAlloc_io_alloc_5_bits_dirty),
    .io_alloc_5_bits_fromProbeHelper(mshrAlloc_io_alloc_5_bits_fromProbeHelper),
    .io_alloc_5_bits_fromCmoHelper(mshrAlloc_io_alloc_5_bits_fromCmoHelper),
    .io_alloc_5_bits_needProbeAckData(mshrAlloc_io_alloc_5_bits_needProbeAckData),
    .io_alloc_6_valid(mshrAlloc_io_alloc_6_valid),
    .io_alloc_6_bits_channel(mshrAlloc_io_alloc_6_bits_channel),
    .io_alloc_6_bits_opcode(mshrAlloc_io_alloc_6_bits_opcode),
    .io_alloc_6_bits_param(mshrAlloc_io_alloc_6_bits_param),
    .io_alloc_6_bits_size(mshrAlloc_io_alloc_6_bits_size),
    .io_alloc_6_bits_source(mshrAlloc_io_alloc_6_bits_source),
    .io_alloc_6_bits_set(mshrAlloc_io_alloc_6_bits_set),
    .io_alloc_6_bits_tag(mshrAlloc_io_alloc_6_bits_tag),
    .io_alloc_6_bits_off(mshrAlloc_io_alloc_6_bits_off),
    .io_alloc_6_bits_mask(mshrAlloc_io_alloc_6_bits_mask),
    .io_alloc_6_bits_bufIdx(mshrAlloc_io_alloc_6_bits_bufIdx),
    .io_alloc_6_bits_preferCache(mshrAlloc_io_alloc_6_bits_preferCache),
    .io_alloc_6_bits_dirty(mshrAlloc_io_alloc_6_bits_dirty),
    .io_alloc_6_bits_fromProbeHelper(mshrAlloc_io_alloc_6_bits_fromProbeHelper),
    .io_alloc_6_bits_fromCmoHelper(mshrAlloc_io_alloc_6_bits_fromCmoHelper),
    .io_alloc_6_bits_needProbeAckData(mshrAlloc_io_alloc_6_bits_needProbeAckData),
    .io_alloc_7_valid(mshrAlloc_io_alloc_7_valid),
    .io_alloc_7_bits_channel(mshrAlloc_io_alloc_7_bits_channel),
    .io_alloc_7_bits_opcode(mshrAlloc_io_alloc_7_bits_opcode),
    .io_alloc_7_bits_param(mshrAlloc_io_alloc_7_bits_param),
    .io_alloc_7_bits_size(mshrAlloc_io_alloc_7_bits_size),
    .io_alloc_7_bits_source(mshrAlloc_io_alloc_7_bits_source),
    .io_alloc_7_bits_set(mshrAlloc_io_alloc_7_bits_set),
    .io_alloc_7_bits_tag(mshrAlloc_io_alloc_7_bits_tag),
    .io_alloc_7_bits_off(mshrAlloc_io_alloc_7_bits_off),
    .io_alloc_7_bits_mask(mshrAlloc_io_alloc_7_bits_mask),
    .io_alloc_7_bits_bufIdx(mshrAlloc_io_alloc_7_bits_bufIdx),
    .io_alloc_7_bits_preferCache(mshrAlloc_io_alloc_7_bits_preferCache),
    .io_alloc_7_bits_dirty(mshrAlloc_io_alloc_7_bits_dirty),
    .io_alloc_7_bits_fromProbeHelper(mshrAlloc_io_alloc_7_bits_fromProbeHelper),
    .io_alloc_7_bits_fromCmoHelper(mshrAlloc_io_alloc_7_bits_fromCmoHelper),
    .io_alloc_7_bits_needProbeAckData(mshrAlloc_io_alloc_7_bits_needProbeAckData),
    .io_alloc_8_valid(mshrAlloc_io_alloc_8_valid),
    .io_alloc_8_bits_channel(mshrAlloc_io_alloc_8_bits_channel),
    .io_alloc_8_bits_opcode(mshrAlloc_io_alloc_8_bits_opcode),
    .io_alloc_8_bits_param(mshrAlloc_io_alloc_8_bits_param),
    .io_alloc_8_bits_size(mshrAlloc_io_alloc_8_bits_size),
    .io_alloc_8_bits_source(mshrAlloc_io_alloc_8_bits_source),
    .io_alloc_8_bits_set(mshrAlloc_io_alloc_8_bits_set),
    .io_alloc_8_bits_tag(mshrAlloc_io_alloc_8_bits_tag),
    .io_alloc_8_bits_off(mshrAlloc_io_alloc_8_bits_off),
    .io_alloc_8_bits_mask(mshrAlloc_io_alloc_8_bits_mask),
    .io_alloc_8_bits_bufIdx(mshrAlloc_io_alloc_8_bits_bufIdx),
    .io_alloc_8_bits_preferCache(mshrAlloc_io_alloc_8_bits_preferCache),
    .io_alloc_8_bits_dirty(mshrAlloc_io_alloc_8_bits_dirty),
    .io_alloc_8_bits_fromProbeHelper(mshrAlloc_io_alloc_8_bits_fromProbeHelper),
    .io_alloc_8_bits_fromCmoHelper(mshrAlloc_io_alloc_8_bits_fromCmoHelper),
    .io_alloc_8_bits_needProbeAckData(mshrAlloc_io_alloc_8_bits_needProbeAckData),
    .io_alloc_9_valid(mshrAlloc_io_alloc_9_valid),
    .io_alloc_9_bits_channel(mshrAlloc_io_alloc_9_bits_channel),
    .io_alloc_9_bits_opcode(mshrAlloc_io_alloc_9_bits_opcode),
    .io_alloc_9_bits_param(mshrAlloc_io_alloc_9_bits_param),
    .io_alloc_9_bits_size(mshrAlloc_io_alloc_9_bits_size),
    .io_alloc_9_bits_source(mshrAlloc_io_alloc_9_bits_source),
    .io_alloc_9_bits_set(mshrAlloc_io_alloc_9_bits_set),
    .io_alloc_9_bits_tag(mshrAlloc_io_alloc_9_bits_tag),
    .io_alloc_9_bits_off(mshrAlloc_io_alloc_9_bits_off),
    .io_alloc_9_bits_mask(mshrAlloc_io_alloc_9_bits_mask),
    .io_alloc_9_bits_bufIdx(mshrAlloc_io_alloc_9_bits_bufIdx),
    .io_alloc_9_bits_preferCache(mshrAlloc_io_alloc_9_bits_preferCache),
    .io_alloc_9_bits_dirty(mshrAlloc_io_alloc_9_bits_dirty),
    .io_alloc_9_bits_fromProbeHelper(mshrAlloc_io_alloc_9_bits_fromProbeHelper),
    .io_alloc_9_bits_fromCmoHelper(mshrAlloc_io_alloc_9_bits_fromCmoHelper),
    .io_alloc_9_bits_needProbeAckData(mshrAlloc_io_alloc_9_bits_needProbeAckData),
    .io_alloc_10_valid(mshrAlloc_io_alloc_10_valid),
    .io_alloc_10_bits_channel(mshrAlloc_io_alloc_10_bits_channel),
    .io_alloc_10_bits_opcode(mshrAlloc_io_alloc_10_bits_opcode),
    .io_alloc_10_bits_param(mshrAlloc_io_alloc_10_bits_param),
    .io_alloc_10_bits_size(mshrAlloc_io_alloc_10_bits_size),
    .io_alloc_10_bits_source(mshrAlloc_io_alloc_10_bits_source),
    .io_alloc_10_bits_set(mshrAlloc_io_alloc_10_bits_set),
    .io_alloc_10_bits_tag(mshrAlloc_io_alloc_10_bits_tag),
    .io_alloc_10_bits_off(mshrAlloc_io_alloc_10_bits_off),
    .io_alloc_10_bits_mask(mshrAlloc_io_alloc_10_bits_mask),
    .io_alloc_10_bits_bufIdx(mshrAlloc_io_alloc_10_bits_bufIdx),
    .io_alloc_10_bits_preferCache(mshrAlloc_io_alloc_10_bits_preferCache),
    .io_alloc_10_bits_dirty(mshrAlloc_io_alloc_10_bits_dirty),
    .io_alloc_10_bits_fromProbeHelper(mshrAlloc_io_alloc_10_bits_fromProbeHelper),
    .io_alloc_10_bits_fromCmoHelper(mshrAlloc_io_alloc_10_bits_fromCmoHelper),
    .io_alloc_10_bits_needProbeAckData(mshrAlloc_io_alloc_10_bits_needProbeAckData),
    .io_alloc_11_valid(mshrAlloc_io_alloc_11_valid),
    .io_alloc_11_bits_channel(mshrAlloc_io_alloc_11_bits_channel),
    .io_alloc_11_bits_opcode(mshrAlloc_io_alloc_11_bits_opcode),
    .io_alloc_11_bits_param(mshrAlloc_io_alloc_11_bits_param),
    .io_alloc_11_bits_size(mshrAlloc_io_alloc_11_bits_size),
    .io_alloc_11_bits_source(mshrAlloc_io_alloc_11_bits_source),
    .io_alloc_11_bits_set(mshrAlloc_io_alloc_11_bits_set),
    .io_alloc_11_bits_tag(mshrAlloc_io_alloc_11_bits_tag),
    .io_alloc_11_bits_off(mshrAlloc_io_alloc_11_bits_off),
    .io_alloc_11_bits_mask(mshrAlloc_io_alloc_11_bits_mask),
    .io_alloc_11_bits_bufIdx(mshrAlloc_io_alloc_11_bits_bufIdx),
    .io_alloc_11_bits_preferCache(mshrAlloc_io_alloc_11_bits_preferCache),
    .io_alloc_11_bits_dirty(mshrAlloc_io_alloc_11_bits_dirty),
    .io_alloc_11_bits_fromProbeHelper(mshrAlloc_io_alloc_11_bits_fromProbeHelper),
    .io_alloc_11_bits_fromCmoHelper(mshrAlloc_io_alloc_11_bits_fromCmoHelper),
    .io_alloc_11_bits_needProbeAckData(mshrAlloc_io_alloc_11_bits_needProbeAckData),
    .io_alloc_12_valid(mshrAlloc_io_alloc_12_valid),
    .io_alloc_12_bits_channel(mshrAlloc_io_alloc_12_bits_channel),
    .io_alloc_12_bits_opcode(mshrAlloc_io_alloc_12_bits_opcode),
    .io_alloc_12_bits_param(mshrAlloc_io_alloc_12_bits_param),
    .io_alloc_12_bits_size(mshrAlloc_io_alloc_12_bits_size),
    .io_alloc_12_bits_source(mshrAlloc_io_alloc_12_bits_source),
    .io_alloc_12_bits_set(mshrAlloc_io_alloc_12_bits_set),
    .io_alloc_12_bits_tag(mshrAlloc_io_alloc_12_bits_tag),
    .io_alloc_12_bits_off(mshrAlloc_io_alloc_12_bits_off),
    .io_alloc_12_bits_mask(mshrAlloc_io_alloc_12_bits_mask),
    .io_alloc_12_bits_bufIdx(mshrAlloc_io_alloc_12_bits_bufIdx),
    .io_alloc_12_bits_preferCache(mshrAlloc_io_alloc_12_bits_preferCache),
    .io_alloc_12_bits_dirty(mshrAlloc_io_alloc_12_bits_dirty),
    .io_alloc_12_bits_fromProbeHelper(mshrAlloc_io_alloc_12_bits_fromProbeHelper),
    .io_alloc_12_bits_fromCmoHelper(mshrAlloc_io_alloc_12_bits_fromCmoHelper),
    .io_alloc_12_bits_needProbeAckData(mshrAlloc_io_alloc_12_bits_needProbeAckData),
    .io_alloc_13_valid(mshrAlloc_io_alloc_13_valid),
    .io_alloc_13_bits_channel(mshrAlloc_io_alloc_13_bits_channel),
    .io_alloc_13_bits_opcode(mshrAlloc_io_alloc_13_bits_opcode),
    .io_alloc_13_bits_param(mshrAlloc_io_alloc_13_bits_param),
    .io_alloc_13_bits_size(mshrAlloc_io_alloc_13_bits_size),
    .io_alloc_13_bits_source(mshrAlloc_io_alloc_13_bits_source),
    .io_alloc_13_bits_set(mshrAlloc_io_alloc_13_bits_set),
    .io_alloc_13_bits_tag(mshrAlloc_io_alloc_13_bits_tag),
    .io_alloc_13_bits_off(mshrAlloc_io_alloc_13_bits_off),
    .io_alloc_13_bits_mask(mshrAlloc_io_alloc_13_bits_mask),
    .io_alloc_13_bits_bufIdx(mshrAlloc_io_alloc_13_bits_bufIdx),
    .io_alloc_13_bits_preferCache(mshrAlloc_io_alloc_13_bits_preferCache),
    .io_alloc_13_bits_dirty(mshrAlloc_io_alloc_13_bits_dirty),
    .io_alloc_13_bits_fromProbeHelper(mshrAlloc_io_alloc_13_bits_fromProbeHelper),
    .io_alloc_13_bits_fromCmoHelper(mshrAlloc_io_alloc_13_bits_fromCmoHelper),
    .io_alloc_13_bits_needProbeAckData(mshrAlloc_io_alloc_13_bits_needProbeAckData),
    .io_alloc_14_valid(mshrAlloc_io_alloc_14_valid),
    .io_alloc_14_bits_channel(mshrAlloc_io_alloc_14_bits_channel),
    .io_alloc_14_bits_opcode(mshrAlloc_io_alloc_14_bits_opcode),
    .io_alloc_14_bits_param(mshrAlloc_io_alloc_14_bits_param),
    .io_alloc_14_bits_size(mshrAlloc_io_alloc_14_bits_size),
    .io_alloc_14_bits_source(mshrAlloc_io_alloc_14_bits_source),
    .io_alloc_14_bits_set(mshrAlloc_io_alloc_14_bits_set),
    .io_alloc_14_bits_tag(mshrAlloc_io_alloc_14_bits_tag),
    .io_alloc_14_bits_off(mshrAlloc_io_alloc_14_bits_off),
    .io_alloc_14_bits_mask(mshrAlloc_io_alloc_14_bits_mask),
    .io_alloc_14_bits_bufIdx(mshrAlloc_io_alloc_14_bits_bufIdx),
    .io_alloc_14_bits_preferCache(mshrAlloc_io_alloc_14_bits_preferCache),
    .io_alloc_14_bits_dirty(mshrAlloc_io_alloc_14_bits_dirty),
    .io_alloc_14_bits_fromProbeHelper(mshrAlloc_io_alloc_14_bits_fromProbeHelper),
    .io_alloc_14_bits_fromCmoHelper(mshrAlloc_io_alloc_14_bits_fromCmoHelper),
    .io_alloc_14_bits_needProbeAckData(mshrAlloc_io_alloc_14_bits_needProbeAckData),
    .io_alloc_15_valid(mshrAlloc_io_alloc_15_valid),
    .io_alloc_15_bits_opcode(mshrAlloc_io_alloc_15_bits_opcode),
    .io_alloc_15_bits_param(mshrAlloc_io_alloc_15_bits_param),
    .io_alloc_15_bits_size(mshrAlloc_io_alloc_15_bits_size),
    .io_alloc_15_bits_source(mshrAlloc_io_alloc_15_bits_source),
    .io_alloc_15_bits_set(mshrAlloc_io_alloc_15_bits_set),
    .io_alloc_15_bits_tag(mshrAlloc_io_alloc_15_bits_tag),
    .io_alloc_15_bits_off(mshrAlloc_io_alloc_15_bits_off),
    .io_alloc_15_bits_bufIdx(mshrAlloc_io_alloc_15_bits_bufIdx),
    .io_alloc_15_bits_dirty(mshrAlloc_io_alloc_15_bits_dirty),
    .io_dirRead_ready(mshrAlloc_io_dirRead_ready),
    .io_dirRead_valid(mshrAlloc_io_dirRead_valid),
    .io_dirRead_bits_idOH(mshrAlloc_io_dirRead_bits_idOH),
    .io_dirRead_bits_tag(mshrAlloc_io_dirRead_bits_tag),
    .io_dirRead_bits_set(mshrAlloc_io_dirRead_bits_set),
    .io_dirRead_bits_replacerInfo_channel(mshrAlloc_io_dirRead_bits_replacerInfo_channel),
    .io_dirRead_bits_replacerInfo_opcode(mshrAlloc_io_dirRead_bits_replacerInfo_opcode),
    .io_dirRead_bits_source(mshrAlloc_io_dirRead_bits_source),
    .io_bc_mask_valid(mshrAlloc_io_bc_mask_valid),
    .io_bc_mask_bits_0(mshrAlloc_io_bc_mask_bits_0),
    .io_bc_mask_bits_1(mshrAlloc_io_bc_mask_bits_1),
    .io_bc_mask_bits_2(mshrAlloc_io_bc_mask_bits_2),
    .io_bc_mask_bits_3(mshrAlloc_io_bc_mask_bits_3),
    .io_bc_mask_bits_4(mshrAlloc_io_bc_mask_bits_4),
    .io_bc_mask_bits_5(mshrAlloc_io_bc_mask_bits_5),
    .io_bc_mask_bits_6(mshrAlloc_io_bc_mask_bits_6),
    .io_bc_mask_bits_7(mshrAlloc_io_bc_mask_bits_7),
    .io_bc_mask_bits_8(mshrAlloc_io_bc_mask_bits_8),
    .io_bc_mask_bits_9(mshrAlloc_io_bc_mask_bits_9),
    .io_bc_mask_bits_10(mshrAlloc_io_bc_mask_bits_10),
    .io_bc_mask_bits_11(mshrAlloc_io_bc_mask_bits_11),
    .io_bc_mask_bits_12(mshrAlloc_io_bc_mask_bits_12),
    .io_bc_mask_bits_13(mshrAlloc_io_bc_mask_bits_13),
    .io_c_mask_valid(mshrAlloc_io_c_mask_valid),
    .io_c_mask_bits_0(mshrAlloc_io_c_mask_bits_0),
    .io_c_mask_bits_1(mshrAlloc_io_c_mask_bits_1),
    .io_c_mask_bits_2(mshrAlloc_io_c_mask_bits_2),
    .io_c_mask_bits_3(mshrAlloc_io_c_mask_bits_3),
    .io_c_mask_bits_4(mshrAlloc_io_c_mask_bits_4),
    .io_c_mask_bits_5(mshrAlloc_io_c_mask_bits_5),
    .io_c_mask_bits_6(mshrAlloc_io_c_mask_bits_6),
    .io_c_mask_bits_7(mshrAlloc_io_c_mask_bits_7),
    .io_c_mask_bits_8(mshrAlloc_io_c_mask_bits_8),
    .io_c_mask_bits_9(mshrAlloc_io_c_mask_bits_9),
    .io_c_mask_bits_10(mshrAlloc_io_c_mask_bits_10),
    .io_c_mask_bits_11(mshrAlloc_io_c_mask_bits_11),
    .io_c_mask_bits_12(mshrAlloc_io_c_mask_bits_12),
    .io_c_mask_bits_13(mshrAlloc_io_c_mask_bits_13),
    .io_c_mask_bits_14(mshrAlloc_io_c_mask_bits_14)
  );
  RequestBuffer a_req_buffer ( // @[Slice.scala 124:28]
    .clock(a_req_buffer_clock),
    .reset(a_req_buffer_reset),
    .io_in_ready(a_req_buffer_io_in_ready),
    .io_in_valid(a_req_buffer_io_in_valid),
    .io_in_bits_opcode(a_req_buffer_io_in_bits_opcode),
    .io_in_bits_param(a_req_buffer_io_in_bits_param),
    .io_in_bits_size(a_req_buffer_io_in_bits_size),
    .io_in_bits_source(a_req_buffer_io_in_bits_source),
    .io_in_bits_set(a_req_buffer_io_in_bits_set),
    .io_in_bits_tag(a_req_buffer_io_in_bits_tag),
    .io_in_bits_off(a_req_buffer_io_in_bits_off),
    .io_in_bits_mask(a_req_buffer_io_in_bits_mask),
    .io_in_bits_bufIdx(a_req_buffer_io_in_bits_bufIdx),
    .io_in_bits_preferCache(a_req_buffer_io_in_bits_preferCache),
    .io_out_ready(a_req_buffer_io_out_ready),
    .io_out_valid(a_req_buffer_io_out_valid),
    .io_out_bits_channel(a_req_buffer_io_out_bits_channel),
    .io_out_bits_opcode(a_req_buffer_io_out_bits_opcode),
    .io_out_bits_param(a_req_buffer_io_out_bits_param),
    .io_out_bits_size(a_req_buffer_io_out_bits_size),
    .io_out_bits_source(a_req_buffer_io_out_bits_source),
    .io_out_bits_set(a_req_buffer_io_out_bits_set),
    .io_out_bits_tag(a_req_buffer_io_out_bits_tag),
    .io_out_bits_off(a_req_buffer_io_out_bits_off),
    .io_out_bits_mask(a_req_buffer_io_out_bits_mask),
    .io_out_bits_bufIdx(a_req_buffer_io_out_bits_bufIdx),
    .io_out_bits_preferCache(a_req_buffer_io_out_bits_preferCache),
    .io_out_bits_dirty(a_req_buffer_io_out_bits_dirty),
    .io_out_bits_fromProbeHelper(a_req_buffer_io_out_bits_fromProbeHelper),
    .io_out_bits_fromCmoHelper(a_req_buffer_io_out_bits_fromCmoHelper),
    .io_out_bits_needProbeAckData(a_req_buffer_io_out_bits_needProbeAckData),
    .io_mshr_status_0_valid(a_req_buffer_io_mshr_status_0_valid),
    .io_mshr_status_0_bits_set(a_req_buffer_io_mshr_status_0_bits_set),
    .io_mshr_status_0_bits_will_free(a_req_buffer_io_mshr_status_0_bits_will_free),
    .io_mshr_status_1_valid(a_req_buffer_io_mshr_status_1_valid),
    .io_mshr_status_1_bits_set(a_req_buffer_io_mshr_status_1_bits_set),
    .io_mshr_status_1_bits_will_free(a_req_buffer_io_mshr_status_1_bits_will_free),
    .io_mshr_status_2_valid(a_req_buffer_io_mshr_status_2_valid),
    .io_mshr_status_2_bits_set(a_req_buffer_io_mshr_status_2_bits_set),
    .io_mshr_status_2_bits_will_free(a_req_buffer_io_mshr_status_2_bits_will_free),
    .io_mshr_status_3_valid(a_req_buffer_io_mshr_status_3_valid),
    .io_mshr_status_3_bits_set(a_req_buffer_io_mshr_status_3_bits_set),
    .io_mshr_status_3_bits_will_free(a_req_buffer_io_mshr_status_3_bits_will_free),
    .io_mshr_status_4_valid(a_req_buffer_io_mshr_status_4_valid),
    .io_mshr_status_4_bits_set(a_req_buffer_io_mshr_status_4_bits_set),
    .io_mshr_status_4_bits_will_free(a_req_buffer_io_mshr_status_4_bits_will_free),
    .io_mshr_status_5_valid(a_req_buffer_io_mshr_status_5_valid),
    .io_mshr_status_5_bits_set(a_req_buffer_io_mshr_status_5_bits_set),
    .io_mshr_status_5_bits_will_free(a_req_buffer_io_mshr_status_5_bits_will_free),
    .io_mshr_status_6_valid(a_req_buffer_io_mshr_status_6_valid),
    .io_mshr_status_6_bits_set(a_req_buffer_io_mshr_status_6_bits_set),
    .io_mshr_status_6_bits_will_free(a_req_buffer_io_mshr_status_6_bits_will_free),
    .io_mshr_status_7_valid(a_req_buffer_io_mshr_status_7_valid),
    .io_mshr_status_7_bits_set(a_req_buffer_io_mshr_status_7_bits_set),
    .io_mshr_status_7_bits_will_free(a_req_buffer_io_mshr_status_7_bits_will_free),
    .io_mshr_status_8_valid(a_req_buffer_io_mshr_status_8_valid),
    .io_mshr_status_8_bits_set(a_req_buffer_io_mshr_status_8_bits_set),
    .io_mshr_status_8_bits_will_free(a_req_buffer_io_mshr_status_8_bits_will_free),
    .io_mshr_status_9_valid(a_req_buffer_io_mshr_status_9_valid),
    .io_mshr_status_9_bits_set(a_req_buffer_io_mshr_status_9_bits_set),
    .io_mshr_status_9_bits_will_free(a_req_buffer_io_mshr_status_9_bits_will_free),
    .io_mshr_status_10_valid(a_req_buffer_io_mshr_status_10_valid),
    .io_mshr_status_10_bits_set(a_req_buffer_io_mshr_status_10_bits_set),
    .io_mshr_status_10_bits_will_free(a_req_buffer_io_mshr_status_10_bits_will_free),
    .io_mshr_status_11_valid(a_req_buffer_io_mshr_status_11_valid),
    .io_mshr_status_11_bits_set(a_req_buffer_io_mshr_status_11_bits_set),
    .io_mshr_status_11_bits_will_free(a_req_buffer_io_mshr_status_11_bits_will_free),
    .io_mshr_status_12_valid(a_req_buffer_io_mshr_status_12_valid),
    .io_mshr_status_12_bits_set(a_req_buffer_io_mshr_status_12_bits_set),
    .io_mshr_status_12_bits_will_free(a_req_buffer_io_mshr_status_12_bits_will_free),
    .io_mshr_status_13_valid(a_req_buffer_io_mshr_status_13_valid),
    .io_mshr_status_13_bits_set(a_req_buffer_io_mshr_status_13_bits_set),
    .io_mshr_status_13_bits_will_free(a_req_buffer_io_mshr_status_13_bits_will_free)
  );
  ProbeHelper probeHelperOpt ( // @[Slice.scala 126:16]
    .clock(probeHelperOpt_clock),
    .reset(probeHelperOpt_reset),
    .io_dirResult_valid(probeHelperOpt_io_dirResult_valid),
    .io_dirResult_bits_clients_states_0_state(probeHelperOpt_io_dirResult_bits_clients_states_0_state),
    .io_dirResult_bits_clients_states_0_hit(probeHelperOpt_io_dirResult_bits_clients_states_0_hit),
    .io_dirResult_bits_clients_states_1_state(probeHelperOpt_io_dirResult_bits_clients_states_1_state),
    .io_dirResult_bits_clients_states_1_hit(probeHelperOpt_io_dirResult_bits_clients_states_1_hit),
    .io_dirResult_bits_clients_tag_match(probeHelperOpt_io_dirResult_bits_clients_tag_match),
    .io_dirResult_bits_clients_tag(probeHelperOpt_io_dirResult_bits_clients_tag),
    .io_dirResult_bits_sourceId(probeHelperOpt_io_dirResult_bits_sourceId),
    .io_dirResult_bits_set(probeHelperOpt_io_dirResult_bits_set),
    .io_dirResult_bits_replacerInfo_channel(probeHelperOpt_io_dirResult_bits_replacerInfo_channel),
    .io_dirResult_bits_replacerInfo_opcode(probeHelperOpt_io_dirResult_bits_replacerInfo_opcode),
    .io_probe_ready(probeHelperOpt_io_probe_ready),
    .io_probe_valid(probeHelperOpt_io_probe_valid),
    .io_probe_bits_channel(probeHelperOpt_io_probe_bits_channel),
    .io_probe_bits_opcode(probeHelperOpt_io_probe_bits_opcode),
    .io_probe_bits_param(probeHelperOpt_io_probe_bits_param),
    .io_probe_bits_size(probeHelperOpt_io_probe_bits_size),
    .io_probe_bits_source(probeHelperOpt_io_probe_bits_source),
    .io_probe_bits_set(probeHelperOpt_io_probe_bits_set),
    .io_probe_bits_tag(probeHelperOpt_io_probe_bits_tag),
    .io_probe_bits_off(probeHelperOpt_io_probe_bits_off),
    .io_probe_bits_mask(probeHelperOpt_io_probe_bits_mask),
    .io_probe_bits_bufIdx(probeHelperOpt_io_probe_bits_bufIdx),
    .io_probe_bits_preferCache(probeHelperOpt_io_probe_bits_preferCache),
    .io_probe_bits_dirty(probeHelperOpt_io_probe_bits_dirty),
    .io_probe_bits_fromProbeHelper(probeHelperOpt_io_probe_bits_fromProbeHelper),
    .io_probe_bits_fromCmoHelper(probeHelperOpt_io_probe_bits_fromCmoHelper),
    .io_probe_bits_needProbeAckData(probeHelperOpt_io_probe_bits_needProbeAckData),
    .io_full(probeHelperOpt_io_full)
  );
  Arbiter_39 b_arb ( // @[Slice.scala 136:23]
    .io_in_0_ready(b_arb_io_in_0_ready),
    .io_in_0_valid(b_arb_io_in_0_valid),
    .io_in_0_bits_channel(b_arb_io_in_0_bits_channel),
    .io_in_0_bits_opcode(b_arb_io_in_0_bits_opcode),
    .io_in_0_bits_param(b_arb_io_in_0_bits_param),
    .io_in_0_bits_size(b_arb_io_in_0_bits_size),
    .io_in_0_bits_source(b_arb_io_in_0_bits_source),
    .io_in_0_bits_set(b_arb_io_in_0_bits_set),
    .io_in_0_bits_tag(b_arb_io_in_0_bits_tag),
    .io_in_0_bits_off(b_arb_io_in_0_bits_off),
    .io_in_0_bits_mask(b_arb_io_in_0_bits_mask),
    .io_in_0_bits_bufIdx(b_arb_io_in_0_bits_bufIdx),
    .io_in_0_bits_preferCache(b_arb_io_in_0_bits_preferCache),
    .io_in_0_bits_dirty(b_arb_io_in_0_bits_dirty),
    .io_in_0_bits_fromProbeHelper(b_arb_io_in_0_bits_fromProbeHelper),
    .io_in_0_bits_fromCmoHelper(b_arb_io_in_0_bits_fromCmoHelper),
    .io_in_0_bits_needProbeAckData(b_arb_io_in_0_bits_needProbeAckData),
    .io_in_1_ready(b_arb_io_in_1_ready),
    .io_in_1_valid(b_arb_io_in_1_valid),
    .io_in_1_bits_opcode(b_arb_io_in_1_bits_opcode),
    .io_in_1_bits_param(b_arb_io_in_1_bits_param),
    .io_in_1_bits_size(b_arb_io_in_1_bits_size),
    .io_in_1_bits_source(b_arb_io_in_1_bits_source),
    .io_in_1_bits_set(b_arb_io_in_1_bits_set),
    .io_in_1_bits_tag(b_arb_io_in_1_bits_tag),
    .io_in_1_bits_off(b_arb_io_in_1_bits_off),
    .io_in_1_bits_mask(b_arb_io_in_1_bits_mask),
    .io_in_1_bits_needProbeAckData(b_arb_io_in_1_bits_needProbeAckData),
    .io_out_ready(b_arb_io_out_ready),
    .io_out_valid(b_arb_io_out_valid),
    .io_out_bits_channel(b_arb_io_out_bits_channel),
    .io_out_bits_opcode(b_arb_io_out_bits_opcode),
    .io_out_bits_param(b_arb_io_out_bits_param),
    .io_out_bits_size(b_arb_io_out_bits_size),
    .io_out_bits_source(b_arb_io_out_bits_source),
    .io_out_bits_set(b_arb_io_out_bits_set),
    .io_out_bits_tag(b_arb_io_out_bits_tag),
    .io_out_bits_off(b_arb_io_out_bits_off),
    .io_out_bits_mask(b_arb_io_out_bits_mask),
    .io_out_bits_bufIdx(b_arb_io_out_bits_bufIdx),
    .io_out_bits_preferCache(b_arb_io_out_bits_preferCache),
    .io_out_bits_dirty(b_arb_io_out_bits_dirty),
    .io_out_bits_fromProbeHelper(b_arb_io_out_bits_fromProbeHelper),
    .io_out_bits_fromCmoHelper(b_arb_io_out_bits_fromCmoHelper),
    .io_out_bits_needProbeAckData(b_arb_io_out_bits_needProbeAckData)
  );
  Directory directory ( // @[Slice.scala 372:25]
    .clock(directory_clock),
    .reset(directory_reset),
    .io_read_ready(directory_io_read_ready),
    .io_read_valid(directory_io_read_valid),
    .io_read_bits_idOH(directory_io_read_bits_idOH),
    .io_read_bits_tag(directory_io_read_bits_tag),
    .io_read_bits_set(directory_io_read_bits_set),
    .io_read_bits_replacerInfo_channel(directory_io_read_bits_replacerInfo_channel),
    .io_read_bits_replacerInfo_opcode(directory_io_read_bits_replacerInfo_opcode),
    .io_read_bits_source(directory_io_read_bits_source),
    .io_result_valid(directory_io_result_valid),
    .io_result_bits_idOH(directory_io_result_bits_idOH),
    .io_result_bits_self_dirty(directory_io_result_bits_self_dirty),
    .io_result_bits_self_state(directory_io_result_bits_self_state),
    .io_result_bits_self_clientStates_0(directory_io_result_bits_self_clientStates_0),
    .io_result_bits_self_clientStates_1(directory_io_result_bits_self_clientStates_1),
    .io_result_bits_self_hit(directory_io_result_bits_self_hit),
    .io_result_bits_self_way(directory_io_result_bits_self_way),
    .io_result_bits_self_tag(directory_io_result_bits_self_tag),
    .io_result_bits_clients_states_0_state(directory_io_result_bits_clients_states_0_state),
    .io_result_bits_clients_states_0_hit(directory_io_result_bits_clients_states_0_hit),
    .io_result_bits_clients_states_1_state(directory_io_result_bits_clients_states_1_state),
    .io_result_bits_clients_states_1_hit(directory_io_result_bits_clients_states_1_hit),
    .io_result_bits_clients_tag_match(directory_io_result_bits_clients_tag_match),
    .io_result_bits_clients_tag(directory_io_result_bits_clients_tag),
    .io_result_bits_clients_way(directory_io_result_bits_clients_way),
    .io_result_bits_sourceId(directory_io_result_bits_sourceId),
    .io_result_bits_set(directory_io_result_bits_set),
    .io_result_bits_replacerInfo_channel(directory_io_result_bits_replacerInfo_channel),
    .io_result_bits_replacerInfo_opcode(directory_io_result_bits_replacerInfo_opcode),
    .io_dirWReq_valid(directory_io_dirWReq_valid),
    .io_dirWReq_bits_set(directory_io_dirWReq_bits_set),
    .io_dirWReq_bits_way(directory_io_dirWReq_bits_way),
    .io_dirWReq_bits_data_dirty(directory_io_dirWReq_bits_data_dirty),
    .io_dirWReq_bits_data_state(directory_io_dirWReq_bits_data_state),
    .io_dirWReq_bits_data_clientStates_0(directory_io_dirWReq_bits_data_clientStates_0),
    .io_dirWReq_bits_data_clientStates_1(directory_io_dirWReq_bits_data_clientStates_1),
    .io_tagWReq_valid(directory_io_tagWReq_valid),
    .io_tagWReq_bits_set(directory_io_tagWReq_bits_set),
    .io_tagWReq_bits_way(directory_io_tagWReq_bits_way),
    .io_tagWReq_bits_tag(directory_io_tagWReq_bits_tag),
    .io_clientDirWReq_valid(directory_io_clientDirWReq_valid),
    .io_clientDirWReq_bits_set(directory_io_clientDirWReq_bits_set),
    .io_clientDirWReq_bits_way(directory_io_clientDirWReq_bits_way),
    .io_clientDirWReq_bits_data_0_state(directory_io_clientDirWReq_bits_data_0_state),
    .io_clientDirWReq_bits_data_1_state(directory_io_clientDirWReq_bits_data_1_state),
    .io_clientTagWreq_valid(directory_io_clientTagWreq_valid),
    .io_clientTagWreq_bits_set(directory_io_clientTagWreq_bits_set),
    .io_clientTagWreq_bits_way(directory_io_clientTagWreq_bits_way),
    .io_clientTagWreq_bits_tag(directory_io_clientTagWreq_bits_tag)
  );
  Pipeline_1 pipeline ( // @[Pipeline.scala 39:26]
    .clock(pipeline_clock),
    .reset(pipeline_reset),
    .io_in_valid(pipeline_io_in_valid),
    .io_in_bits_set(pipeline_io_in_bits_set),
    .io_in_bits_way(pipeline_io_in_bits_way),
    .io_in_bits_data_dirty(pipeline_io_in_bits_data_dirty),
    .io_in_bits_data_state(pipeline_io_in_bits_data_state),
    .io_in_bits_data_clientStates_0(pipeline_io_in_bits_data_clientStates_0),
    .io_in_bits_data_clientStates_1(pipeline_io_in_bits_data_clientStates_1),
    .io_out_valid(pipeline_io_out_valid),
    .io_out_bits_set(pipeline_io_out_bits_set),
    .io_out_bits_way(pipeline_io_out_bits_way),
    .io_out_bits_data_dirty(pipeline_io_out_bits_data_dirty),
    .io_out_bits_data_state(pipeline_io_out_bits_data_state),
    .io_out_bits_data_clientStates_0(pipeline_io_out_bits_data_clientStates_0),
    .io_out_bits_data_clientStates_1(pipeline_io_out_bits_data_clientStates_1)
  );
  FastArbiter_2 arbiter ( // @[Slice.scala 405:25]
    .clock(arbiter_clock),
    .reset(arbiter_reset),
    .io_in_0_ready(arbiter_io_in_0_ready),
    .io_in_0_valid(arbiter_io_in_0_valid),
    .io_in_0_bits_set(arbiter_io_in_0_bits_set),
    .io_in_0_bits_way(arbiter_io_in_0_bits_way),
    .io_in_0_bits_data_dirty(arbiter_io_in_0_bits_data_dirty),
    .io_in_0_bits_data_state(arbiter_io_in_0_bits_data_state),
    .io_in_0_bits_data_clientStates_0(arbiter_io_in_0_bits_data_clientStates_0),
    .io_in_0_bits_data_clientStates_1(arbiter_io_in_0_bits_data_clientStates_1),
    .io_in_1_ready(arbiter_io_in_1_ready),
    .io_in_1_valid(arbiter_io_in_1_valid),
    .io_in_1_bits_set(arbiter_io_in_1_bits_set),
    .io_in_1_bits_way(arbiter_io_in_1_bits_way),
    .io_in_1_bits_data_dirty(arbiter_io_in_1_bits_data_dirty),
    .io_in_1_bits_data_state(arbiter_io_in_1_bits_data_state),
    .io_in_1_bits_data_clientStates_0(arbiter_io_in_1_bits_data_clientStates_0),
    .io_in_1_bits_data_clientStates_1(arbiter_io_in_1_bits_data_clientStates_1),
    .io_in_2_ready(arbiter_io_in_2_ready),
    .io_in_2_valid(arbiter_io_in_2_valid),
    .io_in_2_bits_set(arbiter_io_in_2_bits_set),
    .io_in_2_bits_way(arbiter_io_in_2_bits_way),
    .io_in_2_bits_data_dirty(arbiter_io_in_2_bits_data_dirty),
    .io_in_2_bits_data_state(arbiter_io_in_2_bits_data_state),
    .io_in_2_bits_data_clientStates_0(arbiter_io_in_2_bits_data_clientStates_0),
    .io_in_2_bits_data_clientStates_1(arbiter_io_in_2_bits_data_clientStates_1),
    .io_in_3_ready(arbiter_io_in_3_ready),
    .io_in_3_valid(arbiter_io_in_3_valid),
    .io_in_3_bits_set(arbiter_io_in_3_bits_set),
    .io_in_3_bits_way(arbiter_io_in_3_bits_way),
    .io_in_3_bits_data_dirty(arbiter_io_in_3_bits_data_dirty),
    .io_in_3_bits_data_state(arbiter_io_in_3_bits_data_state),
    .io_in_3_bits_data_clientStates_0(arbiter_io_in_3_bits_data_clientStates_0),
    .io_in_3_bits_data_clientStates_1(arbiter_io_in_3_bits_data_clientStates_1),
    .io_in_4_ready(arbiter_io_in_4_ready),
    .io_in_4_valid(arbiter_io_in_4_valid),
    .io_in_4_bits_set(arbiter_io_in_4_bits_set),
    .io_in_4_bits_way(arbiter_io_in_4_bits_way),
    .io_in_4_bits_data_dirty(arbiter_io_in_4_bits_data_dirty),
    .io_in_4_bits_data_state(arbiter_io_in_4_bits_data_state),
    .io_in_4_bits_data_clientStates_0(arbiter_io_in_4_bits_data_clientStates_0),
    .io_in_4_bits_data_clientStates_1(arbiter_io_in_4_bits_data_clientStates_1),
    .io_in_5_ready(arbiter_io_in_5_ready),
    .io_in_5_valid(arbiter_io_in_5_valid),
    .io_in_5_bits_set(arbiter_io_in_5_bits_set),
    .io_in_5_bits_way(arbiter_io_in_5_bits_way),
    .io_in_5_bits_data_dirty(arbiter_io_in_5_bits_data_dirty),
    .io_in_5_bits_data_state(arbiter_io_in_5_bits_data_state),
    .io_in_5_bits_data_clientStates_0(arbiter_io_in_5_bits_data_clientStates_0),
    .io_in_5_bits_data_clientStates_1(arbiter_io_in_5_bits_data_clientStates_1),
    .io_in_6_ready(arbiter_io_in_6_ready),
    .io_in_6_valid(arbiter_io_in_6_valid),
    .io_in_6_bits_set(arbiter_io_in_6_bits_set),
    .io_in_6_bits_way(arbiter_io_in_6_bits_way),
    .io_in_6_bits_data_dirty(arbiter_io_in_6_bits_data_dirty),
    .io_in_6_bits_data_state(arbiter_io_in_6_bits_data_state),
    .io_in_6_bits_data_clientStates_0(arbiter_io_in_6_bits_data_clientStates_0),
    .io_in_6_bits_data_clientStates_1(arbiter_io_in_6_bits_data_clientStates_1),
    .io_in_7_ready(arbiter_io_in_7_ready),
    .io_in_7_valid(arbiter_io_in_7_valid),
    .io_in_7_bits_set(arbiter_io_in_7_bits_set),
    .io_in_7_bits_way(arbiter_io_in_7_bits_way),
    .io_in_7_bits_data_dirty(arbiter_io_in_7_bits_data_dirty),
    .io_in_7_bits_data_state(arbiter_io_in_7_bits_data_state),
    .io_in_7_bits_data_clientStates_0(arbiter_io_in_7_bits_data_clientStates_0),
    .io_in_7_bits_data_clientStates_1(arbiter_io_in_7_bits_data_clientStates_1),
    .io_in_8_ready(arbiter_io_in_8_ready),
    .io_in_8_valid(arbiter_io_in_8_valid),
    .io_in_8_bits_set(arbiter_io_in_8_bits_set),
    .io_in_8_bits_way(arbiter_io_in_8_bits_way),
    .io_in_8_bits_data_dirty(arbiter_io_in_8_bits_data_dirty),
    .io_in_8_bits_data_state(arbiter_io_in_8_bits_data_state),
    .io_in_8_bits_data_clientStates_0(arbiter_io_in_8_bits_data_clientStates_0),
    .io_in_8_bits_data_clientStates_1(arbiter_io_in_8_bits_data_clientStates_1),
    .io_in_9_ready(arbiter_io_in_9_ready),
    .io_in_9_valid(arbiter_io_in_9_valid),
    .io_in_9_bits_set(arbiter_io_in_9_bits_set),
    .io_in_9_bits_way(arbiter_io_in_9_bits_way),
    .io_in_9_bits_data_dirty(arbiter_io_in_9_bits_data_dirty),
    .io_in_9_bits_data_state(arbiter_io_in_9_bits_data_state),
    .io_in_9_bits_data_clientStates_0(arbiter_io_in_9_bits_data_clientStates_0),
    .io_in_9_bits_data_clientStates_1(arbiter_io_in_9_bits_data_clientStates_1),
    .io_in_10_ready(arbiter_io_in_10_ready),
    .io_in_10_valid(arbiter_io_in_10_valid),
    .io_in_10_bits_set(arbiter_io_in_10_bits_set),
    .io_in_10_bits_way(arbiter_io_in_10_bits_way),
    .io_in_10_bits_data_dirty(arbiter_io_in_10_bits_data_dirty),
    .io_in_10_bits_data_state(arbiter_io_in_10_bits_data_state),
    .io_in_10_bits_data_clientStates_0(arbiter_io_in_10_bits_data_clientStates_0),
    .io_in_10_bits_data_clientStates_1(arbiter_io_in_10_bits_data_clientStates_1),
    .io_in_11_ready(arbiter_io_in_11_ready),
    .io_in_11_valid(arbiter_io_in_11_valid),
    .io_in_11_bits_set(arbiter_io_in_11_bits_set),
    .io_in_11_bits_way(arbiter_io_in_11_bits_way),
    .io_in_11_bits_data_dirty(arbiter_io_in_11_bits_data_dirty),
    .io_in_11_bits_data_state(arbiter_io_in_11_bits_data_state),
    .io_in_11_bits_data_clientStates_0(arbiter_io_in_11_bits_data_clientStates_0),
    .io_in_11_bits_data_clientStates_1(arbiter_io_in_11_bits_data_clientStates_1),
    .io_in_12_ready(arbiter_io_in_12_ready),
    .io_in_12_valid(arbiter_io_in_12_valid),
    .io_in_12_bits_set(arbiter_io_in_12_bits_set),
    .io_in_12_bits_way(arbiter_io_in_12_bits_way),
    .io_in_12_bits_data_dirty(arbiter_io_in_12_bits_data_dirty),
    .io_in_12_bits_data_state(arbiter_io_in_12_bits_data_state),
    .io_in_12_bits_data_clientStates_0(arbiter_io_in_12_bits_data_clientStates_0),
    .io_in_12_bits_data_clientStates_1(arbiter_io_in_12_bits_data_clientStates_1),
    .io_in_13_ready(arbiter_io_in_13_ready),
    .io_in_13_valid(arbiter_io_in_13_valid),
    .io_in_13_bits_set(arbiter_io_in_13_bits_set),
    .io_in_13_bits_way(arbiter_io_in_13_bits_way),
    .io_in_13_bits_data_dirty(arbiter_io_in_13_bits_data_dirty),
    .io_in_13_bits_data_state(arbiter_io_in_13_bits_data_state),
    .io_in_13_bits_data_clientStates_0(arbiter_io_in_13_bits_data_clientStates_0),
    .io_in_13_bits_data_clientStates_1(arbiter_io_in_13_bits_data_clientStates_1),
    .io_in_14_ready(arbiter_io_in_14_ready),
    .io_in_14_valid(arbiter_io_in_14_valid),
    .io_in_14_bits_set(arbiter_io_in_14_bits_set),
    .io_in_14_bits_way(arbiter_io_in_14_bits_way),
    .io_in_14_bits_data_dirty(arbiter_io_in_14_bits_data_dirty),
    .io_in_14_bits_data_state(arbiter_io_in_14_bits_data_state),
    .io_in_14_bits_data_clientStates_0(arbiter_io_in_14_bits_data_clientStates_0),
    .io_in_14_bits_data_clientStates_1(arbiter_io_in_14_bits_data_clientStates_1),
    .io_in_15_ready(arbiter_io_in_15_ready),
    .io_in_15_valid(arbiter_io_in_15_valid),
    .io_in_15_bits_set(arbiter_io_in_15_bits_set),
    .io_in_15_bits_way(arbiter_io_in_15_bits_way),
    .io_in_15_bits_data_dirty(arbiter_io_in_15_bits_data_dirty),
    .io_in_15_bits_data_state(arbiter_io_in_15_bits_data_state),
    .io_in_15_bits_data_clientStates_0(arbiter_io_in_15_bits_data_clientStates_0),
    .io_in_15_bits_data_clientStates_1(arbiter_io_in_15_bits_data_clientStates_1),
    .io_out_valid(arbiter_io_out_valid),
    .io_out_bits_set(arbiter_io_out_bits_set),
    .io_out_bits_way(arbiter_io_out_bits_way),
    .io_out_bits_data_dirty(arbiter_io_out_bits_data_dirty),
    .io_out_bits_data_state(arbiter_io_out_bits_data_state),
    .io_out_bits_data_clientStates_0(arbiter_io_out_bits_data_clientStates_0),
    .io_out_bits_data_clientStates_1(arbiter_io_out_bits_data_clientStates_1)
  );
  LatchFastArbiter sourceA_task_arb ( // @[Slice.scala 468:27]
    .clock(sourceA_task_arb_clock),
    .reset(sourceA_task_arb_reset),
    .io_in_0_ready(sourceA_task_arb_io_in_0_ready),
    .io_in_0_valid(sourceA_task_arb_io_in_0_valid),
    .io_in_0_bits_tag(sourceA_task_arb_io_in_0_bits_tag),
    .io_in_0_bits_set(sourceA_task_arb_io_in_0_bits_set),
    .io_in_0_bits_off(sourceA_task_arb_io_in_0_bits_off),
    .io_in_0_bits_opcode(sourceA_task_arb_io_in_0_bits_opcode),
    .io_in_0_bits_param(sourceA_task_arb_io_in_0_bits_param),
    .io_in_0_bits_source(sourceA_task_arb_io_in_0_bits_source),
    .io_in_0_bits_bufIdx(sourceA_task_arb_io_in_0_bits_bufIdx),
    .io_in_0_bits_size(sourceA_task_arb_io_in_0_bits_size),
    .io_in_0_bits_putData(sourceA_task_arb_io_in_0_bits_putData),
    .io_in_1_ready(sourceA_task_arb_io_in_1_ready),
    .io_in_1_valid(sourceA_task_arb_io_in_1_valid),
    .io_in_1_bits_tag(sourceA_task_arb_io_in_1_bits_tag),
    .io_in_1_bits_set(sourceA_task_arb_io_in_1_bits_set),
    .io_in_1_bits_off(sourceA_task_arb_io_in_1_bits_off),
    .io_in_1_bits_opcode(sourceA_task_arb_io_in_1_bits_opcode),
    .io_in_1_bits_param(sourceA_task_arb_io_in_1_bits_param),
    .io_in_1_bits_source(sourceA_task_arb_io_in_1_bits_source),
    .io_in_1_bits_bufIdx(sourceA_task_arb_io_in_1_bits_bufIdx),
    .io_in_1_bits_size(sourceA_task_arb_io_in_1_bits_size),
    .io_in_1_bits_putData(sourceA_task_arb_io_in_1_bits_putData),
    .io_in_2_ready(sourceA_task_arb_io_in_2_ready),
    .io_in_2_valid(sourceA_task_arb_io_in_2_valid),
    .io_in_2_bits_tag(sourceA_task_arb_io_in_2_bits_tag),
    .io_in_2_bits_set(sourceA_task_arb_io_in_2_bits_set),
    .io_in_2_bits_off(sourceA_task_arb_io_in_2_bits_off),
    .io_in_2_bits_opcode(sourceA_task_arb_io_in_2_bits_opcode),
    .io_in_2_bits_param(sourceA_task_arb_io_in_2_bits_param),
    .io_in_2_bits_source(sourceA_task_arb_io_in_2_bits_source),
    .io_in_2_bits_bufIdx(sourceA_task_arb_io_in_2_bits_bufIdx),
    .io_in_2_bits_size(sourceA_task_arb_io_in_2_bits_size),
    .io_in_2_bits_putData(sourceA_task_arb_io_in_2_bits_putData),
    .io_in_3_ready(sourceA_task_arb_io_in_3_ready),
    .io_in_3_valid(sourceA_task_arb_io_in_3_valid),
    .io_in_3_bits_tag(sourceA_task_arb_io_in_3_bits_tag),
    .io_in_3_bits_set(sourceA_task_arb_io_in_3_bits_set),
    .io_in_3_bits_off(sourceA_task_arb_io_in_3_bits_off),
    .io_in_3_bits_opcode(sourceA_task_arb_io_in_3_bits_opcode),
    .io_in_3_bits_param(sourceA_task_arb_io_in_3_bits_param),
    .io_in_3_bits_source(sourceA_task_arb_io_in_3_bits_source),
    .io_in_3_bits_bufIdx(sourceA_task_arb_io_in_3_bits_bufIdx),
    .io_in_3_bits_size(sourceA_task_arb_io_in_3_bits_size),
    .io_in_3_bits_putData(sourceA_task_arb_io_in_3_bits_putData),
    .io_in_4_ready(sourceA_task_arb_io_in_4_ready),
    .io_in_4_valid(sourceA_task_arb_io_in_4_valid),
    .io_in_4_bits_tag(sourceA_task_arb_io_in_4_bits_tag),
    .io_in_4_bits_set(sourceA_task_arb_io_in_4_bits_set),
    .io_in_4_bits_off(sourceA_task_arb_io_in_4_bits_off),
    .io_in_4_bits_opcode(sourceA_task_arb_io_in_4_bits_opcode),
    .io_in_4_bits_param(sourceA_task_arb_io_in_4_bits_param),
    .io_in_4_bits_source(sourceA_task_arb_io_in_4_bits_source),
    .io_in_4_bits_bufIdx(sourceA_task_arb_io_in_4_bits_bufIdx),
    .io_in_4_bits_size(sourceA_task_arb_io_in_4_bits_size),
    .io_in_4_bits_putData(sourceA_task_arb_io_in_4_bits_putData),
    .io_in_5_ready(sourceA_task_arb_io_in_5_ready),
    .io_in_5_valid(sourceA_task_arb_io_in_5_valid),
    .io_in_5_bits_tag(sourceA_task_arb_io_in_5_bits_tag),
    .io_in_5_bits_set(sourceA_task_arb_io_in_5_bits_set),
    .io_in_5_bits_off(sourceA_task_arb_io_in_5_bits_off),
    .io_in_5_bits_opcode(sourceA_task_arb_io_in_5_bits_opcode),
    .io_in_5_bits_param(sourceA_task_arb_io_in_5_bits_param),
    .io_in_5_bits_source(sourceA_task_arb_io_in_5_bits_source),
    .io_in_5_bits_bufIdx(sourceA_task_arb_io_in_5_bits_bufIdx),
    .io_in_5_bits_size(sourceA_task_arb_io_in_5_bits_size),
    .io_in_5_bits_putData(sourceA_task_arb_io_in_5_bits_putData),
    .io_in_6_ready(sourceA_task_arb_io_in_6_ready),
    .io_in_6_valid(sourceA_task_arb_io_in_6_valid),
    .io_in_6_bits_tag(sourceA_task_arb_io_in_6_bits_tag),
    .io_in_6_bits_set(sourceA_task_arb_io_in_6_bits_set),
    .io_in_6_bits_off(sourceA_task_arb_io_in_6_bits_off),
    .io_in_6_bits_opcode(sourceA_task_arb_io_in_6_bits_opcode),
    .io_in_6_bits_param(sourceA_task_arb_io_in_6_bits_param),
    .io_in_6_bits_source(sourceA_task_arb_io_in_6_bits_source),
    .io_in_6_bits_bufIdx(sourceA_task_arb_io_in_6_bits_bufIdx),
    .io_in_6_bits_size(sourceA_task_arb_io_in_6_bits_size),
    .io_in_6_bits_putData(sourceA_task_arb_io_in_6_bits_putData),
    .io_in_7_ready(sourceA_task_arb_io_in_7_ready),
    .io_in_7_valid(sourceA_task_arb_io_in_7_valid),
    .io_in_7_bits_tag(sourceA_task_arb_io_in_7_bits_tag),
    .io_in_7_bits_set(sourceA_task_arb_io_in_7_bits_set),
    .io_in_7_bits_off(sourceA_task_arb_io_in_7_bits_off),
    .io_in_7_bits_opcode(sourceA_task_arb_io_in_7_bits_opcode),
    .io_in_7_bits_param(sourceA_task_arb_io_in_7_bits_param),
    .io_in_7_bits_source(sourceA_task_arb_io_in_7_bits_source),
    .io_in_7_bits_bufIdx(sourceA_task_arb_io_in_7_bits_bufIdx),
    .io_in_7_bits_size(sourceA_task_arb_io_in_7_bits_size),
    .io_in_7_bits_putData(sourceA_task_arb_io_in_7_bits_putData),
    .io_in_8_ready(sourceA_task_arb_io_in_8_ready),
    .io_in_8_valid(sourceA_task_arb_io_in_8_valid),
    .io_in_8_bits_tag(sourceA_task_arb_io_in_8_bits_tag),
    .io_in_8_bits_set(sourceA_task_arb_io_in_8_bits_set),
    .io_in_8_bits_off(sourceA_task_arb_io_in_8_bits_off),
    .io_in_8_bits_opcode(sourceA_task_arb_io_in_8_bits_opcode),
    .io_in_8_bits_param(sourceA_task_arb_io_in_8_bits_param),
    .io_in_8_bits_source(sourceA_task_arb_io_in_8_bits_source),
    .io_in_8_bits_bufIdx(sourceA_task_arb_io_in_8_bits_bufIdx),
    .io_in_8_bits_size(sourceA_task_arb_io_in_8_bits_size),
    .io_in_8_bits_putData(sourceA_task_arb_io_in_8_bits_putData),
    .io_in_9_ready(sourceA_task_arb_io_in_9_ready),
    .io_in_9_valid(sourceA_task_arb_io_in_9_valid),
    .io_in_9_bits_tag(sourceA_task_arb_io_in_9_bits_tag),
    .io_in_9_bits_set(sourceA_task_arb_io_in_9_bits_set),
    .io_in_9_bits_off(sourceA_task_arb_io_in_9_bits_off),
    .io_in_9_bits_opcode(sourceA_task_arb_io_in_9_bits_opcode),
    .io_in_9_bits_param(sourceA_task_arb_io_in_9_bits_param),
    .io_in_9_bits_source(sourceA_task_arb_io_in_9_bits_source),
    .io_in_9_bits_bufIdx(sourceA_task_arb_io_in_9_bits_bufIdx),
    .io_in_9_bits_size(sourceA_task_arb_io_in_9_bits_size),
    .io_in_9_bits_putData(sourceA_task_arb_io_in_9_bits_putData),
    .io_in_10_ready(sourceA_task_arb_io_in_10_ready),
    .io_in_10_valid(sourceA_task_arb_io_in_10_valid),
    .io_in_10_bits_tag(sourceA_task_arb_io_in_10_bits_tag),
    .io_in_10_bits_set(sourceA_task_arb_io_in_10_bits_set),
    .io_in_10_bits_off(sourceA_task_arb_io_in_10_bits_off),
    .io_in_10_bits_opcode(sourceA_task_arb_io_in_10_bits_opcode),
    .io_in_10_bits_param(sourceA_task_arb_io_in_10_bits_param),
    .io_in_10_bits_source(sourceA_task_arb_io_in_10_bits_source),
    .io_in_10_bits_bufIdx(sourceA_task_arb_io_in_10_bits_bufIdx),
    .io_in_10_bits_size(sourceA_task_arb_io_in_10_bits_size),
    .io_in_10_bits_putData(sourceA_task_arb_io_in_10_bits_putData),
    .io_in_11_ready(sourceA_task_arb_io_in_11_ready),
    .io_in_11_valid(sourceA_task_arb_io_in_11_valid),
    .io_in_11_bits_tag(sourceA_task_arb_io_in_11_bits_tag),
    .io_in_11_bits_set(sourceA_task_arb_io_in_11_bits_set),
    .io_in_11_bits_off(sourceA_task_arb_io_in_11_bits_off),
    .io_in_11_bits_opcode(sourceA_task_arb_io_in_11_bits_opcode),
    .io_in_11_bits_param(sourceA_task_arb_io_in_11_bits_param),
    .io_in_11_bits_source(sourceA_task_arb_io_in_11_bits_source),
    .io_in_11_bits_bufIdx(sourceA_task_arb_io_in_11_bits_bufIdx),
    .io_in_11_bits_size(sourceA_task_arb_io_in_11_bits_size),
    .io_in_11_bits_putData(sourceA_task_arb_io_in_11_bits_putData),
    .io_in_12_ready(sourceA_task_arb_io_in_12_ready),
    .io_in_12_valid(sourceA_task_arb_io_in_12_valid),
    .io_in_12_bits_tag(sourceA_task_arb_io_in_12_bits_tag),
    .io_in_12_bits_set(sourceA_task_arb_io_in_12_bits_set),
    .io_in_12_bits_off(sourceA_task_arb_io_in_12_bits_off),
    .io_in_12_bits_opcode(sourceA_task_arb_io_in_12_bits_opcode),
    .io_in_12_bits_param(sourceA_task_arb_io_in_12_bits_param),
    .io_in_12_bits_source(sourceA_task_arb_io_in_12_bits_source),
    .io_in_12_bits_bufIdx(sourceA_task_arb_io_in_12_bits_bufIdx),
    .io_in_12_bits_size(sourceA_task_arb_io_in_12_bits_size),
    .io_in_12_bits_putData(sourceA_task_arb_io_in_12_bits_putData),
    .io_in_13_ready(sourceA_task_arb_io_in_13_ready),
    .io_in_13_valid(sourceA_task_arb_io_in_13_valid),
    .io_in_13_bits_tag(sourceA_task_arb_io_in_13_bits_tag),
    .io_in_13_bits_set(sourceA_task_arb_io_in_13_bits_set),
    .io_in_13_bits_off(sourceA_task_arb_io_in_13_bits_off),
    .io_in_13_bits_opcode(sourceA_task_arb_io_in_13_bits_opcode),
    .io_in_13_bits_param(sourceA_task_arb_io_in_13_bits_param),
    .io_in_13_bits_source(sourceA_task_arb_io_in_13_bits_source),
    .io_in_13_bits_bufIdx(sourceA_task_arb_io_in_13_bits_bufIdx),
    .io_in_13_bits_size(sourceA_task_arb_io_in_13_bits_size),
    .io_in_13_bits_putData(sourceA_task_arb_io_in_13_bits_putData),
    .io_out_ready(sourceA_task_arb_io_out_ready),
    .io_out_valid(sourceA_task_arb_io_out_valid),
    .io_out_bits_tag(sourceA_task_arb_io_out_bits_tag),
    .io_out_bits_set(sourceA_task_arb_io_out_bits_set),
    .io_out_bits_off(sourceA_task_arb_io_out_bits_off),
    .io_out_bits_opcode(sourceA_task_arb_io_out_bits_opcode),
    .io_out_bits_param(sourceA_task_arb_io_out_bits_param),
    .io_out_bits_source(sourceA_task_arb_io_out_bits_source),
    .io_out_bits_bufIdx(sourceA_task_arb_io_out_bits_bufIdx),
    .io_out_bits_size(sourceA_task_arb_io_out_bits_size),
    .io_out_bits_putData(sourceA_task_arb_io_out_bits_putData)
  );
  LatchFastArbiter_1 sourceB_task_arb ( // @[Slice.scala 468:27]
    .clock(sourceB_task_arb_clock),
    .reset(sourceB_task_arb_reset),
    .io_in_0_ready(sourceB_task_arb_io_in_0_ready),
    .io_in_0_valid(sourceB_task_arb_io_in_0_valid),
    .io_in_0_bits_set(sourceB_task_arb_io_in_0_bits_set),
    .io_in_0_bits_tag(sourceB_task_arb_io_in_0_bits_tag),
    .io_in_0_bits_param(sourceB_task_arb_io_in_0_bits_param),
    .io_in_0_bits_clients(sourceB_task_arb_io_in_0_bits_clients),
    .io_in_0_bits_needData(sourceB_task_arb_io_in_0_bits_needData),
    .io_in_1_ready(sourceB_task_arb_io_in_1_ready),
    .io_in_1_valid(sourceB_task_arb_io_in_1_valid),
    .io_in_1_bits_set(sourceB_task_arb_io_in_1_bits_set),
    .io_in_1_bits_tag(sourceB_task_arb_io_in_1_bits_tag),
    .io_in_1_bits_param(sourceB_task_arb_io_in_1_bits_param),
    .io_in_1_bits_clients(sourceB_task_arb_io_in_1_bits_clients),
    .io_in_1_bits_needData(sourceB_task_arb_io_in_1_bits_needData),
    .io_in_2_ready(sourceB_task_arb_io_in_2_ready),
    .io_in_2_valid(sourceB_task_arb_io_in_2_valid),
    .io_in_2_bits_set(sourceB_task_arb_io_in_2_bits_set),
    .io_in_2_bits_tag(sourceB_task_arb_io_in_2_bits_tag),
    .io_in_2_bits_param(sourceB_task_arb_io_in_2_bits_param),
    .io_in_2_bits_clients(sourceB_task_arb_io_in_2_bits_clients),
    .io_in_2_bits_needData(sourceB_task_arb_io_in_2_bits_needData),
    .io_in_3_ready(sourceB_task_arb_io_in_3_ready),
    .io_in_3_valid(sourceB_task_arb_io_in_3_valid),
    .io_in_3_bits_set(sourceB_task_arb_io_in_3_bits_set),
    .io_in_3_bits_tag(sourceB_task_arb_io_in_3_bits_tag),
    .io_in_3_bits_param(sourceB_task_arb_io_in_3_bits_param),
    .io_in_3_bits_clients(sourceB_task_arb_io_in_3_bits_clients),
    .io_in_3_bits_needData(sourceB_task_arb_io_in_3_bits_needData),
    .io_in_4_ready(sourceB_task_arb_io_in_4_ready),
    .io_in_4_valid(sourceB_task_arb_io_in_4_valid),
    .io_in_4_bits_set(sourceB_task_arb_io_in_4_bits_set),
    .io_in_4_bits_tag(sourceB_task_arb_io_in_4_bits_tag),
    .io_in_4_bits_param(sourceB_task_arb_io_in_4_bits_param),
    .io_in_4_bits_clients(sourceB_task_arb_io_in_4_bits_clients),
    .io_in_4_bits_needData(sourceB_task_arb_io_in_4_bits_needData),
    .io_in_5_ready(sourceB_task_arb_io_in_5_ready),
    .io_in_5_valid(sourceB_task_arb_io_in_5_valid),
    .io_in_5_bits_set(sourceB_task_arb_io_in_5_bits_set),
    .io_in_5_bits_tag(sourceB_task_arb_io_in_5_bits_tag),
    .io_in_5_bits_param(sourceB_task_arb_io_in_5_bits_param),
    .io_in_5_bits_clients(sourceB_task_arb_io_in_5_bits_clients),
    .io_in_5_bits_needData(sourceB_task_arb_io_in_5_bits_needData),
    .io_in_6_ready(sourceB_task_arb_io_in_6_ready),
    .io_in_6_valid(sourceB_task_arb_io_in_6_valid),
    .io_in_6_bits_set(sourceB_task_arb_io_in_6_bits_set),
    .io_in_6_bits_tag(sourceB_task_arb_io_in_6_bits_tag),
    .io_in_6_bits_param(sourceB_task_arb_io_in_6_bits_param),
    .io_in_6_bits_clients(sourceB_task_arb_io_in_6_bits_clients),
    .io_in_6_bits_needData(sourceB_task_arb_io_in_6_bits_needData),
    .io_in_7_ready(sourceB_task_arb_io_in_7_ready),
    .io_in_7_valid(sourceB_task_arb_io_in_7_valid),
    .io_in_7_bits_set(sourceB_task_arb_io_in_7_bits_set),
    .io_in_7_bits_tag(sourceB_task_arb_io_in_7_bits_tag),
    .io_in_7_bits_param(sourceB_task_arb_io_in_7_bits_param),
    .io_in_7_bits_clients(sourceB_task_arb_io_in_7_bits_clients),
    .io_in_7_bits_needData(sourceB_task_arb_io_in_7_bits_needData),
    .io_in_8_ready(sourceB_task_arb_io_in_8_ready),
    .io_in_8_valid(sourceB_task_arb_io_in_8_valid),
    .io_in_8_bits_set(sourceB_task_arb_io_in_8_bits_set),
    .io_in_8_bits_tag(sourceB_task_arb_io_in_8_bits_tag),
    .io_in_8_bits_param(sourceB_task_arb_io_in_8_bits_param),
    .io_in_8_bits_clients(sourceB_task_arb_io_in_8_bits_clients),
    .io_in_8_bits_needData(sourceB_task_arb_io_in_8_bits_needData),
    .io_in_9_ready(sourceB_task_arb_io_in_9_ready),
    .io_in_9_valid(sourceB_task_arb_io_in_9_valid),
    .io_in_9_bits_set(sourceB_task_arb_io_in_9_bits_set),
    .io_in_9_bits_tag(sourceB_task_arb_io_in_9_bits_tag),
    .io_in_9_bits_param(sourceB_task_arb_io_in_9_bits_param),
    .io_in_9_bits_clients(sourceB_task_arb_io_in_9_bits_clients),
    .io_in_9_bits_needData(sourceB_task_arb_io_in_9_bits_needData),
    .io_in_10_ready(sourceB_task_arb_io_in_10_ready),
    .io_in_10_valid(sourceB_task_arb_io_in_10_valid),
    .io_in_10_bits_set(sourceB_task_arb_io_in_10_bits_set),
    .io_in_10_bits_tag(sourceB_task_arb_io_in_10_bits_tag),
    .io_in_10_bits_param(sourceB_task_arb_io_in_10_bits_param),
    .io_in_10_bits_clients(sourceB_task_arb_io_in_10_bits_clients),
    .io_in_10_bits_needData(sourceB_task_arb_io_in_10_bits_needData),
    .io_in_11_ready(sourceB_task_arb_io_in_11_ready),
    .io_in_11_valid(sourceB_task_arb_io_in_11_valid),
    .io_in_11_bits_set(sourceB_task_arb_io_in_11_bits_set),
    .io_in_11_bits_tag(sourceB_task_arb_io_in_11_bits_tag),
    .io_in_11_bits_param(sourceB_task_arb_io_in_11_bits_param),
    .io_in_11_bits_clients(sourceB_task_arb_io_in_11_bits_clients),
    .io_in_11_bits_needData(sourceB_task_arb_io_in_11_bits_needData),
    .io_in_12_ready(sourceB_task_arb_io_in_12_ready),
    .io_in_12_valid(sourceB_task_arb_io_in_12_valid),
    .io_in_12_bits_set(sourceB_task_arb_io_in_12_bits_set),
    .io_in_12_bits_tag(sourceB_task_arb_io_in_12_bits_tag),
    .io_in_12_bits_param(sourceB_task_arb_io_in_12_bits_param),
    .io_in_12_bits_clients(sourceB_task_arb_io_in_12_bits_clients),
    .io_in_12_bits_needData(sourceB_task_arb_io_in_12_bits_needData),
    .io_in_13_ready(sourceB_task_arb_io_in_13_ready),
    .io_in_13_valid(sourceB_task_arb_io_in_13_valid),
    .io_in_13_bits_set(sourceB_task_arb_io_in_13_bits_set),
    .io_in_13_bits_tag(sourceB_task_arb_io_in_13_bits_tag),
    .io_in_13_bits_param(sourceB_task_arb_io_in_13_bits_param),
    .io_in_13_bits_clients(sourceB_task_arb_io_in_13_bits_clients),
    .io_in_13_bits_needData(sourceB_task_arb_io_in_13_bits_needData),
    .io_out_ready(sourceB_task_arb_io_out_ready),
    .io_out_valid(sourceB_task_arb_io_out_valid),
    .io_out_bits_set(sourceB_task_arb_io_out_bits_set),
    .io_out_bits_tag(sourceB_task_arb_io_out_bits_tag),
    .io_out_bits_param(sourceB_task_arb_io_out_bits_param),
    .io_out_bits_clients(sourceB_task_arb_io_out_bits_clients),
    .io_out_bits_needData(sourceB_task_arb_io_out_bits_needData)
  );
  LatchFastArbiter_2 sourceC_task_arb ( // @[Slice.scala 468:27]
    .clock(sourceC_task_arb_clock),
    .reset(sourceC_task_arb_reset),
    .io_in_0_ready(sourceC_task_arb_io_in_0_ready),
    .io_in_0_valid(sourceC_task_arb_io_in_0_valid),
    .io_in_0_bits_opcode(sourceC_task_arb_io_in_0_bits_opcode),
    .io_in_0_bits_tag(sourceC_task_arb_io_in_0_bits_tag),
    .io_in_0_bits_set(sourceC_task_arb_io_in_0_bits_set),
    .io_in_0_bits_source(sourceC_task_arb_io_in_0_bits_source),
    .io_in_0_bits_way(sourceC_task_arb_io_in_0_bits_way),
    .io_in_1_ready(sourceC_task_arb_io_in_1_ready),
    .io_in_1_valid(sourceC_task_arb_io_in_1_valid),
    .io_in_1_bits_opcode(sourceC_task_arb_io_in_1_bits_opcode),
    .io_in_1_bits_tag(sourceC_task_arb_io_in_1_bits_tag),
    .io_in_1_bits_set(sourceC_task_arb_io_in_1_bits_set),
    .io_in_1_bits_source(sourceC_task_arb_io_in_1_bits_source),
    .io_in_1_bits_way(sourceC_task_arb_io_in_1_bits_way),
    .io_in_2_ready(sourceC_task_arb_io_in_2_ready),
    .io_in_2_valid(sourceC_task_arb_io_in_2_valid),
    .io_in_2_bits_opcode(sourceC_task_arb_io_in_2_bits_opcode),
    .io_in_2_bits_tag(sourceC_task_arb_io_in_2_bits_tag),
    .io_in_2_bits_set(sourceC_task_arb_io_in_2_bits_set),
    .io_in_2_bits_source(sourceC_task_arb_io_in_2_bits_source),
    .io_in_2_bits_way(sourceC_task_arb_io_in_2_bits_way),
    .io_in_3_ready(sourceC_task_arb_io_in_3_ready),
    .io_in_3_valid(sourceC_task_arb_io_in_3_valid),
    .io_in_3_bits_opcode(sourceC_task_arb_io_in_3_bits_opcode),
    .io_in_3_bits_tag(sourceC_task_arb_io_in_3_bits_tag),
    .io_in_3_bits_set(sourceC_task_arb_io_in_3_bits_set),
    .io_in_3_bits_source(sourceC_task_arb_io_in_3_bits_source),
    .io_in_3_bits_way(sourceC_task_arb_io_in_3_bits_way),
    .io_in_4_ready(sourceC_task_arb_io_in_4_ready),
    .io_in_4_valid(sourceC_task_arb_io_in_4_valid),
    .io_in_4_bits_opcode(sourceC_task_arb_io_in_4_bits_opcode),
    .io_in_4_bits_tag(sourceC_task_arb_io_in_4_bits_tag),
    .io_in_4_bits_set(sourceC_task_arb_io_in_4_bits_set),
    .io_in_4_bits_source(sourceC_task_arb_io_in_4_bits_source),
    .io_in_4_bits_way(sourceC_task_arb_io_in_4_bits_way),
    .io_in_5_ready(sourceC_task_arb_io_in_5_ready),
    .io_in_5_valid(sourceC_task_arb_io_in_5_valid),
    .io_in_5_bits_opcode(sourceC_task_arb_io_in_5_bits_opcode),
    .io_in_5_bits_tag(sourceC_task_arb_io_in_5_bits_tag),
    .io_in_5_bits_set(sourceC_task_arb_io_in_5_bits_set),
    .io_in_5_bits_source(sourceC_task_arb_io_in_5_bits_source),
    .io_in_5_bits_way(sourceC_task_arb_io_in_5_bits_way),
    .io_in_6_ready(sourceC_task_arb_io_in_6_ready),
    .io_in_6_valid(sourceC_task_arb_io_in_6_valid),
    .io_in_6_bits_opcode(sourceC_task_arb_io_in_6_bits_opcode),
    .io_in_6_bits_tag(sourceC_task_arb_io_in_6_bits_tag),
    .io_in_6_bits_set(sourceC_task_arb_io_in_6_bits_set),
    .io_in_6_bits_source(sourceC_task_arb_io_in_6_bits_source),
    .io_in_6_bits_way(sourceC_task_arb_io_in_6_bits_way),
    .io_in_7_ready(sourceC_task_arb_io_in_7_ready),
    .io_in_7_valid(sourceC_task_arb_io_in_7_valid),
    .io_in_7_bits_opcode(sourceC_task_arb_io_in_7_bits_opcode),
    .io_in_7_bits_tag(sourceC_task_arb_io_in_7_bits_tag),
    .io_in_7_bits_set(sourceC_task_arb_io_in_7_bits_set),
    .io_in_7_bits_source(sourceC_task_arb_io_in_7_bits_source),
    .io_in_7_bits_way(sourceC_task_arb_io_in_7_bits_way),
    .io_in_8_ready(sourceC_task_arb_io_in_8_ready),
    .io_in_8_valid(sourceC_task_arb_io_in_8_valid),
    .io_in_8_bits_opcode(sourceC_task_arb_io_in_8_bits_opcode),
    .io_in_8_bits_tag(sourceC_task_arb_io_in_8_bits_tag),
    .io_in_8_bits_set(sourceC_task_arb_io_in_8_bits_set),
    .io_in_8_bits_source(sourceC_task_arb_io_in_8_bits_source),
    .io_in_8_bits_way(sourceC_task_arb_io_in_8_bits_way),
    .io_in_9_ready(sourceC_task_arb_io_in_9_ready),
    .io_in_9_valid(sourceC_task_arb_io_in_9_valid),
    .io_in_9_bits_opcode(sourceC_task_arb_io_in_9_bits_opcode),
    .io_in_9_bits_tag(sourceC_task_arb_io_in_9_bits_tag),
    .io_in_9_bits_set(sourceC_task_arb_io_in_9_bits_set),
    .io_in_9_bits_source(sourceC_task_arb_io_in_9_bits_source),
    .io_in_9_bits_way(sourceC_task_arb_io_in_9_bits_way),
    .io_in_10_ready(sourceC_task_arb_io_in_10_ready),
    .io_in_10_valid(sourceC_task_arb_io_in_10_valid),
    .io_in_10_bits_opcode(sourceC_task_arb_io_in_10_bits_opcode),
    .io_in_10_bits_tag(sourceC_task_arb_io_in_10_bits_tag),
    .io_in_10_bits_set(sourceC_task_arb_io_in_10_bits_set),
    .io_in_10_bits_source(sourceC_task_arb_io_in_10_bits_source),
    .io_in_10_bits_way(sourceC_task_arb_io_in_10_bits_way),
    .io_in_11_ready(sourceC_task_arb_io_in_11_ready),
    .io_in_11_valid(sourceC_task_arb_io_in_11_valid),
    .io_in_11_bits_opcode(sourceC_task_arb_io_in_11_bits_opcode),
    .io_in_11_bits_tag(sourceC_task_arb_io_in_11_bits_tag),
    .io_in_11_bits_set(sourceC_task_arb_io_in_11_bits_set),
    .io_in_11_bits_source(sourceC_task_arb_io_in_11_bits_source),
    .io_in_11_bits_way(sourceC_task_arb_io_in_11_bits_way),
    .io_in_12_ready(sourceC_task_arb_io_in_12_ready),
    .io_in_12_valid(sourceC_task_arb_io_in_12_valid),
    .io_in_12_bits_opcode(sourceC_task_arb_io_in_12_bits_opcode),
    .io_in_12_bits_tag(sourceC_task_arb_io_in_12_bits_tag),
    .io_in_12_bits_set(sourceC_task_arb_io_in_12_bits_set),
    .io_in_12_bits_source(sourceC_task_arb_io_in_12_bits_source),
    .io_in_12_bits_way(sourceC_task_arb_io_in_12_bits_way),
    .io_in_13_ready(sourceC_task_arb_io_in_13_ready),
    .io_in_13_valid(sourceC_task_arb_io_in_13_valid),
    .io_in_13_bits_opcode(sourceC_task_arb_io_in_13_bits_opcode),
    .io_in_13_bits_tag(sourceC_task_arb_io_in_13_bits_tag),
    .io_in_13_bits_set(sourceC_task_arb_io_in_13_bits_set),
    .io_in_13_bits_source(sourceC_task_arb_io_in_13_bits_source),
    .io_in_13_bits_way(sourceC_task_arb_io_in_13_bits_way),
    .io_out_ready(sourceC_task_arb_io_out_ready),
    .io_out_valid(sourceC_task_arb_io_out_valid),
    .io_out_bits_opcode(sourceC_task_arb_io_out_bits_opcode),
    .io_out_bits_tag(sourceC_task_arb_io_out_bits_tag),
    .io_out_bits_set(sourceC_task_arb_io_out_bits_set),
    .io_out_bits_source(sourceC_task_arb_io_out_bits_source),
    .io_out_bits_way(sourceC_task_arb_io_out_bits_way)
  );
  LatchFastArbiter_3 sourceD_task_arb ( // @[Slice.scala 468:27]
    .clock(sourceD_task_arb_clock),
    .reset(sourceD_task_arb_reset),
    .io_in_0_ready(sourceD_task_arb_io_in_0_ready),
    .io_in_0_valid(sourceD_task_arb_io_in_0_valid),
    .io_in_0_bits_sourceId(sourceD_task_arb_io_in_0_bits_sourceId),
    .io_in_0_bits_set(sourceD_task_arb_io_in_0_bits_set),
    .io_in_0_bits_channel(sourceD_task_arb_io_in_0_bits_channel),
    .io_in_0_bits_opcode(sourceD_task_arb_io_in_0_bits_opcode),
    .io_in_0_bits_param(sourceD_task_arb_io_in_0_bits_param),
    .io_in_0_bits_size(sourceD_task_arb_io_in_0_bits_size),
    .io_in_0_bits_way(sourceD_task_arb_io_in_0_bits_way),
    .io_in_0_bits_off(sourceD_task_arb_io_in_0_bits_off),
    .io_in_0_bits_useBypass(sourceD_task_arb_io_in_0_bits_useBypass),
    .io_in_0_bits_bufIdx(sourceD_task_arb_io_in_0_bits_bufIdx),
    .io_in_0_bits_denied(sourceD_task_arb_io_in_0_bits_denied),
    .io_in_0_bits_sinkId(sourceD_task_arb_io_in_0_bits_sinkId),
    .io_in_0_bits_bypassPut(sourceD_task_arb_io_in_0_bits_bypassPut),
    .io_in_0_bits_dirty(sourceD_task_arb_io_in_0_bits_dirty),
    .io_in_1_ready(sourceD_task_arb_io_in_1_ready),
    .io_in_1_valid(sourceD_task_arb_io_in_1_valid),
    .io_in_1_bits_sourceId(sourceD_task_arb_io_in_1_bits_sourceId),
    .io_in_1_bits_set(sourceD_task_arb_io_in_1_bits_set),
    .io_in_1_bits_channel(sourceD_task_arb_io_in_1_bits_channel),
    .io_in_1_bits_opcode(sourceD_task_arb_io_in_1_bits_opcode),
    .io_in_1_bits_param(sourceD_task_arb_io_in_1_bits_param),
    .io_in_1_bits_size(sourceD_task_arb_io_in_1_bits_size),
    .io_in_1_bits_way(sourceD_task_arb_io_in_1_bits_way),
    .io_in_1_bits_off(sourceD_task_arb_io_in_1_bits_off),
    .io_in_1_bits_useBypass(sourceD_task_arb_io_in_1_bits_useBypass),
    .io_in_1_bits_bufIdx(sourceD_task_arb_io_in_1_bits_bufIdx),
    .io_in_1_bits_denied(sourceD_task_arb_io_in_1_bits_denied),
    .io_in_1_bits_sinkId(sourceD_task_arb_io_in_1_bits_sinkId),
    .io_in_1_bits_bypassPut(sourceD_task_arb_io_in_1_bits_bypassPut),
    .io_in_1_bits_dirty(sourceD_task_arb_io_in_1_bits_dirty),
    .io_in_2_ready(sourceD_task_arb_io_in_2_ready),
    .io_in_2_valid(sourceD_task_arb_io_in_2_valid),
    .io_in_2_bits_sourceId(sourceD_task_arb_io_in_2_bits_sourceId),
    .io_in_2_bits_set(sourceD_task_arb_io_in_2_bits_set),
    .io_in_2_bits_channel(sourceD_task_arb_io_in_2_bits_channel),
    .io_in_2_bits_opcode(sourceD_task_arb_io_in_2_bits_opcode),
    .io_in_2_bits_param(sourceD_task_arb_io_in_2_bits_param),
    .io_in_2_bits_size(sourceD_task_arb_io_in_2_bits_size),
    .io_in_2_bits_way(sourceD_task_arb_io_in_2_bits_way),
    .io_in_2_bits_off(sourceD_task_arb_io_in_2_bits_off),
    .io_in_2_bits_useBypass(sourceD_task_arb_io_in_2_bits_useBypass),
    .io_in_2_bits_bufIdx(sourceD_task_arb_io_in_2_bits_bufIdx),
    .io_in_2_bits_denied(sourceD_task_arb_io_in_2_bits_denied),
    .io_in_2_bits_sinkId(sourceD_task_arb_io_in_2_bits_sinkId),
    .io_in_2_bits_bypassPut(sourceD_task_arb_io_in_2_bits_bypassPut),
    .io_in_2_bits_dirty(sourceD_task_arb_io_in_2_bits_dirty),
    .io_in_3_ready(sourceD_task_arb_io_in_3_ready),
    .io_in_3_valid(sourceD_task_arb_io_in_3_valid),
    .io_in_3_bits_sourceId(sourceD_task_arb_io_in_3_bits_sourceId),
    .io_in_3_bits_set(sourceD_task_arb_io_in_3_bits_set),
    .io_in_3_bits_channel(sourceD_task_arb_io_in_3_bits_channel),
    .io_in_3_bits_opcode(sourceD_task_arb_io_in_3_bits_opcode),
    .io_in_3_bits_param(sourceD_task_arb_io_in_3_bits_param),
    .io_in_3_bits_size(sourceD_task_arb_io_in_3_bits_size),
    .io_in_3_bits_way(sourceD_task_arb_io_in_3_bits_way),
    .io_in_3_bits_off(sourceD_task_arb_io_in_3_bits_off),
    .io_in_3_bits_useBypass(sourceD_task_arb_io_in_3_bits_useBypass),
    .io_in_3_bits_bufIdx(sourceD_task_arb_io_in_3_bits_bufIdx),
    .io_in_3_bits_denied(sourceD_task_arb_io_in_3_bits_denied),
    .io_in_3_bits_sinkId(sourceD_task_arb_io_in_3_bits_sinkId),
    .io_in_3_bits_bypassPut(sourceD_task_arb_io_in_3_bits_bypassPut),
    .io_in_3_bits_dirty(sourceD_task_arb_io_in_3_bits_dirty),
    .io_in_4_ready(sourceD_task_arb_io_in_4_ready),
    .io_in_4_valid(sourceD_task_arb_io_in_4_valid),
    .io_in_4_bits_sourceId(sourceD_task_arb_io_in_4_bits_sourceId),
    .io_in_4_bits_set(sourceD_task_arb_io_in_4_bits_set),
    .io_in_4_bits_channel(sourceD_task_arb_io_in_4_bits_channel),
    .io_in_4_bits_opcode(sourceD_task_arb_io_in_4_bits_opcode),
    .io_in_4_bits_param(sourceD_task_arb_io_in_4_bits_param),
    .io_in_4_bits_size(sourceD_task_arb_io_in_4_bits_size),
    .io_in_4_bits_way(sourceD_task_arb_io_in_4_bits_way),
    .io_in_4_bits_off(sourceD_task_arb_io_in_4_bits_off),
    .io_in_4_bits_useBypass(sourceD_task_arb_io_in_4_bits_useBypass),
    .io_in_4_bits_bufIdx(sourceD_task_arb_io_in_4_bits_bufIdx),
    .io_in_4_bits_denied(sourceD_task_arb_io_in_4_bits_denied),
    .io_in_4_bits_sinkId(sourceD_task_arb_io_in_4_bits_sinkId),
    .io_in_4_bits_bypassPut(sourceD_task_arb_io_in_4_bits_bypassPut),
    .io_in_4_bits_dirty(sourceD_task_arb_io_in_4_bits_dirty),
    .io_in_5_ready(sourceD_task_arb_io_in_5_ready),
    .io_in_5_valid(sourceD_task_arb_io_in_5_valid),
    .io_in_5_bits_sourceId(sourceD_task_arb_io_in_5_bits_sourceId),
    .io_in_5_bits_set(sourceD_task_arb_io_in_5_bits_set),
    .io_in_5_bits_channel(sourceD_task_arb_io_in_5_bits_channel),
    .io_in_5_bits_opcode(sourceD_task_arb_io_in_5_bits_opcode),
    .io_in_5_bits_param(sourceD_task_arb_io_in_5_bits_param),
    .io_in_5_bits_size(sourceD_task_arb_io_in_5_bits_size),
    .io_in_5_bits_way(sourceD_task_arb_io_in_5_bits_way),
    .io_in_5_bits_off(sourceD_task_arb_io_in_5_bits_off),
    .io_in_5_bits_useBypass(sourceD_task_arb_io_in_5_bits_useBypass),
    .io_in_5_bits_bufIdx(sourceD_task_arb_io_in_5_bits_bufIdx),
    .io_in_5_bits_denied(sourceD_task_arb_io_in_5_bits_denied),
    .io_in_5_bits_sinkId(sourceD_task_arb_io_in_5_bits_sinkId),
    .io_in_5_bits_bypassPut(sourceD_task_arb_io_in_5_bits_bypassPut),
    .io_in_5_bits_dirty(sourceD_task_arb_io_in_5_bits_dirty),
    .io_in_6_ready(sourceD_task_arb_io_in_6_ready),
    .io_in_6_valid(sourceD_task_arb_io_in_6_valid),
    .io_in_6_bits_sourceId(sourceD_task_arb_io_in_6_bits_sourceId),
    .io_in_6_bits_set(sourceD_task_arb_io_in_6_bits_set),
    .io_in_6_bits_channel(sourceD_task_arb_io_in_6_bits_channel),
    .io_in_6_bits_opcode(sourceD_task_arb_io_in_6_bits_opcode),
    .io_in_6_bits_param(sourceD_task_arb_io_in_6_bits_param),
    .io_in_6_bits_size(sourceD_task_arb_io_in_6_bits_size),
    .io_in_6_bits_way(sourceD_task_arb_io_in_6_bits_way),
    .io_in_6_bits_off(sourceD_task_arb_io_in_6_bits_off),
    .io_in_6_bits_useBypass(sourceD_task_arb_io_in_6_bits_useBypass),
    .io_in_6_bits_bufIdx(sourceD_task_arb_io_in_6_bits_bufIdx),
    .io_in_6_bits_denied(sourceD_task_arb_io_in_6_bits_denied),
    .io_in_6_bits_sinkId(sourceD_task_arb_io_in_6_bits_sinkId),
    .io_in_6_bits_bypassPut(sourceD_task_arb_io_in_6_bits_bypassPut),
    .io_in_6_bits_dirty(sourceD_task_arb_io_in_6_bits_dirty),
    .io_in_7_ready(sourceD_task_arb_io_in_7_ready),
    .io_in_7_valid(sourceD_task_arb_io_in_7_valid),
    .io_in_7_bits_sourceId(sourceD_task_arb_io_in_7_bits_sourceId),
    .io_in_7_bits_set(sourceD_task_arb_io_in_7_bits_set),
    .io_in_7_bits_channel(sourceD_task_arb_io_in_7_bits_channel),
    .io_in_7_bits_opcode(sourceD_task_arb_io_in_7_bits_opcode),
    .io_in_7_bits_param(sourceD_task_arb_io_in_7_bits_param),
    .io_in_7_bits_size(sourceD_task_arb_io_in_7_bits_size),
    .io_in_7_bits_way(sourceD_task_arb_io_in_7_bits_way),
    .io_in_7_bits_off(sourceD_task_arb_io_in_7_bits_off),
    .io_in_7_bits_useBypass(sourceD_task_arb_io_in_7_bits_useBypass),
    .io_in_7_bits_bufIdx(sourceD_task_arb_io_in_7_bits_bufIdx),
    .io_in_7_bits_denied(sourceD_task_arb_io_in_7_bits_denied),
    .io_in_7_bits_sinkId(sourceD_task_arb_io_in_7_bits_sinkId),
    .io_in_7_bits_bypassPut(sourceD_task_arb_io_in_7_bits_bypassPut),
    .io_in_7_bits_dirty(sourceD_task_arb_io_in_7_bits_dirty),
    .io_in_8_ready(sourceD_task_arb_io_in_8_ready),
    .io_in_8_valid(sourceD_task_arb_io_in_8_valid),
    .io_in_8_bits_sourceId(sourceD_task_arb_io_in_8_bits_sourceId),
    .io_in_8_bits_set(sourceD_task_arb_io_in_8_bits_set),
    .io_in_8_bits_channel(sourceD_task_arb_io_in_8_bits_channel),
    .io_in_8_bits_opcode(sourceD_task_arb_io_in_8_bits_opcode),
    .io_in_8_bits_param(sourceD_task_arb_io_in_8_bits_param),
    .io_in_8_bits_size(sourceD_task_arb_io_in_8_bits_size),
    .io_in_8_bits_way(sourceD_task_arb_io_in_8_bits_way),
    .io_in_8_bits_off(sourceD_task_arb_io_in_8_bits_off),
    .io_in_8_bits_useBypass(sourceD_task_arb_io_in_8_bits_useBypass),
    .io_in_8_bits_bufIdx(sourceD_task_arb_io_in_8_bits_bufIdx),
    .io_in_8_bits_denied(sourceD_task_arb_io_in_8_bits_denied),
    .io_in_8_bits_sinkId(sourceD_task_arb_io_in_8_bits_sinkId),
    .io_in_8_bits_bypassPut(sourceD_task_arb_io_in_8_bits_bypassPut),
    .io_in_8_bits_dirty(sourceD_task_arb_io_in_8_bits_dirty),
    .io_in_9_ready(sourceD_task_arb_io_in_9_ready),
    .io_in_9_valid(sourceD_task_arb_io_in_9_valid),
    .io_in_9_bits_sourceId(sourceD_task_arb_io_in_9_bits_sourceId),
    .io_in_9_bits_set(sourceD_task_arb_io_in_9_bits_set),
    .io_in_9_bits_channel(sourceD_task_arb_io_in_9_bits_channel),
    .io_in_9_bits_opcode(sourceD_task_arb_io_in_9_bits_opcode),
    .io_in_9_bits_param(sourceD_task_arb_io_in_9_bits_param),
    .io_in_9_bits_size(sourceD_task_arb_io_in_9_bits_size),
    .io_in_9_bits_way(sourceD_task_arb_io_in_9_bits_way),
    .io_in_9_bits_off(sourceD_task_arb_io_in_9_bits_off),
    .io_in_9_bits_useBypass(sourceD_task_arb_io_in_9_bits_useBypass),
    .io_in_9_bits_bufIdx(sourceD_task_arb_io_in_9_bits_bufIdx),
    .io_in_9_bits_denied(sourceD_task_arb_io_in_9_bits_denied),
    .io_in_9_bits_sinkId(sourceD_task_arb_io_in_9_bits_sinkId),
    .io_in_9_bits_bypassPut(sourceD_task_arb_io_in_9_bits_bypassPut),
    .io_in_9_bits_dirty(sourceD_task_arb_io_in_9_bits_dirty),
    .io_in_10_ready(sourceD_task_arb_io_in_10_ready),
    .io_in_10_valid(sourceD_task_arb_io_in_10_valid),
    .io_in_10_bits_sourceId(sourceD_task_arb_io_in_10_bits_sourceId),
    .io_in_10_bits_set(sourceD_task_arb_io_in_10_bits_set),
    .io_in_10_bits_channel(sourceD_task_arb_io_in_10_bits_channel),
    .io_in_10_bits_opcode(sourceD_task_arb_io_in_10_bits_opcode),
    .io_in_10_bits_param(sourceD_task_arb_io_in_10_bits_param),
    .io_in_10_bits_size(sourceD_task_arb_io_in_10_bits_size),
    .io_in_10_bits_way(sourceD_task_arb_io_in_10_bits_way),
    .io_in_10_bits_off(sourceD_task_arb_io_in_10_bits_off),
    .io_in_10_bits_useBypass(sourceD_task_arb_io_in_10_bits_useBypass),
    .io_in_10_bits_bufIdx(sourceD_task_arb_io_in_10_bits_bufIdx),
    .io_in_10_bits_denied(sourceD_task_arb_io_in_10_bits_denied),
    .io_in_10_bits_sinkId(sourceD_task_arb_io_in_10_bits_sinkId),
    .io_in_10_bits_bypassPut(sourceD_task_arb_io_in_10_bits_bypassPut),
    .io_in_10_bits_dirty(sourceD_task_arb_io_in_10_bits_dirty),
    .io_in_11_ready(sourceD_task_arb_io_in_11_ready),
    .io_in_11_valid(sourceD_task_arb_io_in_11_valid),
    .io_in_11_bits_sourceId(sourceD_task_arb_io_in_11_bits_sourceId),
    .io_in_11_bits_set(sourceD_task_arb_io_in_11_bits_set),
    .io_in_11_bits_channel(sourceD_task_arb_io_in_11_bits_channel),
    .io_in_11_bits_opcode(sourceD_task_arb_io_in_11_bits_opcode),
    .io_in_11_bits_param(sourceD_task_arb_io_in_11_bits_param),
    .io_in_11_bits_size(sourceD_task_arb_io_in_11_bits_size),
    .io_in_11_bits_way(sourceD_task_arb_io_in_11_bits_way),
    .io_in_11_bits_off(sourceD_task_arb_io_in_11_bits_off),
    .io_in_11_bits_useBypass(sourceD_task_arb_io_in_11_bits_useBypass),
    .io_in_11_bits_bufIdx(sourceD_task_arb_io_in_11_bits_bufIdx),
    .io_in_11_bits_denied(sourceD_task_arb_io_in_11_bits_denied),
    .io_in_11_bits_sinkId(sourceD_task_arb_io_in_11_bits_sinkId),
    .io_in_11_bits_bypassPut(sourceD_task_arb_io_in_11_bits_bypassPut),
    .io_in_11_bits_dirty(sourceD_task_arb_io_in_11_bits_dirty),
    .io_in_12_ready(sourceD_task_arb_io_in_12_ready),
    .io_in_12_valid(sourceD_task_arb_io_in_12_valid),
    .io_in_12_bits_sourceId(sourceD_task_arb_io_in_12_bits_sourceId),
    .io_in_12_bits_set(sourceD_task_arb_io_in_12_bits_set),
    .io_in_12_bits_channel(sourceD_task_arb_io_in_12_bits_channel),
    .io_in_12_bits_opcode(sourceD_task_arb_io_in_12_bits_opcode),
    .io_in_12_bits_param(sourceD_task_arb_io_in_12_bits_param),
    .io_in_12_bits_size(sourceD_task_arb_io_in_12_bits_size),
    .io_in_12_bits_way(sourceD_task_arb_io_in_12_bits_way),
    .io_in_12_bits_off(sourceD_task_arb_io_in_12_bits_off),
    .io_in_12_bits_useBypass(sourceD_task_arb_io_in_12_bits_useBypass),
    .io_in_12_bits_bufIdx(sourceD_task_arb_io_in_12_bits_bufIdx),
    .io_in_12_bits_denied(sourceD_task_arb_io_in_12_bits_denied),
    .io_in_12_bits_sinkId(sourceD_task_arb_io_in_12_bits_sinkId),
    .io_in_12_bits_bypassPut(sourceD_task_arb_io_in_12_bits_bypassPut),
    .io_in_12_bits_dirty(sourceD_task_arb_io_in_12_bits_dirty),
    .io_in_13_ready(sourceD_task_arb_io_in_13_ready),
    .io_in_13_valid(sourceD_task_arb_io_in_13_valid),
    .io_in_13_bits_sourceId(sourceD_task_arb_io_in_13_bits_sourceId),
    .io_in_13_bits_set(sourceD_task_arb_io_in_13_bits_set),
    .io_in_13_bits_channel(sourceD_task_arb_io_in_13_bits_channel),
    .io_in_13_bits_opcode(sourceD_task_arb_io_in_13_bits_opcode),
    .io_in_13_bits_param(sourceD_task_arb_io_in_13_bits_param),
    .io_in_13_bits_size(sourceD_task_arb_io_in_13_bits_size),
    .io_in_13_bits_way(sourceD_task_arb_io_in_13_bits_way),
    .io_in_13_bits_off(sourceD_task_arb_io_in_13_bits_off),
    .io_in_13_bits_useBypass(sourceD_task_arb_io_in_13_bits_useBypass),
    .io_in_13_bits_bufIdx(sourceD_task_arb_io_in_13_bits_bufIdx),
    .io_in_13_bits_denied(sourceD_task_arb_io_in_13_bits_denied),
    .io_in_13_bits_sinkId(sourceD_task_arb_io_in_13_bits_sinkId),
    .io_in_13_bits_bypassPut(sourceD_task_arb_io_in_13_bits_bypassPut),
    .io_in_13_bits_dirty(sourceD_task_arb_io_in_13_bits_dirty),
    .io_out_ready(sourceD_task_arb_io_out_ready),
    .io_out_valid(sourceD_task_arb_io_out_valid),
    .io_out_bits_sourceId(sourceD_task_arb_io_out_bits_sourceId),
    .io_out_bits_set(sourceD_task_arb_io_out_bits_set),
    .io_out_bits_channel(sourceD_task_arb_io_out_bits_channel),
    .io_out_bits_opcode(sourceD_task_arb_io_out_bits_opcode),
    .io_out_bits_param(sourceD_task_arb_io_out_bits_param),
    .io_out_bits_size(sourceD_task_arb_io_out_bits_size),
    .io_out_bits_way(sourceD_task_arb_io_out_bits_way),
    .io_out_bits_off(sourceD_task_arb_io_out_bits_off),
    .io_out_bits_useBypass(sourceD_task_arb_io_out_bits_useBypass),
    .io_out_bits_bufIdx(sourceD_task_arb_io_out_bits_bufIdx),
    .io_out_bits_denied(sourceD_task_arb_io_out_bits_denied),
    .io_out_bits_sinkId(sourceD_task_arb_io_out_bits_sinkId),
    .io_out_bits_bypassPut(sourceD_task_arb_io_out_bits_bypassPut),
    .io_out_bits_dirty(sourceD_task_arb_io_out_bits_dirty)
  );
  LatchFastArbiter_4 sourceE_task_arb ( // @[Slice.scala 468:27]
    .clock(sourceE_task_arb_clock),
    .reset(sourceE_task_arb_reset),
    .io_in_0_ready(sourceE_task_arb_io_in_0_ready),
    .io_in_0_valid(sourceE_task_arb_io_in_0_valid),
    .io_in_0_bits_sink(sourceE_task_arb_io_in_0_bits_sink),
    .io_in_1_ready(sourceE_task_arb_io_in_1_ready),
    .io_in_1_valid(sourceE_task_arb_io_in_1_valid),
    .io_in_1_bits_sink(sourceE_task_arb_io_in_1_bits_sink),
    .io_in_2_ready(sourceE_task_arb_io_in_2_ready),
    .io_in_2_valid(sourceE_task_arb_io_in_2_valid),
    .io_in_2_bits_sink(sourceE_task_arb_io_in_2_bits_sink),
    .io_in_3_ready(sourceE_task_arb_io_in_3_ready),
    .io_in_3_valid(sourceE_task_arb_io_in_3_valid),
    .io_in_3_bits_sink(sourceE_task_arb_io_in_3_bits_sink),
    .io_in_4_ready(sourceE_task_arb_io_in_4_ready),
    .io_in_4_valid(sourceE_task_arb_io_in_4_valid),
    .io_in_4_bits_sink(sourceE_task_arb_io_in_4_bits_sink),
    .io_in_5_ready(sourceE_task_arb_io_in_5_ready),
    .io_in_5_valid(sourceE_task_arb_io_in_5_valid),
    .io_in_5_bits_sink(sourceE_task_arb_io_in_5_bits_sink),
    .io_in_6_ready(sourceE_task_arb_io_in_6_ready),
    .io_in_6_valid(sourceE_task_arb_io_in_6_valid),
    .io_in_6_bits_sink(sourceE_task_arb_io_in_6_bits_sink),
    .io_in_7_ready(sourceE_task_arb_io_in_7_ready),
    .io_in_7_valid(sourceE_task_arb_io_in_7_valid),
    .io_in_7_bits_sink(sourceE_task_arb_io_in_7_bits_sink),
    .io_in_8_ready(sourceE_task_arb_io_in_8_ready),
    .io_in_8_valid(sourceE_task_arb_io_in_8_valid),
    .io_in_8_bits_sink(sourceE_task_arb_io_in_8_bits_sink),
    .io_in_9_ready(sourceE_task_arb_io_in_9_ready),
    .io_in_9_valid(sourceE_task_arb_io_in_9_valid),
    .io_in_9_bits_sink(sourceE_task_arb_io_in_9_bits_sink),
    .io_in_10_ready(sourceE_task_arb_io_in_10_ready),
    .io_in_10_valid(sourceE_task_arb_io_in_10_valid),
    .io_in_10_bits_sink(sourceE_task_arb_io_in_10_bits_sink),
    .io_in_11_ready(sourceE_task_arb_io_in_11_ready),
    .io_in_11_valid(sourceE_task_arb_io_in_11_valid),
    .io_in_11_bits_sink(sourceE_task_arb_io_in_11_bits_sink),
    .io_in_12_ready(sourceE_task_arb_io_in_12_ready),
    .io_in_12_valid(sourceE_task_arb_io_in_12_valid),
    .io_in_12_bits_sink(sourceE_task_arb_io_in_12_bits_sink),
    .io_in_13_ready(sourceE_task_arb_io_in_13_ready),
    .io_in_13_valid(sourceE_task_arb_io_in_13_valid),
    .io_in_13_bits_sink(sourceE_task_arb_io_in_13_bits_sink),
    .io_out_ready(sourceE_task_arb_io_out_ready),
    .io_out_valid(sourceE_task_arb_io_out_valid),
    .io_out_bits_sink(sourceE_task_arb_io_out_bits_sink)
  );
  LatchFastArbiter_6 sinkC_task_arb ( // @[Slice.scala 468:27]
    .clock(sinkC_task_arb_clock),
    .reset(sinkC_task_arb_reset),
    .io_in_0_ready(sinkC_task_arb_io_in_0_ready),
    .io_in_0_valid(sinkC_task_arb_io_in_0_valid),
    .io_in_0_bits_set(sinkC_task_arb_io_in_0_bits_set),
    .io_in_0_bits_tag(sinkC_task_arb_io_in_0_bits_tag),
    .io_in_0_bits_way(sinkC_task_arb_io_in_0_bits_way),
    .io_in_0_bits_bufIdx(sinkC_task_arb_io_in_0_bits_bufIdx),
    .io_in_0_bits_opcode(sinkC_task_arb_io_in_0_bits_opcode),
    .io_in_0_bits_source(sinkC_task_arb_io_in_0_bits_source),
    .io_in_0_bits_save(sinkC_task_arb_io_in_0_bits_save),
    .io_in_0_bits_drop(sinkC_task_arb_io_in_0_bits_drop),
    .io_in_0_bits_release(sinkC_task_arb_io_in_0_bits_release),
    .io_in_1_ready(sinkC_task_arb_io_in_1_ready),
    .io_in_1_valid(sinkC_task_arb_io_in_1_valid),
    .io_in_1_bits_set(sinkC_task_arb_io_in_1_bits_set),
    .io_in_1_bits_tag(sinkC_task_arb_io_in_1_bits_tag),
    .io_in_1_bits_way(sinkC_task_arb_io_in_1_bits_way),
    .io_in_1_bits_bufIdx(sinkC_task_arb_io_in_1_bits_bufIdx),
    .io_in_1_bits_opcode(sinkC_task_arb_io_in_1_bits_opcode),
    .io_in_1_bits_source(sinkC_task_arb_io_in_1_bits_source),
    .io_in_1_bits_save(sinkC_task_arb_io_in_1_bits_save),
    .io_in_1_bits_drop(sinkC_task_arb_io_in_1_bits_drop),
    .io_in_1_bits_release(sinkC_task_arb_io_in_1_bits_release),
    .io_in_2_ready(sinkC_task_arb_io_in_2_ready),
    .io_in_2_valid(sinkC_task_arb_io_in_2_valid),
    .io_in_2_bits_set(sinkC_task_arb_io_in_2_bits_set),
    .io_in_2_bits_tag(sinkC_task_arb_io_in_2_bits_tag),
    .io_in_2_bits_way(sinkC_task_arb_io_in_2_bits_way),
    .io_in_2_bits_bufIdx(sinkC_task_arb_io_in_2_bits_bufIdx),
    .io_in_2_bits_opcode(sinkC_task_arb_io_in_2_bits_opcode),
    .io_in_2_bits_source(sinkC_task_arb_io_in_2_bits_source),
    .io_in_2_bits_save(sinkC_task_arb_io_in_2_bits_save),
    .io_in_2_bits_drop(sinkC_task_arb_io_in_2_bits_drop),
    .io_in_2_bits_release(sinkC_task_arb_io_in_2_bits_release),
    .io_in_3_ready(sinkC_task_arb_io_in_3_ready),
    .io_in_3_valid(sinkC_task_arb_io_in_3_valid),
    .io_in_3_bits_set(sinkC_task_arb_io_in_3_bits_set),
    .io_in_3_bits_tag(sinkC_task_arb_io_in_3_bits_tag),
    .io_in_3_bits_way(sinkC_task_arb_io_in_3_bits_way),
    .io_in_3_bits_bufIdx(sinkC_task_arb_io_in_3_bits_bufIdx),
    .io_in_3_bits_opcode(sinkC_task_arb_io_in_3_bits_opcode),
    .io_in_3_bits_source(sinkC_task_arb_io_in_3_bits_source),
    .io_in_3_bits_save(sinkC_task_arb_io_in_3_bits_save),
    .io_in_3_bits_drop(sinkC_task_arb_io_in_3_bits_drop),
    .io_in_3_bits_release(sinkC_task_arb_io_in_3_bits_release),
    .io_in_4_ready(sinkC_task_arb_io_in_4_ready),
    .io_in_4_valid(sinkC_task_arb_io_in_4_valid),
    .io_in_4_bits_set(sinkC_task_arb_io_in_4_bits_set),
    .io_in_4_bits_tag(sinkC_task_arb_io_in_4_bits_tag),
    .io_in_4_bits_way(sinkC_task_arb_io_in_4_bits_way),
    .io_in_4_bits_bufIdx(sinkC_task_arb_io_in_4_bits_bufIdx),
    .io_in_4_bits_opcode(sinkC_task_arb_io_in_4_bits_opcode),
    .io_in_4_bits_source(sinkC_task_arb_io_in_4_bits_source),
    .io_in_4_bits_save(sinkC_task_arb_io_in_4_bits_save),
    .io_in_4_bits_drop(sinkC_task_arb_io_in_4_bits_drop),
    .io_in_4_bits_release(sinkC_task_arb_io_in_4_bits_release),
    .io_in_5_ready(sinkC_task_arb_io_in_5_ready),
    .io_in_5_valid(sinkC_task_arb_io_in_5_valid),
    .io_in_5_bits_set(sinkC_task_arb_io_in_5_bits_set),
    .io_in_5_bits_tag(sinkC_task_arb_io_in_5_bits_tag),
    .io_in_5_bits_way(sinkC_task_arb_io_in_5_bits_way),
    .io_in_5_bits_bufIdx(sinkC_task_arb_io_in_5_bits_bufIdx),
    .io_in_5_bits_opcode(sinkC_task_arb_io_in_5_bits_opcode),
    .io_in_5_bits_source(sinkC_task_arb_io_in_5_bits_source),
    .io_in_5_bits_save(sinkC_task_arb_io_in_5_bits_save),
    .io_in_5_bits_drop(sinkC_task_arb_io_in_5_bits_drop),
    .io_in_5_bits_release(sinkC_task_arb_io_in_5_bits_release),
    .io_in_6_ready(sinkC_task_arb_io_in_6_ready),
    .io_in_6_valid(sinkC_task_arb_io_in_6_valid),
    .io_in_6_bits_set(sinkC_task_arb_io_in_6_bits_set),
    .io_in_6_bits_tag(sinkC_task_arb_io_in_6_bits_tag),
    .io_in_6_bits_way(sinkC_task_arb_io_in_6_bits_way),
    .io_in_6_bits_bufIdx(sinkC_task_arb_io_in_6_bits_bufIdx),
    .io_in_6_bits_opcode(sinkC_task_arb_io_in_6_bits_opcode),
    .io_in_6_bits_source(sinkC_task_arb_io_in_6_bits_source),
    .io_in_6_bits_save(sinkC_task_arb_io_in_6_bits_save),
    .io_in_6_bits_drop(sinkC_task_arb_io_in_6_bits_drop),
    .io_in_6_bits_release(sinkC_task_arb_io_in_6_bits_release),
    .io_in_7_ready(sinkC_task_arb_io_in_7_ready),
    .io_in_7_valid(sinkC_task_arb_io_in_7_valid),
    .io_in_7_bits_set(sinkC_task_arb_io_in_7_bits_set),
    .io_in_7_bits_tag(sinkC_task_arb_io_in_7_bits_tag),
    .io_in_7_bits_way(sinkC_task_arb_io_in_7_bits_way),
    .io_in_7_bits_bufIdx(sinkC_task_arb_io_in_7_bits_bufIdx),
    .io_in_7_bits_opcode(sinkC_task_arb_io_in_7_bits_opcode),
    .io_in_7_bits_source(sinkC_task_arb_io_in_7_bits_source),
    .io_in_7_bits_save(sinkC_task_arb_io_in_7_bits_save),
    .io_in_7_bits_drop(sinkC_task_arb_io_in_7_bits_drop),
    .io_in_7_bits_release(sinkC_task_arb_io_in_7_bits_release),
    .io_in_8_ready(sinkC_task_arb_io_in_8_ready),
    .io_in_8_valid(sinkC_task_arb_io_in_8_valid),
    .io_in_8_bits_set(sinkC_task_arb_io_in_8_bits_set),
    .io_in_8_bits_tag(sinkC_task_arb_io_in_8_bits_tag),
    .io_in_8_bits_way(sinkC_task_arb_io_in_8_bits_way),
    .io_in_8_bits_bufIdx(sinkC_task_arb_io_in_8_bits_bufIdx),
    .io_in_8_bits_opcode(sinkC_task_arb_io_in_8_bits_opcode),
    .io_in_8_bits_source(sinkC_task_arb_io_in_8_bits_source),
    .io_in_8_bits_save(sinkC_task_arb_io_in_8_bits_save),
    .io_in_8_bits_drop(sinkC_task_arb_io_in_8_bits_drop),
    .io_in_8_bits_release(sinkC_task_arb_io_in_8_bits_release),
    .io_in_9_ready(sinkC_task_arb_io_in_9_ready),
    .io_in_9_valid(sinkC_task_arb_io_in_9_valid),
    .io_in_9_bits_set(sinkC_task_arb_io_in_9_bits_set),
    .io_in_9_bits_tag(sinkC_task_arb_io_in_9_bits_tag),
    .io_in_9_bits_way(sinkC_task_arb_io_in_9_bits_way),
    .io_in_9_bits_bufIdx(sinkC_task_arb_io_in_9_bits_bufIdx),
    .io_in_9_bits_opcode(sinkC_task_arb_io_in_9_bits_opcode),
    .io_in_9_bits_source(sinkC_task_arb_io_in_9_bits_source),
    .io_in_9_bits_save(sinkC_task_arb_io_in_9_bits_save),
    .io_in_9_bits_drop(sinkC_task_arb_io_in_9_bits_drop),
    .io_in_9_bits_release(sinkC_task_arb_io_in_9_bits_release),
    .io_in_10_ready(sinkC_task_arb_io_in_10_ready),
    .io_in_10_valid(sinkC_task_arb_io_in_10_valid),
    .io_in_10_bits_set(sinkC_task_arb_io_in_10_bits_set),
    .io_in_10_bits_tag(sinkC_task_arb_io_in_10_bits_tag),
    .io_in_10_bits_way(sinkC_task_arb_io_in_10_bits_way),
    .io_in_10_bits_bufIdx(sinkC_task_arb_io_in_10_bits_bufIdx),
    .io_in_10_bits_opcode(sinkC_task_arb_io_in_10_bits_opcode),
    .io_in_10_bits_source(sinkC_task_arb_io_in_10_bits_source),
    .io_in_10_bits_save(sinkC_task_arb_io_in_10_bits_save),
    .io_in_10_bits_drop(sinkC_task_arb_io_in_10_bits_drop),
    .io_in_10_bits_release(sinkC_task_arb_io_in_10_bits_release),
    .io_in_11_ready(sinkC_task_arb_io_in_11_ready),
    .io_in_11_valid(sinkC_task_arb_io_in_11_valid),
    .io_in_11_bits_set(sinkC_task_arb_io_in_11_bits_set),
    .io_in_11_bits_tag(sinkC_task_arb_io_in_11_bits_tag),
    .io_in_11_bits_way(sinkC_task_arb_io_in_11_bits_way),
    .io_in_11_bits_bufIdx(sinkC_task_arb_io_in_11_bits_bufIdx),
    .io_in_11_bits_opcode(sinkC_task_arb_io_in_11_bits_opcode),
    .io_in_11_bits_source(sinkC_task_arb_io_in_11_bits_source),
    .io_in_11_bits_save(sinkC_task_arb_io_in_11_bits_save),
    .io_in_11_bits_drop(sinkC_task_arb_io_in_11_bits_drop),
    .io_in_11_bits_release(sinkC_task_arb_io_in_11_bits_release),
    .io_in_12_ready(sinkC_task_arb_io_in_12_ready),
    .io_in_12_valid(sinkC_task_arb_io_in_12_valid),
    .io_in_12_bits_set(sinkC_task_arb_io_in_12_bits_set),
    .io_in_12_bits_tag(sinkC_task_arb_io_in_12_bits_tag),
    .io_in_12_bits_way(sinkC_task_arb_io_in_12_bits_way),
    .io_in_12_bits_bufIdx(sinkC_task_arb_io_in_12_bits_bufIdx),
    .io_in_12_bits_opcode(sinkC_task_arb_io_in_12_bits_opcode),
    .io_in_12_bits_source(sinkC_task_arb_io_in_12_bits_source),
    .io_in_12_bits_save(sinkC_task_arb_io_in_12_bits_save),
    .io_in_12_bits_drop(sinkC_task_arb_io_in_12_bits_drop),
    .io_in_12_bits_release(sinkC_task_arb_io_in_12_bits_release),
    .io_in_13_ready(sinkC_task_arb_io_in_13_ready),
    .io_in_13_valid(sinkC_task_arb_io_in_13_valid),
    .io_in_13_bits_set(sinkC_task_arb_io_in_13_bits_set),
    .io_in_13_bits_tag(sinkC_task_arb_io_in_13_bits_tag),
    .io_in_13_bits_way(sinkC_task_arb_io_in_13_bits_way),
    .io_in_13_bits_bufIdx(sinkC_task_arb_io_in_13_bits_bufIdx),
    .io_in_13_bits_opcode(sinkC_task_arb_io_in_13_bits_opcode),
    .io_in_13_bits_source(sinkC_task_arb_io_in_13_bits_source),
    .io_in_13_bits_save(sinkC_task_arb_io_in_13_bits_save),
    .io_in_13_bits_drop(sinkC_task_arb_io_in_13_bits_drop),
    .io_in_13_bits_release(sinkC_task_arb_io_in_13_bits_release),
    .io_out_ready(sinkC_task_arb_io_out_ready),
    .io_out_valid(sinkC_task_arb_io_out_valid),
    .io_out_bits_set(sinkC_task_arb_io_out_bits_set),
    .io_out_bits_tag(sinkC_task_arb_io_out_bits_tag),
    .io_out_bits_way(sinkC_task_arb_io_out_bits_way),
    .io_out_bits_bufIdx(sinkC_task_arb_io_out_bits_bufIdx),
    .io_out_bits_opcode(sinkC_task_arb_io_out_bits_opcode),
    .io_out_bits_source(sinkC_task_arb_io_out_bits_source),
    .io_out_bits_save(sinkC_task_arb_io_out_bits_save),
    .io_out_bits_drop(sinkC_task_arb_io_out_bits_drop),
    .io_out_bits_release(sinkC_task_arb_io_out_bits_release)
  );
  Pipeline_2 pipeline_1 ( // @[Pipeline.scala 39:26]
    .clock(pipeline_1_clock),
    .reset(pipeline_1_reset),
    .io_in_valid(pipeline_1_io_in_valid),
    .io_in_bits_set(pipeline_1_io_in_bits_set),
    .io_in_bits_way(pipeline_1_io_in_bits_way),
    .io_in_bits_tag(pipeline_1_io_in_bits_tag),
    .io_out_valid(pipeline_1_io_out_valid),
    .io_out_bits_set(pipeline_1_io_out_bits_set),
    .io_out_bits_way(pipeline_1_io_out_bits_way),
    .io_out_bits_tag(pipeline_1_io_out_bits_tag)
  );
  FastArbiter_3 tagWrite_task_arb ( // @[Slice.scala 468:27]
    .clock(tagWrite_task_arb_clock),
    .reset(tagWrite_task_arb_reset),
    .io_in_0_ready(tagWrite_task_arb_io_in_0_ready),
    .io_in_0_valid(tagWrite_task_arb_io_in_0_valid),
    .io_in_0_bits_set(tagWrite_task_arb_io_in_0_bits_set),
    .io_in_0_bits_way(tagWrite_task_arb_io_in_0_bits_way),
    .io_in_0_bits_tag(tagWrite_task_arb_io_in_0_bits_tag),
    .io_in_1_ready(tagWrite_task_arb_io_in_1_ready),
    .io_in_1_valid(tagWrite_task_arb_io_in_1_valid),
    .io_in_1_bits_set(tagWrite_task_arb_io_in_1_bits_set),
    .io_in_1_bits_way(tagWrite_task_arb_io_in_1_bits_way),
    .io_in_1_bits_tag(tagWrite_task_arb_io_in_1_bits_tag),
    .io_in_2_ready(tagWrite_task_arb_io_in_2_ready),
    .io_in_2_valid(tagWrite_task_arb_io_in_2_valid),
    .io_in_2_bits_set(tagWrite_task_arb_io_in_2_bits_set),
    .io_in_2_bits_way(tagWrite_task_arb_io_in_2_bits_way),
    .io_in_2_bits_tag(tagWrite_task_arb_io_in_2_bits_tag),
    .io_in_3_ready(tagWrite_task_arb_io_in_3_ready),
    .io_in_3_valid(tagWrite_task_arb_io_in_3_valid),
    .io_in_3_bits_set(tagWrite_task_arb_io_in_3_bits_set),
    .io_in_3_bits_way(tagWrite_task_arb_io_in_3_bits_way),
    .io_in_3_bits_tag(tagWrite_task_arb_io_in_3_bits_tag),
    .io_in_4_ready(tagWrite_task_arb_io_in_4_ready),
    .io_in_4_valid(tagWrite_task_arb_io_in_4_valid),
    .io_in_4_bits_set(tagWrite_task_arb_io_in_4_bits_set),
    .io_in_4_bits_way(tagWrite_task_arb_io_in_4_bits_way),
    .io_in_4_bits_tag(tagWrite_task_arb_io_in_4_bits_tag),
    .io_in_5_ready(tagWrite_task_arb_io_in_5_ready),
    .io_in_5_valid(tagWrite_task_arb_io_in_5_valid),
    .io_in_5_bits_set(tagWrite_task_arb_io_in_5_bits_set),
    .io_in_5_bits_way(tagWrite_task_arb_io_in_5_bits_way),
    .io_in_5_bits_tag(tagWrite_task_arb_io_in_5_bits_tag),
    .io_in_6_ready(tagWrite_task_arb_io_in_6_ready),
    .io_in_6_valid(tagWrite_task_arb_io_in_6_valid),
    .io_in_6_bits_set(tagWrite_task_arb_io_in_6_bits_set),
    .io_in_6_bits_way(tagWrite_task_arb_io_in_6_bits_way),
    .io_in_6_bits_tag(tagWrite_task_arb_io_in_6_bits_tag),
    .io_in_7_ready(tagWrite_task_arb_io_in_7_ready),
    .io_in_7_valid(tagWrite_task_arb_io_in_7_valid),
    .io_in_7_bits_set(tagWrite_task_arb_io_in_7_bits_set),
    .io_in_7_bits_way(tagWrite_task_arb_io_in_7_bits_way),
    .io_in_7_bits_tag(tagWrite_task_arb_io_in_7_bits_tag),
    .io_in_8_ready(tagWrite_task_arb_io_in_8_ready),
    .io_in_8_valid(tagWrite_task_arb_io_in_8_valid),
    .io_in_8_bits_set(tagWrite_task_arb_io_in_8_bits_set),
    .io_in_8_bits_way(tagWrite_task_arb_io_in_8_bits_way),
    .io_in_8_bits_tag(tagWrite_task_arb_io_in_8_bits_tag),
    .io_in_9_ready(tagWrite_task_arb_io_in_9_ready),
    .io_in_9_valid(tagWrite_task_arb_io_in_9_valid),
    .io_in_9_bits_set(tagWrite_task_arb_io_in_9_bits_set),
    .io_in_9_bits_way(tagWrite_task_arb_io_in_9_bits_way),
    .io_in_9_bits_tag(tagWrite_task_arb_io_in_9_bits_tag),
    .io_in_10_ready(tagWrite_task_arb_io_in_10_ready),
    .io_in_10_valid(tagWrite_task_arb_io_in_10_valid),
    .io_in_10_bits_set(tagWrite_task_arb_io_in_10_bits_set),
    .io_in_10_bits_way(tagWrite_task_arb_io_in_10_bits_way),
    .io_in_10_bits_tag(tagWrite_task_arb_io_in_10_bits_tag),
    .io_in_11_ready(tagWrite_task_arb_io_in_11_ready),
    .io_in_11_valid(tagWrite_task_arb_io_in_11_valid),
    .io_in_11_bits_set(tagWrite_task_arb_io_in_11_bits_set),
    .io_in_11_bits_way(tagWrite_task_arb_io_in_11_bits_way),
    .io_in_11_bits_tag(tagWrite_task_arb_io_in_11_bits_tag),
    .io_in_12_ready(tagWrite_task_arb_io_in_12_ready),
    .io_in_12_valid(tagWrite_task_arb_io_in_12_valid),
    .io_in_12_bits_set(tagWrite_task_arb_io_in_12_bits_set),
    .io_in_12_bits_way(tagWrite_task_arb_io_in_12_bits_way),
    .io_in_12_bits_tag(tagWrite_task_arb_io_in_12_bits_tag),
    .io_in_13_ready(tagWrite_task_arb_io_in_13_ready),
    .io_in_13_valid(tagWrite_task_arb_io_in_13_valid),
    .io_in_13_bits_set(tagWrite_task_arb_io_in_13_bits_set),
    .io_in_13_bits_way(tagWrite_task_arb_io_in_13_bits_way),
    .io_in_13_bits_tag(tagWrite_task_arb_io_in_13_bits_tag),
    .io_out_ready(tagWrite_task_arb_io_out_ready),
    .io_out_valid(tagWrite_task_arb_io_out_valid),
    .io_out_bits_set(tagWrite_task_arb_io_out_bits_set),
    .io_out_bits_way(tagWrite_task_arb_io_out_bits_way),
    .io_out_bits_tag(tagWrite_task_arb_io_out_bits_tag)
  );
  Pipeline_3 pipeline_2 ( // @[Pipeline.scala 39:26]
    .clock(pipeline_2_clock),
    .reset(pipeline_2_reset),
    .io_in_valid(pipeline_2_io_in_valid),
    .io_in_bits_set(pipeline_2_io_in_bits_set),
    .io_in_bits_way(pipeline_2_io_in_bits_way),
    .io_in_bits_data_0_state(pipeline_2_io_in_bits_data_0_state),
    .io_in_bits_data_1_state(pipeline_2_io_in_bits_data_1_state),
    .io_out_valid(pipeline_2_io_out_valid),
    .io_out_bits_set(pipeline_2_io_out_bits_set),
    .io_out_bits_way(pipeline_2_io_out_bits_way),
    .io_out_bits_data_0_state(pipeline_2_io_out_bits_data_0_state),
    .io_out_bits_data_1_state(pipeline_2_io_out_bits_data_1_state)
  );
  FastArbiter_4 arbiter_1 ( // @[Slice.scala 405:25]
    .clock(arbiter_1_clock),
    .reset(arbiter_1_reset),
    .io_in_0_ready(arbiter_1_io_in_0_ready),
    .io_in_0_valid(arbiter_1_io_in_0_valid),
    .io_in_0_bits_set(arbiter_1_io_in_0_bits_set),
    .io_in_0_bits_way(arbiter_1_io_in_0_bits_way),
    .io_in_0_bits_data_0_state(arbiter_1_io_in_0_bits_data_0_state),
    .io_in_0_bits_data_1_state(arbiter_1_io_in_0_bits_data_1_state),
    .io_in_1_ready(arbiter_1_io_in_1_ready),
    .io_in_1_valid(arbiter_1_io_in_1_valid),
    .io_in_1_bits_set(arbiter_1_io_in_1_bits_set),
    .io_in_1_bits_way(arbiter_1_io_in_1_bits_way),
    .io_in_1_bits_data_0_state(arbiter_1_io_in_1_bits_data_0_state),
    .io_in_1_bits_data_1_state(arbiter_1_io_in_1_bits_data_1_state),
    .io_in_2_ready(arbiter_1_io_in_2_ready),
    .io_in_2_valid(arbiter_1_io_in_2_valid),
    .io_in_2_bits_set(arbiter_1_io_in_2_bits_set),
    .io_in_2_bits_way(arbiter_1_io_in_2_bits_way),
    .io_in_2_bits_data_0_state(arbiter_1_io_in_2_bits_data_0_state),
    .io_in_2_bits_data_1_state(arbiter_1_io_in_2_bits_data_1_state),
    .io_in_3_ready(arbiter_1_io_in_3_ready),
    .io_in_3_valid(arbiter_1_io_in_3_valid),
    .io_in_3_bits_set(arbiter_1_io_in_3_bits_set),
    .io_in_3_bits_way(arbiter_1_io_in_3_bits_way),
    .io_in_3_bits_data_0_state(arbiter_1_io_in_3_bits_data_0_state),
    .io_in_3_bits_data_1_state(arbiter_1_io_in_3_bits_data_1_state),
    .io_in_4_ready(arbiter_1_io_in_4_ready),
    .io_in_4_valid(arbiter_1_io_in_4_valid),
    .io_in_4_bits_set(arbiter_1_io_in_4_bits_set),
    .io_in_4_bits_way(arbiter_1_io_in_4_bits_way),
    .io_in_4_bits_data_0_state(arbiter_1_io_in_4_bits_data_0_state),
    .io_in_4_bits_data_1_state(arbiter_1_io_in_4_bits_data_1_state),
    .io_in_5_ready(arbiter_1_io_in_5_ready),
    .io_in_5_valid(arbiter_1_io_in_5_valid),
    .io_in_5_bits_set(arbiter_1_io_in_5_bits_set),
    .io_in_5_bits_way(arbiter_1_io_in_5_bits_way),
    .io_in_5_bits_data_0_state(arbiter_1_io_in_5_bits_data_0_state),
    .io_in_5_bits_data_1_state(arbiter_1_io_in_5_bits_data_1_state),
    .io_in_6_ready(arbiter_1_io_in_6_ready),
    .io_in_6_valid(arbiter_1_io_in_6_valid),
    .io_in_6_bits_set(arbiter_1_io_in_6_bits_set),
    .io_in_6_bits_way(arbiter_1_io_in_6_bits_way),
    .io_in_6_bits_data_0_state(arbiter_1_io_in_6_bits_data_0_state),
    .io_in_6_bits_data_1_state(arbiter_1_io_in_6_bits_data_1_state),
    .io_in_7_ready(arbiter_1_io_in_7_ready),
    .io_in_7_valid(arbiter_1_io_in_7_valid),
    .io_in_7_bits_set(arbiter_1_io_in_7_bits_set),
    .io_in_7_bits_way(arbiter_1_io_in_7_bits_way),
    .io_in_7_bits_data_0_state(arbiter_1_io_in_7_bits_data_0_state),
    .io_in_7_bits_data_1_state(arbiter_1_io_in_7_bits_data_1_state),
    .io_in_8_ready(arbiter_1_io_in_8_ready),
    .io_in_8_valid(arbiter_1_io_in_8_valid),
    .io_in_8_bits_set(arbiter_1_io_in_8_bits_set),
    .io_in_8_bits_way(arbiter_1_io_in_8_bits_way),
    .io_in_8_bits_data_0_state(arbiter_1_io_in_8_bits_data_0_state),
    .io_in_8_bits_data_1_state(arbiter_1_io_in_8_bits_data_1_state),
    .io_in_9_ready(arbiter_1_io_in_9_ready),
    .io_in_9_valid(arbiter_1_io_in_9_valid),
    .io_in_9_bits_set(arbiter_1_io_in_9_bits_set),
    .io_in_9_bits_way(arbiter_1_io_in_9_bits_way),
    .io_in_9_bits_data_0_state(arbiter_1_io_in_9_bits_data_0_state),
    .io_in_9_bits_data_1_state(arbiter_1_io_in_9_bits_data_1_state),
    .io_in_10_ready(arbiter_1_io_in_10_ready),
    .io_in_10_valid(arbiter_1_io_in_10_valid),
    .io_in_10_bits_set(arbiter_1_io_in_10_bits_set),
    .io_in_10_bits_way(arbiter_1_io_in_10_bits_way),
    .io_in_10_bits_data_0_state(arbiter_1_io_in_10_bits_data_0_state),
    .io_in_10_bits_data_1_state(arbiter_1_io_in_10_bits_data_1_state),
    .io_in_11_ready(arbiter_1_io_in_11_ready),
    .io_in_11_valid(arbiter_1_io_in_11_valid),
    .io_in_11_bits_set(arbiter_1_io_in_11_bits_set),
    .io_in_11_bits_way(arbiter_1_io_in_11_bits_way),
    .io_in_11_bits_data_0_state(arbiter_1_io_in_11_bits_data_0_state),
    .io_in_11_bits_data_1_state(arbiter_1_io_in_11_bits_data_1_state),
    .io_in_12_ready(arbiter_1_io_in_12_ready),
    .io_in_12_valid(arbiter_1_io_in_12_valid),
    .io_in_12_bits_set(arbiter_1_io_in_12_bits_set),
    .io_in_12_bits_way(arbiter_1_io_in_12_bits_way),
    .io_in_12_bits_data_0_state(arbiter_1_io_in_12_bits_data_0_state),
    .io_in_12_bits_data_1_state(arbiter_1_io_in_12_bits_data_1_state),
    .io_in_13_ready(arbiter_1_io_in_13_ready),
    .io_in_13_valid(arbiter_1_io_in_13_valid),
    .io_in_13_bits_set(arbiter_1_io_in_13_bits_set),
    .io_in_13_bits_way(arbiter_1_io_in_13_bits_way),
    .io_in_13_bits_data_0_state(arbiter_1_io_in_13_bits_data_0_state),
    .io_in_13_bits_data_1_state(arbiter_1_io_in_13_bits_data_1_state),
    .io_in_14_ready(arbiter_1_io_in_14_ready),
    .io_in_14_valid(arbiter_1_io_in_14_valid),
    .io_in_14_bits_set(arbiter_1_io_in_14_bits_set),
    .io_in_14_bits_way(arbiter_1_io_in_14_bits_way),
    .io_in_14_bits_data_0_state(arbiter_1_io_in_14_bits_data_0_state),
    .io_in_14_bits_data_1_state(arbiter_1_io_in_14_bits_data_1_state),
    .io_in_15_ready(arbiter_1_io_in_15_ready),
    .io_in_15_valid(arbiter_1_io_in_15_valid),
    .io_in_15_bits_set(arbiter_1_io_in_15_bits_set),
    .io_in_15_bits_way(arbiter_1_io_in_15_bits_way),
    .io_in_15_bits_data_0_state(arbiter_1_io_in_15_bits_data_0_state),
    .io_in_15_bits_data_1_state(arbiter_1_io_in_15_bits_data_1_state),
    .io_out_valid(arbiter_1_io_out_valid),
    .io_out_bits_set(arbiter_1_io_out_bits_set),
    .io_out_bits_way(arbiter_1_io_out_bits_way),
    .io_out_bits_data_0_state(arbiter_1_io_out_bits_data_0_state),
    .io_out_bits_data_1_state(arbiter_1_io_out_bits_data_1_state)
  );
  Pipeline_4 pipeline_3 ( // @[Pipeline.scala 39:26]
    .clock(pipeline_3_clock),
    .reset(pipeline_3_reset),
    .io_in_valid(pipeline_3_io_in_valid),
    .io_in_bits_set(pipeline_3_io_in_bits_set),
    .io_in_bits_way(pipeline_3_io_in_bits_way),
    .io_in_bits_tag(pipeline_3_io_in_bits_tag),
    .io_out_valid(pipeline_3_io_out_valid),
    .io_out_bits_set(pipeline_3_io_out_bits_set),
    .io_out_bits_way(pipeline_3_io_out_bits_way),
    .io_out_bits_tag(pipeline_3_io_out_bits_tag)
  );
  FastArbiter_5 arbiter_2 ( // @[Slice.scala 468:27]
    .clock(arbiter_2_clock),
    .reset(arbiter_2_reset),
    .io_in_0_ready(arbiter_2_io_in_0_ready),
    .io_in_0_valid(arbiter_2_io_in_0_valid),
    .io_in_0_bits_set(arbiter_2_io_in_0_bits_set),
    .io_in_0_bits_way(arbiter_2_io_in_0_bits_way),
    .io_in_0_bits_tag(arbiter_2_io_in_0_bits_tag),
    .io_in_1_ready(arbiter_2_io_in_1_ready),
    .io_in_1_valid(arbiter_2_io_in_1_valid),
    .io_in_1_bits_set(arbiter_2_io_in_1_bits_set),
    .io_in_1_bits_way(arbiter_2_io_in_1_bits_way),
    .io_in_1_bits_tag(arbiter_2_io_in_1_bits_tag),
    .io_in_2_ready(arbiter_2_io_in_2_ready),
    .io_in_2_valid(arbiter_2_io_in_2_valid),
    .io_in_2_bits_set(arbiter_2_io_in_2_bits_set),
    .io_in_2_bits_way(arbiter_2_io_in_2_bits_way),
    .io_in_2_bits_tag(arbiter_2_io_in_2_bits_tag),
    .io_in_3_ready(arbiter_2_io_in_3_ready),
    .io_in_3_valid(arbiter_2_io_in_3_valid),
    .io_in_3_bits_set(arbiter_2_io_in_3_bits_set),
    .io_in_3_bits_way(arbiter_2_io_in_3_bits_way),
    .io_in_3_bits_tag(arbiter_2_io_in_3_bits_tag),
    .io_in_4_ready(arbiter_2_io_in_4_ready),
    .io_in_4_valid(arbiter_2_io_in_4_valid),
    .io_in_4_bits_set(arbiter_2_io_in_4_bits_set),
    .io_in_4_bits_way(arbiter_2_io_in_4_bits_way),
    .io_in_4_bits_tag(arbiter_2_io_in_4_bits_tag),
    .io_in_5_ready(arbiter_2_io_in_5_ready),
    .io_in_5_valid(arbiter_2_io_in_5_valid),
    .io_in_5_bits_set(arbiter_2_io_in_5_bits_set),
    .io_in_5_bits_way(arbiter_2_io_in_5_bits_way),
    .io_in_5_bits_tag(arbiter_2_io_in_5_bits_tag),
    .io_in_6_ready(arbiter_2_io_in_6_ready),
    .io_in_6_valid(arbiter_2_io_in_6_valid),
    .io_in_6_bits_set(arbiter_2_io_in_6_bits_set),
    .io_in_6_bits_way(arbiter_2_io_in_6_bits_way),
    .io_in_6_bits_tag(arbiter_2_io_in_6_bits_tag),
    .io_in_7_ready(arbiter_2_io_in_7_ready),
    .io_in_7_valid(arbiter_2_io_in_7_valid),
    .io_in_7_bits_set(arbiter_2_io_in_7_bits_set),
    .io_in_7_bits_way(arbiter_2_io_in_7_bits_way),
    .io_in_7_bits_tag(arbiter_2_io_in_7_bits_tag),
    .io_in_8_ready(arbiter_2_io_in_8_ready),
    .io_in_8_valid(arbiter_2_io_in_8_valid),
    .io_in_8_bits_set(arbiter_2_io_in_8_bits_set),
    .io_in_8_bits_way(arbiter_2_io_in_8_bits_way),
    .io_in_8_bits_tag(arbiter_2_io_in_8_bits_tag),
    .io_in_9_ready(arbiter_2_io_in_9_ready),
    .io_in_9_valid(arbiter_2_io_in_9_valid),
    .io_in_9_bits_set(arbiter_2_io_in_9_bits_set),
    .io_in_9_bits_way(arbiter_2_io_in_9_bits_way),
    .io_in_9_bits_tag(arbiter_2_io_in_9_bits_tag),
    .io_in_10_ready(arbiter_2_io_in_10_ready),
    .io_in_10_valid(arbiter_2_io_in_10_valid),
    .io_in_10_bits_set(arbiter_2_io_in_10_bits_set),
    .io_in_10_bits_way(arbiter_2_io_in_10_bits_way),
    .io_in_10_bits_tag(arbiter_2_io_in_10_bits_tag),
    .io_in_11_ready(arbiter_2_io_in_11_ready),
    .io_in_11_valid(arbiter_2_io_in_11_valid),
    .io_in_11_bits_set(arbiter_2_io_in_11_bits_set),
    .io_in_11_bits_way(arbiter_2_io_in_11_bits_way),
    .io_in_11_bits_tag(arbiter_2_io_in_11_bits_tag),
    .io_in_12_ready(arbiter_2_io_in_12_ready),
    .io_in_12_valid(arbiter_2_io_in_12_valid),
    .io_in_12_bits_set(arbiter_2_io_in_12_bits_set),
    .io_in_12_bits_way(arbiter_2_io_in_12_bits_way),
    .io_in_12_bits_tag(arbiter_2_io_in_12_bits_tag),
    .io_in_13_ready(arbiter_2_io_in_13_ready),
    .io_in_13_valid(arbiter_2_io_in_13_valid),
    .io_in_13_bits_set(arbiter_2_io_in_13_bits_set),
    .io_in_13_bits_way(arbiter_2_io_in_13_bits_way),
    .io_in_13_bits_tag(arbiter_2_io_in_13_bits_tag),
    .io_out_ready(arbiter_2_io_out_ready),
    .io_out_valid(arbiter_2_io_out_valid),
    .io_out_bits_set(arbiter_2_io_out_bits_set),
    .io_out_bits_way(arbiter_2_io_out_bits_way),
    .io_out_bits_tag(arbiter_2_io_out_bits_tag)
  );
  assign io_in_a_ready = sinkA_io_a_ready; // @[Slice.scala 63:14]
  assign io_in_bvalid = sourceB_io_bvalid; // @[Slice.scala 64:11]
  assign io_in_bparam = sourceB_io_bparam; // @[Slice.scala 64:11]
  assign io_in_bsource = sourceB_io_bsource; // @[Slice.scala 64:11]
  assign io_in_baddress = sourceB_io_baddress; // @[Slice.scala 64:11]
  assign io_in_bdata = sourceB_io_bdata; // @[Slice.scala 64:11]
  assign io_in_c_ready = sinkC_io_c_ready; // @[Slice.scala 65:14]
  assign io_in_d_valid = sourceD_io_d_valid; // @[Slice.scala 66:11]
  assign io_in_d_bits_opcode = sourceD_io_d_bits_opcode; // @[Slice.scala 66:11]
  assign io_in_d_bits_param = sourceD_io_d_bits_param; // @[Slice.scala 66:11]
  assign io_in_d_bits_size = sourceD_io_d_bits_size; // @[Slice.scala 66:11]
  assign io_in_d_bits_source = sourceD_io_d_bits_source; // @[Slice.scala 66:11]
  assign io_in_d_bits_sink = sourceD_io_d_bits_sink; // @[Slice.scala 66:11]
  assign io_in_d_bits_denied = sourceD_io_d_bits_denied; // @[Slice.scala 66:11]
  assign io_in_d_bits_echo_blockisdirty = sourceD_io_d_bits_echo_blockisdirty; // @[Slice.scala 66:11]
  assign io_in_d_bits_data = sourceD_io_d_bits_data; // @[Slice.scala 66:11]
  assign io_in_d_bits_corrupt = sourceD_io_d_bits_corrupt; // @[Slice.scala 66:11]
  assign io_out_a_valid = io_out_a_q_io_deq_valid; // @[Slice.scala 82:12]
  assign io_out_a_bits_opcode = io_out_a_q_io_deq_bits_opcode; // @[Slice.scala 82:12]
  assign io_out_a_bits_param = io_out_a_q_io_deq_bits_param; // @[Slice.scala 82:12]
  assign io_out_a_bits_size = io_out_a_q_io_deq_bits_size; // @[Slice.scala 82:12]
  assign io_out_a_bits_source = io_out_a_q_io_deq_bits_source; // @[Slice.scala 82:12]
  assign io_out_a_bits_address = io_out_a_q_io_deq_bits_address; // @[Slice.scala 82:12]
  assign io_out_a_bits_mask = io_out_a_q_io_deq_bits_mask; // @[Slice.scala 82:12]
  assign io_out_a_bits_data = io_out_a_q_io_deq_bits_data; // @[Slice.scala 82:12]
  assign io_out_c_valid = io_out_c_q_io_deq_valid; // @[Slice.scala 86:12]
  assign io_out_c_bits_opcode = io_out_c_q_io_deq_bits_opcode; // @[Slice.scala 86:12]
  assign io_out_c_bits_size = io_out_c_q_io_deq_bits_size; // @[Slice.scala 86:12]
  assign io_out_c_bits_source = io_out_c_q_io_deq_bits_source; // @[Slice.scala 86:12]
  assign io_out_c_bits_address = io_out_c_q_io_deq_bits_address; // @[Slice.scala 86:12]
  assign io_out_c_bits_data = io_out_c_q_io_deq_bits_data; // @[Slice.scala 86:12]
  assign io_out_d_ready = sinkD_io_d_q_io_enq_ready; // @[Decoupled.scala 365:17]
  assign io_out_e_valid = io_out_e_q_io_deq_valid; // @[Slice.scala 88:12]
  assign io_out_e_bits_sink = io_out_e_q_io_deq_bits_sink; // @[Slice.scala 88:12]
  assign sinkA_clock = clock;
  assign sinkA_reset = reset;
  assign sinkA_io_a_valid = io_in_a_valid; // @[Slice.scala 63:14]
  assign sinkA_io_a_bits_opcode = io_in_a_bits_opcode; // @[Slice.scala 63:14]
  assign sinkA_io_a_bits_param = io_in_a_bits_param; // @[Slice.scala 63:14]
  assign sinkA_io_a_bits_size = io_in_a_bits_size; // @[Slice.scala 63:14]
  assign sinkA_io_a_bits_source = io_in_a_bits_source; // @[Slice.scala 63:14]
  assign sinkA_io_a_bits_address = io_in_a_bits_address; // @[Slice.scala 63:14]
  assign sinkA_io_a_bits_user_preferCache = io_in_a_bits_user_preferCache; // @[Slice.scala 63:14]
  assign sinkA_io_a_bits_mask = io_in_a_bits_mask; // @[Slice.scala 63:14]
  assign sinkA_io_a_bits_data = io_in_a_bits_data; // @[Slice.scala 63:14]
  assign sinkA_io_alloc_ready = _a_req_valid_T & a_req_ready; // @[Slice.scala 391:28]
  assign sinkA_io_d_pb_pop_valid = sourceD_io_pb_pop_valid; // @[Slice.scala 586:21]
  assign sinkA_io_d_pb_pop_bits_bufIdx = sourceD_io_pb_pop_bits_bufIdx; // @[Slice.scala 586:21]
  assign sinkA_io_d_pb_pop_bits_count = sourceD_io_pb_pop_bits_count; // @[Slice.scala 586:21]
  assign sinkA_io_d_pb_pop_bits_last = sourceD_io_pb_pop_bits_last; // @[Slice.scala 586:21]
  assign sinkA_io_a_pb_pop_valid = sourceA_io_pb_pop_valid; // @[Slice.scala 589:21]
  assign sinkA_io_a_pb_pop_bits_bufIdx = sourceA_io_pb_pop_bits_bufIdx; // @[Slice.scala 589:21]
  assign sinkA_io_a_pb_pop_bits_count = sourceA_io_pb_pop_bits_count; // @[Slice.scala 589:21]
  assign sinkA_io_a_pb_pop_bits_last = sourceA_io_pb_pop_bits_last; // @[Slice.scala 589:21]
  assign sourceB_clock = clock;
  assign sourceB_reset = reset;
  assign sourceB_io_bready = io_in_bready; // @[Slice.scala 64:11]
  assign sourceB_io_task_valid = c_real_valid_1 | bc_real_valid_1 | sourceB_task_arb_io_out_valid; // @[Slice.scala 489:52]
  assign sourceB_io_task_bits_set = c_real_valid_1 ? c_bits_latch_1_set : _sourceB_io_task_bits_T_set; // @[Slice.scala 490:24]
  assign sourceB_io_task_bits_tag = c_real_valid_1 ? c_bits_latch_1_tag : _sourceB_io_task_bits_T_tag; // @[Slice.scala 490:24]
  assign sourceB_io_task_bits_param = c_real_valid_1 ? c_bits_latch_1_param : _sourceB_io_task_bits_T_param; // @[Slice.scala 490:24]
  assign sourceB_io_task_bits_clients = c_real_valid_1 ? c_bits_latch_1_clients : _sourceB_io_task_bits_T_clients; // @[Slice.scala 490:24]
  assign sourceB_io_task_bits_needData = c_real_valid_1 ? c_bits_latch_1_needData : _sourceB_io_task_bits_T_needData; // @[Slice.scala 490:24]
  assign sinkC_clock = clock;
  assign sinkC_reset = reset;
  assign sinkC_io_c_valid = io_in_c_valid; // @[Slice.scala 65:14]
  assign sinkC_io_c_bits_opcode = io_in_c_bits_opcode; // @[Slice.scala 65:14]
  assign sinkC_io_c_bits_param = io_in_c_bits_param; // @[Slice.scala 65:14]
  assign sinkC_io_c_bits_size = io_in_c_bits_size; // @[Slice.scala 65:14]
  assign sinkC_io_c_bits_source = io_in_c_bits_source; // @[Slice.scala 65:14]
  assign sinkC_io_c_bits_address = io_in_c_bits_address; // @[Slice.scala 65:14]
  assign sinkC_io_c_bits_echo_blockisdirty = io_in_c_bits_echo_blockisdirty; // @[Slice.scala 65:14]
  assign sinkC_io_c_bits_data = io_in_c_bits_data; // @[Slice.scala 65:14]
  assign sinkC_io_alloc_ready = mshrAlloc_io_c_req_ready; // @[Slice.scala 161:24]
  assign sinkC_io_task_valid = c_real_valid_6 | bc_real_valid_6 | sinkC_task_arb_io_out_valid; // @[Slice.scala 489:52]
  assign sinkC_io_task_bits_set = c_real_valid_6 ? c_bits_latch_6_set : _sinkC_io_task_bits_T_set; // @[Slice.scala 490:24]
  assign sinkC_io_task_bits_tag = c_real_valid_6 ? c_bits_latch_6_tag : _sinkC_io_task_bits_T_tag; // @[Slice.scala 490:24]
  assign sinkC_io_task_bits_way = c_real_valid_6 ? c_bits_latch_6_way : _sinkC_io_task_bits_T_way; // @[Slice.scala 490:24]
  assign sinkC_io_task_bits_bufIdx = c_real_valid_6 ? c_bits_latch_6_bufIdx : _sinkC_io_task_bits_T_bufIdx; // @[Slice.scala 490:24]
  assign sinkC_io_task_bits_opcode = c_real_valid_6 ? c_bits_latch_6_opcode : _sinkC_io_task_bits_T_opcode; // @[Slice.scala 490:24]
  assign sinkC_io_task_bits_source = c_real_valid_6 ? c_bits_latch_6_source : _sinkC_io_task_bits_T_source; // @[Slice.scala 490:24]
  assign sinkC_io_task_bits_save = c_real_valid_6 ? c_bits_latch_6_save : _sinkC_io_task_bits_T_save; // @[Slice.scala 490:24]
  assign sinkC_io_task_bits_drop = c_real_valid_6 ? c_bits_latch_6_drop : _sinkC_io_task_bits_T_drop; // @[Slice.scala 490:24]
  assign sinkC_io_task_bits_release = c_real_valid_6 ? c_bits_latch_6_release : _sinkC_io_task_bits_T_release; // @[Slice.scala 490:24]
  assign sinkC_io_bs_waddr_ready = dataStorage_io_sinkC_waddr_ready; // @[Slice.scala 114:30]
  assign sinkC_io_sourceD_rhazard_valid = sourceD_io_sourceD_rhazard_valid; // @[Slice.scala 583:29]
  assign sinkC_io_sourceD_rhazard_bits_way = sourceD_io_sourceD_rhazard_bits_way; // @[Slice.scala 583:29]
  assign sinkC_io_sourceD_rhazard_bits_set = sourceD_io_sourceD_rhazard_bits_set; // @[Slice.scala 583:29]
  assign sinkC_io_release_ready = out_c_ready & allowed_0; // @[Arbiter.scala 123:31]
  assign sourceD_clock = clock;
  assign sourceD_reset = reset;
  assign sourceD_io_d_ready = io_in_d_ready; // @[Slice.scala 66:11]
  assign sourceD_io_task_valid = c_real_valid_3 | bc_real_valid_3 | sourceD_task_arb_io_out_valid; // @[Slice.scala 489:52]
  assign sourceD_io_task_bits_sourceId = c_real_valid_3 ? c_bits_latch_3_sourceId : _sourceD_io_task_bits_T_sourceId; // @[Slice.scala 490:24]
  assign sourceD_io_task_bits_set = c_real_valid_3 ? c_bits_latch_3_set : _sourceD_io_task_bits_T_set; // @[Slice.scala 490:24]
  assign sourceD_io_task_bits_channel = c_real_valid_3 ? c_bits_latch_3_channel : _sourceD_io_task_bits_T_channel; // @[Slice.scala 490:24]
  assign sourceD_io_task_bits_opcode = c_real_valid_3 ? c_bits_latch_3_opcode : _sourceD_io_task_bits_T_opcode; // @[Slice.scala 490:24]
  assign sourceD_io_task_bits_param = c_real_valid_3 ? c_bits_latch_3_param : _sourceD_io_task_bits_T_param; // @[Slice.scala 490:24]
  assign sourceD_io_task_bits_size = c_real_valid_3 ? c_bits_latch_3_size : _sourceD_io_task_bits_T_size; // @[Slice.scala 490:24]
  assign sourceD_io_task_bits_way = c_real_valid_3 ? c_bits_latch_3_way : _sourceD_io_task_bits_T_way; // @[Slice.scala 490:24]
  assign sourceD_io_task_bits_off = c_real_valid_3 ? c_bits_latch_3_off : _sourceD_io_task_bits_T_off; // @[Slice.scala 490:24]
  assign sourceD_io_task_bits_useBypass = c_real_valid_3 ? c_bits_latch_3_useBypass : _sourceD_io_task_bits_T_useBypass; // @[Slice.scala 490:24]
  assign sourceD_io_task_bits_bufIdx = c_real_valid_3 ? c_bits_latch_3_bufIdx : _sourceD_io_task_bits_T_bufIdx; // @[Slice.scala 490:24]
  assign sourceD_io_task_bits_denied = c_real_valid_3 ? c_bits_latch_3_denied : _sourceD_io_task_bits_T_denied; // @[Slice.scala 490:24]
  assign sourceD_io_task_bits_sinkId = c_real_valid_3 ? c_bits_latch_3_sinkId : _sourceD_io_task_bits_T_sinkId; // @[Slice.scala 490:24]
  assign sourceD_io_task_bits_bypassPut = c_real_valid_3 ? c_bits_latch_3_bypassPut : _sourceD_io_task_bits_T_bypassPut; // @[Slice.scala 490:24]
  assign sourceD_io_task_bits_dirty = c_real_valid_3 ? c_bits_latch_3_dirty : _sourceD_io_task_bits_T_dirty; // @[Slice.scala 490:24]
  assign sourceD_io_bs_raddr_ready = dataStorage_io_sourceD_raddr_ready; // @[Slice.scala 110:32]
  assign sourceD_io_bs_rdata_data = dataStorage_io_sourceD_rdata_data; // @[Slice.scala 109:23]
  assign sourceD_io_bypass_read_ready = refillBuffer_io_rready; // @[Slice.scala 78:21]
  assign sourceD_io_bypass_read_buffer_data_data = refillBuffer_io_rbuffer_data_data; // @[Slice.scala 78:21]
  assign sourceD_io_bs_waddr_ready = dataStorage_io_sourceD_waddr_ready; // @[Slice.scala 111:32]
  assign sourceD_io_pb_pop_ready = sinkA_io_d_pb_pop_ready; // @[Slice.scala 586:21]
  assign sourceD_io_pb_beat_data = sinkA_io_d_pb_beat_data; // @[Slice.scala 587:22]
  assign sourceD_io_pb_beat_mask = sinkA_io_d_pb_beat_mask; // @[Slice.scala 587:22]
  assign sinkE_io_e_valid = io_in_e_valid; // @[Slice.scala 67:14]
  assign sinkE_io_e_bits_sink = io_in_e_bits_sink; // @[Slice.scala 67:14]
  assign sourceA_clock = clock;
  assign sourceA_reset = reset;
  assign sourceA_io_a_ready = io_out_a_q_io_enq_ready; // @[Decoupled.scala 365:17]
  assign sourceA_io_task_valid = c_real_valid | bc_real_valid | sourceA_task_arb_io_out_valid; // @[Slice.scala 489:52]
  assign sourceA_io_task_bits_tag = c_real_valid ? c_bits_latch_tag : _sourceA_io_task_bits_T_tag; // @[Slice.scala 490:24]
  assign sourceA_io_task_bits_set = c_real_valid ? c_bits_latch_set : _sourceA_io_task_bits_T_set; // @[Slice.scala 490:24]
  assign sourceA_io_task_bits_off = c_real_valid ? c_bits_latch_off : _sourceA_io_task_bits_T_off; // @[Slice.scala 490:24]
  assign sourceA_io_task_bits_opcode = c_real_valid ? c_bits_latch_opcode : _sourceA_io_task_bits_T_opcode; // @[Slice.scala 490:24]
  assign sourceA_io_task_bits_param = c_real_valid ? c_bits_latch_param : _sourceA_io_task_bits_T_param; // @[Slice.scala 490:24]
  assign sourceA_io_task_bits_source = c_real_valid ? c_bits_latch_source : _sourceA_io_task_bits_T_source; // @[Slice.scala 490:24]
  assign sourceA_io_task_bits_bufIdx = c_real_valid ? c_bits_latch_bufIdx : _sourceA_io_task_bits_T_bufIdx; // @[Slice.scala 490:24]
  assign sourceA_io_task_bits_size = c_real_valid ? c_bits_latch_size : _sourceA_io_task_bits_T_size; // @[Slice.scala 490:24]
  assign sourceA_io_task_bits_putData = c_real_valid ? c_bits_latch_putData : _sourceA_io_task_bits_T_putData; // @[Slice.scala 490:24]
  assign sourceA_io_pb_pop_ready = sinkA_io_a_pb_pop_ready; // @[Slice.scala 589:21]
  assign sourceA_io_pb_beat_data = sinkA_io_a_pb_beat_data; // @[Slice.scala 590:22]
  assign sourceA_io_pb_beat_mask = sinkA_io_a_pb_beat_mask; // @[Slice.scala 590:22]
  assign sinkB_io_bvalid = sinkB_io_bq_io_deq_valid; // @[Slice.scala 83:14]
  assign sinkB_io_bopcode = sinkB_io_bq_io_deq_bits_opcode; // @[Slice.scala 83:14]
  assign sinkB_io_bparam = sinkB_io_bq_io_deq_bits_param; // @[Slice.scala 83:14]
  assign sinkB_io_bsize = sinkB_io_bq_io_deq_bits_size; // @[Slice.scala 83:14]
  assign sinkB_io_bsource = sinkB_io_bq_io_deq_bits_source; // @[Slice.scala 83:14]
  assign sinkB_io_baddress = sinkB_io_bq_io_deq_bits_address; // @[Slice.scala 83:14]
  assign sinkB_io_bmask = sinkB_io_bq_io_deq_bits_mask; // @[Slice.scala 83:14]
  assign sinkB_io_bdata = sinkB_io_bq_io_deq_bits_data; // @[Slice.scala 83:14]
  assign sinkB_io_alloc_ready = b_arb_io_in_1_ready; // @[Slice.scala 138:20]
  assign sourceC_clock = clock;
  assign sourceC_reset = reset;
  assign sourceC_io_c_ready = out_c_ready & allowed_1; // @[Arbiter.scala 123:31]
  assign sourceC_io_bs_raddr_ready = dataStorage_io_sourceC_raddr_ready; // @[Slice.scala 113:32]
  assign sourceC_io_bs_rdata_data = dataStorage_io_sourceC_rdata_data; // @[Slice.scala 105:23]
  assign sourceC_io_task_valid = c_real_valid_2 | bc_real_valid_2 | sourceC_task_arb_io_out_valid; // @[Slice.scala 489:52]
  assign sourceC_io_task_bits_opcode = c_real_valid_2 ? c_bits_latch_2_opcode : _sourceC_io_task_bits_T_opcode; // @[Slice.scala 490:24]
  assign sourceC_io_task_bits_tag = c_real_valid_2 ? c_bits_latch_2_tag : _sourceC_io_task_bits_T_tag; // @[Slice.scala 490:24]
  assign sourceC_io_task_bits_set = c_real_valid_2 ? c_bits_latch_2_set : _sourceC_io_task_bits_T_set; // @[Slice.scala 490:24]
  assign sourceC_io_task_bits_source = c_real_valid_2 ? c_bits_latch_2_source : _sourceC_io_task_bits_T_source; // @[Slice.scala 490:24]
  assign sourceC_io_task_bits_way = c_real_valid_2 ? c_bits_latch_2_way : _sourceC_io_task_bits_T_way; // @[Slice.scala 490:24]
  assign sinkD_clock = clock;
  assign sinkD_reset = reset;
  assign sinkD_io_d_valid = sinkD_io_d_q_io_deq_valid; // @[Slice.scala 87:14]
  assign sinkD_io_d_bits_opcode = sinkD_io_d_q_io_deq_bits_opcode; // @[Slice.scala 87:14]
  assign sinkD_io_d_bits_param = sinkD_io_d_q_io_deq_bits_param; // @[Slice.scala 87:14]
  assign sinkD_io_d_bits_size = sinkD_io_d_q_io_deq_bits_size; // @[Slice.scala 87:14]
  assign sinkD_io_d_bits_source = sinkD_io_d_q_io_deq_bits_source; // @[Slice.scala 87:14]
  assign sinkD_io_d_bits_sink = sinkD_io_d_q_io_deq_bits_sink; // @[Slice.scala 87:14]
  assign sinkD_io_d_bits_denied = sinkD_io_d_q_io_deq_bits_denied; // @[Slice.scala 87:14]
  assign sinkD_io_d_bits_data = sinkD_io_d_q_io_deq_bits_data; // @[Slice.scala 87:14]
  assign sinkD_io_bs_waddr_ready = dataStorage_io_sinkD_waddr_ready; // @[Slice.scala 104:30]
  assign sinkD_io_bypass_write_ready = refillBuffer_io_wready; // @[Slice.scala 79:21]
  assign sinkD_io_bypass_write_id = refillBuffer_io_wid; // @[Slice.scala 79:21]
  assign sinkD_io_way = _sinkD_status_T_324 | _sinkD_status_T_310; // @[Mux.scala 27:73]
  assign sinkD_io_set = _sinkD_status_T_417 | _sinkD_status_T_403; // @[Mux.scala 27:73]
  assign sinkD_io_inner_grant = _sinkD_status_T & abc_mshr_0_io_status_bits_will_grant_data | _sinkD_status_T_1 &
    abc_mshr_1_io_status_bits_will_grant_data | _sinkD_status_T_2 & abc_mshr_2_io_status_bits_will_grant_data |
    _sinkD_status_T_3 & abc_mshr_3_io_status_bits_will_grant_data | _sinkD_status_T_4 &
    abc_mshr_4_io_status_bits_will_grant_data | _sinkD_status_T_5 & abc_mshr_5_io_status_bits_will_grant_data |
    _sinkD_status_T_6 & abc_mshr_6_io_status_bits_will_grant_data | _sinkD_status_T_7 &
    abc_mshr_7_io_status_bits_will_grant_data | _sinkD_status_T_8 & abc_mshr_8_io_status_bits_will_grant_data |
    _sinkD_status_T_9 & abc_mshr_9_io_status_bits_will_grant_data | _sinkD_status_T_10 &
    abc_mshr_10_io_status_bits_will_grant_data | _sinkD_status_T_11 & abc_mshr_11_io_status_bits_will_grant_data |
    _sinkD_status_T_12 & abc_mshr_12_io_status_bits_will_grant_data | _sinkD_status_T_13 &
    abc_mshr_13_io_status_bits_will_grant_data | _sinkD_status_T_14 & bc_mshr_io_status_bits_will_grant_data |
    _sinkD_status_T_124; // @[Mux.scala 27:73]
  assign sinkD_io_save_data_in_bs = _sinkD_status_T & abc_mshr_0_io_status_bits_will_save_data | _sinkD_status_T_1 &
    abc_mshr_1_io_status_bits_will_save_data | _sinkD_status_T_2 & abc_mshr_2_io_status_bits_will_save_data |
    _sinkD_status_T_3 & abc_mshr_3_io_status_bits_will_save_data | _sinkD_status_T_4 &
    abc_mshr_4_io_status_bits_will_save_data | _sinkD_status_T_5 & abc_mshr_5_io_status_bits_will_save_data |
    _sinkD_status_T_6 & abc_mshr_6_io_status_bits_will_save_data | _sinkD_status_T_7 &
    abc_mshr_7_io_status_bits_will_save_data | _sinkD_status_T_8 & abc_mshr_8_io_status_bits_will_save_data |
    _sinkD_status_T_9 & abc_mshr_9_io_status_bits_will_save_data | _sinkD_status_T_10 &
    abc_mshr_10_io_status_bits_will_save_data | _sinkD_status_T_11 & abc_mshr_11_io_status_bits_will_save_data |
    _sinkD_status_T_12 & abc_mshr_12_io_status_bits_will_save_data | _sinkD_status_T_13 &
    abc_mshr_13_io_status_bits_will_save_data | _sinkD_status_T_14 & bc_mshr_io_status_bits_will_save_data |
    _sinkD_status_T_93; // @[Mux.scala 27:73]
  assign sinkD_io_sourceD_rhazard_valid = sourceD_io_sourceD_rhazard_valid; // @[Slice.scala 584:29]
  assign sinkD_io_sourceD_rhazard_bits_way = sourceD_io_sourceD_rhazard_bits_way; // @[Slice.scala 584:29]
  assign sinkD_io_sourceD_rhazard_bits_set = sourceD_io_sourceD_rhazard_bits_set; // @[Slice.scala 584:29]
  assign sourceE_io_e_ready = io_out_e_q_io_enq_ready; // @[Decoupled.scala 365:17]
  assign sourceE_io_task_valid = c_real_valid_4 | bc_real_valid_4 | sourceE_task_arb_io_out_valid; // @[Slice.scala 489:52]
  assign sourceE_io_task_bits_sink = c_real_valid_4 ? c_bits_latch_4_sink : _sourceE_io_task_bits_T_sink; // @[Slice.scala 490:24]
  assign refillBuffer_clock = clock;
  assign refillBuffer_reset = reset;
  assign refillBuffer_io_rvalid = sourceD_io_bypass_read_valid; // @[Slice.scala 78:21]
  assign refillBuffer_io_rbeat = sourceD_io_bypass_read_beat; // @[Slice.scala 78:21]
  assign refillBuffer_io_rid = sourceD_io_bypass_read_id; // @[Slice.scala 78:21]
  assign refillBuffer_io_rlast = sourceD_io_bypass_read_last; // @[Slice.scala 78:21]
  assign refillBuffer_io_wvalid = sinkD_io_bypass_write_valid; // @[Slice.scala 79:21]
  assign refillBuffer_io_wbeat = sinkD_io_bypass_write_beat; // @[Slice.scala 79:21]
  assign refillBuffer_io_wdata_data = sinkD_io_bypass_write_data_data; // @[Slice.scala 79:21]
  assign io_out_a_q_clock = clock;
  assign io_out_a_q_reset = reset;
  assign io_out_a_q_io_enq_valid = sourceA_io_a_valid; // @[Decoupled.scala 363:22]
  assign io_out_a_q_io_enq_bits_opcode = sourceA_io_a_bits_opcode; // @[Decoupled.scala 364:21]
  assign io_out_a_q_io_enq_bits_param = sourceA_io_a_bits_param; // @[Decoupled.scala 364:21]
  assign io_out_a_q_io_enq_bits_size = sourceA_io_a_bits_size; // @[Decoupled.scala 364:21]
  assign io_out_a_q_io_enq_bits_source = sourceA_io_a_bits_source; // @[Decoupled.scala 364:21]
  assign io_out_a_q_io_enq_bits_address = sourceA_io_a_bits_address; // @[Decoupled.scala 364:21]
  assign io_out_a_q_io_enq_bits_mask = sourceA_io_a_bits_mask; // @[Decoupled.scala 364:21]
  assign io_out_a_q_io_enq_bits_data = sourceA_io_a_bits_data; // @[Decoupled.scala 364:21]
  assign io_out_a_q_io_deq_ready = io_out_a_ready; // @[Slice.scala 82:12]
  assign sinkB_io_bq_clock = clock;
  assign sinkB_io_bq_reset = reset;
  assign sinkB_io_bq_io_enq_valid = 1'h0; // @[Decoupled.scala 363:22]
  assign sinkB_io_bq_io_enq_bits_opcode = 3'h0; // @[Decoupled.scala 364:21]
  assign sinkB_io_bq_io_enq_bits_param = 2'h0; // @[Decoupled.scala 364:21]
  assign sinkB_io_bq_io_enq_bits_size = 3'h0; // @[Decoupled.scala 364:21]
  assign sinkB_io_bq_io_enq_bits_source = 4'h0; // @[Decoupled.scala 364:21]
  assign sinkB_io_bq_io_enq_bits_address = 36'h0; // @[Decoupled.scala 364:21]
  assign sinkB_io_bq_io_enq_bits_mask = 32'h0; // @[Decoupled.scala 364:21]
  assign sinkB_io_bq_io_enq_bits_data = 256'h0; // @[Decoupled.scala 364:21]
  assign sinkB_io_bq_io_deq_ready = sinkB_io_bready; // @[Slice.scala 83:14]
  assign io_out_c_q_clock = clock;
  assign io_out_c_q_reset = reset;
  assign io_out_c_q_io_enq_valid = idle ? _T_12 : _sink_ACancel_earlyValid_T_3; // @[Arbiter.scala 125:29]
  assign io_out_c_q_io_enq_bits_opcode = _T_44 | _T_45; // @[Mux.scala 27:73]
  assign io_out_c_q_io_enq_bits_size = _T_38 | _T_39; // @[Mux.scala 27:73]
  assign io_out_c_q_io_enq_bits_source = _T_35 | _T_36; // @[Mux.scala 27:73]
  assign io_out_c_q_io_enq_bits_address = _T_32 | _T_33; // @[Mux.scala 27:73]
  assign io_out_c_q_io_enq_bits_data = _T_29 | _T_30; // @[Mux.scala 27:73]
  assign io_out_c_q_io_deq_ready = io_out_c_ready; // @[Slice.scala 86:12]
  assign sinkD_io_d_q_clock = clock;
  assign sinkD_io_d_q_reset = reset;
  assign sinkD_io_d_q_io_enq_valid = io_out_d_valid; // @[Decoupled.scala 363:22]
  assign sinkD_io_d_q_io_enq_bits_opcode = io_out_d_bits_opcode; // @[Decoupled.scala 364:21]
  assign sinkD_io_d_q_io_enq_bits_param = io_out_d_bits_param; // @[Decoupled.scala 364:21]
  assign sinkD_io_d_q_io_enq_bits_size = io_out_d_bits_size; // @[Decoupled.scala 364:21]
  assign sinkD_io_d_q_io_enq_bits_source = io_out_d_bits_source; // @[Decoupled.scala 364:21]
  assign sinkD_io_d_q_io_enq_bits_sink = io_out_d_bits_sink; // @[Decoupled.scala 364:21]
  assign sinkD_io_d_q_io_enq_bits_denied = io_out_d_bits_denied; // @[Decoupled.scala 364:21]
  assign sinkD_io_d_q_io_enq_bits_data = io_out_d_bits_data; // @[Decoupled.scala 364:21]
  assign sinkD_io_d_q_io_deq_ready = sinkD_io_d_ready; // @[Slice.scala 87:14]
  assign io_out_e_q_clock = clock;
  assign io_out_e_q_reset = reset;
  assign io_out_e_q_io_enq_valid = sourceE_io_e_valid; // @[Decoupled.scala 363:22]
  assign io_out_e_q_io_enq_bits_sink = sourceE_io_e_bits_sink; // @[Decoupled.scala 364:21]
  assign abc_mshr_0_clock = clock;
  assign abc_mshr_0_reset = reset;
  assign abc_mshr_0_io_id = 4'h0; // @[Slice.scala 166:18]
  assign abc_mshr_0_io_enable = ~(bc_disable | c_disable); // @[Slice.scala 198:25]
  assign abc_mshr_0_io_alloc_valid = mshrAlloc_io_alloc_0_valid; // @[Slice.scala 167:21]
  assign abc_mshr_0_io_alloc_bits_channel = mshrAlloc_io_alloc_0_bits_channel; // @[Slice.scala 167:21]
  assign abc_mshr_0_io_alloc_bits_opcode = mshrAlloc_io_alloc_0_bits_opcode; // @[Slice.scala 167:21]
  assign abc_mshr_0_io_alloc_bits_param = mshrAlloc_io_alloc_0_bits_param; // @[Slice.scala 167:21]
  assign abc_mshr_0_io_alloc_bits_size = mshrAlloc_io_alloc_0_bits_size; // @[Slice.scala 167:21]
  assign abc_mshr_0_io_alloc_bits_source = mshrAlloc_io_alloc_0_bits_source; // @[Slice.scala 167:21]
  assign abc_mshr_0_io_alloc_bits_set = mshrAlloc_io_alloc_0_bits_set; // @[Slice.scala 167:21]
  assign abc_mshr_0_io_alloc_bits_tag = mshrAlloc_io_alloc_0_bits_tag; // @[Slice.scala 167:21]
  assign abc_mshr_0_io_alloc_bits_off = mshrAlloc_io_alloc_0_bits_off; // @[Slice.scala 167:21]
  assign abc_mshr_0_io_alloc_bits_mask = mshrAlloc_io_alloc_0_bits_mask; // @[Slice.scala 167:21]
  assign abc_mshr_0_io_alloc_bits_bufIdx = mshrAlloc_io_alloc_0_bits_bufIdx; // @[Slice.scala 167:21]
  assign abc_mshr_0_io_alloc_bits_preferCache = mshrAlloc_io_alloc_0_bits_preferCache; // @[Slice.scala 167:21]
  assign abc_mshr_0_io_alloc_bits_dirty = mshrAlloc_io_alloc_0_bits_dirty; // @[Slice.scala 167:21]
  assign abc_mshr_0_io_alloc_bits_fromProbeHelper = mshrAlloc_io_alloc_0_bits_fromProbeHelper; // @[Slice.scala 167:21]
  assign abc_mshr_0_io_alloc_bits_fromCmoHelper = mshrAlloc_io_alloc_0_bits_fromCmoHelper; // @[Slice.scala 167:21]
  assign abc_mshr_0_io_alloc_bits_needProbeAckData = mshrAlloc_io_alloc_0_bits_needProbeAckData; // @[Slice.scala 167:21]
  assign abc_mshr_0_io_resps_sink_c_valid = sinkC_io_resp_valid & sinkC_io_resp_bits_set ==
    abc_mshr_0_io_status_bits_set; // @[Slice.scala 527:57]
  assign abc_mshr_0_io_resps_sink_c_bits_hasData = sinkC_io_resp_bits_hasData; // @[Slice.scala 531:33]
  assign abc_mshr_0_io_resps_sink_c_bits_param = sinkC_io_resp_bits_param; // @[Slice.scala 531:33]
  assign abc_mshr_0_io_resps_sink_c_bits_source = sinkC_io_resp_bits_source; // @[Slice.scala 531:33]
  assign abc_mshr_0_io_resps_sink_c_bits_last = sinkC_io_resp_bits_last; // @[Slice.scala 531:33]
  assign abc_mshr_0_io_resps_sink_c_bits_bufIdx = sinkC_io_resp_bits_bufIdx; // @[Slice.scala 531:33]
  assign abc_mshr_0_io_resps_sink_d_valid = sinkD_io_resp_valid & sinkD_io_resp_bits_source == 4'h0; // @[Slice.scala 528:57]
  assign abc_mshr_0_io_resps_sink_d_bits_opcode = sinkD_io_resp_bits_opcode; // @[Slice.scala 532:33]
  assign abc_mshr_0_io_resps_sink_d_bits_param = sinkD_io_resp_bits_param; // @[Slice.scala 532:33]
  assign abc_mshr_0_io_resps_sink_d_bits_sink = sinkD_io_resp_bits_sink; // @[Slice.scala 532:33]
  assign abc_mshr_0_io_resps_sink_d_bits_last = sinkD_io_resp_bits_last; // @[Slice.scala 532:33]
  assign abc_mshr_0_io_resps_sink_d_bits_denied = sinkD_io_resp_bits_denied; // @[Slice.scala 532:33]
  assign abc_mshr_0_io_resps_sink_d_bits_bufIdx = sinkD_io_resp_bits_bufIdx; // @[Slice.scala 532:33]
  assign abc_mshr_0_io_resps_sink_e_valid = sinkE_io_resp_valid & sinkE_io_resp_bits_sink == 4'h0; // @[Slice.scala 529:57]
  assign abc_mshr_0_io_resps_source_d_valid = sourceD_io_resp_valid & sourceD_io_resp_bits_sink == 4'h0; // @[Slice.scala 530:61]
  assign abc_mshr_0_io_nestedwb_set = c_mshr_io_status_valid ? c_mshr_io_status_bits_set : bc_mshr_io_status_bits_set; // @[Slice.scala 258:22]
  assign abc_mshr_0_io_nestedwb_tag = c_mshr_io_status_valid ? c_mshr_io_status_bits_tag : bc_mshr_io_status_bits_tag; // @[Slice.scala 259:22]
  assign abc_mshr_0_io_nestedwb_btoN = _nestedWb_btoN_T_2 & _nestedWb_btoN_T_3; // @[Slice.scala 280:38]
  assign abc_mshr_0_io_nestedwb_btoB = _nestedWb_btoN_T_2 & _nestedWb_btoB_T_3; // @[Slice.scala 283:38]
  assign abc_mshr_0_io_nestedwb_bclr_dirty = _nestedWb_btoN_T_2 & _nestedWb_bclr_dirty_T_4; // @[Slice.scala 286:38]
  assign abc_mshr_0_io_nestedwb_bset_dirty = _nestedWb_btoN_T_2 & bc_mshr_io_tasks_dir_write_bits_data_dirty; // @[Slice.scala 289:38]
  assign abc_mshr_0_io_nestedwb_c_set_dirty = _nestedWb_c_set_dirty_T & c_mshr_io_tasks_dir_write_bits_data_dirty; // @[Slice.scala 292:37]
  assign abc_mshr_0_io_nestedwb_c_set_hit = c_mshr_io_status_valid & c_mshr_io_tasks_tag_write_valid &
    _nestedWb_c_set_hit_T_1; // @[Slice.scala 304:50]
  assign abc_mshr_0_io_nestedwb_clients_0_isToN = c_mshr_io_status_valid ? _nestedWb_clients_0_isToN_T_1 :
    _nestedWb_clients_0_isToN_T_3; // @[Slice.scala 314:25]
  assign abc_mshr_0_io_nestedwb_clients_1_isToN = c_mshr_io_status_valid ? _nestedWb_clients_1_isToN_T_1 :
    _nestedWb_clients_1_isToN_T_3; // @[Slice.scala 314:25]
  assign abc_mshr_0_io_tasks_sink_a_ready = 1'h0; // @[Slice.scala 472:13]
  assign abc_mshr_0_io_tasks_source_bready = sourceB_task_arb_io_in_0_ready; // @[Slice.scala 472:13]
  assign abc_mshr_0_io_tasks_sink_c_ready = sinkC_task_arb_io_in_0_ready; // @[Slice.scala 472:13]
  assign abc_mshr_0_io_tasks_source_d_ready = sourceD_task_arb_io_in_0_ready; // @[Slice.scala 472:13]
  assign abc_mshr_0_io_tasks_source_a_ready = sourceA_task_arb_io_in_0_ready; // @[Slice.scala 472:13]
  assign abc_mshr_0_io_tasks_source_c_ready = sourceC_task_arb_io_in_0_ready; // @[Slice.scala 472:13]
  assign abc_mshr_0_io_tasks_source_e_ready = sourceE_task_arb_io_in_0_ready; // @[Slice.scala 472:13]
  assign abc_mshr_0_io_tasks_dir_write_ready = arbiter_io_in_0_ready; // @[Slice.scala 406:60]
  assign abc_mshr_0_io_tasks_tag_write_ready = tagWrite_task_arb_io_in_0_ready; // @[Slice.scala 472:13]
  assign abc_mshr_0_io_tasks_client_dir_write_ready = arbiter_1_io_in_0_ready; // @[Slice.scala 406:60]
  assign abc_mshr_0_io_tasks_client_tag_write_ready = arbiter_2_io_in_0_ready; // @[Slice.scala 472:13]
  assign abc_mshr_0_io_dirResult_valid = ms_0_io_dirResult_valid_REG; // @[Slice.scala 556:31]
  assign abc_mshr_0_io_dirResult_bits_self_dirty = directory_io_result_bits_self_dirty; // @[Slice.scala 555:30]
  assign abc_mshr_0_io_dirResult_bits_self_state = directory_io_result_bits_self_state; // @[Slice.scala 555:30]
  assign abc_mshr_0_io_dirResult_bits_self_clientStates_0 = directory_io_result_bits_self_clientStates_0; // @[Slice.scala 555:30]
  assign abc_mshr_0_io_dirResult_bits_self_clientStates_1 = directory_io_result_bits_self_clientStates_1; // @[Slice.scala 555:30]
  assign abc_mshr_0_io_dirResult_bits_self_hit = directory_io_result_bits_self_hit; // @[Slice.scala 555:30]
  assign abc_mshr_0_io_dirResult_bits_self_way = directory_io_result_bits_self_way; // @[Slice.scala 555:30]
  assign abc_mshr_0_io_dirResult_bits_self_tag = directory_io_result_bits_self_tag; // @[Slice.scala 555:30]
  assign abc_mshr_0_io_dirResult_bits_clients_states_0_state = directory_io_result_bits_clients_states_0_state; // @[Slice.scala 555:30]
  assign abc_mshr_0_io_dirResult_bits_clients_states_0_hit = directory_io_result_bits_clients_states_0_hit; // @[Slice.scala 555:30]
  assign abc_mshr_0_io_dirResult_bits_clients_states_1_state = directory_io_result_bits_clients_states_1_state; // @[Slice.scala 555:30]
  assign abc_mshr_0_io_dirResult_bits_clients_states_1_hit = directory_io_result_bits_clients_states_1_hit; // @[Slice.scala 555:30]
  assign abc_mshr_0_io_dirResult_bits_clients_tag = directory_io_result_bits_clients_tag; // @[Slice.scala 555:30]
  assign abc_mshr_0_io_dirResult_bits_clients_way = directory_io_result_bits_clients_way; // @[Slice.scala 555:30]
  assign abc_mshr_0_io_c_status_set = c_mshr_io_status_bits_set; // @[Slice.scala 209:28]
  assign abc_mshr_0_io_c_status_tag = c_mshr_io_status_bits_tag; // @[Slice.scala 210:28]
  assign abc_mshr_0_io_c_status_way = c_mshr_io_status_bits_way; // @[Slice.scala 211:28]
  assign abc_mshr_0_io_c_status_nestedReleaseData = c_mshr_io_status_valid & c_mshr_io_is_nestedReleaseData; // @[Slice.scala 213:32]
  assign abc_mshr_0_io_bstatus_set = bc_mshr_io_status_bits_set; // @[Slice.scala 214:28]
  assign abc_mshr_0_io_bstatus_tag = bc_mshr_io_status_bits_tag; // @[Slice.scala 215:28]
  assign abc_mshr_0_io_bstatus_way = bc_mshr_io_status_bits_way; // @[Slice.scala 216:28]
  assign abc_mshr_0_io_bstatus_nestedProbeAckData = bc_mshr_io_status_valid & bc_mshr_io_is_nestedProbeAckData; // @[Slice.scala 218:33]
  assign abc_mshr_0_io_bstatus_probeHelperFinish = bc_mshr_io_status_valid & bc_mshr_io_probeHelperFinish; // @[Slice.scala 220:33]
  assign abc_mshr_0_io_releaseThrough = 1'h0; // @[Slice.scala 221:30]
  assign abc_mshr_0_io_probeAckDataThrough = 1'h0; // @[Slice.scala 222:35]
  assign abc_mshr_1_clock = clock;
  assign abc_mshr_1_reset = reset;
  assign abc_mshr_1_io_id = 4'h1; // @[Slice.scala 166:18]
  assign abc_mshr_1_io_enable = ~(bc_disable_1 | c_disable_1); // @[Slice.scala 198:25]
  assign abc_mshr_1_io_alloc_valid = mshrAlloc_io_alloc_1_valid; // @[Slice.scala 167:21]
  assign abc_mshr_1_io_alloc_bits_channel = mshrAlloc_io_alloc_1_bits_channel; // @[Slice.scala 167:21]
  assign abc_mshr_1_io_alloc_bits_opcode = mshrAlloc_io_alloc_1_bits_opcode; // @[Slice.scala 167:21]
  assign abc_mshr_1_io_alloc_bits_param = mshrAlloc_io_alloc_1_bits_param; // @[Slice.scala 167:21]
  assign abc_mshr_1_io_alloc_bits_size = mshrAlloc_io_alloc_1_bits_size; // @[Slice.scala 167:21]
  assign abc_mshr_1_io_alloc_bits_source = mshrAlloc_io_alloc_1_bits_source; // @[Slice.scala 167:21]
  assign abc_mshr_1_io_alloc_bits_set = mshrAlloc_io_alloc_1_bits_set; // @[Slice.scala 167:21]
  assign abc_mshr_1_io_alloc_bits_tag = mshrAlloc_io_alloc_1_bits_tag; // @[Slice.scala 167:21]
  assign abc_mshr_1_io_alloc_bits_off = mshrAlloc_io_alloc_1_bits_off; // @[Slice.scala 167:21]
  assign abc_mshr_1_io_alloc_bits_mask = mshrAlloc_io_alloc_1_bits_mask; // @[Slice.scala 167:21]
  assign abc_mshr_1_io_alloc_bits_bufIdx = mshrAlloc_io_alloc_1_bits_bufIdx; // @[Slice.scala 167:21]
  assign abc_mshr_1_io_alloc_bits_preferCache = mshrAlloc_io_alloc_1_bits_preferCache; // @[Slice.scala 167:21]
  assign abc_mshr_1_io_alloc_bits_dirty = mshrAlloc_io_alloc_1_bits_dirty; // @[Slice.scala 167:21]
  assign abc_mshr_1_io_alloc_bits_fromProbeHelper = mshrAlloc_io_alloc_1_bits_fromProbeHelper; // @[Slice.scala 167:21]
  assign abc_mshr_1_io_alloc_bits_fromCmoHelper = mshrAlloc_io_alloc_1_bits_fromCmoHelper; // @[Slice.scala 167:21]
  assign abc_mshr_1_io_alloc_bits_needProbeAckData = mshrAlloc_io_alloc_1_bits_needProbeAckData; // @[Slice.scala 167:21]
  assign abc_mshr_1_io_resps_sink_c_valid = sinkC_io_resp_valid & sinkC_io_resp_bits_set ==
    abc_mshr_1_io_status_bits_set; // @[Slice.scala 527:57]
  assign abc_mshr_1_io_resps_sink_c_bits_hasData = sinkC_io_resp_bits_hasData; // @[Slice.scala 531:33]
  assign abc_mshr_1_io_resps_sink_c_bits_param = sinkC_io_resp_bits_param; // @[Slice.scala 531:33]
  assign abc_mshr_1_io_resps_sink_c_bits_source = sinkC_io_resp_bits_source; // @[Slice.scala 531:33]
  assign abc_mshr_1_io_resps_sink_c_bits_last = sinkC_io_resp_bits_last; // @[Slice.scala 531:33]
  assign abc_mshr_1_io_resps_sink_c_bits_bufIdx = sinkC_io_resp_bits_bufIdx; // @[Slice.scala 531:33]
  assign abc_mshr_1_io_resps_sink_d_valid = sinkD_io_resp_valid & sinkD_io_resp_bits_source == 4'h1; // @[Slice.scala 528:57]
  assign abc_mshr_1_io_resps_sink_d_bits_opcode = sinkD_io_resp_bits_opcode; // @[Slice.scala 532:33]
  assign abc_mshr_1_io_resps_sink_d_bits_param = sinkD_io_resp_bits_param; // @[Slice.scala 532:33]
  assign abc_mshr_1_io_resps_sink_d_bits_sink = sinkD_io_resp_bits_sink; // @[Slice.scala 532:33]
  assign abc_mshr_1_io_resps_sink_d_bits_last = sinkD_io_resp_bits_last; // @[Slice.scala 532:33]
  assign abc_mshr_1_io_resps_sink_d_bits_denied = sinkD_io_resp_bits_denied; // @[Slice.scala 532:33]
  assign abc_mshr_1_io_resps_sink_d_bits_bufIdx = sinkD_io_resp_bits_bufIdx; // @[Slice.scala 532:33]
  assign abc_mshr_1_io_resps_sink_e_valid = sinkE_io_resp_valid & sinkE_io_resp_bits_sink == 4'h1; // @[Slice.scala 529:57]
  assign abc_mshr_1_io_resps_source_d_valid = sourceD_io_resp_valid & sourceD_io_resp_bits_sink == 4'h1; // @[Slice.scala 530:61]
  assign abc_mshr_1_io_nestedwb_set = c_mshr_io_status_valid ? c_mshr_io_status_bits_set : bc_mshr_io_status_bits_set; // @[Slice.scala 258:22]
  assign abc_mshr_1_io_nestedwb_tag = c_mshr_io_status_valid ? c_mshr_io_status_bits_tag : bc_mshr_io_status_bits_tag; // @[Slice.scala 259:22]
  assign abc_mshr_1_io_nestedwb_btoN = _nestedWb_btoN_T_2 & _nestedWb_btoN_T_3; // @[Slice.scala 280:38]
  assign abc_mshr_1_io_nestedwb_btoB = _nestedWb_btoN_T_2 & _nestedWb_btoB_T_3; // @[Slice.scala 283:38]
  assign abc_mshr_1_io_nestedwb_bclr_dirty = _nestedWb_btoN_T_2 & _nestedWb_bclr_dirty_T_4; // @[Slice.scala 286:38]
  assign abc_mshr_1_io_nestedwb_bset_dirty = _nestedWb_btoN_T_2 & bc_mshr_io_tasks_dir_write_bits_data_dirty; // @[Slice.scala 289:38]
  assign abc_mshr_1_io_nestedwb_c_set_dirty = _nestedWb_c_set_dirty_T & c_mshr_io_tasks_dir_write_bits_data_dirty; // @[Slice.scala 292:37]
  assign abc_mshr_1_io_nestedwb_c_set_hit = c_mshr_io_status_valid & c_mshr_io_tasks_tag_write_valid &
    _nestedWb_c_set_hit_T_3; // @[Slice.scala 304:50]
  assign abc_mshr_1_io_nestedwb_clients_0_isToN = c_mshr_io_status_valid ? _nestedWb_clients_0_isToN_T_1 :
    _nestedWb_clients_0_isToN_T_3; // @[Slice.scala 314:25]
  assign abc_mshr_1_io_nestedwb_clients_1_isToN = c_mshr_io_status_valid ? _nestedWb_clients_1_isToN_T_1 :
    _nestedWb_clients_1_isToN_T_3; // @[Slice.scala 314:25]
  assign abc_mshr_1_io_tasks_sink_a_ready = 1'h0; // @[Slice.scala 472:13]
  assign abc_mshr_1_io_tasks_source_bready = sourceB_task_arb_io_in_1_ready; // @[Slice.scala 472:13]
  assign abc_mshr_1_io_tasks_sink_c_ready = sinkC_task_arb_io_in_1_ready; // @[Slice.scala 472:13]
  assign abc_mshr_1_io_tasks_source_d_ready = sourceD_task_arb_io_in_1_ready; // @[Slice.scala 472:13]
  assign abc_mshr_1_io_tasks_source_a_ready = sourceA_task_arb_io_in_1_ready; // @[Slice.scala 472:13]
  assign abc_mshr_1_io_tasks_source_c_ready = sourceC_task_arb_io_in_1_ready; // @[Slice.scala 472:13]
  assign abc_mshr_1_io_tasks_source_e_ready = sourceE_task_arb_io_in_1_ready; // @[Slice.scala 472:13]
  assign abc_mshr_1_io_tasks_dir_write_ready = arbiter_io_in_1_ready; // @[Slice.scala 406:60]
  assign abc_mshr_1_io_tasks_tag_write_ready = tagWrite_task_arb_io_in_1_ready; // @[Slice.scala 472:13]
  assign abc_mshr_1_io_tasks_client_dir_write_ready = arbiter_1_io_in_1_ready; // @[Slice.scala 406:60]
  assign abc_mshr_1_io_tasks_client_tag_write_ready = arbiter_2_io_in_1_ready; // @[Slice.scala 472:13]
  assign abc_mshr_1_io_dirResult_valid = ms_1_io_dirResult_valid_REG; // @[Slice.scala 556:31]
  assign abc_mshr_1_io_dirResult_bits_self_dirty = directory_io_result_bits_self_dirty; // @[Slice.scala 555:30]
  assign abc_mshr_1_io_dirResult_bits_self_state = directory_io_result_bits_self_state; // @[Slice.scala 555:30]
  assign abc_mshr_1_io_dirResult_bits_self_clientStates_0 = directory_io_result_bits_self_clientStates_0; // @[Slice.scala 555:30]
  assign abc_mshr_1_io_dirResult_bits_self_clientStates_1 = directory_io_result_bits_self_clientStates_1; // @[Slice.scala 555:30]
  assign abc_mshr_1_io_dirResult_bits_self_hit = directory_io_result_bits_self_hit; // @[Slice.scala 555:30]
  assign abc_mshr_1_io_dirResult_bits_self_way = directory_io_result_bits_self_way; // @[Slice.scala 555:30]
  assign abc_mshr_1_io_dirResult_bits_self_tag = directory_io_result_bits_self_tag; // @[Slice.scala 555:30]
  assign abc_mshr_1_io_dirResult_bits_clients_states_0_state = directory_io_result_bits_clients_states_0_state; // @[Slice.scala 555:30]
  assign abc_mshr_1_io_dirResult_bits_clients_states_0_hit = directory_io_result_bits_clients_states_0_hit; // @[Slice.scala 555:30]
  assign abc_mshr_1_io_dirResult_bits_clients_states_1_state = directory_io_result_bits_clients_states_1_state; // @[Slice.scala 555:30]
  assign abc_mshr_1_io_dirResult_bits_clients_states_1_hit = directory_io_result_bits_clients_states_1_hit; // @[Slice.scala 555:30]
  assign abc_mshr_1_io_dirResult_bits_clients_tag = directory_io_result_bits_clients_tag; // @[Slice.scala 555:30]
  assign abc_mshr_1_io_dirResult_bits_clients_way = directory_io_result_bits_clients_way; // @[Slice.scala 555:30]
  assign abc_mshr_1_io_c_status_set = c_mshr_io_status_bits_set; // @[Slice.scala 209:28]
  assign abc_mshr_1_io_c_status_tag = c_mshr_io_status_bits_tag; // @[Slice.scala 210:28]
  assign abc_mshr_1_io_c_status_way = c_mshr_io_status_bits_way; // @[Slice.scala 211:28]
  assign abc_mshr_1_io_c_status_nestedReleaseData = c_mshr_io_status_valid & c_mshr_io_is_nestedReleaseData; // @[Slice.scala 213:32]
  assign abc_mshr_1_io_bstatus_set = bc_mshr_io_status_bits_set; // @[Slice.scala 214:28]
  assign abc_mshr_1_io_bstatus_tag = bc_mshr_io_status_bits_tag; // @[Slice.scala 215:28]
  assign abc_mshr_1_io_bstatus_way = bc_mshr_io_status_bits_way; // @[Slice.scala 216:28]
  assign abc_mshr_1_io_bstatus_nestedProbeAckData = bc_mshr_io_status_valid & bc_mshr_io_is_nestedProbeAckData; // @[Slice.scala 218:33]
  assign abc_mshr_1_io_bstatus_probeHelperFinish = bc_mshr_io_status_valid & bc_mshr_io_probeHelperFinish; // @[Slice.scala 220:33]
  assign abc_mshr_1_io_releaseThrough = 1'h0; // @[Slice.scala 221:30]
  assign abc_mshr_1_io_probeAckDataThrough = 1'h0; // @[Slice.scala 222:35]
  assign abc_mshr_2_clock = clock;
  assign abc_mshr_2_reset = reset;
  assign abc_mshr_2_io_id = 4'h2; // @[Slice.scala 166:18]
  assign abc_mshr_2_io_enable = ~(bc_disable_2 | c_disable_2); // @[Slice.scala 198:25]
  assign abc_mshr_2_io_alloc_valid = mshrAlloc_io_alloc_2_valid; // @[Slice.scala 167:21]
  assign abc_mshr_2_io_alloc_bits_channel = mshrAlloc_io_alloc_2_bits_channel; // @[Slice.scala 167:21]
  assign abc_mshr_2_io_alloc_bits_opcode = mshrAlloc_io_alloc_2_bits_opcode; // @[Slice.scala 167:21]
  assign abc_mshr_2_io_alloc_bits_param = mshrAlloc_io_alloc_2_bits_param; // @[Slice.scala 167:21]
  assign abc_mshr_2_io_alloc_bits_size = mshrAlloc_io_alloc_2_bits_size; // @[Slice.scala 167:21]
  assign abc_mshr_2_io_alloc_bits_source = mshrAlloc_io_alloc_2_bits_source; // @[Slice.scala 167:21]
  assign abc_mshr_2_io_alloc_bits_set = mshrAlloc_io_alloc_2_bits_set; // @[Slice.scala 167:21]
  assign abc_mshr_2_io_alloc_bits_tag = mshrAlloc_io_alloc_2_bits_tag; // @[Slice.scala 167:21]
  assign abc_mshr_2_io_alloc_bits_off = mshrAlloc_io_alloc_2_bits_off; // @[Slice.scala 167:21]
  assign abc_mshr_2_io_alloc_bits_mask = mshrAlloc_io_alloc_2_bits_mask; // @[Slice.scala 167:21]
  assign abc_mshr_2_io_alloc_bits_bufIdx = mshrAlloc_io_alloc_2_bits_bufIdx; // @[Slice.scala 167:21]
  assign abc_mshr_2_io_alloc_bits_preferCache = mshrAlloc_io_alloc_2_bits_preferCache; // @[Slice.scala 167:21]
  assign abc_mshr_2_io_alloc_bits_dirty = mshrAlloc_io_alloc_2_bits_dirty; // @[Slice.scala 167:21]
  assign abc_mshr_2_io_alloc_bits_fromProbeHelper = mshrAlloc_io_alloc_2_bits_fromProbeHelper; // @[Slice.scala 167:21]
  assign abc_mshr_2_io_alloc_bits_fromCmoHelper = mshrAlloc_io_alloc_2_bits_fromCmoHelper; // @[Slice.scala 167:21]
  assign abc_mshr_2_io_alloc_bits_needProbeAckData = mshrAlloc_io_alloc_2_bits_needProbeAckData; // @[Slice.scala 167:21]
  assign abc_mshr_2_io_resps_sink_c_valid = sinkC_io_resp_valid & sinkC_io_resp_bits_set ==
    abc_mshr_2_io_status_bits_set; // @[Slice.scala 527:57]
  assign abc_mshr_2_io_resps_sink_c_bits_hasData = sinkC_io_resp_bits_hasData; // @[Slice.scala 531:33]
  assign abc_mshr_2_io_resps_sink_c_bits_param = sinkC_io_resp_bits_param; // @[Slice.scala 531:33]
  assign abc_mshr_2_io_resps_sink_c_bits_source = sinkC_io_resp_bits_source; // @[Slice.scala 531:33]
  assign abc_mshr_2_io_resps_sink_c_bits_last = sinkC_io_resp_bits_last; // @[Slice.scala 531:33]
  assign abc_mshr_2_io_resps_sink_c_bits_bufIdx = sinkC_io_resp_bits_bufIdx; // @[Slice.scala 531:33]
  assign abc_mshr_2_io_resps_sink_d_valid = sinkD_io_resp_valid & sinkD_io_resp_bits_source == 4'h2; // @[Slice.scala 528:57]
  assign abc_mshr_2_io_resps_sink_d_bits_opcode = sinkD_io_resp_bits_opcode; // @[Slice.scala 532:33]
  assign abc_mshr_2_io_resps_sink_d_bits_param = sinkD_io_resp_bits_param; // @[Slice.scala 532:33]
  assign abc_mshr_2_io_resps_sink_d_bits_sink = sinkD_io_resp_bits_sink; // @[Slice.scala 532:33]
  assign abc_mshr_2_io_resps_sink_d_bits_last = sinkD_io_resp_bits_last; // @[Slice.scala 532:33]
  assign abc_mshr_2_io_resps_sink_d_bits_denied = sinkD_io_resp_bits_denied; // @[Slice.scala 532:33]
  assign abc_mshr_2_io_resps_sink_d_bits_bufIdx = sinkD_io_resp_bits_bufIdx; // @[Slice.scala 532:33]
  assign abc_mshr_2_io_resps_sink_e_valid = sinkE_io_resp_valid & sinkE_io_resp_bits_sink == 4'h2; // @[Slice.scala 529:57]
  assign abc_mshr_2_io_resps_source_d_valid = sourceD_io_resp_valid & sourceD_io_resp_bits_sink == 4'h2; // @[Slice.scala 530:61]
  assign abc_mshr_2_io_nestedwb_set = c_mshr_io_status_valid ? c_mshr_io_status_bits_set : bc_mshr_io_status_bits_set; // @[Slice.scala 258:22]
  assign abc_mshr_2_io_nestedwb_tag = c_mshr_io_status_valid ? c_mshr_io_status_bits_tag : bc_mshr_io_status_bits_tag; // @[Slice.scala 259:22]
  assign abc_mshr_2_io_nestedwb_btoN = _nestedWb_btoN_T_2 & _nestedWb_btoN_T_3; // @[Slice.scala 280:38]
  assign abc_mshr_2_io_nestedwb_btoB = _nestedWb_btoN_T_2 & _nestedWb_btoB_T_3; // @[Slice.scala 283:38]
  assign abc_mshr_2_io_nestedwb_bclr_dirty = _nestedWb_btoN_T_2 & _nestedWb_bclr_dirty_T_4; // @[Slice.scala 286:38]
  assign abc_mshr_2_io_nestedwb_bset_dirty = _nestedWb_btoN_T_2 & bc_mshr_io_tasks_dir_write_bits_data_dirty; // @[Slice.scala 289:38]
  assign abc_mshr_2_io_nestedwb_c_set_dirty = _nestedWb_c_set_dirty_T & c_mshr_io_tasks_dir_write_bits_data_dirty; // @[Slice.scala 292:37]
  assign abc_mshr_2_io_nestedwb_c_set_hit = c_mshr_io_status_valid & c_mshr_io_tasks_tag_write_valid &
    _nestedWb_c_set_hit_T_5; // @[Slice.scala 304:50]
  assign abc_mshr_2_io_nestedwb_clients_0_isToN = c_mshr_io_status_valid ? _nestedWb_clients_0_isToN_T_1 :
    _nestedWb_clients_0_isToN_T_3; // @[Slice.scala 314:25]
  assign abc_mshr_2_io_nestedwb_clients_1_isToN = c_mshr_io_status_valid ? _nestedWb_clients_1_isToN_T_1 :
    _nestedWb_clients_1_isToN_T_3; // @[Slice.scala 314:25]
  assign abc_mshr_2_io_tasks_sink_a_ready = 1'h0; // @[Slice.scala 472:13]
  assign abc_mshr_2_io_tasks_source_bready = sourceB_task_arb_io_in_2_ready; // @[Slice.scala 472:13]
  assign abc_mshr_2_io_tasks_sink_c_ready = sinkC_task_arb_io_in_2_ready; // @[Slice.scala 472:13]
  assign abc_mshr_2_io_tasks_source_d_ready = sourceD_task_arb_io_in_2_ready; // @[Slice.scala 472:13]
  assign abc_mshr_2_io_tasks_source_a_ready = sourceA_task_arb_io_in_2_ready; // @[Slice.scala 472:13]
  assign abc_mshr_2_io_tasks_source_c_ready = sourceC_task_arb_io_in_2_ready; // @[Slice.scala 472:13]
  assign abc_mshr_2_io_tasks_source_e_ready = sourceE_task_arb_io_in_2_ready; // @[Slice.scala 472:13]
  assign abc_mshr_2_io_tasks_dir_write_ready = arbiter_io_in_2_ready; // @[Slice.scala 406:60]
  assign abc_mshr_2_io_tasks_tag_write_ready = tagWrite_task_arb_io_in_2_ready; // @[Slice.scala 472:13]
  assign abc_mshr_2_io_tasks_client_dir_write_ready = arbiter_1_io_in_2_ready; // @[Slice.scala 406:60]
  assign abc_mshr_2_io_tasks_client_tag_write_ready = arbiter_2_io_in_2_ready; // @[Slice.scala 472:13]
  assign abc_mshr_2_io_dirResult_valid = ms_2_io_dirResult_valid_REG; // @[Slice.scala 556:31]
  assign abc_mshr_2_io_dirResult_bits_self_dirty = directory_io_result_bits_self_dirty; // @[Slice.scala 555:30]
  assign abc_mshr_2_io_dirResult_bits_self_state = directory_io_result_bits_self_state; // @[Slice.scala 555:30]
  assign abc_mshr_2_io_dirResult_bits_self_clientStates_0 = directory_io_result_bits_self_clientStates_0; // @[Slice.scala 555:30]
  assign abc_mshr_2_io_dirResult_bits_self_clientStates_1 = directory_io_result_bits_self_clientStates_1; // @[Slice.scala 555:30]
  assign abc_mshr_2_io_dirResult_bits_self_hit = directory_io_result_bits_self_hit; // @[Slice.scala 555:30]
  assign abc_mshr_2_io_dirResult_bits_self_way = directory_io_result_bits_self_way; // @[Slice.scala 555:30]
  assign abc_mshr_2_io_dirResult_bits_self_tag = directory_io_result_bits_self_tag; // @[Slice.scala 555:30]
  assign abc_mshr_2_io_dirResult_bits_clients_states_0_state = directory_io_result_bits_clients_states_0_state; // @[Slice.scala 555:30]
  assign abc_mshr_2_io_dirResult_bits_clients_states_0_hit = directory_io_result_bits_clients_states_0_hit; // @[Slice.scala 555:30]
  assign abc_mshr_2_io_dirResult_bits_clients_states_1_state = directory_io_result_bits_clients_states_1_state; // @[Slice.scala 555:30]
  assign abc_mshr_2_io_dirResult_bits_clients_states_1_hit = directory_io_result_bits_clients_states_1_hit; // @[Slice.scala 555:30]
  assign abc_mshr_2_io_dirResult_bits_clients_tag = directory_io_result_bits_clients_tag; // @[Slice.scala 555:30]
  assign abc_mshr_2_io_dirResult_bits_clients_way = directory_io_result_bits_clients_way; // @[Slice.scala 555:30]
  assign abc_mshr_2_io_c_status_set = c_mshr_io_status_bits_set; // @[Slice.scala 209:28]
  assign abc_mshr_2_io_c_status_tag = c_mshr_io_status_bits_tag; // @[Slice.scala 210:28]
  assign abc_mshr_2_io_c_status_way = c_mshr_io_status_bits_way; // @[Slice.scala 211:28]
  assign abc_mshr_2_io_c_status_nestedReleaseData = c_mshr_io_status_valid & c_mshr_io_is_nestedReleaseData; // @[Slice.scala 213:32]
  assign abc_mshr_2_io_bstatus_set = bc_mshr_io_status_bits_set; // @[Slice.scala 214:28]
  assign abc_mshr_2_io_bstatus_tag = bc_mshr_io_status_bits_tag; // @[Slice.scala 215:28]
  assign abc_mshr_2_io_bstatus_way = bc_mshr_io_status_bits_way; // @[Slice.scala 216:28]
  assign abc_mshr_2_io_bstatus_nestedProbeAckData = bc_mshr_io_status_valid & bc_mshr_io_is_nestedProbeAckData; // @[Slice.scala 218:33]
  assign abc_mshr_2_io_bstatus_probeHelperFinish = bc_mshr_io_status_valid & bc_mshr_io_probeHelperFinish; // @[Slice.scala 220:33]
  assign abc_mshr_2_io_releaseThrough = 1'h0; // @[Slice.scala 221:30]
  assign abc_mshr_2_io_probeAckDataThrough = 1'h0; // @[Slice.scala 222:35]
  assign abc_mshr_3_clock = clock;
  assign abc_mshr_3_reset = reset;
  assign abc_mshr_3_io_id = 4'h3; // @[Slice.scala 166:18]
  assign abc_mshr_3_io_enable = ~(bc_disable_3 | c_disable_3); // @[Slice.scala 198:25]
  assign abc_mshr_3_io_alloc_valid = mshrAlloc_io_alloc_3_valid; // @[Slice.scala 167:21]
  assign abc_mshr_3_io_alloc_bits_channel = mshrAlloc_io_alloc_3_bits_channel; // @[Slice.scala 167:21]
  assign abc_mshr_3_io_alloc_bits_opcode = mshrAlloc_io_alloc_3_bits_opcode; // @[Slice.scala 167:21]
  assign abc_mshr_3_io_alloc_bits_param = mshrAlloc_io_alloc_3_bits_param; // @[Slice.scala 167:21]
  assign abc_mshr_3_io_alloc_bits_size = mshrAlloc_io_alloc_3_bits_size; // @[Slice.scala 167:21]
  assign abc_mshr_3_io_alloc_bits_source = mshrAlloc_io_alloc_3_bits_source; // @[Slice.scala 167:21]
  assign abc_mshr_3_io_alloc_bits_set = mshrAlloc_io_alloc_3_bits_set; // @[Slice.scala 167:21]
  assign abc_mshr_3_io_alloc_bits_tag = mshrAlloc_io_alloc_3_bits_tag; // @[Slice.scala 167:21]
  assign abc_mshr_3_io_alloc_bits_off = mshrAlloc_io_alloc_3_bits_off; // @[Slice.scala 167:21]
  assign abc_mshr_3_io_alloc_bits_mask = mshrAlloc_io_alloc_3_bits_mask; // @[Slice.scala 167:21]
  assign abc_mshr_3_io_alloc_bits_bufIdx = mshrAlloc_io_alloc_3_bits_bufIdx; // @[Slice.scala 167:21]
  assign abc_mshr_3_io_alloc_bits_preferCache = mshrAlloc_io_alloc_3_bits_preferCache; // @[Slice.scala 167:21]
  assign abc_mshr_3_io_alloc_bits_dirty = mshrAlloc_io_alloc_3_bits_dirty; // @[Slice.scala 167:21]
  assign abc_mshr_3_io_alloc_bits_fromProbeHelper = mshrAlloc_io_alloc_3_bits_fromProbeHelper; // @[Slice.scala 167:21]
  assign abc_mshr_3_io_alloc_bits_fromCmoHelper = mshrAlloc_io_alloc_3_bits_fromCmoHelper; // @[Slice.scala 167:21]
  assign abc_mshr_3_io_alloc_bits_needProbeAckData = mshrAlloc_io_alloc_3_bits_needProbeAckData; // @[Slice.scala 167:21]
  assign abc_mshr_3_io_resps_sink_c_valid = sinkC_io_resp_valid & sinkC_io_resp_bits_set ==
    abc_mshr_3_io_status_bits_set; // @[Slice.scala 527:57]
  assign abc_mshr_3_io_resps_sink_c_bits_hasData = sinkC_io_resp_bits_hasData; // @[Slice.scala 531:33]
  assign abc_mshr_3_io_resps_sink_c_bits_param = sinkC_io_resp_bits_param; // @[Slice.scala 531:33]
  assign abc_mshr_3_io_resps_sink_c_bits_source = sinkC_io_resp_bits_source; // @[Slice.scala 531:33]
  assign abc_mshr_3_io_resps_sink_c_bits_last = sinkC_io_resp_bits_last; // @[Slice.scala 531:33]
  assign abc_mshr_3_io_resps_sink_c_bits_bufIdx = sinkC_io_resp_bits_bufIdx; // @[Slice.scala 531:33]
  assign abc_mshr_3_io_resps_sink_d_valid = sinkD_io_resp_valid & sinkD_io_resp_bits_source == 4'h3; // @[Slice.scala 528:57]
  assign abc_mshr_3_io_resps_sink_d_bits_opcode = sinkD_io_resp_bits_opcode; // @[Slice.scala 532:33]
  assign abc_mshr_3_io_resps_sink_d_bits_param = sinkD_io_resp_bits_param; // @[Slice.scala 532:33]
  assign abc_mshr_3_io_resps_sink_d_bits_sink = sinkD_io_resp_bits_sink; // @[Slice.scala 532:33]
  assign abc_mshr_3_io_resps_sink_d_bits_last = sinkD_io_resp_bits_last; // @[Slice.scala 532:33]
  assign abc_mshr_3_io_resps_sink_d_bits_denied = sinkD_io_resp_bits_denied; // @[Slice.scala 532:33]
  assign abc_mshr_3_io_resps_sink_d_bits_bufIdx = sinkD_io_resp_bits_bufIdx; // @[Slice.scala 532:33]
  assign abc_mshr_3_io_resps_sink_e_valid = sinkE_io_resp_valid & sinkE_io_resp_bits_sink == 4'h3; // @[Slice.scala 529:57]
  assign abc_mshr_3_io_resps_source_d_valid = sourceD_io_resp_valid & sourceD_io_resp_bits_sink == 4'h3; // @[Slice.scala 530:61]
  assign abc_mshr_3_io_nestedwb_set = c_mshr_io_status_valid ? c_mshr_io_status_bits_set : bc_mshr_io_status_bits_set; // @[Slice.scala 258:22]
  assign abc_mshr_3_io_nestedwb_tag = c_mshr_io_status_valid ? c_mshr_io_status_bits_tag : bc_mshr_io_status_bits_tag; // @[Slice.scala 259:22]
  assign abc_mshr_3_io_nestedwb_btoN = _nestedWb_btoN_T_2 & _nestedWb_btoN_T_3; // @[Slice.scala 280:38]
  assign abc_mshr_3_io_nestedwb_btoB = _nestedWb_btoN_T_2 & _nestedWb_btoB_T_3; // @[Slice.scala 283:38]
  assign abc_mshr_3_io_nestedwb_bclr_dirty = _nestedWb_btoN_T_2 & _nestedWb_bclr_dirty_T_4; // @[Slice.scala 286:38]
  assign abc_mshr_3_io_nestedwb_bset_dirty = _nestedWb_btoN_T_2 & bc_mshr_io_tasks_dir_write_bits_data_dirty; // @[Slice.scala 289:38]
  assign abc_mshr_3_io_nestedwb_c_set_dirty = _nestedWb_c_set_dirty_T & c_mshr_io_tasks_dir_write_bits_data_dirty; // @[Slice.scala 292:37]
  assign abc_mshr_3_io_nestedwb_c_set_hit = c_mshr_io_status_valid & c_mshr_io_tasks_tag_write_valid &
    _nestedWb_c_set_hit_T_7; // @[Slice.scala 304:50]
  assign abc_mshr_3_io_nestedwb_clients_0_isToN = c_mshr_io_status_valid ? _nestedWb_clients_0_isToN_T_1 :
    _nestedWb_clients_0_isToN_T_3; // @[Slice.scala 314:25]
  assign abc_mshr_3_io_nestedwb_clients_1_isToN = c_mshr_io_status_valid ? _nestedWb_clients_1_isToN_T_1 :
    _nestedWb_clients_1_isToN_T_3; // @[Slice.scala 314:25]
  assign abc_mshr_3_io_tasks_sink_a_ready = 1'h0; // @[Slice.scala 472:13]
  assign abc_mshr_3_io_tasks_source_bready = sourceB_task_arb_io_in_3_ready; // @[Slice.scala 472:13]
  assign abc_mshr_3_io_tasks_sink_c_ready = sinkC_task_arb_io_in_3_ready; // @[Slice.scala 472:13]
  assign abc_mshr_3_io_tasks_source_d_ready = sourceD_task_arb_io_in_3_ready; // @[Slice.scala 472:13]
  assign abc_mshr_3_io_tasks_source_a_ready = sourceA_task_arb_io_in_3_ready; // @[Slice.scala 472:13]
  assign abc_mshr_3_io_tasks_source_c_ready = sourceC_task_arb_io_in_3_ready; // @[Slice.scala 472:13]
  assign abc_mshr_3_io_tasks_source_e_ready = sourceE_task_arb_io_in_3_ready; // @[Slice.scala 472:13]
  assign abc_mshr_3_io_tasks_dir_write_ready = arbiter_io_in_3_ready; // @[Slice.scala 406:60]
  assign abc_mshr_3_io_tasks_tag_write_ready = tagWrite_task_arb_io_in_3_ready; // @[Slice.scala 472:13]
  assign abc_mshr_3_io_tasks_client_dir_write_ready = arbiter_1_io_in_3_ready; // @[Slice.scala 406:60]
  assign abc_mshr_3_io_tasks_client_tag_write_ready = arbiter_2_io_in_3_ready; // @[Slice.scala 472:13]
  assign abc_mshr_3_io_dirResult_valid = ms_3_io_dirResult_valid_REG; // @[Slice.scala 556:31]
  assign abc_mshr_3_io_dirResult_bits_self_dirty = directory_io_result_bits_self_dirty; // @[Slice.scala 555:30]
  assign abc_mshr_3_io_dirResult_bits_self_state = directory_io_result_bits_self_state; // @[Slice.scala 555:30]
  assign abc_mshr_3_io_dirResult_bits_self_clientStates_0 = directory_io_result_bits_self_clientStates_0; // @[Slice.scala 555:30]
  assign abc_mshr_3_io_dirResult_bits_self_clientStates_1 = directory_io_result_bits_self_clientStates_1; // @[Slice.scala 555:30]
  assign abc_mshr_3_io_dirResult_bits_self_hit = directory_io_result_bits_self_hit; // @[Slice.scala 555:30]
  assign abc_mshr_3_io_dirResult_bits_self_way = directory_io_result_bits_self_way; // @[Slice.scala 555:30]
  assign abc_mshr_3_io_dirResult_bits_self_tag = directory_io_result_bits_self_tag; // @[Slice.scala 555:30]
  assign abc_mshr_3_io_dirResult_bits_clients_states_0_state = directory_io_result_bits_clients_states_0_state; // @[Slice.scala 555:30]
  assign abc_mshr_3_io_dirResult_bits_clients_states_0_hit = directory_io_result_bits_clients_states_0_hit; // @[Slice.scala 555:30]
  assign abc_mshr_3_io_dirResult_bits_clients_states_1_state = directory_io_result_bits_clients_states_1_state; // @[Slice.scala 555:30]
  assign abc_mshr_3_io_dirResult_bits_clients_states_1_hit = directory_io_result_bits_clients_states_1_hit; // @[Slice.scala 555:30]
  assign abc_mshr_3_io_dirResult_bits_clients_tag = directory_io_result_bits_clients_tag; // @[Slice.scala 555:30]
  assign abc_mshr_3_io_dirResult_bits_clients_way = directory_io_result_bits_clients_way; // @[Slice.scala 555:30]
  assign abc_mshr_3_io_c_status_set = c_mshr_io_status_bits_set; // @[Slice.scala 209:28]
  assign abc_mshr_3_io_c_status_tag = c_mshr_io_status_bits_tag; // @[Slice.scala 210:28]
  assign abc_mshr_3_io_c_status_way = c_mshr_io_status_bits_way; // @[Slice.scala 211:28]
  assign abc_mshr_3_io_c_status_nestedReleaseData = c_mshr_io_status_valid & c_mshr_io_is_nestedReleaseData; // @[Slice.scala 213:32]
  assign abc_mshr_3_io_bstatus_set = bc_mshr_io_status_bits_set; // @[Slice.scala 214:28]
  assign abc_mshr_3_io_bstatus_tag = bc_mshr_io_status_bits_tag; // @[Slice.scala 215:28]
  assign abc_mshr_3_io_bstatus_way = bc_mshr_io_status_bits_way; // @[Slice.scala 216:28]
  assign abc_mshr_3_io_bstatus_nestedProbeAckData = bc_mshr_io_status_valid & bc_mshr_io_is_nestedProbeAckData; // @[Slice.scala 218:33]
  assign abc_mshr_3_io_bstatus_probeHelperFinish = bc_mshr_io_status_valid & bc_mshr_io_probeHelperFinish; // @[Slice.scala 220:33]
  assign abc_mshr_3_io_releaseThrough = 1'h0; // @[Slice.scala 221:30]
  assign abc_mshr_3_io_probeAckDataThrough = 1'h0; // @[Slice.scala 222:35]
  assign abc_mshr_4_clock = clock;
  assign abc_mshr_4_reset = reset;
  assign abc_mshr_4_io_id = 4'h4; // @[Slice.scala 166:18]
  assign abc_mshr_4_io_enable = ~(bc_disable_4 | c_disable_4); // @[Slice.scala 198:25]
  assign abc_mshr_4_io_alloc_valid = mshrAlloc_io_alloc_4_valid; // @[Slice.scala 167:21]
  assign abc_mshr_4_io_alloc_bits_channel = mshrAlloc_io_alloc_4_bits_channel; // @[Slice.scala 167:21]
  assign abc_mshr_4_io_alloc_bits_opcode = mshrAlloc_io_alloc_4_bits_opcode; // @[Slice.scala 167:21]
  assign abc_mshr_4_io_alloc_bits_param = mshrAlloc_io_alloc_4_bits_param; // @[Slice.scala 167:21]
  assign abc_mshr_4_io_alloc_bits_size = mshrAlloc_io_alloc_4_bits_size; // @[Slice.scala 167:21]
  assign abc_mshr_4_io_alloc_bits_source = mshrAlloc_io_alloc_4_bits_source; // @[Slice.scala 167:21]
  assign abc_mshr_4_io_alloc_bits_set = mshrAlloc_io_alloc_4_bits_set; // @[Slice.scala 167:21]
  assign abc_mshr_4_io_alloc_bits_tag = mshrAlloc_io_alloc_4_bits_tag; // @[Slice.scala 167:21]
  assign abc_mshr_4_io_alloc_bits_off = mshrAlloc_io_alloc_4_bits_off; // @[Slice.scala 167:21]
  assign abc_mshr_4_io_alloc_bits_mask = mshrAlloc_io_alloc_4_bits_mask; // @[Slice.scala 167:21]
  assign abc_mshr_4_io_alloc_bits_bufIdx = mshrAlloc_io_alloc_4_bits_bufIdx; // @[Slice.scala 167:21]
  assign abc_mshr_4_io_alloc_bits_preferCache = mshrAlloc_io_alloc_4_bits_preferCache; // @[Slice.scala 167:21]
  assign abc_mshr_4_io_alloc_bits_dirty = mshrAlloc_io_alloc_4_bits_dirty; // @[Slice.scala 167:21]
  assign abc_mshr_4_io_alloc_bits_fromProbeHelper = mshrAlloc_io_alloc_4_bits_fromProbeHelper; // @[Slice.scala 167:21]
  assign abc_mshr_4_io_alloc_bits_fromCmoHelper = mshrAlloc_io_alloc_4_bits_fromCmoHelper; // @[Slice.scala 167:21]
  assign abc_mshr_4_io_alloc_bits_needProbeAckData = mshrAlloc_io_alloc_4_bits_needProbeAckData; // @[Slice.scala 167:21]
  assign abc_mshr_4_io_resps_sink_c_valid = sinkC_io_resp_valid & sinkC_io_resp_bits_set ==
    abc_mshr_4_io_status_bits_set; // @[Slice.scala 527:57]
  assign abc_mshr_4_io_resps_sink_c_bits_hasData = sinkC_io_resp_bits_hasData; // @[Slice.scala 531:33]
  assign abc_mshr_4_io_resps_sink_c_bits_param = sinkC_io_resp_bits_param; // @[Slice.scala 531:33]
  assign abc_mshr_4_io_resps_sink_c_bits_source = sinkC_io_resp_bits_source; // @[Slice.scala 531:33]
  assign abc_mshr_4_io_resps_sink_c_bits_last = sinkC_io_resp_bits_last; // @[Slice.scala 531:33]
  assign abc_mshr_4_io_resps_sink_c_bits_bufIdx = sinkC_io_resp_bits_bufIdx; // @[Slice.scala 531:33]
  assign abc_mshr_4_io_resps_sink_d_valid = sinkD_io_resp_valid & sinkD_io_resp_bits_source == 4'h4; // @[Slice.scala 528:57]
  assign abc_mshr_4_io_resps_sink_d_bits_opcode = sinkD_io_resp_bits_opcode; // @[Slice.scala 532:33]
  assign abc_mshr_4_io_resps_sink_d_bits_param = sinkD_io_resp_bits_param; // @[Slice.scala 532:33]
  assign abc_mshr_4_io_resps_sink_d_bits_sink = sinkD_io_resp_bits_sink; // @[Slice.scala 532:33]
  assign abc_mshr_4_io_resps_sink_d_bits_last = sinkD_io_resp_bits_last; // @[Slice.scala 532:33]
  assign abc_mshr_4_io_resps_sink_d_bits_denied = sinkD_io_resp_bits_denied; // @[Slice.scala 532:33]
  assign abc_mshr_4_io_resps_sink_d_bits_bufIdx = sinkD_io_resp_bits_bufIdx; // @[Slice.scala 532:33]
  assign abc_mshr_4_io_resps_sink_e_valid = sinkE_io_resp_valid & sinkE_io_resp_bits_sink == 4'h4; // @[Slice.scala 529:57]
  assign abc_mshr_4_io_resps_source_d_valid = sourceD_io_resp_valid & sourceD_io_resp_bits_sink == 4'h4; // @[Slice.scala 530:61]
  assign abc_mshr_4_io_nestedwb_set = c_mshr_io_status_valid ? c_mshr_io_status_bits_set : bc_mshr_io_status_bits_set; // @[Slice.scala 258:22]
  assign abc_mshr_4_io_nestedwb_tag = c_mshr_io_status_valid ? c_mshr_io_status_bits_tag : bc_mshr_io_status_bits_tag; // @[Slice.scala 259:22]
  assign abc_mshr_4_io_nestedwb_btoN = _nestedWb_btoN_T_2 & _nestedWb_btoN_T_3; // @[Slice.scala 280:38]
  assign abc_mshr_4_io_nestedwb_btoB = _nestedWb_btoN_T_2 & _nestedWb_btoB_T_3; // @[Slice.scala 283:38]
  assign abc_mshr_4_io_nestedwb_bclr_dirty = _nestedWb_btoN_T_2 & _nestedWb_bclr_dirty_T_4; // @[Slice.scala 286:38]
  assign abc_mshr_4_io_nestedwb_bset_dirty = _nestedWb_btoN_T_2 & bc_mshr_io_tasks_dir_write_bits_data_dirty; // @[Slice.scala 289:38]
  assign abc_mshr_4_io_nestedwb_c_set_dirty = _nestedWb_c_set_dirty_T & c_mshr_io_tasks_dir_write_bits_data_dirty; // @[Slice.scala 292:37]
  assign abc_mshr_4_io_nestedwb_c_set_hit = c_mshr_io_status_valid & c_mshr_io_tasks_tag_write_valid &
    _nestedWb_c_set_hit_T_9; // @[Slice.scala 304:50]
  assign abc_mshr_4_io_nestedwb_clients_0_isToN = c_mshr_io_status_valid ? _nestedWb_clients_0_isToN_T_1 :
    _nestedWb_clients_0_isToN_T_3; // @[Slice.scala 314:25]
  assign abc_mshr_4_io_nestedwb_clients_1_isToN = c_mshr_io_status_valid ? _nestedWb_clients_1_isToN_T_1 :
    _nestedWb_clients_1_isToN_T_3; // @[Slice.scala 314:25]
  assign abc_mshr_4_io_tasks_sink_a_ready = 1'h0; // @[Slice.scala 472:13]
  assign abc_mshr_4_io_tasks_source_bready = sourceB_task_arb_io_in_4_ready; // @[Slice.scala 472:13]
  assign abc_mshr_4_io_tasks_sink_c_ready = sinkC_task_arb_io_in_4_ready; // @[Slice.scala 472:13]
  assign abc_mshr_4_io_tasks_source_d_ready = sourceD_task_arb_io_in_4_ready; // @[Slice.scala 472:13]
  assign abc_mshr_4_io_tasks_source_a_ready = sourceA_task_arb_io_in_4_ready; // @[Slice.scala 472:13]
  assign abc_mshr_4_io_tasks_source_c_ready = sourceC_task_arb_io_in_4_ready; // @[Slice.scala 472:13]
  assign abc_mshr_4_io_tasks_source_e_ready = sourceE_task_arb_io_in_4_ready; // @[Slice.scala 472:13]
  assign abc_mshr_4_io_tasks_dir_write_ready = arbiter_io_in_4_ready; // @[Slice.scala 406:60]
  assign abc_mshr_4_io_tasks_tag_write_ready = tagWrite_task_arb_io_in_4_ready; // @[Slice.scala 472:13]
  assign abc_mshr_4_io_tasks_client_dir_write_ready = arbiter_1_io_in_4_ready; // @[Slice.scala 406:60]
  assign abc_mshr_4_io_tasks_client_tag_write_ready = arbiter_2_io_in_4_ready; // @[Slice.scala 472:13]
  assign abc_mshr_4_io_dirResult_valid = ms_4_io_dirResult_valid_REG; // @[Slice.scala 556:31]
  assign abc_mshr_4_io_dirResult_bits_self_dirty = directory_io_result_bits_self_dirty; // @[Slice.scala 555:30]
  assign abc_mshr_4_io_dirResult_bits_self_state = directory_io_result_bits_self_state; // @[Slice.scala 555:30]
  assign abc_mshr_4_io_dirResult_bits_self_clientStates_0 = directory_io_result_bits_self_clientStates_0; // @[Slice.scala 555:30]
  assign abc_mshr_4_io_dirResult_bits_self_clientStates_1 = directory_io_result_bits_self_clientStates_1; // @[Slice.scala 555:30]
  assign abc_mshr_4_io_dirResult_bits_self_hit = directory_io_result_bits_self_hit; // @[Slice.scala 555:30]
  assign abc_mshr_4_io_dirResult_bits_self_way = directory_io_result_bits_self_way; // @[Slice.scala 555:30]
  assign abc_mshr_4_io_dirResult_bits_self_tag = directory_io_result_bits_self_tag; // @[Slice.scala 555:30]
  assign abc_mshr_4_io_dirResult_bits_clients_states_0_state = directory_io_result_bits_clients_states_0_state; // @[Slice.scala 555:30]
  assign abc_mshr_4_io_dirResult_bits_clients_states_0_hit = directory_io_result_bits_clients_states_0_hit; // @[Slice.scala 555:30]
  assign abc_mshr_4_io_dirResult_bits_clients_states_1_state = directory_io_result_bits_clients_states_1_state; // @[Slice.scala 555:30]
  assign abc_mshr_4_io_dirResult_bits_clients_states_1_hit = directory_io_result_bits_clients_states_1_hit; // @[Slice.scala 555:30]
  assign abc_mshr_4_io_dirResult_bits_clients_tag = directory_io_result_bits_clients_tag; // @[Slice.scala 555:30]
  assign abc_mshr_4_io_dirResult_bits_clients_way = directory_io_result_bits_clients_way; // @[Slice.scala 555:30]
  assign abc_mshr_4_io_c_status_set = c_mshr_io_status_bits_set; // @[Slice.scala 209:28]
  assign abc_mshr_4_io_c_status_tag = c_mshr_io_status_bits_tag; // @[Slice.scala 210:28]
  assign abc_mshr_4_io_c_status_way = c_mshr_io_status_bits_way; // @[Slice.scala 211:28]
  assign abc_mshr_4_io_c_status_nestedReleaseData = c_mshr_io_status_valid & c_mshr_io_is_nestedReleaseData; // @[Slice.scala 213:32]
  assign abc_mshr_4_io_bstatus_set = bc_mshr_io_status_bits_set; // @[Slice.scala 214:28]
  assign abc_mshr_4_io_bstatus_tag = bc_mshr_io_status_bits_tag; // @[Slice.scala 215:28]
  assign abc_mshr_4_io_bstatus_way = bc_mshr_io_status_bits_way; // @[Slice.scala 216:28]
  assign abc_mshr_4_io_bstatus_nestedProbeAckData = bc_mshr_io_status_valid & bc_mshr_io_is_nestedProbeAckData; // @[Slice.scala 218:33]
  assign abc_mshr_4_io_bstatus_probeHelperFinish = bc_mshr_io_status_valid & bc_mshr_io_probeHelperFinish; // @[Slice.scala 220:33]
  assign abc_mshr_4_io_releaseThrough = 1'h0; // @[Slice.scala 221:30]
  assign abc_mshr_4_io_probeAckDataThrough = 1'h0; // @[Slice.scala 222:35]
  assign abc_mshr_5_clock = clock;
  assign abc_mshr_5_reset = reset;
  assign abc_mshr_5_io_id = 4'h5; // @[Slice.scala 166:18]
  assign abc_mshr_5_io_enable = ~(bc_disable_5 | c_disable_5); // @[Slice.scala 198:25]
  assign abc_mshr_5_io_alloc_valid = mshrAlloc_io_alloc_5_valid; // @[Slice.scala 167:21]
  assign abc_mshr_5_io_alloc_bits_channel = mshrAlloc_io_alloc_5_bits_channel; // @[Slice.scala 167:21]
  assign abc_mshr_5_io_alloc_bits_opcode = mshrAlloc_io_alloc_5_bits_opcode; // @[Slice.scala 167:21]
  assign abc_mshr_5_io_alloc_bits_param = mshrAlloc_io_alloc_5_bits_param; // @[Slice.scala 167:21]
  assign abc_mshr_5_io_alloc_bits_size = mshrAlloc_io_alloc_5_bits_size; // @[Slice.scala 167:21]
  assign abc_mshr_5_io_alloc_bits_source = mshrAlloc_io_alloc_5_bits_source; // @[Slice.scala 167:21]
  assign abc_mshr_5_io_alloc_bits_set = mshrAlloc_io_alloc_5_bits_set; // @[Slice.scala 167:21]
  assign abc_mshr_5_io_alloc_bits_tag = mshrAlloc_io_alloc_5_bits_tag; // @[Slice.scala 167:21]
  assign abc_mshr_5_io_alloc_bits_off = mshrAlloc_io_alloc_5_bits_off; // @[Slice.scala 167:21]
  assign abc_mshr_5_io_alloc_bits_mask = mshrAlloc_io_alloc_5_bits_mask; // @[Slice.scala 167:21]
  assign abc_mshr_5_io_alloc_bits_bufIdx = mshrAlloc_io_alloc_5_bits_bufIdx; // @[Slice.scala 167:21]
  assign abc_mshr_5_io_alloc_bits_preferCache = mshrAlloc_io_alloc_5_bits_preferCache; // @[Slice.scala 167:21]
  assign abc_mshr_5_io_alloc_bits_dirty = mshrAlloc_io_alloc_5_bits_dirty; // @[Slice.scala 167:21]
  assign abc_mshr_5_io_alloc_bits_fromProbeHelper = mshrAlloc_io_alloc_5_bits_fromProbeHelper; // @[Slice.scala 167:21]
  assign abc_mshr_5_io_alloc_bits_fromCmoHelper = mshrAlloc_io_alloc_5_bits_fromCmoHelper; // @[Slice.scala 167:21]
  assign abc_mshr_5_io_alloc_bits_needProbeAckData = mshrAlloc_io_alloc_5_bits_needProbeAckData; // @[Slice.scala 167:21]
  assign abc_mshr_5_io_resps_sink_c_valid = sinkC_io_resp_valid & sinkC_io_resp_bits_set ==
    abc_mshr_5_io_status_bits_set; // @[Slice.scala 527:57]
  assign abc_mshr_5_io_resps_sink_c_bits_hasData = sinkC_io_resp_bits_hasData; // @[Slice.scala 531:33]
  assign abc_mshr_5_io_resps_sink_c_bits_param = sinkC_io_resp_bits_param; // @[Slice.scala 531:33]
  assign abc_mshr_5_io_resps_sink_c_bits_source = sinkC_io_resp_bits_source; // @[Slice.scala 531:33]
  assign abc_mshr_5_io_resps_sink_c_bits_last = sinkC_io_resp_bits_last; // @[Slice.scala 531:33]
  assign abc_mshr_5_io_resps_sink_c_bits_bufIdx = sinkC_io_resp_bits_bufIdx; // @[Slice.scala 531:33]
  assign abc_mshr_5_io_resps_sink_d_valid = sinkD_io_resp_valid & sinkD_io_resp_bits_source == 4'h5; // @[Slice.scala 528:57]
  assign abc_mshr_5_io_resps_sink_d_bits_opcode = sinkD_io_resp_bits_opcode; // @[Slice.scala 532:33]
  assign abc_mshr_5_io_resps_sink_d_bits_param = sinkD_io_resp_bits_param; // @[Slice.scala 532:33]
  assign abc_mshr_5_io_resps_sink_d_bits_sink = sinkD_io_resp_bits_sink; // @[Slice.scala 532:33]
  assign abc_mshr_5_io_resps_sink_d_bits_last = sinkD_io_resp_bits_last; // @[Slice.scala 532:33]
  assign abc_mshr_5_io_resps_sink_d_bits_denied = sinkD_io_resp_bits_denied; // @[Slice.scala 532:33]
  assign abc_mshr_5_io_resps_sink_d_bits_bufIdx = sinkD_io_resp_bits_bufIdx; // @[Slice.scala 532:33]
  assign abc_mshr_5_io_resps_sink_e_valid = sinkE_io_resp_valid & sinkE_io_resp_bits_sink == 4'h5; // @[Slice.scala 529:57]
  assign abc_mshr_5_io_resps_source_d_valid = sourceD_io_resp_valid & sourceD_io_resp_bits_sink == 4'h5; // @[Slice.scala 530:61]
  assign abc_mshr_5_io_nestedwb_set = c_mshr_io_status_valid ? c_mshr_io_status_bits_set : bc_mshr_io_status_bits_set; // @[Slice.scala 258:22]
  assign abc_mshr_5_io_nestedwb_tag = c_mshr_io_status_valid ? c_mshr_io_status_bits_tag : bc_mshr_io_status_bits_tag; // @[Slice.scala 259:22]
  assign abc_mshr_5_io_nestedwb_btoN = _nestedWb_btoN_T_2 & _nestedWb_btoN_T_3; // @[Slice.scala 280:38]
  assign abc_mshr_5_io_nestedwb_btoB = _nestedWb_btoN_T_2 & _nestedWb_btoB_T_3; // @[Slice.scala 283:38]
  assign abc_mshr_5_io_nestedwb_bclr_dirty = _nestedWb_btoN_T_2 & _nestedWb_bclr_dirty_T_4; // @[Slice.scala 286:38]
  assign abc_mshr_5_io_nestedwb_bset_dirty = _nestedWb_btoN_T_2 & bc_mshr_io_tasks_dir_write_bits_data_dirty; // @[Slice.scala 289:38]
  assign abc_mshr_5_io_nestedwb_c_set_dirty = _nestedWb_c_set_dirty_T & c_mshr_io_tasks_dir_write_bits_data_dirty; // @[Slice.scala 292:37]
  assign abc_mshr_5_io_nestedwb_c_set_hit = c_mshr_io_status_valid & c_mshr_io_tasks_tag_write_valid &
    _nestedWb_c_set_hit_T_11; // @[Slice.scala 304:50]
  assign abc_mshr_5_io_nestedwb_clients_0_isToN = c_mshr_io_status_valid ? _nestedWb_clients_0_isToN_T_1 :
    _nestedWb_clients_0_isToN_T_3; // @[Slice.scala 314:25]
  assign abc_mshr_5_io_nestedwb_clients_1_isToN = c_mshr_io_status_valid ? _nestedWb_clients_1_isToN_T_1 :
    _nestedWb_clients_1_isToN_T_3; // @[Slice.scala 314:25]
  assign abc_mshr_5_io_tasks_sink_a_ready = 1'h0; // @[Slice.scala 472:13]
  assign abc_mshr_5_io_tasks_source_bready = sourceB_task_arb_io_in_5_ready; // @[Slice.scala 472:13]
  assign abc_mshr_5_io_tasks_sink_c_ready = sinkC_task_arb_io_in_5_ready; // @[Slice.scala 472:13]
  assign abc_mshr_5_io_tasks_source_d_ready = sourceD_task_arb_io_in_5_ready; // @[Slice.scala 472:13]
  assign abc_mshr_5_io_tasks_source_a_ready = sourceA_task_arb_io_in_5_ready; // @[Slice.scala 472:13]
  assign abc_mshr_5_io_tasks_source_c_ready = sourceC_task_arb_io_in_5_ready; // @[Slice.scala 472:13]
  assign abc_mshr_5_io_tasks_source_e_ready = sourceE_task_arb_io_in_5_ready; // @[Slice.scala 472:13]
  assign abc_mshr_5_io_tasks_dir_write_ready = arbiter_io_in_5_ready; // @[Slice.scala 406:60]
  assign abc_mshr_5_io_tasks_tag_write_ready = tagWrite_task_arb_io_in_5_ready; // @[Slice.scala 472:13]
  assign abc_mshr_5_io_tasks_client_dir_write_ready = arbiter_1_io_in_5_ready; // @[Slice.scala 406:60]
  assign abc_mshr_5_io_tasks_client_tag_write_ready = arbiter_2_io_in_5_ready; // @[Slice.scala 472:13]
  assign abc_mshr_5_io_dirResult_valid = ms_5_io_dirResult_valid_REG; // @[Slice.scala 556:31]
  assign abc_mshr_5_io_dirResult_bits_self_dirty = directory_io_result_bits_self_dirty; // @[Slice.scala 555:30]
  assign abc_mshr_5_io_dirResult_bits_self_state = directory_io_result_bits_self_state; // @[Slice.scala 555:30]
  assign abc_mshr_5_io_dirResult_bits_self_clientStates_0 = directory_io_result_bits_self_clientStates_0; // @[Slice.scala 555:30]
  assign abc_mshr_5_io_dirResult_bits_self_clientStates_1 = directory_io_result_bits_self_clientStates_1; // @[Slice.scala 555:30]
  assign abc_mshr_5_io_dirResult_bits_self_hit = directory_io_result_bits_self_hit; // @[Slice.scala 555:30]
  assign abc_mshr_5_io_dirResult_bits_self_way = directory_io_result_bits_self_way; // @[Slice.scala 555:30]
  assign abc_mshr_5_io_dirResult_bits_self_tag = directory_io_result_bits_self_tag; // @[Slice.scala 555:30]
  assign abc_mshr_5_io_dirResult_bits_clients_states_0_state = directory_io_result_bits_clients_states_0_state; // @[Slice.scala 555:30]
  assign abc_mshr_5_io_dirResult_bits_clients_states_0_hit = directory_io_result_bits_clients_states_0_hit; // @[Slice.scala 555:30]
  assign abc_mshr_5_io_dirResult_bits_clients_states_1_state = directory_io_result_bits_clients_states_1_state; // @[Slice.scala 555:30]
  assign abc_mshr_5_io_dirResult_bits_clients_states_1_hit = directory_io_result_bits_clients_states_1_hit; // @[Slice.scala 555:30]
  assign abc_mshr_5_io_dirResult_bits_clients_tag = directory_io_result_bits_clients_tag; // @[Slice.scala 555:30]
  assign abc_mshr_5_io_dirResult_bits_clients_way = directory_io_result_bits_clients_way; // @[Slice.scala 555:30]
  assign abc_mshr_5_io_c_status_set = c_mshr_io_status_bits_set; // @[Slice.scala 209:28]
  assign abc_mshr_5_io_c_status_tag = c_mshr_io_status_bits_tag; // @[Slice.scala 210:28]
  assign abc_mshr_5_io_c_status_way = c_mshr_io_status_bits_way; // @[Slice.scala 211:28]
  assign abc_mshr_5_io_c_status_nestedReleaseData = c_mshr_io_status_valid & c_mshr_io_is_nestedReleaseData; // @[Slice.scala 213:32]
  assign abc_mshr_5_io_bstatus_set = bc_mshr_io_status_bits_set; // @[Slice.scala 214:28]
  assign abc_mshr_5_io_bstatus_tag = bc_mshr_io_status_bits_tag; // @[Slice.scala 215:28]
  assign abc_mshr_5_io_bstatus_way = bc_mshr_io_status_bits_way; // @[Slice.scala 216:28]
  assign abc_mshr_5_io_bstatus_nestedProbeAckData = bc_mshr_io_status_valid & bc_mshr_io_is_nestedProbeAckData; // @[Slice.scala 218:33]
  assign abc_mshr_5_io_bstatus_probeHelperFinish = bc_mshr_io_status_valid & bc_mshr_io_probeHelperFinish; // @[Slice.scala 220:33]
  assign abc_mshr_5_io_releaseThrough = 1'h0; // @[Slice.scala 221:30]
  assign abc_mshr_5_io_probeAckDataThrough = 1'h0; // @[Slice.scala 222:35]
  assign abc_mshr_6_clock = clock;
  assign abc_mshr_6_reset = reset;
  assign abc_mshr_6_io_id = 4'h6; // @[Slice.scala 166:18]
  assign abc_mshr_6_io_enable = ~(bc_disable_6 | c_disable_6); // @[Slice.scala 198:25]
  assign abc_mshr_6_io_alloc_valid = mshrAlloc_io_alloc_6_valid; // @[Slice.scala 167:21]
  assign abc_mshr_6_io_alloc_bits_channel = mshrAlloc_io_alloc_6_bits_channel; // @[Slice.scala 167:21]
  assign abc_mshr_6_io_alloc_bits_opcode = mshrAlloc_io_alloc_6_bits_opcode; // @[Slice.scala 167:21]
  assign abc_mshr_6_io_alloc_bits_param = mshrAlloc_io_alloc_6_bits_param; // @[Slice.scala 167:21]
  assign abc_mshr_6_io_alloc_bits_size = mshrAlloc_io_alloc_6_bits_size; // @[Slice.scala 167:21]
  assign abc_mshr_6_io_alloc_bits_source = mshrAlloc_io_alloc_6_bits_source; // @[Slice.scala 167:21]
  assign abc_mshr_6_io_alloc_bits_set = mshrAlloc_io_alloc_6_bits_set; // @[Slice.scala 167:21]
  assign abc_mshr_6_io_alloc_bits_tag = mshrAlloc_io_alloc_6_bits_tag; // @[Slice.scala 167:21]
  assign abc_mshr_6_io_alloc_bits_off = mshrAlloc_io_alloc_6_bits_off; // @[Slice.scala 167:21]
  assign abc_mshr_6_io_alloc_bits_mask = mshrAlloc_io_alloc_6_bits_mask; // @[Slice.scala 167:21]
  assign abc_mshr_6_io_alloc_bits_bufIdx = mshrAlloc_io_alloc_6_bits_bufIdx; // @[Slice.scala 167:21]
  assign abc_mshr_6_io_alloc_bits_preferCache = mshrAlloc_io_alloc_6_bits_preferCache; // @[Slice.scala 167:21]
  assign abc_mshr_6_io_alloc_bits_dirty = mshrAlloc_io_alloc_6_bits_dirty; // @[Slice.scala 167:21]
  assign abc_mshr_6_io_alloc_bits_fromProbeHelper = mshrAlloc_io_alloc_6_bits_fromProbeHelper; // @[Slice.scala 167:21]
  assign abc_mshr_6_io_alloc_bits_fromCmoHelper = mshrAlloc_io_alloc_6_bits_fromCmoHelper; // @[Slice.scala 167:21]
  assign abc_mshr_6_io_alloc_bits_needProbeAckData = mshrAlloc_io_alloc_6_bits_needProbeAckData; // @[Slice.scala 167:21]
  assign abc_mshr_6_io_resps_sink_c_valid = sinkC_io_resp_valid & sinkC_io_resp_bits_set ==
    abc_mshr_6_io_status_bits_set; // @[Slice.scala 527:57]
  assign abc_mshr_6_io_resps_sink_c_bits_hasData = sinkC_io_resp_bits_hasData; // @[Slice.scala 531:33]
  assign abc_mshr_6_io_resps_sink_c_bits_param = sinkC_io_resp_bits_param; // @[Slice.scala 531:33]
  assign abc_mshr_6_io_resps_sink_c_bits_source = sinkC_io_resp_bits_source; // @[Slice.scala 531:33]
  assign abc_mshr_6_io_resps_sink_c_bits_last = sinkC_io_resp_bits_last; // @[Slice.scala 531:33]
  assign abc_mshr_6_io_resps_sink_c_bits_bufIdx = sinkC_io_resp_bits_bufIdx; // @[Slice.scala 531:33]
  assign abc_mshr_6_io_resps_sink_d_valid = sinkD_io_resp_valid & sinkD_io_resp_bits_source == 4'h6; // @[Slice.scala 528:57]
  assign abc_mshr_6_io_resps_sink_d_bits_opcode = sinkD_io_resp_bits_opcode; // @[Slice.scala 532:33]
  assign abc_mshr_6_io_resps_sink_d_bits_param = sinkD_io_resp_bits_param; // @[Slice.scala 532:33]
  assign abc_mshr_6_io_resps_sink_d_bits_sink = sinkD_io_resp_bits_sink; // @[Slice.scala 532:33]
  assign abc_mshr_6_io_resps_sink_d_bits_last = sinkD_io_resp_bits_last; // @[Slice.scala 532:33]
  assign abc_mshr_6_io_resps_sink_d_bits_denied = sinkD_io_resp_bits_denied; // @[Slice.scala 532:33]
  assign abc_mshr_6_io_resps_sink_d_bits_bufIdx = sinkD_io_resp_bits_bufIdx; // @[Slice.scala 532:33]
  assign abc_mshr_6_io_resps_sink_e_valid = sinkE_io_resp_valid & sinkE_io_resp_bits_sink == 4'h6; // @[Slice.scala 529:57]
  assign abc_mshr_6_io_resps_source_d_valid = sourceD_io_resp_valid & sourceD_io_resp_bits_sink == 4'h6; // @[Slice.scala 530:61]
  assign abc_mshr_6_io_nestedwb_set = c_mshr_io_status_valid ? c_mshr_io_status_bits_set : bc_mshr_io_status_bits_set; // @[Slice.scala 258:22]
  assign abc_mshr_6_io_nestedwb_tag = c_mshr_io_status_valid ? c_mshr_io_status_bits_tag : bc_mshr_io_status_bits_tag; // @[Slice.scala 259:22]
  assign abc_mshr_6_io_nestedwb_btoN = _nestedWb_btoN_T_2 & _nestedWb_btoN_T_3; // @[Slice.scala 280:38]
  assign abc_mshr_6_io_nestedwb_btoB = _nestedWb_btoN_T_2 & _nestedWb_btoB_T_3; // @[Slice.scala 283:38]
  assign abc_mshr_6_io_nestedwb_bclr_dirty = _nestedWb_btoN_T_2 & _nestedWb_bclr_dirty_T_4; // @[Slice.scala 286:38]
  assign abc_mshr_6_io_nestedwb_bset_dirty = _nestedWb_btoN_T_2 & bc_mshr_io_tasks_dir_write_bits_data_dirty; // @[Slice.scala 289:38]
  assign abc_mshr_6_io_nestedwb_c_set_dirty = _nestedWb_c_set_dirty_T & c_mshr_io_tasks_dir_write_bits_data_dirty; // @[Slice.scala 292:37]
  assign abc_mshr_6_io_nestedwb_c_set_hit = c_mshr_io_status_valid & c_mshr_io_tasks_tag_write_valid &
    _nestedWb_c_set_hit_T_13; // @[Slice.scala 304:50]
  assign abc_mshr_6_io_nestedwb_clients_0_isToN = c_mshr_io_status_valid ? _nestedWb_clients_0_isToN_T_1 :
    _nestedWb_clients_0_isToN_T_3; // @[Slice.scala 314:25]
  assign abc_mshr_6_io_nestedwb_clients_1_isToN = c_mshr_io_status_valid ? _nestedWb_clients_1_isToN_T_1 :
    _nestedWb_clients_1_isToN_T_3; // @[Slice.scala 314:25]
  assign abc_mshr_6_io_tasks_sink_a_ready = 1'h0; // @[Slice.scala 472:13]
  assign abc_mshr_6_io_tasks_source_bready = sourceB_task_arb_io_in_6_ready; // @[Slice.scala 472:13]
  assign abc_mshr_6_io_tasks_sink_c_ready = sinkC_task_arb_io_in_6_ready; // @[Slice.scala 472:13]
  assign abc_mshr_6_io_tasks_source_d_ready = sourceD_task_arb_io_in_6_ready; // @[Slice.scala 472:13]
  assign abc_mshr_6_io_tasks_source_a_ready = sourceA_task_arb_io_in_6_ready; // @[Slice.scala 472:13]
  assign abc_mshr_6_io_tasks_source_c_ready = sourceC_task_arb_io_in_6_ready; // @[Slice.scala 472:13]
  assign abc_mshr_6_io_tasks_source_e_ready = sourceE_task_arb_io_in_6_ready; // @[Slice.scala 472:13]
  assign abc_mshr_6_io_tasks_dir_write_ready = arbiter_io_in_6_ready; // @[Slice.scala 406:60]
  assign abc_mshr_6_io_tasks_tag_write_ready = tagWrite_task_arb_io_in_6_ready; // @[Slice.scala 472:13]
  assign abc_mshr_6_io_tasks_client_dir_write_ready = arbiter_1_io_in_6_ready; // @[Slice.scala 406:60]
  assign abc_mshr_6_io_tasks_client_tag_write_ready = arbiter_2_io_in_6_ready; // @[Slice.scala 472:13]
  assign abc_mshr_6_io_dirResult_valid = ms_6_io_dirResult_valid_REG; // @[Slice.scala 556:31]
  assign abc_mshr_6_io_dirResult_bits_self_dirty = directory_io_result_bits_self_dirty; // @[Slice.scala 555:30]
  assign abc_mshr_6_io_dirResult_bits_self_state = directory_io_result_bits_self_state; // @[Slice.scala 555:30]
  assign abc_mshr_6_io_dirResult_bits_self_clientStates_0 = directory_io_result_bits_self_clientStates_0; // @[Slice.scala 555:30]
  assign abc_mshr_6_io_dirResult_bits_self_clientStates_1 = directory_io_result_bits_self_clientStates_1; // @[Slice.scala 555:30]
  assign abc_mshr_6_io_dirResult_bits_self_hit = directory_io_result_bits_self_hit; // @[Slice.scala 555:30]
  assign abc_mshr_6_io_dirResult_bits_self_way = directory_io_result_bits_self_way; // @[Slice.scala 555:30]
  assign abc_mshr_6_io_dirResult_bits_self_tag = directory_io_result_bits_self_tag; // @[Slice.scala 555:30]
  assign abc_mshr_6_io_dirResult_bits_clients_states_0_state = directory_io_result_bits_clients_states_0_state; // @[Slice.scala 555:30]
  assign abc_mshr_6_io_dirResult_bits_clients_states_0_hit = directory_io_result_bits_clients_states_0_hit; // @[Slice.scala 555:30]
  assign abc_mshr_6_io_dirResult_bits_clients_states_1_state = directory_io_result_bits_clients_states_1_state; // @[Slice.scala 555:30]
  assign abc_mshr_6_io_dirResult_bits_clients_states_1_hit = directory_io_result_bits_clients_states_1_hit; // @[Slice.scala 555:30]
  assign abc_mshr_6_io_dirResult_bits_clients_tag = directory_io_result_bits_clients_tag; // @[Slice.scala 555:30]
  assign abc_mshr_6_io_dirResult_bits_clients_way = directory_io_result_bits_clients_way; // @[Slice.scala 555:30]
  assign abc_mshr_6_io_c_status_set = c_mshr_io_status_bits_set; // @[Slice.scala 209:28]
  assign abc_mshr_6_io_c_status_tag = c_mshr_io_status_bits_tag; // @[Slice.scala 210:28]
  assign abc_mshr_6_io_c_status_way = c_mshr_io_status_bits_way; // @[Slice.scala 211:28]
  assign abc_mshr_6_io_c_status_nestedReleaseData = c_mshr_io_status_valid & c_mshr_io_is_nestedReleaseData; // @[Slice.scala 213:32]
  assign abc_mshr_6_io_bstatus_set = bc_mshr_io_status_bits_set; // @[Slice.scala 214:28]
  assign abc_mshr_6_io_bstatus_tag = bc_mshr_io_status_bits_tag; // @[Slice.scala 215:28]
  assign abc_mshr_6_io_bstatus_way = bc_mshr_io_status_bits_way; // @[Slice.scala 216:28]
  assign abc_mshr_6_io_bstatus_nestedProbeAckData = bc_mshr_io_status_valid & bc_mshr_io_is_nestedProbeAckData; // @[Slice.scala 218:33]
  assign abc_mshr_6_io_bstatus_probeHelperFinish = bc_mshr_io_status_valid & bc_mshr_io_probeHelperFinish; // @[Slice.scala 220:33]
  assign abc_mshr_6_io_releaseThrough = 1'h0; // @[Slice.scala 221:30]
  assign abc_mshr_6_io_probeAckDataThrough = 1'h0; // @[Slice.scala 222:35]
  assign abc_mshr_7_clock = clock;
  assign abc_mshr_7_reset = reset;
  assign abc_mshr_7_io_id = 4'h7; // @[Slice.scala 166:18]
  assign abc_mshr_7_io_enable = ~(bc_disable_7 | c_disable_7); // @[Slice.scala 198:25]
  assign abc_mshr_7_io_alloc_valid = mshrAlloc_io_alloc_7_valid; // @[Slice.scala 167:21]
  assign abc_mshr_7_io_alloc_bits_channel = mshrAlloc_io_alloc_7_bits_channel; // @[Slice.scala 167:21]
  assign abc_mshr_7_io_alloc_bits_opcode = mshrAlloc_io_alloc_7_bits_opcode; // @[Slice.scala 167:21]
  assign abc_mshr_7_io_alloc_bits_param = mshrAlloc_io_alloc_7_bits_param; // @[Slice.scala 167:21]
  assign abc_mshr_7_io_alloc_bits_size = mshrAlloc_io_alloc_7_bits_size; // @[Slice.scala 167:21]
  assign abc_mshr_7_io_alloc_bits_source = mshrAlloc_io_alloc_7_bits_source; // @[Slice.scala 167:21]
  assign abc_mshr_7_io_alloc_bits_set = mshrAlloc_io_alloc_7_bits_set; // @[Slice.scala 167:21]
  assign abc_mshr_7_io_alloc_bits_tag = mshrAlloc_io_alloc_7_bits_tag; // @[Slice.scala 167:21]
  assign abc_mshr_7_io_alloc_bits_off = mshrAlloc_io_alloc_7_bits_off; // @[Slice.scala 167:21]
  assign abc_mshr_7_io_alloc_bits_mask = mshrAlloc_io_alloc_7_bits_mask; // @[Slice.scala 167:21]
  assign abc_mshr_7_io_alloc_bits_bufIdx = mshrAlloc_io_alloc_7_bits_bufIdx; // @[Slice.scala 167:21]
  assign abc_mshr_7_io_alloc_bits_preferCache = mshrAlloc_io_alloc_7_bits_preferCache; // @[Slice.scala 167:21]
  assign abc_mshr_7_io_alloc_bits_dirty = mshrAlloc_io_alloc_7_bits_dirty; // @[Slice.scala 167:21]
  assign abc_mshr_7_io_alloc_bits_fromProbeHelper = mshrAlloc_io_alloc_7_bits_fromProbeHelper; // @[Slice.scala 167:21]
  assign abc_mshr_7_io_alloc_bits_fromCmoHelper = mshrAlloc_io_alloc_7_bits_fromCmoHelper; // @[Slice.scala 167:21]
  assign abc_mshr_7_io_alloc_bits_needProbeAckData = mshrAlloc_io_alloc_7_bits_needProbeAckData; // @[Slice.scala 167:21]
  assign abc_mshr_7_io_resps_sink_c_valid = sinkC_io_resp_valid & sinkC_io_resp_bits_set ==
    abc_mshr_7_io_status_bits_set; // @[Slice.scala 527:57]
  assign abc_mshr_7_io_resps_sink_c_bits_hasData = sinkC_io_resp_bits_hasData; // @[Slice.scala 531:33]
  assign abc_mshr_7_io_resps_sink_c_bits_param = sinkC_io_resp_bits_param; // @[Slice.scala 531:33]
  assign abc_mshr_7_io_resps_sink_c_bits_source = sinkC_io_resp_bits_source; // @[Slice.scala 531:33]
  assign abc_mshr_7_io_resps_sink_c_bits_last = sinkC_io_resp_bits_last; // @[Slice.scala 531:33]
  assign abc_mshr_7_io_resps_sink_c_bits_bufIdx = sinkC_io_resp_bits_bufIdx; // @[Slice.scala 531:33]
  assign abc_mshr_7_io_resps_sink_d_valid = sinkD_io_resp_valid & sinkD_io_resp_bits_source == 4'h7; // @[Slice.scala 528:57]
  assign abc_mshr_7_io_resps_sink_d_bits_opcode = sinkD_io_resp_bits_opcode; // @[Slice.scala 532:33]
  assign abc_mshr_7_io_resps_sink_d_bits_param = sinkD_io_resp_bits_param; // @[Slice.scala 532:33]
  assign abc_mshr_7_io_resps_sink_d_bits_sink = sinkD_io_resp_bits_sink; // @[Slice.scala 532:33]
  assign abc_mshr_7_io_resps_sink_d_bits_last = sinkD_io_resp_bits_last; // @[Slice.scala 532:33]
  assign abc_mshr_7_io_resps_sink_d_bits_denied = sinkD_io_resp_bits_denied; // @[Slice.scala 532:33]
  assign abc_mshr_7_io_resps_sink_d_bits_bufIdx = sinkD_io_resp_bits_bufIdx; // @[Slice.scala 532:33]
  assign abc_mshr_7_io_resps_sink_e_valid = sinkE_io_resp_valid & sinkE_io_resp_bits_sink == 4'h7; // @[Slice.scala 529:57]
  assign abc_mshr_7_io_resps_source_d_valid = sourceD_io_resp_valid & sourceD_io_resp_bits_sink == 4'h7; // @[Slice.scala 530:61]
  assign abc_mshr_7_io_nestedwb_set = c_mshr_io_status_valid ? c_mshr_io_status_bits_set : bc_mshr_io_status_bits_set; // @[Slice.scala 258:22]
  assign abc_mshr_7_io_nestedwb_tag = c_mshr_io_status_valid ? c_mshr_io_status_bits_tag : bc_mshr_io_status_bits_tag; // @[Slice.scala 259:22]
  assign abc_mshr_7_io_nestedwb_btoN = _nestedWb_btoN_T_2 & _nestedWb_btoN_T_3; // @[Slice.scala 280:38]
  assign abc_mshr_7_io_nestedwb_btoB = _nestedWb_btoN_T_2 & _nestedWb_btoB_T_3; // @[Slice.scala 283:38]
  assign abc_mshr_7_io_nestedwb_bclr_dirty = _nestedWb_btoN_T_2 & _nestedWb_bclr_dirty_T_4; // @[Slice.scala 286:38]
  assign abc_mshr_7_io_nestedwb_bset_dirty = _nestedWb_btoN_T_2 & bc_mshr_io_tasks_dir_write_bits_data_dirty; // @[Slice.scala 289:38]
  assign abc_mshr_7_io_nestedwb_c_set_dirty = _nestedWb_c_set_dirty_T & c_mshr_io_tasks_dir_write_bits_data_dirty; // @[Slice.scala 292:37]
  assign abc_mshr_7_io_nestedwb_c_set_hit = c_mshr_io_status_valid & c_mshr_io_tasks_tag_write_valid &
    _nestedWb_c_set_hit_T_15; // @[Slice.scala 304:50]
  assign abc_mshr_7_io_nestedwb_clients_0_isToN = c_mshr_io_status_valid ? _nestedWb_clients_0_isToN_T_1 :
    _nestedWb_clients_0_isToN_T_3; // @[Slice.scala 314:25]
  assign abc_mshr_7_io_nestedwb_clients_1_isToN = c_mshr_io_status_valid ? _nestedWb_clients_1_isToN_T_1 :
    _nestedWb_clients_1_isToN_T_3; // @[Slice.scala 314:25]
  assign abc_mshr_7_io_tasks_sink_a_ready = 1'h0; // @[Slice.scala 472:13]
  assign abc_mshr_7_io_tasks_source_bready = sourceB_task_arb_io_in_7_ready; // @[Slice.scala 472:13]
  assign abc_mshr_7_io_tasks_sink_c_ready = sinkC_task_arb_io_in_7_ready; // @[Slice.scala 472:13]
  assign abc_mshr_7_io_tasks_source_d_ready = sourceD_task_arb_io_in_7_ready; // @[Slice.scala 472:13]
  assign abc_mshr_7_io_tasks_source_a_ready = sourceA_task_arb_io_in_7_ready; // @[Slice.scala 472:13]
  assign abc_mshr_7_io_tasks_source_c_ready = sourceC_task_arb_io_in_7_ready; // @[Slice.scala 472:13]
  assign abc_mshr_7_io_tasks_source_e_ready = sourceE_task_arb_io_in_7_ready; // @[Slice.scala 472:13]
  assign abc_mshr_7_io_tasks_dir_write_ready = arbiter_io_in_7_ready; // @[Slice.scala 406:60]
  assign abc_mshr_7_io_tasks_tag_write_ready = tagWrite_task_arb_io_in_7_ready; // @[Slice.scala 472:13]
  assign abc_mshr_7_io_tasks_client_dir_write_ready = arbiter_1_io_in_7_ready; // @[Slice.scala 406:60]
  assign abc_mshr_7_io_tasks_client_tag_write_ready = arbiter_2_io_in_7_ready; // @[Slice.scala 472:13]
  assign abc_mshr_7_io_dirResult_valid = ms_7_io_dirResult_valid_REG; // @[Slice.scala 556:31]
  assign abc_mshr_7_io_dirResult_bits_self_dirty = directory_io_result_bits_self_dirty; // @[Slice.scala 555:30]
  assign abc_mshr_7_io_dirResult_bits_self_state = directory_io_result_bits_self_state; // @[Slice.scala 555:30]
  assign abc_mshr_7_io_dirResult_bits_self_clientStates_0 = directory_io_result_bits_self_clientStates_0; // @[Slice.scala 555:30]
  assign abc_mshr_7_io_dirResult_bits_self_clientStates_1 = directory_io_result_bits_self_clientStates_1; // @[Slice.scala 555:30]
  assign abc_mshr_7_io_dirResult_bits_self_hit = directory_io_result_bits_self_hit; // @[Slice.scala 555:30]
  assign abc_mshr_7_io_dirResult_bits_self_way = directory_io_result_bits_self_way; // @[Slice.scala 555:30]
  assign abc_mshr_7_io_dirResult_bits_self_tag = directory_io_result_bits_self_tag; // @[Slice.scala 555:30]
  assign abc_mshr_7_io_dirResult_bits_clients_states_0_state = directory_io_result_bits_clients_states_0_state; // @[Slice.scala 555:30]
  assign abc_mshr_7_io_dirResult_bits_clients_states_0_hit = directory_io_result_bits_clients_states_0_hit; // @[Slice.scala 555:30]
  assign abc_mshr_7_io_dirResult_bits_clients_states_1_state = directory_io_result_bits_clients_states_1_state; // @[Slice.scala 555:30]
  assign abc_mshr_7_io_dirResult_bits_clients_states_1_hit = directory_io_result_bits_clients_states_1_hit; // @[Slice.scala 555:30]
  assign abc_mshr_7_io_dirResult_bits_clients_tag = directory_io_result_bits_clients_tag; // @[Slice.scala 555:30]
  assign abc_mshr_7_io_dirResult_bits_clients_way = directory_io_result_bits_clients_way; // @[Slice.scala 555:30]
  assign abc_mshr_7_io_c_status_set = c_mshr_io_status_bits_set; // @[Slice.scala 209:28]
  assign abc_mshr_7_io_c_status_tag = c_mshr_io_status_bits_tag; // @[Slice.scala 210:28]
  assign abc_mshr_7_io_c_status_way = c_mshr_io_status_bits_way; // @[Slice.scala 211:28]
  assign abc_mshr_7_io_c_status_nestedReleaseData = c_mshr_io_status_valid & c_mshr_io_is_nestedReleaseData; // @[Slice.scala 213:32]
  assign abc_mshr_7_io_bstatus_set = bc_mshr_io_status_bits_set; // @[Slice.scala 214:28]
  assign abc_mshr_7_io_bstatus_tag = bc_mshr_io_status_bits_tag; // @[Slice.scala 215:28]
  assign abc_mshr_7_io_bstatus_way = bc_mshr_io_status_bits_way; // @[Slice.scala 216:28]
  assign abc_mshr_7_io_bstatus_nestedProbeAckData = bc_mshr_io_status_valid & bc_mshr_io_is_nestedProbeAckData; // @[Slice.scala 218:33]
  assign abc_mshr_7_io_bstatus_probeHelperFinish = bc_mshr_io_status_valid & bc_mshr_io_probeHelperFinish; // @[Slice.scala 220:33]
  assign abc_mshr_7_io_releaseThrough = 1'h0; // @[Slice.scala 221:30]
  assign abc_mshr_7_io_probeAckDataThrough = 1'h0; // @[Slice.scala 222:35]
  assign abc_mshr_8_clock = clock;
  assign abc_mshr_8_reset = reset;
  assign abc_mshr_8_io_id = 4'h8; // @[Slice.scala 166:18]
  assign abc_mshr_8_io_enable = ~(bc_disable_8 | c_disable_8); // @[Slice.scala 198:25]
  assign abc_mshr_8_io_alloc_valid = mshrAlloc_io_alloc_8_valid; // @[Slice.scala 167:21]
  assign abc_mshr_8_io_alloc_bits_channel = mshrAlloc_io_alloc_8_bits_channel; // @[Slice.scala 167:21]
  assign abc_mshr_8_io_alloc_bits_opcode = mshrAlloc_io_alloc_8_bits_opcode; // @[Slice.scala 167:21]
  assign abc_mshr_8_io_alloc_bits_param = mshrAlloc_io_alloc_8_bits_param; // @[Slice.scala 167:21]
  assign abc_mshr_8_io_alloc_bits_size = mshrAlloc_io_alloc_8_bits_size; // @[Slice.scala 167:21]
  assign abc_mshr_8_io_alloc_bits_source = mshrAlloc_io_alloc_8_bits_source; // @[Slice.scala 167:21]
  assign abc_mshr_8_io_alloc_bits_set = mshrAlloc_io_alloc_8_bits_set; // @[Slice.scala 167:21]
  assign abc_mshr_8_io_alloc_bits_tag = mshrAlloc_io_alloc_8_bits_tag; // @[Slice.scala 167:21]
  assign abc_mshr_8_io_alloc_bits_off = mshrAlloc_io_alloc_8_bits_off; // @[Slice.scala 167:21]
  assign abc_mshr_8_io_alloc_bits_mask = mshrAlloc_io_alloc_8_bits_mask; // @[Slice.scala 167:21]
  assign abc_mshr_8_io_alloc_bits_bufIdx = mshrAlloc_io_alloc_8_bits_bufIdx; // @[Slice.scala 167:21]
  assign abc_mshr_8_io_alloc_bits_preferCache = mshrAlloc_io_alloc_8_bits_preferCache; // @[Slice.scala 167:21]
  assign abc_mshr_8_io_alloc_bits_dirty = mshrAlloc_io_alloc_8_bits_dirty; // @[Slice.scala 167:21]
  assign abc_mshr_8_io_alloc_bits_fromProbeHelper = mshrAlloc_io_alloc_8_bits_fromProbeHelper; // @[Slice.scala 167:21]
  assign abc_mshr_8_io_alloc_bits_fromCmoHelper = mshrAlloc_io_alloc_8_bits_fromCmoHelper; // @[Slice.scala 167:21]
  assign abc_mshr_8_io_alloc_bits_needProbeAckData = mshrAlloc_io_alloc_8_bits_needProbeAckData; // @[Slice.scala 167:21]
  assign abc_mshr_8_io_resps_sink_c_valid = sinkC_io_resp_valid & sinkC_io_resp_bits_set ==
    abc_mshr_8_io_status_bits_set; // @[Slice.scala 527:57]
  assign abc_mshr_8_io_resps_sink_c_bits_hasData = sinkC_io_resp_bits_hasData; // @[Slice.scala 531:33]
  assign abc_mshr_8_io_resps_sink_c_bits_param = sinkC_io_resp_bits_param; // @[Slice.scala 531:33]
  assign abc_mshr_8_io_resps_sink_c_bits_source = sinkC_io_resp_bits_source; // @[Slice.scala 531:33]
  assign abc_mshr_8_io_resps_sink_c_bits_last = sinkC_io_resp_bits_last; // @[Slice.scala 531:33]
  assign abc_mshr_8_io_resps_sink_c_bits_bufIdx = sinkC_io_resp_bits_bufIdx; // @[Slice.scala 531:33]
  assign abc_mshr_8_io_resps_sink_d_valid = sinkD_io_resp_valid & sinkD_io_resp_bits_source == 4'h8; // @[Slice.scala 528:57]
  assign abc_mshr_8_io_resps_sink_d_bits_opcode = sinkD_io_resp_bits_opcode; // @[Slice.scala 532:33]
  assign abc_mshr_8_io_resps_sink_d_bits_param = sinkD_io_resp_bits_param; // @[Slice.scala 532:33]
  assign abc_mshr_8_io_resps_sink_d_bits_sink = sinkD_io_resp_bits_sink; // @[Slice.scala 532:33]
  assign abc_mshr_8_io_resps_sink_d_bits_last = sinkD_io_resp_bits_last; // @[Slice.scala 532:33]
  assign abc_mshr_8_io_resps_sink_d_bits_denied = sinkD_io_resp_bits_denied; // @[Slice.scala 532:33]
  assign abc_mshr_8_io_resps_sink_d_bits_bufIdx = sinkD_io_resp_bits_bufIdx; // @[Slice.scala 532:33]
  assign abc_mshr_8_io_resps_sink_e_valid = sinkE_io_resp_valid & sinkE_io_resp_bits_sink == 4'h8; // @[Slice.scala 529:57]
  assign abc_mshr_8_io_resps_source_d_valid = sourceD_io_resp_valid & sourceD_io_resp_bits_sink == 4'h8; // @[Slice.scala 530:61]
  assign abc_mshr_8_io_nestedwb_set = c_mshr_io_status_valid ? c_mshr_io_status_bits_set : bc_mshr_io_status_bits_set; // @[Slice.scala 258:22]
  assign abc_mshr_8_io_nestedwb_tag = c_mshr_io_status_valid ? c_mshr_io_status_bits_tag : bc_mshr_io_status_bits_tag; // @[Slice.scala 259:22]
  assign abc_mshr_8_io_nestedwb_btoN = _nestedWb_btoN_T_2 & _nestedWb_btoN_T_3; // @[Slice.scala 280:38]
  assign abc_mshr_8_io_nestedwb_btoB = _nestedWb_btoN_T_2 & _nestedWb_btoB_T_3; // @[Slice.scala 283:38]
  assign abc_mshr_8_io_nestedwb_bclr_dirty = _nestedWb_btoN_T_2 & _nestedWb_bclr_dirty_T_4; // @[Slice.scala 286:38]
  assign abc_mshr_8_io_nestedwb_bset_dirty = _nestedWb_btoN_T_2 & bc_mshr_io_tasks_dir_write_bits_data_dirty; // @[Slice.scala 289:38]
  assign abc_mshr_8_io_nestedwb_c_set_dirty = _nestedWb_c_set_dirty_T & c_mshr_io_tasks_dir_write_bits_data_dirty; // @[Slice.scala 292:37]
  assign abc_mshr_8_io_nestedwb_c_set_hit = c_mshr_io_status_valid & c_mshr_io_tasks_tag_write_valid &
    _nestedWb_c_set_hit_T_17; // @[Slice.scala 304:50]
  assign abc_mshr_8_io_nestedwb_clients_0_isToN = c_mshr_io_status_valid ? _nestedWb_clients_0_isToN_T_1 :
    _nestedWb_clients_0_isToN_T_3; // @[Slice.scala 314:25]
  assign abc_mshr_8_io_nestedwb_clients_1_isToN = c_mshr_io_status_valid ? _nestedWb_clients_1_isToN_T_1 :
    _nestedWb_clients_1_isToN_T_3; // @[Slice.scala 314:25]
  assign abc_mshr_8_io_tasks_sink_a_ready = 1'h0; // @[Slice.scala 472:13]
  assign abc_mshr_8_io_tasks_source_bready = sourceB_task_arb_io_in_8_ready; // @[Slice.scala 472:13]
  assign abc_mshr_8_io_tasks_sink_c_ready = sinkC_task_arb_io_in_8_ready; // @[Slice.scala 472:13]
  assign abc_mshr_8_io_tasks_source_d_ready = sourceD_task_arb_io_in_8_ready; // @[Slice.scala 472:13]
  assign abc_mshr_8_io_tasks_source_a_ready = sourceA_task_arb_io_in_8_ready; // @[Slice.scala 472:13]
  assign abc_mshr_8_io_tasks_source_c_ready = sourceC_task_arb_io_in_8_ready; // @[Slice.scala 472:13]
  assign abc_mshr_8_io_tasks_source_e_ready = sourceE_task_arb_io_in_8_ready; // @[Slice.scala 472:13]
  assign abc_mshr_8_io_tasks_dir_write_ready = arbiter_io_in_8_ready; // @[Slice.scala 406:60]
  assign abc_mshr_8_io_tasks_tag_write_ready = tagWrite_task_arb_io_in_8_ready; // @[Slice.scala 472:13]
  assign abc_mshr_8_io_tasks_client_dir_write_ready = arbiter_1_io_in_8_ready; // @[Slice.scala 406:60]
  assign abc_mshr_8_io_tasks_client_tag_write_ready = arbiter_2_io_in_8_ready; // @[Slice.scala 472:13]
  assign abc_mshr_8_io_dirResult_valid = ms_8_io_dirResult_valid_REG; // @[Slice.scala 556:31]
  assign abc_mshr_8_io_dirResult_bits_self_dirty = directory_io_result_bits_self_dirty; // @[Slice.scala 555:30]
  assign abc_mshr_8_io_dirResult_bits_self_state = directory_io_result_bits_self_state; // @[Slice.scala 555:30]
  assign abc_mshr_8_io_dirResult_bits_self_clientStates_0 = directory_io_result_bits_self_clientStates_0; // @[Slice.scala 555:30]
  assign abc_mshr_8_io_dirResult_bits_self_clientStates_1 = directory_io_result_bits_self_clientStates_1; // @[Slice.scala 555:30]
  assign abc_mshr_8_io_dirResult_bits_self_hit = directory_io_result_bits_self_hit; // @[Slice.scala 555:30]
  assign abc_mshr_8_io_dirResult_bits_self_way = directory_io_result_bits_self_way; // @[Slice.scala 555:30]
  assign abc_mshr_8_io_dirResult_bits_self_tag = directory_io_result_bits_self_tag; // @[Slice.scala 555:30]
  assign abc_mshr_8_io_dirResult_bits_clients_states_0_state = directory_io_result_bits_clients_states_0_state; // @[Slice.scala 555:30]
  assign abc_mshr_8_io_dirResult_bits_clients_states_0_hit = directory_io_result_bits_clients_states_0_hit; // @[Slice.scala 555:30]
  assign abc_mshr_8_io_dirResult_bits_clients_states_1_state = directory_io_result_bits_clients_states_1_state; // @[Slice.scala 555:30]
  assign abc_mshr_8_io_dirResult_bits_clients_states_1_hit = directory_io_result_bits_clients_states_1_hit; // @[Slice.scala 555:30]
  assign abc_mshr_8_io_dirResult_bits_clients_tag = directory_io_result_bits_clients_tag; // @[Slice.scala 555:30]
  assign abc_mshr_8_io_dirResult_bits_clients_way = directory_io_result_bits_clients_way; // @[Slice.scala 555:30]
  assign abc_mshr_8_io_c_status_set = c_mshr_io_status_bits_set; // @[Slice.scala 209:28]
  assign abc_mshr_8_io_c_status_tag = c_mshr_io_status_bits_tag; // @[Slice.scala 210:28]
  assign abc_mshr_8_io_c_status_way = c_mshr_io_status_bits_way; // @[Slice.scala 211:28]
  assign abc_mshr_8_io_c_status_nestedReleaseData = c_mshr_io_status_valid & c_mshr_io_is_nestedReleaseData; // @[Slice.scala 213:32]
  assign abc_mshr_8_io_bstatus_set = bc_mshr_io_status_bits_set; // @[Slice.scala 214:28]
  assign abc_mshr_8_io_bstatus_tag = bc_mshr_io_status_bits_tag; // @[Slice.scala 215:28]
  assign abc_mshr_8_io_bstatus_way = bc_mshr_io_status_bits_way; // @[Slice.scala 216:28]
  assign abc_mshr_8_io_bstatus_nestedProbeAckData = bc_mshr_io_status_valid & bc_mshr_io_is_nestedProbeAckData; // @[Slice.scala 218:33]
  assign abc_mshr_8_io_bstatus_probeHelperFinish = bc_mshr_io_status_valid & bc_mshr_io_probeHelperFinish; // @[Slice.scala 220:33]
  assign abc_mshr_8_io_releaseThrough = 1'h0; // @[Slice.scala 221:30]
  assign abc_mshr_8_io_probeAckDataThrough = 1'h0; // @[Slice.scala 222:35]
  assign abc_mshr_9_clock = clock;
  assign abc_mshr_9_reset = reset;
  assign abc_mshr_9_io_id = 4'h9; // @[Slice.scala 166:18]
  assign abc_mshr_9_io_enable = ~(bc_disable_9 | c_disable_9); // @[Slice.scala 198:25]
  assign abc_mshr_9_io_alloc_valid = mshrAlloc_io_alloc_9_valid; // @[Slice.scala 167:21]
  assign abc_mshr_9_io_alloc_bits_channel = mshrAlloc_io_alloc_9_bits_channel; // @[Slice.scala 167:21]
  assign abc_mshr_9_io_alloc_bits_opcode = mshrAlloc_io_alloc_9_bits_opcode; // @[Slice.scala 167:21]
  assign abc_mshr_9_io_alloc_bits_param = mshrAlloc_io_alloc_9_bits_param; // @[Slice.scala 167:21]
  assign abc_mshr_9_io_alloc_bits_size = mshrAlloc_io_alloc_9_bits_size; // @[Slice.scala 167:21]
  assign abc_mshr_9_io_alloc_bits_source = mshrAlloc_io_alloc_9_bits_source; // @[Slice.scala 167:21]
  assign abc_mshr_9_io_alloc_bits_set = mshrAlloc_io_alloc_9_bits_set; // @[Slice.scala 167:21]
  assign abc_mshr_9_io_alloc_bits_tag = mshrAlloc_io_alloc_9_bits_tag; // @[Slice.scala 167:21]
  assign abc_mshr_9_io_alloc_bits_off = mshrAlloc_io_alloc_9_bits_off; // @[Slice.scala 167:21]
  assign abc_mshr_9_io_alloc_bits_mask = mshrAlloc_io_alloc_9_bits_mask; // @[Slice.scala 167:21]
  assign abc_mshr_9_io_alloc_bits_bufIdx = mshrAlloc_io_alloc_9_bits_bufIdx; // @[Slice.scala 167:21]
  assign abc_mshr_9_io_alloc_bits_preferCache = mshrAlloc_io_alloc_9_bits_preferCache; // @[Slice.scala 167:21]
  assign abc_mshr_9_io_alloc_bits_dirty = mshrAlloc_io_alloc_9_bits_dirty; // @[Slice.scala 167:21]
  assign abc_mshr_9_io_alloc_bits_fromProbeHelper = mshrAlloc_io_alloc_9_bits_fromProbeHelper; // @[Slice.scala 167:21]
  assign abc_mshr_9_io_alloc_bits_fromCmoHelper = mshrAlloc_io_alloc_9_bits_fromCmoHelper; // @[Slice.scala 167:21]
  assign abc_mshr_9_io_alloc_bits_needProbeAckData = mshrAlloc_io_alloc_9_bits_needProbeAckData; // @[Slice.scala 167:21]
  assign abc_mshr_9_io_resps_sink_c_valid = sinkC_io_resp_valid & sinkC_io_resp_bits_set ==
    abc_mshr_9_io_status_bits_set; // @[Slice.scala 527:57]
  assign abc_mshr_9_io_resps_sink_c_bits_hasData = sinkC_io_resp_bits_hasData; // @[Slice.scala 531:33]
  assign abc_mshr_9_io_resps_sink_c_bits_param = sinkC_io_resp_bits_param; // @[Slice.scala 531:33]
  assign abc_mshr_9_io_resps_sink_c_bits_source = sinkC_io_resp_bits_source; // @[Slice.scala 531:33]
  assign abc_mshr_9_io_resps_sink_c_bits_last = sinkC_io_resp_bits_last; // @[Slice.scala 531:33]
  assign abc_mshr_9_io_resps_sink_c_bits_bufIdx = sinkC_io_resp_bits_bufIdx; // @[Slice.scala 531:33]
  assign abc_mshr_9_io_resps_sink_d_valid = sinkD_io_resp_valid & sinkD_io_resp_bits_source == 4'h9; // @[Slice.scala 528:57]
  assign abc_mshr_9_io_resps_sink_d_bits_opcode = sinkD_io_resp_bits_opcode; // @[Slice.scala 532:33]
  assign abc_mshr_9_io_resps_sink_d_bits_param = sinkD_io_resp_bits_param; // @[Slice.scala 532:33]
  assign abc_mshr_9_io_resps_sink_d_bits_sink = sinkD_io_resp_bits_sink; // @[Slice.scala 532:33]
  assign abc_mshr_9_io_resps_sink_d_bits_last = sinkD_io_resp_bits_last; // @[Slice.scala 532:33]
  assign abc_mshr_9_io_resps_sink_d_bits_denied = sinkD_io_resp_bits_denied; // @[Slice.scala 532:33]
  assign abc_mshr_9_io_resps_sink_d_bits_bufIdx = sinkD_io_resp_bits_bufIdx; // @[Slice.scala 532:33]
  assign abc_mshr_9_io_resps_sink_e_valid = sinkE_io_resp_valid & sinkE_io_resp_bits_sink == 4'h9; // @[Slice.scala 529:57]
  assign abc_mshr_9_io_resps_source_d_valid = sourceD_io_resp_valid & sourceD_io_resp_bits_sink == 4'h9; // @[Slice.scala 530:61]
  assign abc_mshr_9_io_nestedwb_set = c_mshr_io_status_valid ? c_mshr_io_status_bits_set : bc_mshr_io_status_bits_set; // @[Slice.scala 258:22]
  assign abc_mshr_9_io_nestedwb_tag = c_mshr_io_status_valid ? c_mshr_io_status_bits_tag : bc_mshr_io_status_bits_tag; // @[Slice.scala 259:22]
  assign abc_mshr_9_io_nestedwb_btoN = _nestedWb_btoN_T_2 & _nestedWb_btoN_T_3; // @[Slice.scala 280:38]
  assign abc_mshr_9_io_nestedwb_btoB = _nestedWb_btoN_T_2 & _nestedWb_btoB_T_3; // @[Slice.scala 283:38]
  assign abc_mshr_9_io_nestedwb_bclr_dirty = _nestedWb_btoN_T_2 & _nestedWb_bclr_dirty_T_4; // @[Slice.scala 286:38]
  assign abc_mshr_9_io_nestedwb_bset_dirty = _nestedWb_btoN_T_2 & bc_mshr_io_tasks_dir_write_bits_data_dirty; // @[Slice.scala 289:38]
  assign abc_mshr_9_io_nestedwb_c_set_dirty = _nestedWb_c_set_dirty_T & c_mshr_io_tasks_dir_write_bits_data_dirty; // @[Slice.scala 292:37]
  assign abc_mshr_9_io_nestedwb_c_set_hit = c_mshr_io_status_valid & c_mshr_io_tasks_tag_write_valid &
    _nestedWb_c_set_hit_T_19; // @[Slice.scala 304:50]
  assign abc_mshr_9_io_nestedwb_clients_0_isToN = c_mshr_io_status_valid ? _nestedWb_clients_0_isToN_T_1 :
    _nestedWb_clients_0_isToN_T_3; // @[Slice.scala 314:25]
  assign abc_mshr_9_io_nestedwb_clients_1_isToN = c_mshr_io_status_valid ? _nestedWb_clients_1_isToN_T_1 :
    _nestedWb_clients_1_isToN_T_3; // @[Slice.scala 314:25]
  assign abc_mshr_9_io_tasks_sink_a_ready = 1'h0; // @[Slice.scala 472:13]
  assign abc_mshr_9_io_tasks_source_bready = sourceB_task_arb_io_in_9_ready; // @[Slice.scala 472:13]
  assign abc_mshr_9_io_tasks_sink_c_ready = sinkC_task_arb_io_in_9_ready; // @[Slice.scala 472:13]
  assign abc_mshr_9_io_tasks_source_d_ready = sourceD_task_arb_io_in_9_ready; // @[Slice.scala 472:13]
  assign abc_mshr_9_io_tasks_source_a_ready = sourceA_task_arb_io_in_9_ready; // @[Slice.scala 472:13]
  assign abc_mshr_9_io_tasks_source_c_ready = sourceC_task_arb_io_in_9_ready; // @[Slice.scala 472:13]
  assign abc_mshr_9_io_tasks_source_e_ready = sourceE_task_arb_io_in_9_ready; // @[Slice.scala 472:13]
  assign abc_mshr_9_io_tasks_dir_write_ready = arbiter_io_in_9_ready; // @[Slice.scala 406:60]
  assign abc_mshr_9_io_tasks_tag_write_ready = tagWrite_task_arb_io_in_9_ready; // @[Slice.scala 472:13]
  assign abc_mshr_9_io_tasks_client_dir_write_ready = arbiter_1_io_in_9_ready; // @[Slice.scala 406:60]
  assign abc_mshr_9_io_tasks_client_tag_write_ready = arbiter_2_io_in_9_ready; // @[Slice.scala 472:13]
  assign abc_mshr_9_io_dirResult_valid = ms_9_io_dirResult_valid_REG; // @[Slice.scala 556:31]
  assign abc_mshr_9_io_dirResult_bits_self_dirty = directory_io_result_bits_self_dirty; // @[Slice.scala 555:30]
  assign abc_mshr_9_io_dirResult_bits_self_state = directory_io_result_bits_self_state; // @[Slice.scala 555:30]
  assign abc_mshr_9_io_dirResult_bits_self_clientStates_0 = directory_io_result_bits_self_clientStates_0; // @[Slice.scala 555:30]
  assign abc_mshr_9_io_dirResult_bits_self_clientStates_1 = directory_io_result_bits_self_clientStates_1; // @[Slice.scala 555:30]
  assign abc_mshr_9_io_dirResult_bits_self_hit = directory_io_result_bits_self_hit; // @[Slice.scala 555:30]
  assign abc_mshr_9_io_dirResult_bits_self_way = directory_io_result_bits_self_way; // @[Slice.scala 555:30]
  assign abc_mshr_9_io_dirResult_bits_self_tag = directory_io_result_bits_self_tag; // @[Slice.scala 555:30]
  assign abc_mshr_9_io_dirResult_bits_clients_states_0_state = directory_io_result_bits_clients_states_0_state; // @[Slice.scala 555:30]
  assign abc_mshr_9_io_dirResult_bits_clients_states_0_hit = directory_io_result_bits_clients_states_0_hit; // @[Slice.scala 555:30]
  assign abc_mshr_9_io_dirResult_bits_clients_states_1_state = directory_io_result_bits_clients_states_1_state; // @[Slice.scala 555:30]
  assign abc_mshr_9_io_dirResult_bits_clients_states_1_hit = directory_io_result_bits_clients_states_1_hit; // @[Slice.scala 555:30]
  assign abc_mshr_9_io_dirResult_bits_clients_tag = directory_io_result_bits_clients_tag; // @[Slice.scala 555:30]
  assign abc_mshr_9_io_dirResult_bits_clients_way = directory_io_result_bits_clients_way; // @[Slice.scala 555:30]
  assign abc_mshr_9_io_c_status_set = c_mshr_io_status_bits_set; // @[Slice.scala 209:28]
  assign abc_mshr_9_io_c_status_tag = c_mshr_io_status_bits_tag; // @[Slice.scala 210:28]
  assign abc_mshr_9_io_c_status_way = c_mshr_io_status_bits_way; // @[Slice.scala 211:28]
  assign abc_mshr_9_io_c_status_nestedReleaseData = c_mshr_io_status_valid & c_mshr_io_is_nestedReleaseData; // @[Slice.scala 213:32]
  assign abc_mshr_9_io_bstatus_set = bc_mshr_io_status_bits_set; // @[Slice.scala 214:28]
  assign abc_mshr_9_io_bstatus_tag = bc_mshr_io_status_bits_tag; // @[Slice.scala 215:28]
  assign abc_mshr_9_io_bstatus_way = bc_mshr_io_status_bits_way; // @[Slice.scala 216:28]
  assign abc_mshr_9_io_bstatus_nestedProbeAckData = bc_mshr_io_status_valid & bc_mshr_io_is_nestedProbeAckData; // @[Slice.scala 218:33]
  assign abc_mshr_9_io_bstatus_probeHelperFinish = bc_mshr_io_status_valid & bc_mshr_io_probeHelperFinish; // @[Slice.scala 220:33]
  assign abc_mshr_9_io_releaseThrough = 1'h0; // @[Slice.scala 221:30]
  assign abc_mshr_9_io_probeAckDataThrough = 1'h0; // @[Slice.scala 222:35]
  assign abc_mshr_10_clock = clock;
  assign abc_mshr_10_reset = reset;
  assign abc_mshr_10_io_id = 4'ha; // @[Slice.scala 166:18]
  assign abc_mshr_10_io_enable = ~(bc_disable_10 | c_disable_10); // @[Slice.scala 198:25]
  assign abc_mshr_10_io_alloc_valid = mshrAlloc_io_alloc_10_valid; // @[Slice.scala 167:21]
  assign abc_mshr_10_io_alloc_bits_channel = mshrAlloc_io_alloc_10_bits_channel; // @[Slice.scala 167:21]
  assign abc_mshr_10_io_alloc_bits_opcode = mshrAlloc_io_alloc_10_bits_opcode; // @[Slice.scala 167:21]
  assign abc_mshr_10_io_alloc_bits_param = mshrAlloc_io_alloc_10_bits_param; // @[Slice.scala 167:21]
  assign abc_mshr_10_io_alloc_bits_size = mshrAlloc_io_alloc_10_bits_size; // @[Slice.scala 167:21]
  assign abc_mshr_10_io_alloc_bits_source = mshrAlloc_io_alloc_10_bits_source; // @[Slice.scala 167:21]
  assign abc_mshr_10_io_alloc_bits_set = mshrAlloc_io_alloc_10_bits_set; // @[Slice.scala 167:21]
  assign abc_mshr_10_io_alloc_bits_tag = mshrAlloc_io_alloc_10_bits_tag; // @[Slice.scala 167:21]
  assign abc_mshr_10_io_alloc_bits_off = mshrAlloc_io_alloc_10_bits_off; // @[Slice.scala 167:21]
  assign abc_mshr_10_io_alloc_bits_mask = mshrAlloc_io_alloc_10_bits_mask; // @[Slice.scala 167:21]
  assign abc_mshr_10_io_alloc_bits_bufIdx = mshrAlloc_io_alloc_10_bits_bufIdx; // @[Slice.scala 167:21]
  assign abc_mshr_10_io_alloc_bits_preferCache = mshrAlloc_io_alloc_10_bits_preferCache; // @[Slice.scala 167:21]
  assign abc_mshr_10_io_alloc_bits_dirty = mshrAlloc_io_alloc_10_bits_dirty; // @[Slice.scala 167:21]
  assign abc_mshr_10_io_alloc_bits_fromProbeHelper = mshrAlloc_io_alloc_10_bits_fromProbeHelper; // @[Slice.scala 167:21]
  assign abc_mshr_10_io_alloc_bits_fromCmoHelper = mshrAlloc_io_alloc_10_bits_fromCmoHelper; // @[Slice.scala 167:21]
  assign abc_mshr_10_io_alloc_bits_needProbeAckData = mshrAlloc_io_alloc_10_bits_needProbeAckData; // @[Slice.scala 167:21]
  assign abc_mshr_10_io_resps_sink_c_valid = sinkC_io_resp_valid & sinkC_io_resp_bits_set ==
    abc_mshr_10_io_status_bits_set; // @[Slice.scala 527:57]
  assign abc_mshr_10_io_resps_sink_c_bits_hasData = sinkC_io_resp_bits_hasData; // @[Slice.scala 531:33]
  assign abc_mshr_10_io_resps_sink_c_bits_param = sinkC_io_resp_bits_param; // @[Slice.scala 531:33]
  assign abc_mshr_10_io_resps_sink_c_bits_source = sinkC_io_resp_bits_source; // @[Slice.scala 531:33]
  assign abc_mshr_10_io_resps_sink_c_bits_last = sinkC_io_resp_bits_last; // @[Slice.scala 531:33]
  assign abc_mshr_10_io_resps_sink_c_bits_bufIdx = sinkC_io_resp_bits_bufIdx; // @[Slice.scala 531:33]
  assign abc_mshr_10_io_resps_sink_d_valid = sinkD_io_resp_valid & sinkD_io_resp_bits_source == 4'ha; // @[Slice.scala 528:57]
  assign abc_mshr_10_io_resps_sink_d_bits_opcode = sinkD_io_resp_bits_opcode; // @[Slice.scala 532:33]
  assign abc_mshr_10_io_resps_sink_d_bits_param = sinkD_io_resp_bits_param; // @[Slice.scala 532:33]
  assign abc_mshr_10_io_resps_sink_d_bits_sink = sinkD_io_resp_bits_sink; // @[Slice.scala 532:33]
  assign abc_mshr_10_io_resps_sink_d_bits_last = sinkD_io_resp_bits_last; // @[Slice.scala 532:33]
  assign abc_mshr_10_io_resps_sink_d_bits_denied = sinkD_io_resp_bits_denied; // @[Slice.scala 532:33]
  assign abc_mshr_10_io_resps_sink_d_bits_bufIdx = sinkD_io_resp_bits_bufIdx; // @[Slice.scala 532:33]
  assign abc_mshr_10_io_resps_sink_e_valid = sinkE_io_resp_valid & sinkE_io_resp_bits_sink == 4'ha; // @[Slice.scala 529:57]
  assign abc_mshr_10_io_resps_source_d_valid = sourceD_io_resp_valid & sourceD_io_resp_bits_sink == 4'ha; // @[Slice.scala 530:61]
  assign abc_mshr_10_io_nestedwb_set = c_mshr_io_status_valid ? c_mshr_io_status_bits_set : bc_mshr_io_status_bits_set; // @[Slice.scala 258:22]
  assign abc_mshr_10_io_nestedwb_tag = c_mshr_io_status_valid ? c_mshr_io_status_bits_tag : bc_mshr_io_status_bits_tag; // @[Slice.scala 259:22]
  assign abc_mshr_10_io_nestedwb_btoN = _nestedWb_btoN_T_2 & _nestedWb_btoN_T_3; // @[Slice.scala 280:38]
  assign abc_mshr_10_io_nestedwb_btoB = _nestedWb_btoN_T_2 & _nestedWb_btoB_T_3; // @[Slice.scala 283:38]
  assign abc_mshr_10_io_nestedwb_bclr_dirty = _nestedWb_btoN_T_2 & _nestedWb_bclr_dirty_T_4; // @[Slice.scala 286:38]
  assign abc_mshr_10_io_nestedwb_bset_dirty = _nestedWb_btoN_T_2 & bc_mshr_io_tasks_dir_write_bits_data_dirty; // @[Slice.scala 289:38]
  assign abc_mshr_10_io_nestedwb_c_set_dirty = _nestedWb_c_set_dirty_T & c_mshr_io_tasks_dir_write_bits_data_dirty; // @[Slice.scala 292:37]
  assign abc_mshr_10_io_nestedwb_c_set_hit = c_mshr_io_status_valid & c_mshr_io_tasks_tag_write_valid &
    _nestedWb_c_set_hit_T_21; // @[Slice.scala 304:50]
  assign abc_mshr_10_io_nestedwb_clients_0_isToN = c_mshr_io_status_valid ? _nestedWb_clients_0_isToN_T_1 :
    _nestedWb_clients_0_isToN_T_3; // @[Slice.scala 314:25]
  assign abc_mshr_10_io_nestedwb_clients_1_isToN = c_mshr_io_status_valid ? _nestedWb_clients_1_isToN_T_1 :
    _nestedWb_clients_1_isToN_T_3; // @[Slice.scala 314:25]
  assign abc_mshr_10_io_tasks_sink_a_ready = 1'h0; // @[Slice.scala 472:13]
  assign abc_mshr_10_io_tasks_source_bready = sourceB_task_arb_io_in_10_ready; // @[Slice.scala 472:13]
  assign abc_mshr_10_io_tasks_sink_c_ready = sinkC_task_arb_io_in_10_ready; // @[Slice.scala 472:13]
  assign abc_mshr_10_io_tasks_source_d_ready = sourceD_task_arb_io_in_10_ready; // @[Slice.scala 472:13]
  assign abc_mshr_10_io_tasks_source_a_ready = sourceA_task_arb_io_in_10_ready; // @[Slice.scala 472:13]
  assign abc_mshr_10_io_tasks_source_c_ready = sourceC_task_arb_io_in_10_ready; // @[Slice.scala 472:13]
  assign abc_mshr_10_io_tasks_source_e_ready = sourceE_task_arb_io_in_10_ready; // @[Slice.scala 472:13]
  assign abc_mshr_10_io_tasks_dir_write_ready = arbiter_io_in_10_ready; // @[Slice.scala 406:60]
  assign abc_mshr_10_io_tasks_tag_write_ready = tagWrite_task_arb_io_in_10_ready; // @[Slice.scala 472:13]
  assign abc_mshr_10_io_tasks_client_dir_write_ready = arbiter_1_io_in_10_ready; // @[Slice.scala 406:60]
  assign abc_mshr_10_io_tasks_client_tag_write_ready = arbiter_2_io_in_10_ready; // @[Slice.scala 472:13]
  assign abc_mshr_10_io_dirResult_valid = ms_10_io_dirResult_valid_REG; // @[Slice.scala 556:31]
  assign abc_mshr_10_io_dirResult_bits_self_dirty = directory_io_result_bits_self_dirty; // @[Slice.scala 555:30]
  assign abc_mshr_10_io_dirResult_bits_self_state = directory_io_result_bits_self_state; // @[Slice.scala 555:30]
  assign abc_mshr_10_io_dirResult_bits_self_clientStates_0 = directory_io_result_bits_self_clientStates_0; // @[Slice.scala 555:30]
  assign abc_mshr_10_io_dirResult_bits_self_clientStates_1 = directory_io_result_bits_self_clientStates_1; // @[Slice.scala 555:30]
  assign abc_mshr_10_io_dirResult_bits_self_hit = directory_io_result_bits_self_hit; // @[Slice.scala 555:30]
  assign abc_mshr_10_io_dirResult_bits_self_way = directory_io_result_bits_self_way; // @[Slice.scala 555:30]
  assign abc_mshr_10_io_dirResult_bits_self_tag = directory_io_result_bits_self_tag; // @[Slice.scala 555:30]
  assign abc_mshr_10_io_dirResult_bits_clients_states_0_state = directory_io_result_bits_clients_states_0_state; // @[Slice.scala 555:30]
  assign abc_mshr_10_io_dirResult_bits_clients_states_0_hit = directory_io_result_bits_clients_states_0_hit; // @[Slice.scala 555:30]
  assign abc_mshr_10_io_dirResult_bits_clients_states_1_state = directory_io_result_bits_clients_states_1_state; // @[Slice.scala 555:30]
  assign abc_mshr_10_io_dirResult_bits_clients_states_1_hit = directory_io_result_bits_clients_states_1_hit; // @[Slice.scala 555:30]
  assign abc_mshr_10_io_dirResult_bits_clients_tag = directory_io_result_bits_clients_tag; // @[Slice.scala 555:30]
  assign abc_mshr_10_io_dirResult_bits_clients_way = directory_io_result_bits_clients_way; // @[Slice.scala 555:30]
  assign abc_mshr_10_io_c_status_set = c_mshr_io_status_bits_set; // @[Slice.scala 209:28]
  assign abc_mshr_10_io_c_status_tag = c_mshr_io_status_bits_tag; // @[Slice.scala 210:28]
  assign abc_mshr_10_io_c_status_way = c_mshr_io_status_bits_way; // @[Slice.scala 211:28]
  assign abc_mshr_10_io_c_status_nestedReleaseData = c_mshr_io_status_valid & c_mshr_io_is_nestedReleaseData; // @[Slice.scala 213:32]
  assign abc_mshr_10_io_bstatus_set = bc_mshr_io_status_bits_set; // @[Slice.scala 214:28]
  assign abc_mshr_10_io_bstatus_tag = bc_mshr_io_status_bits_tag; // @[Slice.scala 215:28]
  assign abc_mshr_10_io_bstatus_way = bc_mshr_io_status_bits_way; // @[Slice.scala 216:28]
  assign abc_mshr_10_io_bstatus_nestedProbeAckData = bc_mshr_io_status_valid & bc_mshr_io_is_nestedProbeAckData; // @[Slice.scala 218:33]
  assign abc_mshr_10_io_bstatus_probeHelperFinish = bc_mshr_io_status_valid & bc_mshr_io_probeHelperFinish; // @[Slice.scala 220:33]
  assign abc_mshr_10_io_releaseThrough = 1'h0; // @[Slice.scala 221:30]
  assign abc_mshr_10_io_probeAckDataThrough = 1'h0; // @[Slice.scala 222:35]
  assign abc_mshr_11_clock = clock;
  assign abc_mshr_11_reset = reset;
  assign abc_mshr_11_io_id = 4'hb; // @[Slice.scala 166:18]
  assign abc_mshr_11_io_enable = ~(bc_disable_11 | c_disable_11); // @[Slice.scala 198:25]
  assign abc_mshr_11_io_alloc_valid = mshrAlloc_io_alloc_11_valid; // @[Slice.scala 167:21]
  assign abc_mshr_11_io_alloc_bits_channel = mshrAlloc_io_alloc_11_bits_channel; // @[Slice.scala 167:21]
  assign abc_mshr_11_io_alloc_bits_opcode = mshrAlloc_io_alloc_11_bits_opcode; // @[Slice.scala 167:21]
  assign abc_mshr_11_io_alloc_bits_param = mshrAlloc_io_alloc_11_bits_param; // @[Slice.scala 167:21]
  assign abc_mshr_11_io_alloc_bits_size = mshrAlloc_io_alloc_11_bits_size; // @[Slice.scala 167:21]
  assign abc_mshr_11_io_alloc_bits_source = mshrAlloc_io_alloc_11_bits_source; // @[Slice.scala 167:21]
  assign abc_mshr_11_io_alloc_bits_set = mshrAlloc_io_alloc_11_bits_set; // @[Slice.scala 167:21]
  assign abc_mshr_11_io_alloc_bits_tag = mshrAlloc_io_alloc_11_bits_tag; // @[Slice.scala 167:21]
  assign abc_mshr_11_io_alloc_bits_off = mshrAlloc_io_alloc_11_bits_off; // @[Slice.scala 167:21]
  assign abc_mshr_11_io_alloc_bits_mask = mshrAlloc_io_alloc_11_bits_mask; // @[Slice.scala 167:21]
  assign abc_mshr_11_io_alloc_bits_bufIdx = mshrAlloc_io_alloc_11_bits_bufIdx; // @[Slice.scala 167:21]
  assign abc_mshr_11_io_alloc_bits_preferCache = mshrAlloc_io_alloc_11_bits_preferCache; // @[Slice.scala 167:21]
  assign abc_mshr_11_io_alloc_bits_dirty = mshrAlloc_io_alloc_11_bits_dirty; // @[Slice.scala 167:21]
  assign abc_mshr_11_io_alloc_bits_fromProbeHelper = mshrAlloc_io_alloc_11_bits_fromProbeHelper; // @[Slice.scala 167:21]
  assign abc_mshr_11_io_alloc_bits_fromCmoHelper = mshrAlloc_io_alloc_11_bits_fromCmoHelper; // @[Slice.scala 167:21]
  assign abc_mshr_11_io_alloc_bits_needProbeAckData = mshrAlloc_io_alloc_11_bits_needProbeAckData; // @[Slice.scala 167:21]
  assign abc_mshr_11_io_resps_sink_c_valid = sinkC_io_resp_valid & sinkC_io_resp_bits_set ==
    abc_mshr_11_io_status_bits_set; // @[Slice.scala 527:57]
  assign abc_mshr_11_io_resps_sink_c_bits_hasData = sinkC_io_resp_bits_hasData; // @[Slice.scala 531:33]
  assign abc_mshr_11_io_resps_sink_c_bits_param = sinkC_io_resp_bits_param; // @[Slice.scala 531:33]
  assign abc_mshr_11_io_resps_sink_c_bits_source = sinkC_io_resp_bits_source; // @[Slice.scala 531:33]
  assign abc_mshr_11_io_resps_sink_c_bits_last = sinkC_io_resp_bits_last; // @[Slice.scala 531:33]
  assign abc_mshr_11_io_resps_sink_c_bits_bufIdx = sinkC_io_resp_bits_bufIdx; // @[Slice.scala 531:33]
  assign abc_mshr_11_io_resps_sink_d_valid = sinkD_io_resp_valid & sinkD_io_resp_bits_source == 4'hb; // @[Slice.scala 528:57]
  assign abc_mshr_11_io_resps_sink_d_bits_opcode = sinkD_io_resp_bits_opcode; // @[Slice.scala 532:33]
  assign abc_mshr_11_io_resps_sink_d_bits_param = sinkD_io_resp_bits_param; // @[Slice.scala 532:33]
  assign abc_mshr_11_io_resps_sink_d_bits_sink = sinkD_io_resp_bits_sink; // @[Slice.scala 532:33]
  assign abc_mshr_11_io_resps_sink_d_bits_last = sinkD_io_resp_bits_last; // @[Slice.scala 532:33]
  assign abc_mshr_11_io_resps_sink_d_bits_denied = sinkD_io_resp_bits_denied; // @[Slice.scala 532:33]
  assign abc_mshr_11_io_resps_sink_d_bits_bufIdx = sinkD_io_resp_bits_bufIdx; // @[Slice.scala 532:33]
  assign abc_mshr_11_io_resps_sink_e_valid = sinkE_io_resp_valid & sinkE_io_resp_bits_sink == 4'hb; // @[Slice.scala 529:57]
  assign abc_mshr_11_io_resps_source_d_valid = sourceD_io_resp_valid & sourceD_io_resp_bits_sink == 4'hb; // @[Slice.scala 530:61]
  assign abc_mshr_11_io_nestedwb_set = c_mshr_io_status_valid ? c_mshr_io_status_bits_set : bc_mshr_io_status_bits_set; // @[Slice.scala 258:22]
  assign abc_mshr_11_io_nestedwb_tag = c_mshr_io_status_valid ? c_mshr_io_status_bits_tag : bc_mshr_io_status_bits_tag; // @[Slice.scala 259:22]
  assign abc_mshr_11_io_nestedwb_btoN = _nestedWb_btoN_T_2 & _nestedWb_btoN_T_3; // @[Slice.scala 280:38]
  assign abc_mshr_11_io_nestedwb_btoB = _nestedWb_btoN_T_2 & _nestedWb_btoB_T_3; // @[Slice.scala 283:38]
  assign abc_mshr_11_io_nestedwb_bclr_dirty = _nestedWb_btoN_T_2 & _nestedWb_bclr_dirty_T_4; // @[Slice.scala 286:38]
  assign abc_mshr_11_io_nestedwb_bset_dirty = _nestedWb_btoN_T_2 & bc_mshr_io_tasks_dir_write_bits_data_dirty; // @[Slice.scala 289:38]
  assign abc_mshr_11_io_nestedwb_c_set_dirty = _nestedWb_c_set_dirty_T & c_mshr_io_tasks_dir_write_bits_data_dirty; // @[Slice.scala 292:37]
  assign abc_mshr_11_io_nestedwb_c_set_hit = c_mshr_io_status_valid & c_mshr_io_tasks_tag_write_valid &
    _nestedWb_c_set_hit_T_23; // @[Slice.scala 304:50]
  assign abc_mshr_11_io_nestedwb_clients_0_isToN = c_mshr_io_status_valid ? _nestedWb_clients_0_isToN_T_1 :
    _nestedWb_clients_0_isToN_T_3; // @[Slice.scala 314:25]
  assign abc_mshr_11_io_nestedwb_clients_1_isToN = c_mshr_io_status_valid ? _nestedWb_clients_1_isToN_T_1 :
    _nestedWb_clients_1_isToN_T_3; // @[Slice.scala 314:25]
  assign abc_mshr_11_io_tasks_sink_a_ready = 1'h0; // @[Slice.scala 472:13]
  assign abc_mshr_11_io_tasks_source_bready = sourceB_task_arb_io_in_11_ready; // @[Slice.scala 472:13]
  assign abc_mshr_11_io_tasks_sink_c_ready = sinkC_task_arb_io_in_11_ready; // @[Slice.scala 472:13]
  assign abc_mshr_11_io_tasks_source_d_ready = sourceD_task_arb_io_in_11_ready; // @[Slice.scala 472:13]
  assign abc_mshr_11_io_tasks_source_a_ready = sourceA_task_arb_io_in_11_ready; // @[Slice.scala 472:13]
  assign abc_mshr_11_io_tasks_source_c_ready = sourceC_task_arb_io_in_11_ready; // @[Slice.scala 472:13]
  assign abc_mshr_11_io_tasks_source_e_ready = sourceE_task_arb_io_in_11_ready; // @[Slice.scala 472:13]
  assign abc_mshr_11_io_tasks_dir_write_ready = arbiter_io_in_11_ready; // @[Slice.scala 406:60]
  assign abc_mshr_11_io_tasks_tag_write_ready = tagWrite_task_arb_io_in_11_ready; // @[Slice.scala 472:13]
  assign abc_mshr_11_io_tasks_client_dir_write_ready = arbiter_1_io_in_11_ready; // @[Slice.scala 406:60]
  assign abc_mshr_11_io_tasks_client_tag_write_ready = arbiter_2_io_in_11_ready; // @[Slice.scala 472:13]
  assign abc_mshr_11_io_dirResult_valid = ms_11_io_dirResult_valid_REG; // @[Slice.scala 556:31]
  assign abc_mshr_11_io_dirResult_bits_self_dirty = directory_io_result_bits_self_dirty; // @[Slice.scala 555:30]
  assign abc_mshr_11_io_dirResult_bits_self_state = directory_io_result_bits_self_state; // @[Slice.scala 555:30]
  assign abc_mshr_11_io_dirResult_bits_self_clientStates_0 = directory_io_result_bits_self_clientStates_0; // @[Slice.scala 555:30]
  assign abc_mshr_11_io_dirResult_bits_self_clientStates_1 = directory_io_result_bits_self_clientStates_1; // @[Slice.scala 555:30]
  assign abc_mshr_11_io_dirResult_bits_self_hit = directory_io_result_bits_self_hit; // @[Slice.scala 555:30]
  assign abc_mshr_11_io_dirResult_bits_self_way = directory_io_result_bits_self_way; // @[Slice.scala 555:30]
  assign abc_mshr_11_io_dirResult_bits_self_tag = directory_io_result_bits_self_tag; // @[Slice.scala 555:30]
  assign abc_mshr_11_io_dirResult_bits_clients_states_0_state = directory_io_result_bits_clients_states_0_state; // @[Slice.scala 555:30]
  assign abc_mshr_11_io_dirResult_bits_clients_states_0_hit = directory_io_result_bits_clients_states_0_hit; // @[Slice.scala 555:30]
  assign abc_mshr_11_io_dirResult_bits_clients_states_1_state = directory_io_result_bits_clients_states_1_state; // @[Slice.scala 555:30]
  assign abc_mshr_11_io_dirResult_bits_clients_states_1_hit = directory_io_result_bits_clients_states_1_hit; // @[Slice.scala 555:30]
  assign abc_mshr_11_io_dirResult_bits_clients_tag = directory_io_result_bits_clients_tag; // @[Slice.scala 555:30]
  assign abc_mshr_11_io_dirResult_bits_clients_way = directory_io_result_bits_clients_way; // @[Slice.scala 555:30]
  assign abc_mshr_11_io_c_status_set = c_mshr_io_status_bits_set; // @[Slice.scala 209:28]
  assign abc_mshr_11_io_c_status_tag = c_mshr_io_status_bits_tag; // @[Slice.scala 210:28]
  assign abc_mshr_11_io_c_status_way = c_mshr_io_status_bits_way; // @[Slice.scala 211:28]
  assign abc_mshr_11_io_c_status_nestedReleaseData = c_mshr_io_status_valid & c_mshr_io_is_nestedReleaseData; // @[Slice.scala 213:32]
  assign abc_mshr_11_io_bstatus_set = bc_mshr_io_status_bits_set; // @[Slice.scala 214:28]
  assign abc_mshr_11_io_bstatus_tag = bc_mshr_io_status_bits_tag; // @[Slice.scala 215:28]
  assign abc_mshr_11_io_bstatus_way = bc_mshr_io_status_bits_way; // @[Slice.scala 216:28]
  assign abc_mshr_11_io_bstatus_nestedProbeAckData = bc_mshr_io_status_valid & bc_mshr_io_is_nestedProbeAckData; // @[Slice.scala 218:33]
  assign abc_mshr_11_io_bstatus_probeHelperFinish = bc_mshr_io_status_valid & bc_mshr_io_probeHelperFinish; // @[Slice.scala 220:33]
  assign abc_mshr_11_io_releaseThrough = 1'h0; // @[Slice.scala 221:30]
  assign abc_mshr_11_io_probeAckDataThrough = 1'h0; // @[Slice.scala 222:35]
  assign abc_mshr_12_clock = clock;
  assign abc_mshr_12_reset = reset;
  assign abc_mshr_12_io_id = 4'hc; // @[Slice.scala 166:18]
  assign abc_mshr_12_io_enable = ~(bc_disable_12 | c_disable_12); // @[Slice.scala 198:25]
  assign abc_mshr_12_io_alloc_valid = mshrAlloc_io_alloc_12_valid; // @[Slice.scala 167:21]
  assign abc_mshr_12_io_alloc_bits_channel = mshrAlloc_io_alloc_12_bits_channel; // @[Slice.scala 167:21]
  assign abc_mshr_12_io_alloc_bits_opcode = mshrAlloc_io_alloc_12_bits_opcode; // @[Slice.scala 167:21]
  assign abc_mshr_12_io_alloc_bits_param = mshrAlloc_io_alloc_12_bits_param; // @[Slice.scala 167:21]
  assign abc_mshr_12_io_alloc_bits_size = mshrAlloc_io_alloc_12_bits_size; // @[Slice.scala 167:21]
  assign abc_mshr_12_io_alloc_bits_source = mshrAlloc_io_alloc_12_bits_source; // @[Slice.scala 167:21]
  assign abc_mshr_12_io_alloc_bits_set = mshrAlloc_io_alloc_12_bits_set; // @[Slice.scala 167:21]
  assign abc_mshr_12_io_alloc_bits_tag = mshrAlloc_io_alloc_12_bits_tag; // @[Slice.scala 167:21]
  assign abc_mshr_12_io_alloc_bits_off = mshrAlloc_io_alloc_12_bits_off; // @[Slice.scala 167:21]
  assign abc_mshr_12_io_alloc_bits_mask = mshrAlloc_io_alloc_12_bits_mask; // @[Slice.scala 167:21]
  assign abc_mshr_12_io_alloc_bits_bufIdx = mshrAlloc_io_alloc_12_bits_bufIdx; // @[Slice.scala 167:21]
  assign abc_mshr_12_io_alloc_bits_preferCache = mshrAlloc_io_alloc_12_bits_preferCache; // @[Slice.scala 167:21]
  assign abc_mshr_12_io_alloc_bits_dirty = mshrAlloc_io_alloc_12_bits_dirty; // @[Slice.scala 167:21]
  assign abc_mshr_12_io_alloc_bits_fromProbeHelper = mshrAlloc_io_alloc_12_bits_fromProbeHelper; // @[Slice.scala 167:21]
  assign abc_mshr_12_io_alloc_bits_fromCmoHelper = mshrAlloc_io_alloc_12_bits_fromCmoHelper; // @[Slice.scala 167:21]
  assign abc_mshr_12_io_alloc_bits_needProbeAckData = mshrAlloc_io_alloc_12_bits_needProbeAckData; // @[Slice.scala 167:21]
  assign abc_mshr_12_io_resps_sink_c_valid = sinkC_io_resp_valid & sinkC_io_resp_bits_set ==
    abc_mshr_12_io_status_bits_set; // @[Slice.scala 527:57]
  assign abc_mshr_12_io_resps_sink_c_bits_hasData = sinkC_io_resp_bits_hasData; // @[Slice.scala 531:33]
  assign abc_mshr_12_io_resps_sink_c_bits_param = sinkC_io_resp_bits_param; // @[Slice.scala 531:33]
  assign abc_mshr_12_io_resps_sink_c_bits_source = sinkC_io_resp_bits_source; // @[Slice.scala 531:33]
  assign abc_mshr_12_io_resps_sink_c_bits_last = sinkC_io_resp_bits_last; // @[Slice.scala 531:33]
  assign abc_mshr_12_io_resps_sink_c_bits_bufIdx = sinkC_io_resp_bits_bufIdx; // @[Slice.scala 531:33]
  assign abc_mshr_12_io_resps_sink_d_valid = sinkD_io_resp_valid & sinkD_io_resp_bits_source == 4'hc; // @[Slice.scala 528:57]
  assign abc_mshr_12_io_resps_sink_d_bits_opcode = sinkD_io_resp_bits_opcode; // @[Slice.scala 532:33]
  assign abc_mshr_12_io_resps_sink_d_bits_param = sinkD_io_resp_bits_param; // @[Slice.scala 532:33]
  assign abc_mshr_12_io_resps_sink_d_bits_sink = sinkD_io_resp_bits_sink; // @[Slice.scala 532:33]
  assign abc_mshr_12_io_resps_sink_d_bits_last = sinkD_io_resp_bits_last; // @[Slice.scala 532:33]
  assign abc_mshr_12_io_resps_sink_d_bits_denied = sinkD_io_resp_bits_denied; // @[Slice.scala 532:33]
  assign abc_mshr_12_io_resps_sink_d_bits_bufIdx = sinkD_io_resp_bits_bufIdx; // @[Slice.scala 532:33]
  assign abc_mshr_12_io_resps_sink_e_valid = sinkE_io_resp_valid & sinkE_io_resp_bits_sink == 4'hc; // @[Slice.scala 529:57]
  assign abc_mshr_12_io_resps_source_d_valid = sourceD_io_resp_valid & sourceD_io_resp_bits_sink == 4'hc; // @[Slice.scala 530:61]
  assign abc_mshr_12_io_nestedwb_set = c_mshr_io_status_valid ? c_mshr_io_status_bits_set : bc_mshr_io_status_bits_set; // @[Slice.scala 258:22]
  assign abc_mshr_12_io_nestedwb_tag = c_mshr_io_status_valid ? c_mshr_io_status_bits_tag : bc_mshr_io_status_bits_tag; // @[Slice.scala 259:22]
  assign abc_mshr_12_io_nestedwb_btoN = _nestedWb_btoN_T_2 & _nestedWb_btoN_T_3; // @[Slice.scala 280:38]
  assign abc_mshr_12_io_nestedwb_btoB = _nestedWb_btoN_T_2 & _nestedWb_btoB_T_3; // @[Slice.scala 283:38]
  assign abc_mshr_12_io_nestedwb_bclr_dirty = _nestedWb_btoN_T_2 & _nestedWb_bclr_dirty_T_4; // @[Slice.scala 286:38]
  assign abc_mshr_12_io_nestedwb_bset_dirty = _nestedWb_btoN_T_2 & bc_mshr_io_tasks_dir_write_bits_data_dirty; // @[Slice.scala 289:38]
  assign abc_mshr_12_io_nestedwb_c_set_dirty = _nestedWb_c_set_dirty_T & c_mshr_io_tasks_dir_write_bits_data_dirty; // @[Slice.scala 292:37]
  assign abc_mshr_12_io_nestedwb_c_set_hit = c_mshr_io_status_valid & c_mshr_io_tasks_tag_write_valid &
    _nestedWb_c_set_hit_T_25; // @[Slice.scala 304:50]
  assign abc_mshr_12_io_nestedwb_clients_0_isToN = c_mshr_io_status_valid ? _nestedWb_clients_0_isToN_T_1 :
    _nestedWb_clients_0_isToN_T_3; // @[Slice.scala 314:25]
  assign abc_mshr_12_io_nestedwb_clients_1_isToN = c_mshr_io_status_valid ? _nestedWb_clients_1_isToN_T_1 :
    _nestedWb_clients_1_isToN_T_3; // @[Slice.scala 314:25]
  assign abc_mshr_12_io_tasks_sink_a_ready = 1'h0; // @[Slice.scala 472:13]
  assign abc_mshr_12_io_tasks_source_bready = sourceB_task_arb_io_in_12_ready; // @[Slice.scala 472:13]
  assign abc_mshr_12_io_tasks_sink_c_ready = sinkC_task_arb_io_in_12_ready; // @[Slice.scala 472:13]
  assign abc_mshr_12_io_tasks_source_d_ready = sourceD_task_arb_io_in_12_ready; // @[Slice.scala 472:13]
  assign abc_mshr_12_io_tasks_source_a_ready = sourceA_task_arb_io_in_12_ready; // @[Slice.scala 472:13]
  assign abc_mshr_12_io_tasks_source_c_ready = sourceC_task_arb_io_in_12_ready; // @[Slice.scala 472:13]
  assign abc_mshr_12_io_tasks_source_e_ready = sourceE_task_arb_io_in_12_ready; // @[Slice.scala 472:13]
  assign abc_mshr_12_io_tasks_dir_write_ready = arbiter_io_in_12_ready; // @[Slice.scala 406:60]
  assign abc_mshr_12_io_tasks_tag_write_ready = tagWrite_task_arb_io_in_12_ready; // @[Slice.scala 472:13]
  assign abc_mshr_12_io_tasks_client_dir_write_ready = arbiter_1_io_in_12_ready; // @[Slice.scala 406:60]
  assign abc_mshr_12_io_tasks_client_tag_write_ready = arbiter_2_io_in_12_ready; // @[Slice.scala 472:13]
  assign abc_mshr_12_io_dirResult_valid = ms_12_io_dirResult_valid_REG; // @[Slice.scala 556:31]
  assign abc_mshr_12_io_dirResult_bits_self_dirty = directory_io_result_bits_self_dirty; // @[Slice.scala 555:30]
  assign abc_mshr_12_io_dirResult_bits_self_state = directory_io_result_bits_self_state; // @[Slice.scala 555:30]
  assign abc_mshr_12_io_dirResult_bits_self_clientStates_0 = directory_io_result_bits_self_clientStates_0; // @[Slice.scala 555:30]
  assign abc_mshr_12_io_dirResult_bits_self_clientStates_1 = directory_io_result_bits_self_clientStates_1; // @[Slice.scala 555:30]
  assign abc_mshr_12_io_dirResult_bits_self_hit = directory_io_result_bits_self_hit; // @[Slice.scala 555:30]
  assign abc_mshr_12_io_dirResult_bits_self_way = directory_io_result_bits_self_way; // @[Slice.scala 555:30]
  assign abc_mshr_12_io_dirResult_bits_self_tag = directory_io_result_bits_self_tag; // @[Slice.scala 555:30]
  assign abc_mshr_12_io_dirResult_bits_clients_states_0_state = directory_io_result_bits_clients_states_0_state; // @[Slice.scala 555:30]
  assign abc_mshr_12_io_dirResult_bits_clients_states_0_hit = directory_io_result_bits_clients_states_0_hit; // @[Slice.scala 555:30]
  assign abc_mshr_12_io_dirResult_bits_clients_states_1_state = directory_io_result_bits_clients_states_1_state; // @[Slice.scala 555:30]
  assign abc_mshr_12_io_dirResult_bits_clients_states_1_hit = directory_io_result_bits_clients_states_1_hit; // @[Slice.scala 555:30]
  assign abc_mshr_12_io_dirResult_bits_clients_tag = directory_io_result_bits_clients_tag; // @[Slice.scala 555:30]
  assign abc_mshr_12_io_dirResult_bits_clients_way = directory_io_result_bits_clients_way; // @[Slice.scala 555:30]
  assign abc_mshr_12_io_c_status_set = c_mshr_io_status_bits_set; // @[Slice.scala 209:28]
  assign abc_mshr_12_io_c_status_tag = c_mshr_io_status_bits_tag; // @[Slice.scala 210:28]
  assign abc_mshr_12_io_c_status_way = c_mshr_io_status_bits_way; // @[Slice.scala 211:28]
  assign abc_mshr_12_io_c_status_nestedReleaseData = c_mshr_io_status_valid & c_mshr_io_is_nestedReleaseData; // @[Slice.scala 213:32]
  assign abc_mshr_12_io_bstatus_set = bc_mshr_io_status_bits_set; // @[Slice.scala 214:28]
  assign abc_mshr_12_io_bstatus_tag = bc_mshr_io_status_bits_tag; // @[Slice.scala 215:28]
  assign abc_mshr_12_io_bstatus_way = bc_mshr_io_status_bits_way; // @[Slice.scala 216:28]
  assign abc_mshr_12_io_bstatus_nestedProbeAckData = bc_mshr_io_status_valid & bc_mshr_io_is_nestedProbeAckData; // @[Slice.scala 218:33]
  assign abc_mshr_12_io_bstatus_probeHelperFinish = bc_mshr_io_status_valid & bc_mshr_io_probeHelperFinish; // @[Slice.scala 220:33]
  assign abc_mshr_12_io_releaseThrough = 1'h0; // @[Slice.scala 221:30]
  assign abc_mshr_12_io_probeAckDataThrough = 1'h0; // @[Slice.scala 222:35]
  assign abc_mshr_13_clock = clock;
  assign abc_mshr_13_reset = reset;
  assign abc_mshr_13_io_id = 4'hd; // @[Slice.scala 166:18]
  assign abc_mshr_13_io_enable = ~(bc_disable_13 | c_disable_13); // @[Slice.scala 198:25]
  assign abc_mshr_13_io_alloc_valid = mshrAlloc_io_alloc_13_valid; // @[Slice.scala 167:21]
  assign abc_mshr_13_io_alloc_bits_channel = mshrAlloc_io_alloc_13_bits_channel; // @[Slice.scala 167:21]
  assign abc_mshr_13_io_alloc_bits_opcode = mshrAlloc_io_alloc_13_bits_opcode; // @[Slice.scala 167:21]
  assign abc_mshr_13_io_alloc_bits_param = mshrAlloc_io_alloc_13_bits_param; // @[Slice.scala 167:21]
  assign abc_mshr_13_io_alloc_bits_size = mshrAlloc_io_alloc_13_bits_size; // @[Slice.scala 167:21]
  assign abc_mshr_13_io_alloc_bits_source = mshrAlloc_io_alloc_13_bits_source; // @[Slice.scala 167:21]
  assign abc_mshr_13_io_alloc_bits_set = mshrAlloc_io_alloc_13_bits_set; // @[Slice.scala 167:21]
  assign abc_mshr_13_io_alloc_bits_tag = mshrAlloc_io_alloc_13_bits_tag; // @[Slice.scala 167:21]
  assign abc_mshr_13_io_alloc_bits_off = mshrAlloc_io_alloc_13_bits_off; // @[Slice.scala 167:21]
  assign abc_mshr_13_io_alloc_bits_mask = mshrAlloc_io_alloc_13_bits_mask; // @[Slice.scala 167:21]
  assign abc_mshr_13_io_alloc_bits_bufIdx = mshrAlloc_io_alloc_13_bits_bufIdx; // @[Slice.scala 167:21]
  assign abc_mshr_13_io_alloc_bits_preferCache = mshrAlloc_io_alloc_13_bits_preferCache; // @[Slice.scala 167:21]
  assign abc_mshr_13_io_alloc_bits_dirty = mshrAlloc_io_alloc_13_bits_dirty; // @[Slice.scala 167:21]
  assign abc_mshr_13_io_alloc_bits_fromProbeHelper = mshrAlloc_io_alloc_13_bits_fromProbeHelper; // @[Slice.scala 167:21]
  assign abc_mshr_13_io_alloc_bits_fromCmoHelper = mshrAlloc_io_alloc_13_bits_fromCmoHelper; // @[Slice.scala 167:21]
  assign abc_mshr_13_io_alloc_bits_needProbeAckData = mshrAlloc_io_alloc_13_bits_needProbeAckData; // @[Slice.scala 167:21]
  assign abc_mshr_13_io_resps_sink_c_valid = sinkC_io_resp_valid & sinkC_io_resp_bits_set ==
    abc_mshr_13_io_status_bits_set; // @[Slice.scala 527:57]
  assign abc_mshr_13_io_resps_sink_c_bits_hasData = sinkC_io_resp_bits_hasData; // @[Slice.scala 531:33]
  assign abc_mshr_13_io_resps_sink_c_bits_param = sinkC_io_resp_bits_param; // @[Slice.scala 531:33]
  assign abc_mshr_13_io_resps_sink_c_bits_source = sinkC_io_resp_bits_source; // @[Slice.scala 531:33]
  assign abc_mshr_13_io_resps_sink_c_bits_last = sinkC_io_resp_bits_last; // @[Slice.scala 531:33]
  assign abc_mshr_13_io_resps_sink_c_bits_bufIdx = sinkC_io_resp_bits_bufIdx; // @[Slice.scala 531:33]
  assign abc_mshr_13_io_resps_sink_d_valid = sinkD_io_resp_valid & sinkD_io_resp_bits_source == 4'hd; // @[Slice.scala 528:57]
  assign abc_mshr_13_io_resps_sink_d_bits_opcode = sinkD_io_resp_bits_opcode; // @[Slice.scala 532:33]
  assign abc_mshr_13_io_resps_sink_d_bits_param = sinkD_io_resp_bits_param; // @[Slice.scala 532:33]
  assign abc_mshr_13_io_resps_sink_d_bits_sink = sinkD_io_resp_bits_sink; // @[Slice.scala 532:33]
  assign abc_mshr_13_io_resps_sink_d_bits_last = sinkD_io_resp_bits_last; // @[Slice.scala 532:33]
  assign abc_mshr_13_io_resps_sink_d_bits_denied = sinkD_io_resp_bits_denied; // @[Slice.scala 532:33]
  assign abc_mshr_13_io_resps_sink_d_bits_bufIdx = sinkD_io_resp_bits_bufIdx; // @[Slice.scala 532:33]
  assign abc_mshr_13_io_resps_sink_e_valid = sinkE_io_resp_valid & sinkE_io_resp_bits_sink == 4'hd; // @[Slice.scala 529:57]
  assign abc_mshr_13_io_resps_source_d_valid = sourceD_io_resp_valid & sourceD_io_resp_bits_sink == 4'hd; // @[Slice.scala 530:61]
  assign abc_mshr_13_io_nestedwb_set = c_mshr_io_status_valid ? c_mshr_io_status_bits_set : bc_mshr_io_status_bits_set; // @[Slice.scala 258:22]
  assign abc_mshr_13_io_nestedwb_tag = c_mshr_io_status_valid ? c_mshr_io_status_bits_tag : bc_mshr_io_status_bits_tag; // @[Slice.scala 259:22]
  assign abc_mshr_13_io_nestedwb_btoN = _nestedWb_btoN_T_2 & _nestedWb_btoN_T_3; // @[Slice.scala 280:38]
  assign abc_mshr_13_io_nestedwb_btoB = _nestedWb_btoN_T_2 & _nestedWb_btoB_T_3; // @[Slice.scala 283:38]
  assign abc_mshr_13_io_nestedwb_bclr_dirty = _nestedWb_btoN_T_2 & _nestedWb_bclr_dirty_T_4; // @[Slice.scala 286:38]
  assign abc_mshr_13_io_nestedwb_bset_dirty = _nestedWb_btoN_T_2 & bc_mshr_io_tasks_dir_write_bits_data_dirty; // @[Slice.scala 289:38]
  assign abc_mshr_13_io_nestedwb_c_set_dirty = _nestedWb_c_set_dirty_T & c_mshr_io_tasks_dir_write_bits_data_dirty; // @[Slice.scala 292:37]
  assign abc_mshr_13_io_nestedwb_c_set_hit = c_mshr_io_status_valid & c_mshr_io_tasks_tag_write_valid &
    _nestedWb_c_set_hit_T_27; // @[Slice.scala 304:50]
  assign abc_mshr_13_io_nestedwb_clients_0_isToN = c_mshr_io_status_valid ? _nestedWb_clients_0_isToN_T_1 :
    _nestedWb_clients_0_isToN_T_3; // @[Slice.scala 314:25]
  assign abc_mshr_13_io_nestedwb_clients_1_isToN = c_mshr_io_status_valid ? _nestedWb_clients_1_isToN_T_1 :
    _nestedWb_clients_1_isToN_T_3; // @[Slice.scala 314:25]
  assign abc_mshr_13_io_tasks_sink_a_ready = 1'h0; // @[Slice.scala 472:13]
  assign abc_mshr_13_io_tasks_source_bready = sourceB_task_arb_io_in_13_ready; // @[Slice.scala 472:13]
  assign abc_mshr_13_io_tasks_sink_c_ready = sinkC_task_arb_io_in_13_ready; // @[Slice.scala 472:13]
  assign abc_mshr_13_io_tasks_source_d_ready = sourceD_task_arb_io_in_13_ready; // @[Slice.scala 472:13]
  assign abc_mshr_13_io_tasks_source_a_ready = sourceA_task_arb_io_in_13_ready; // @[Slice.scala 472:13]
  assign abc_mshr_13_io_tasks_source_c_ready = sourceC_task_arb_io_in_13_ready; // @[Slice.scala 472:13]
  assign abc_mshr_13_io_tasks_source_e_ready = sourceE_task_arb_io_in_13_ready; // @[Slice.scala 472:13]
  assign abc_mshr_13_io_tasks_dir_write_ready = arbiter_io_in_13_ready; // @[Slice.scala 406:60]
  assign abc_mshr_13_io_tasks_tag_write_ready = tagWrite_task_arb_io_in_13_ready; // @[Slice.scala 472:13]
  assign abc_mshr_13_io_tasks_client_dir_write_ready = arbiter_1_io_in_13_ready; // @[Slice.scala 406:60]
  assign abc_mshr_13_io_tasks_client_tag_write_ready = arbiter_2_io_in_13_ready; // @[Slice.scala 472:13]
  assign abc_mshr_13_io_dirResult_valid = ms_13_io_dirResult_valid_REG; // @[Slice.scala 556:31]
  assign abc_mshr_13_io_dirResult_bits_self_dirty = directory_io_result_bits_self_dirty; // @[Slice.scala 555:30]
  assign abc_mshr_13_io_dirResult_bits_self_state = directory_io_result_bits_self_state; // @[Slice.scala 555:30]
  assign abc_mshr_13_io_dirResult_bits_self_clientStates_0 = directory_io_result_bits_self_clientStates_0; // @[Slice.scala 555:30]
  assign abc_mshr_13_io_dirResult_bits_self_clientStates_1 = directory_io_result_bits_self_clientStates_1; // @[Slice.scala 555:30]
  assign abc_mshr_13_io_dirResult_bits_self_hit = directory_io_result_bits_self_hit; // @[Slice.scala 555:30]
  assign abc_mshr_13_io_dirResult_bits_self_way = directory_io_result_bits_self_way; // @[Slice.scala 555:30]
  assign abc_mshr_13_io_dirResult_bits_self_tag = directory_io_result_bits_self_tag; // @[Slice.scala 555:30]
  assign abc_mshr_13_io_dirResult_bits_clients_states_0_state = directory_io_result_bits_clients_states_0_state; // @[Slice.scala 555:30]
  assign abc_mshr_13_io_dirResult_bits_clients_states_0_hit = directory_io_result_bits_clients_states_0_hit; // @[Slice.scala 555:30]
  assign abc_mshr_13_io_dirResult_bits_clients_states_1_state = directory_io_result_bits_clients_states_1_state; // @[Slice.scala 555:30]
  assign abc_mshr_13_io_dirResult_bits_clients_states_1_hit = directory_io_result_bits_clients_states_1_hit; // @[Slice.scala 555:30]
  assign abc_mshr_13_io_dirResult_bits_clients_tag = directory_io_result_bits_clients_tag; // @[Slice.scala 555:30]
  assign abc_mshr_13_io_dirResult_bits_clients_way = directory_io_result_bits_clients_way; // @[Slice.scala 555:30]
  assign abc_mshr_13_io_c_status_set = c_mshr_io_status_bits_set; // @[Slice.scala 209:28]
  assign abc_mshr_13_io_c_status_tag = c_mshr_io_status_bits_tag; // @[Slice.scala 210:28]
  assign abc_mshr_13_io_c_status_way = c_mshr_io_status_bits_way; // @[Slice.scala 211:28]
  assign abc_mshr_13_io_c_status_nestedReleaseData = c_mshr_io_status_valid & c_mshr_io_is_nestedReleaseData; // @[Slice.scala 213:32]
  assign abc_mshr_13_io_bstatus_set = bc_mshr_io_status_bits_set; // @[Slice.scala 214:28]
  assign abc_mshr_13_io_bstatus_tag = bc_mshr_io_status_bits_tag; // @[Slice.scala 215:28]
  assign abc_mshr_13_io_bstatus_way = bc_mshr_io_status_bits_way; // @[Slice.scala 216:28]
  assign abc_mshr_13_io_bstatus_nestedProbeAckData = bc_mshr_io_status_valid & bc_mshr_io_is_nestedProbeAckData; // @[Slice.scala 218:33]
  assign abc_mshr_13_io_bstatus_probeHelperFinish = bc_mshr_io_status_valid & bc_mshr_io_probeHelperFinish; // @[Slice.scala 220:33]
  assign abc_mshr_13_io_releaseThrough = 1'h0; // @[Slice.scala 221:30]
  assign abc_mshr_13_io_probeAckDataThrough = 1'h0; // @[Slice.scala 222:35]
  assign bc_mshr_clock = clock;
  assign bc_mshr_reset = reset;
  assign bc_mshr_io_id = 4'he; // @[Slice.scala 166:18]
  assign bc_mshr_io_enable = ~(c_mask_latch_14 & c_mshr_io_status_valid); // @[Slice.scala 200:24]
  assign bc_mshr_io_alloc_valid = mshrAlloc_io_alloc_14_valid; // @[Slice.scala 167:21]
  assign bc_mshr_io_alloc_bits_channel = mshrAlloc_io_alloc_14_bits_channel; // @[Slice.scala 167:21]
  assign bc_mshr_io_alloc_bits_opcode = mshrAlloc_io_alloc_14_bits_opcode; // @[Slice.scala 167:21]
  assign bc_mshr_io_alloc_bits_param = mshrAlloc_io_alloc_14_bits_param; // @[Slice.scala 167:21]
  assign bc_mshr_io_alloc_bits_size = mshrAlloc_io_alloc_14_bits_size; // @[Slice.scala 167:21]
  assign bc_mshr_io_alloc_bits_source = mshrAlloc_io_alloc_14_bits_source; // @[Slice.scala 167:21]
  assign bc_mshr_io_alloc_bits_set = mshrAlloc_io_alloc_14_bits_set; // @[Slice.scala 167:21]
  assign bc_mshr_io_alloc_bits_tag = mshrAlloc_io_alloc_14_bits_tag; // @[Slice.scala 167:21]
  assign bc_mshr_io_alloc_bits_off = mshrAlloc_io_alloc_14_bits_off; // @[Slice.scala 167:21]
  assign bc_mshr_io_alloc_bits_mask = mshrAlloc_io_alloc_14_bits_mask; // @[Slice.scala 167:21]
  assign bc_mshr_io_alloc_bits_bufIdx = mshrAlloc_io_alloc_14_bits_bufIdx; // @[Slice.scala 167:21]
  assign bc_mshr_io_alloc_bits_preferCache = mshrAlloc_io_alloc_14_bits_preferCache; // @[Slice.scala 167:21]
  assign bc_mshr_io_alloc_bits_dirty = mshrAlloc_io_alloc_14_bits_dirty; // @[Slice.scala 167:21]
  assign bc_mshr_io_alloc_bits_fromProbeHelper = mshrAlloc_io_alloc_14_bits_fromProbeHelper; // @[Slice.scala 167:21]
  assign bc_mshr_io_alloc_bits_fromCmoHelper = mshrAlloc_io_alloc_14_bits_fromCmoHelper; // @[Slice.scala 167:21]
  assign bc_mshr_io_alloc_bits_needProbeAckData = mshrAlloc_io_alloc_14_bits_needProbeAckData; // @[Slice.scala 167:21]
  assign bc_mshr_io_resps_sink_c_valid = sinkC_io_resp_valid & sinkC_io_resp_bits_set == bc_mshr_io_status_bits_set; // @[Slice.scala 527:57]
  assign bc_mshr_io_resps_sink_c_bits_hasData = sinkC_io_resp_bits_hasData; // @[Slice.scala 531:33]
  assign bc_mshr_io_resps_sink_c_bits_param = sinkC_io_resp_bits_param; // @[Slice.scala 531:33]
  assign bc_mshr_io_resps_sink_c_bits_source = sinkC_io_resp_bits_source; // @[Slice.scala 531:33]
  assign bc_mshr_io_resps_sink_c_bits_last = sinkC_io_resp_bits_last; // @[Slice.scala 531:33]
  assign bc_mshr_io_resps_sink_c_bits_bufIdx = sinkC_io_resp_bits_bufIdx; // @[Slice.scala 531:33]
  assign bc_mshr_io_resps_sink_d_valid = sinkD_io_resp_valid & sinkD_io_resp_bits_source == 4'he; // @[Slice.scala 528:57]
  assign bc_mshr_io_resps_sink_d_bits_opcode = sinkD_io_resp_bits_opcode; // @[Slice.scala 532:33]
  assign bc_mshr_io_resps_sink_d_bits_param = sinkD_io_resp_bits_param; // @[Slice.scala 532:33]
  assign bc_mshr_io_resps_sink_d_bits_sink = sinkD_io_resp_bits_sink; // @[Slice.scala 532:33]
  assign bc_mshr_io_resps_sink_d_bits_last = sinkD_io_resp_bits_last; // @[Slice.scala 532:33]
  assign bc_mshr_io_resps_sink_d_bits_denied = sinkD_io_resp_bits_denied; // @[Slice.scala 532:33]
  assign bc_mshr_io_resps_sink_d_bits_bufIdx = sinkD_io_resp_bits_bufIdx; // @[Slice.scala 532:33]
  assign bc_mshr_io_resps_sink_e_valid = sinkE_io_resp_valid & sinkE_io_resp_bits_sink == 4'he; // @[Slice.scala 529:57]
  assign bc_mshr_io_resps_source_d_valid = sourceD_io_resp_valid & sourceD_io_resp_bits_sink == 4'he; // @[Slice.scala 530:61]
  assign bc_mshr_io_nestedwb_set = c_mshr_io_status_bits_set; // @[Slice.scala 342:27]
  assign bc_mshr_io_nestedwb_tag = c_mshr_io_status_bits_tag; // @[Slice.scala 343:27]
  assign bc_mshr_io_nestedwb_btoN = 1'h0; // @[Slice.scala 341:{38,38}]
  assign bc_mshr_io_nestedwb_btoB = 1'h0; // @[Slice.scala 341:{38,38}]
  assign bc_mshr_io_nestedwb_bclr_dirty = 1'h0; // @[Slice.scala 341:{38,38}]
  assign bc_mshr_io_nestedwb_bset_dirty = 1'h0; // @[Slice.scala 341:{38,38}]
  assign bc_mshr_io_nestedwb_c_set_dirty = _nestedWb_c_set_dirty_T & c_mshr_io_tasks_dir_write_bits_data_dirty; // @[Slice.scala 292:37]
  assign bc_mshr_io_nestedwb_c_set_hit = c_mshr_io_status_valid & c_mshr_io_tasks_tag_write_valid &
    _nestedWb_c_set_hit_T_29; // @[Slice.scala 304:50]
  assign bc_mshr_io_nestedwb_clients_0_isToN = c_mshr_io_status_valid & nestedWb_clients_0_isToN; // @[Slice.scala 355:18 358:11 341:23]
  assign bc_mshr_io_nestedwb_clients_1_isToN = c_mshr_io_status_valid & nestedWb_clients_1_isToN; // @[Slice.scala 355:18 358:11 341:23]
  assign bc_mshr_io_tasks_sink_a_ready = 1'h0; // @[Slice.scala 492:49]
  assign bc_mshr_io_tasks_source_bready = sourceB_io_task_ready & bc_valid_latch_1 & ~c_real_valid_1; // @[Slice.scala 492:49]
  assign bc_mshr_io_tasks_sink_c_ready = sinkC_io_task_ready & bc_valid_latch_6 & ~c_real_valid_6; // @[Slice.scala 492:49]
  assign bc_mshr_io_tasks_source_d_ready = sourceD_io_task_ready & bc_valid_latch_3 & ~c_real_valid_3; // @[Slice.scala 492:49]
  assign bc_mshr_io_tasks_source_a_ready = sourceA_io_task_ready & bc_valid_latch & ~c_real_valid; // @[Slice.scala 492:49]
  assign bc_mshr_io_tasks_source_c_ready = sourceC_io_task_ready & bc_valid_latch_2 & ~c_real_valid_2; // @[Slice.scala 492:49]
  assign bc_mshr_io_tasks_source_e_ready = sourceE_io_task_ready & bc_valid_latch_4 & ~c_real_valid_4; // @[Slice.scala 492:49]
  assign bc_mshr_io_tasks_dir_write_ready = _nestedWb_btoN_T & arbiter_io_in_14_ready; // @[Slice.scala 391:28]
  assign bc_mshr_io_tasks_tag_write_ready = bc_valid_latch_7 & ~c_real_valid_7; // @[Slice.scala 492:49]
  assign bc_mshr_io_tasks_client_dir_write_ready = _nestedWb_btoN_T & arbiter_1_io_in_14_ready; // @[Slice.scala 391:28]
  assign bc_mshr_io_tasks_client_tag_write_ready = bc_valid_latch_8 & ~c_real_valid_8; // @[Slice.scala 492:49]
  assign bc_mshr_io_dirResult_valid = ms_14_io_dirResult_valid_REG; // @[Slice.scala 556:31]
  assign bc_mshr_io_dirResult_bits_self_dirty = directory_io_result_bits_self_dirty; // @[Slice.scala 555:30]
  assign bc_mshr_io_dirResult_bits_self_state = directory_io_result_bits_self_state; // @[Slice.scala 555:30]
  assign bc_mshr_io_dirResult_bits_self_clientStates_0 = directory_io_result_bits_self_clientStates_0; // @[Slice.scala 555:30]
  assign bc_mshr_io_dirResult_bits_self_clientStates_1 = directory_io_result_bits_self_clientStates_1; // @[Slice.scala 555:30]
  assign bc_mshr_io_dirResult_bits_self_hit = directory_io_result_bits_self_hit; // @[Slice.scala 555:30]
  assign bc_mshr_io_dirResult_bits_self_way = directory_io_result_bits_self_way; // @[Slice.scala 555:30]
  assign bc_mshr_io_dirResult_bits_self_tag = directory_io_result_bits_self_tag; // @[Slice.scala 555:30]
  assign bc_mshr_io_dirResult_bits_clients_states_0_state = directory_io_result_bits_clients_states_0_state; // @[Slice.scala 555:30]
  assign bc_mshr_io_dirResult_bits_clients_states_0_hit = directory_io_result_bits_clients_states_0_hit; // @[Slice.scala 555:30]
  assign bc_mshr_io_dirResult_bits_clients_states_1_state = directory_io_result_bits_clients_states_1_state; // @[Slice.scala 555:30]
  assign bc_mshr_io_dirResult_bits_clients_states_1_hit = directory_io_result_bits_clients_states_1_hit; // @[Slice.scala 555:30]
  assign bc_mshr_io_dirResult_bits_clients_tag = directory_io_result_bits_clients_tag; // @[Slice.scala 555:30]
  assign bc_mshr_io_dirResult_bits_clients_way = directory_io_result_bits_clients_way; // @[Slice.scala 555:30]
  assign bc_mshr_io_c_status_set = c_mshr_io_status_bits_set; // @[Slice.scala 228:28]
  assign bc_mshr_io_c_status_tag = c_mshr_io_status_bits_tag; // @[Slice.scala 229:28]
  assign bc_mshr_io_c_status_way = c_mshr_io_status_bits_way; // @[Slice.scala 230:28]
  assign bc_mshr_io_c_status_nestedReleaseData = c_mshr_io_status_valid & c_mshr_io_is_nestedReleaseData; // @[Slice.scala 232:32]
  assign bc_mshr_io_bstatus_set = 10'h0; // @[Slice.scala 233:28]
  assign bc_mshr_io_bstatus_tag = 20'h0; // @[Slice.scala 234:28]
  assign bc_mshr_io_bstatus_way = 3'h0; // @[Slice.scala 235:28]
  assign bc_mshr_io_bstatus_nestedProbeAckData = 1'h0; // @[Slice.scala 236:43]
  assign bc_mshr_io_bstatus_probeHelperFinish = 1'h0; // @[Slice.scala 237:42]
  assign bc_mshr_io_releaseThrough = 1'h0; // @[Slice.scala 348:30]
  assign bc_mshr_io_probeAckDataThrough = |_ms_14_io_probeAckDataThrough_T; // @[Slice.scala 351:12]
  assign c_mshr_clock = clock;
  assign c_mshr_reset = reset;
  assign c_mshr_io_id = 4'hf; // @[Slice.scala 166:18]
  assign c_mshr_io_enable = 1'h1; // @[Slice.scala 201:20]
  assign c_mshr_io_alloc_valid = mshrAlloc_io_alloc_15_valid; // @[Slice.scala 167:21]
  assign c_mshr_io_alloc_bits_channel = 3'h4; // @[Slice.scala 167:21]
  assign c_mshr_io_alloc_bits_opcode = mshrAlloc_io_alloc_15_bits_opcode; // @[Slice.scala 167:21]
  assign c_mshr_io_alloc_bits_param = mshrAlloc_io_alloc_15_bits_param; // @[Slice.scala 167:21]
  assign c_mshr_io_alloc_bits_size = mshrAlloc_io_alloc_15_bits_size; // @[Slice.scala 167:21]
  assign c_mshr_io_alloc_bits_source = mshrAlloc_io_alloc_15_bits_source; // @[Slice.scala 167:21]
  assign c_mshr_io_alloc_bits_set = mshrAlloc_io_alloc_15_bits_set; // @[Slice.scala 167:21]
  assign c_mshr_io_alloc_bits_tag = mshrAlloc_io_alloc_15_bits_tag; // @[Slice.scala 167:21]
  assign c_mshr_io_alloc_bits_off = mshrAlloc_io_alloc_15_bits_off; // @[Slice.scala 167:21]
  assign c_mshr_io_alloc_bits_mask = 32'h0; // @[Slice.scala 167:21]
  assign c_mshr_io_alloc_bits_bufIdx = mshrAlloc_io_alloc_15_bits_bufIdx; // @[Slice.scala 167:21]
  assign c_mshr_io_alloc_bits_preferCache = 1'h1; // @[Slice.scala 167:21]
  assign c_mshr_io_alloc_bits_dirty = mshrAlloc_io_alloc_15_bits_dirty; // @[Slice.scala 167:21]
  assign c_mshr_io_alloc_bits_fromProbeHelper = 1'h0; // @[Slice.scala 167:21]
  assign c_mshr_io_alloc_bits_fromCmoHelper = 1'h0; // @[Slice.scala 167:21]
  assign c_mshr_io_alloc_bits_needProbeAckData = 1'h0; // @[Slice.scala 167:21]
  assign c_mshr_io_resps_sink_c_valid = 1'h0; // @[Slice.scala 536:32]
  assign c_mshr_io_resps_sink_c_bits_hasData = sinkC_io_resp_bits_hasData; // @[Slice.scala 531:33]
  assign c_mshr_io_resps_sink_c_bits_param = sinkC_io_resp_bits_param; // @[Slice.scala 531:33]
  assign c_mshr_io_resps_sink_c_bits_source = sinkC_io_resp_bits_source; // @[Slice.scala 531:33]
  assign c_mshr_io_resps_sink_c_bits_last = sinkC_io_resp_bits_last; // @[Slice.scala 531:33]
  assign c_mshr_io_resps_sink_c_bits_bufIdx = sinkC_io_resp_bits_bufIdx; // @[Slice.scala 531:33]
  assign c_mshr_io_resps_sink_d_valid = sinkD_io_resp_valid & sinkD_io_resp_bits_source == 4'hf; // @[Slice.scala 528:57]
  assign c_mshr_io_resps_sink_d_bits_opcode = sinkD_io_resp_bits_opcode; // @[Slice.scala 532:33]
  assign c_mshr_io_resps_sink_d_bits_param = sinkD_io_resp_bits_param; // @[Slice.scala 532:33]
  assign c_mshr_io_resps_sink_d_bits_sink = sinkD_io_resp_bits_sink; // @[Slice.scala 532:33]
  assign c_mshr_io_resps_sink_d_bits_last = sinkD_io_resp_bits_last; // @[Slice.scala 532:33]
  assign c_mshr_io_resps_sink_d_bits_denied = sinkD_io_resp_bits_denied; // @[Slice.scala 532:33]
  assign c_mshr_io_resps_sink_d_bits_bufIdx = sinkD_io_resp_bits_bufIdx; // @[Slice.scala 532:33]
  assign c_mshr_io_resps_sink_e_valid = sinkE_io_resp_valid & sinkE_io_resp_bits_sink == 4'hf; // @[Slice.scala 529:57]
  assign c_mshr_io_resps_source_d_valid = sourceD_io_resp_valid & sourceD_io_resp_bits_sink == 4'hf; // @[Slice.scala 530:61]
  assign c_mshr_io_nestedwb_set = 10'h0; // @[Slice.scala 362:{37,37}]
  assign c_mshr_io_nestedwb_tag = 20'h0; // @[Slice.scala 362:{37,37}]
  assign c_mshr_io_nestedwb_btoN = 1'h0; // @[Slice.scala 362:{37,37}]
  assign c_mshr_io_nestedwb_btoB = 1'h0; // @[Slice.scala 362:{37,37}]
  assign c_mshr_io_nestedwb_bclr_dirty = 1'h0; // @[Slice.scala 362:{37,37}]
  assign c_mshr_io_nestedwb_bset_dirty = 1'h0; // @[Slice.scala 362:{37,37}]
  assign c_mshr_io_nestedwb_c_set_dirty = 1'h0; // @[Slice.scala 362:{37,37}]
  assign c_mshr_io_nestedwb_c_set_hit = 1'h0; // @[Slice.scala 362:{37,37}]
  assign c_mshr_io_nestedwb_clients_0_isToN = 1'h0; // @[Slice.scala 362:{37,37}]
  assign c_mshr_io_nestedwb_clients_1_isToN = 1'h0; // @[Slice.scala 362:{37,37}]
  assign c_mshr_io_tasks_sink_a_ready = 1'h0; // @[Slice.scala 491:30]
  assign c_mshr_io_tasks_source_bready = sourceB_io_task_ready & c_valid_latch_1; // @[Slice.scala 491:30]
  assign c_mshr_io_tasks_sink_c_ready = sinkC_io_task_ready & c_valid_latch_6; // @[Slice.scala 491:30]
  assign c_mshr_io_tasks_source_d_ready = sourceD_io_task_ready & c_valid_latch_3; // @[Slice.scala 491:30]
  assign c_mshr_io_tasks_source_a_ready = sourceA_io_task_ready & c_valid_latch; // @[Slice.scala 491:30]
  assign c_mshr_io_tasks_source_c_ready = sourceC_io_task_ready & c_valid_latch_2; // @[Slice.scala 491:30]
  assign c_mshr_io_tasks_source_e_ready = sourceE_io_task_ready & c_valid_latch_4; // @[Slice.scala 491:30]
  assign c_mshr_io_tasks_dir_write_ready = arbiter_io_in_15_ready; // @[Slice.scala 408:24]
  assign c_mshr_io_tasks_tag_write_ready = c_valid_latch_7; // @[Slice.scala 491:30]
  assign c_mshr_io_tasks_client_dir_write_ready = arbiter_1_io_in_15_ready; // @[Slice.scala 408:24]
  assign c_mshr_io_tasks_client_tag_write_ready = c_valid_latch_8; // @[Slice.scala 491:30]
  assign c_mshr_io_dirResult_valid = ms_15_io_dirResult_valid_REG; // @[Slice.scala 556:31]
  assign c_mshr_io_dirResult_bits_self_dirty = directory_io_result_bits_self_dirty; // @[Slice.scala 555:30]
  assign c_mshr_io_dirResult_bits_self_state = directory_io_result_bits_self_state; // @[Slice.scala 555:30]
  assign c_mshr_io_dirResult_bits_self_clientStates_0 = directory_io_result_bits_self_clientStates_0; // @[Slice.scala 555:30]
  assign c_mshr_io_dirResult_bits_self_clientStates_1 = directory_io_result_bits_self_clientStates_1; // @[Slice.scala 555:30]
  assign c_mshr_io_dirResult_bits_self_hit = directory_io_result_bits_self_hit; // @[Slice.scala 555:30]
  assign c_mshr_io_dirResult_bits_self_way = directory_io_result_bits_self_way; // @[Slice.scala 555:30]
  assign c_mshr_io_dirResult_bits_self_tag = directory_io_result_bits_self_tag; // @[Slice.scala 555:30]
  assign c_mshr_io_dirResult_bits_clients_states_0_state = directory_io_result_bits_clients_states_0_state; // @[Slice.scala 555:30]
  assign c_mshr_io_dirResult_bits_clients_states_0_hit = directory_io_result_bits_clients_states_0_hit; // @[Slice.scala 555:30]
  assign c_mshr_io_dirResult_bits_clients_states_1_state = directory_io_result_bits_clients_states_1_state; // @[Slice.scala 555:30]
  assign c_mshr_io_dirResult_bits_clients_states_1_hit = directory_io_result_bits_clients_states_1_hit; // @[Slice.scala 555:30]
  assign c_mshr_io_dirResult_bits_clients_tag = directory_io_result_bits_clients_tag; // @[Slice.scala 555:30]
  assign c_mshr_io_dirResult_bits_clients_way = directory_io_result_bits_clients_way; // @[Slice.scala 555:30]
  assign c_mshr_io_c_status_set = 10'h0; // @[Slice.scala 244:28]
  assign c_mshr_io_c_status_tag = 20'h0; // @[Slice.scala 245:28]
  assign c_mshr_io_c_status_way = 3'h0; // @[Slice.scala 246:28]
  assign c_mshr_io_c_status_nestedReleaseData = 1'h0; // @[Slice.scala 247:42]
  assign c_mshr_io_bstatus_set = 10'h0; // @[Slice.scala 248:28]
  assign c_mshr_io_bstatus_tag = 20'h0; // @[Slice.scala 249:28]
  assign c_mshr_io_bstatus_way = 3'h0; // @[Slice.scala 250:28]
  assign c_mshr_io_bstatus_nestedProbeAckData = 1'h0; // @[Slice.scala 251:43]
  assign c_mshr_io_bstatus_probeHelperFinish = 1'h0; // @[Slice.scala 252:42]
  assign c_mshr_io_releaseThrough = |_ms_15_io_releaseThrough_T; // @[Slice.scala 368:12]
  assign c_mshr_io_probeAckDataThrough = 1'h0; // @[Slice.scala 365:35]
  assign dataStorage_clock = clock;
  assign dataStorage_reset = reset;
  assign dataStorage_io_sourceC_raddr_valid = sourceC_io_bs_raddr_valid; // @[Slice.scala 113:32]
  assign dataStorage_io_sourceC_raddr_bits_way = sourceC_io_bs_raddr_bits_way; // @[Slice.scala 113:32]
  assign dataStorage_io_sourceC_raddr_bits_set = sourceC_io_bs_raddr_bits_set; // @[Slice.scala 113:32]
  assign dataStorage_io_sourceC_raddr_bits_beat = sourceC_io_bs_raddr_bits_beat; // @[Slice.scala 113:32]
  assign dataStorage_io_sinkD_waddr_valid = sinkD_io_bs_waddr_valid; // @[Slice.scala 104:30]
  assign dataStorage_io_sinkD_waddr_bits_way = sinkD_io_bs_waddr_bits_way; // @[Slice.scala 104:30]
  assign dataStorage_io_sinkD_waddr_bits_set = sinkD_io_bs_waddr_bits_set; // @[Slice.scala 104:30]
  assign dataStorage_io_sinkD_waddr_bits_beat = sinkD_io_bs_waddr_bits_beat; // @[Slice.scala 104:30]
  assign dataStorage_io_sinkD_waddr_bits_noop = sinkD_io_bs_waddr_bits_noop; // @[Slice.scala 104:30]
  assign dataStorage_io_sinkD_wdata_data = sinkD_io_bs_wdata_data; // @[Slice.scala 103:30]
  assign dataStorage_io_sourceD_raddr_valid = sourceD_io_bs_raddr_valid; // @[Slice.scala 110:32]
  assign dataStorage_io_sourceD_raddr_bits_way = sourceD_io_bs_raddr_bits_way; // @[Slice.scala 110:32]
  assign dataStorage_io_sourceD_raddr_bits_set = sourceD_io_bs_raddr_bits_set; // @[Slice.scala 110:32]
  assign dataStorage_io_sourceD_raddr_bits_beat = sourceD_io_bs_raddr_bits_beat; // @[Slice.scala 110:32]
  assign dataStorage_io_sourceD_waddr_valid = sourceD_io_bs_waddr_valid; // @[Slice.scala 111:32]
  assign dataStorage_io_sourceD_waddr_bits_way = sourceD_io_bs_waddr_bits_way; // @[Slice.scala 111:32]
  assign dataStorage_io_sourceD_waddr_bits_set = sourceD_io_bs_waddr_bits_set; // @[Slice.scala 111:32]
  assign dataStorage_io_sourceD_waddr_bits_beat = sourceD_io_bs_waddr_bits_beat; // @[Slice.scala 111:32]
  assign dataStorage_io_sourceD_wdata_data = sourceD_io_bs_wdata_data; // @[Slice.scala 112:32]
  assign dataStorage_io_sinkC_waddr_valid = sinkC_io_bs_waddr_valid; // @[Slice.scala 114:30]
  assign dataStorage_io_sinkC_waddr_bits_way = sinkC_io_bs_waddr_bits_way; // @[Slice.scala 114:30]
  assign dataStorage_io_sinkC_waddr_bits_set = sinkC_io_bs_waddr_bits_set; // @[Slice.scala 114:30]
  assign dataStorage_io_sinkC_waddr_bits_beat = sinkC_io_bs_waddr_bits_beat; // @[Slice.scala 114:30]
  assign dataStorage_io_sinkC_waddr_bits_noop = sinkC_io_bs_waddr_bits_noop; // @[Slice.scala 114:30]
  assign dataStorage_io_sinkC_wdata_data = sinkC_io_bs_wdata_data; // @[Slice.scala 115:30]
  assign mshrAlloc_io_a_req_valid = a_req_buffer_io_out_valid; // @[Slice.scala 150:22]
  assign mshrAlloc_io_a_req_bits_channel = a_req_buffer_io_out_bits_channel; // @[Slice.scala 150:22]
  assign mshrAlloc_io_a_req_bits_opcode = a_req_buffer_io_out_bits_opcode; // @[Slice.scala 150:22]
  assign mshrAlloc_io_a_req_bits_param = a_req_buffer_io_out_bits_param; // @[Slice.scala 150:22]
  assign mshrAlloc_io_a_req_bits_size = a_req_buffer_io_out_bits_size; // @[Slice.scala 150:22]
  assign mshrAlloc_io_a_req_bits_source = a_req_buffer_io_out_bits_source; // @[Slice.scala 150:22]
  assign mshrAlloc_io_a_req_bits_set = a_req_buffer_io_out_bits_set; // @[Slice.scala 150:22]
  assign mshrAlloc_io_a_req_bits_tag = a_req_buffer_io_out_bits_tag; // @[Slice.scala 150:22]
  assign mshrAlloc_io_a_req_bits_off = a_req_buffer_io_out_bits_off; // @[Slice.scala 150:22]
  assign mshrAlloc_io_a_req_bits_mask = a_req_buffer_io_out_bits_mask; // @[Slice.scala 150:22]
  assign mshrAlloc_io_a_req_bits_bufIdx = a_req_buffer_io_out_bits_bufIdx; // @[Slice.scala 150:22]
  assign mshrAlloc_io_a_req_bits_preferCache = a_req_buffer_io_out_bits_preferCache; // @[Slice.scala 150:22]
  assign mshrAlloc_io_a_req_bits_dirty = a_req_buffer_io_out_bits_dirty; // @[Slice.scala 150:22]
  assign mshrAlloc_io_a_req_bits_fromProbeHelper = a_req_buffer_io_out_bits_fromProbeHelper; // @[Slice.scala 150:22]
  assign mshrAlloc_io_a_req_bits_fromCmoHelper = a_req_buffer_io_out_bits_fromCmoHelper; // @[Slice.scala 150:22]
  assign mshrAlloc_io_a_req_bits_needProbeAckData = a_req_buffer_io_out_bits_needProbeAckData; // @[Slice.scala 150:22]
  assign mshrAlloc_io_breq_valid = b_arb_io_out_valid; // @[Slice.scala 139:24]
  assign mshrAlloc_io_breq_bits_channel = b_arb_io_out_bits_channel; // @[Slice.scala 139:24]
  assign mshrAlloc_io_breq_bits_opcode = b_arb_io_out_bits_opcode; // @[Slice.scala 139:24]
  assign mshrAlloc_io_breq_bits_param = b_arb_io_out_bits_param; // @[Slice.scala 139:24]
  assign mshrAlloc_io_breq_bits_size = b_arb_io_out_bits_size; // @[Slice.scala 139:24]
  assign mshrAlloc_io_breq_bits_source = b_arb_io_out_bits_source; // @[Slice.scala 139:24]
  assign mshrAlloc_io_breq_bits_set = b_arb_io_out_bits_set; // @[Slice.scala 139:24]
  assign mshrAlloc_io_breq_bits_tag = b_arb_io_out_bits_tag; // @[Slice.scala 139:24]
  assign mshrAlloc_io_breq_bits_off = b_arb_io_out_bits_off; // @[Slice.scala 139:24]
  assign mshrAlloc_io_breq_bits_mask = b_arb_io_out_bits_mask; // @[Slice.scala 139:24]
  assign mshrAlloc_io_breq_bits_bufIdx = b_arb_io_out_bits_bufIdx; // @[Slice.scala 139:24]
  assign mshrAlloc_io_breq_bits_preferCache = b_arb_io_out_bits_preferCache; // @[Slice.scala 139:24]
  assign mshrAlloc_io_breq_bits_dirty = b_arb_io_out_bits_dirty; // @[Slice.scala 139:24]
  assign mshrAlloc_io_breq_bits_fromProbeHelper = b_arb_io_out_bits_fromProbeHelper; // @[Slice.scala 139:24]
  assign mshrAlloc_io_breq_bits_fromCmoHelper = b_arb_io_out_bits_fromCmoHelper; // @[Slice.scala 139:24]
  assign mshrAlloc_io_breq_bits_needProbeAckData = b_arb_io_out_bits_needProbeAckData; // @[Slice.scala 139:24]
  assign mshrAlloc_io_c_req_valid = sinkC_io_alloc_valid; // @[Slice.scala 161:24]
  assign mshrAlloc_io_c_req_bits_opcode = sinkC_io_alloc_bits_opcode; // @[Slice.scala 161:24]
  assign mshrAlloc_io_c_req_bits_param = sinkC_io_alloc_bits_param; // @[Slice.scala 161:24]
  assign mshrAlloc_io_c_req_bits_size = sinkC_io_alloc_bits_size; // @[Slice.scala 161:24]
  assign mshrAlloc_io_c_req_bits_source = sinkC_io_alloc_bits_source; // @[Slice.scala 161:24]
  assign mshrAlloc_io_c_req_bits_set = sinkC_io_alloc_bits_set; // @[Slice.scala 161:24]
  assign mshrAlloc_io_c_req_bits_tag = sinkC_io_alloc_bits_tag; // @[Slice.scala 161:24]
  assign mshrAlloc_io_c_req_bits_off = sinkC_io_alloc_bits_off; // @[Slice.scala 161:24]
  assign mshrAlloc_io_c_req_bits_bufIdx = sinkC_io_alloc_bits_bufIdx; // @[Slice.scala 161:24]
  assign mshrAlloc_io_c_req_bits_dirty = sinkC_io_alloc_bits_dirty; // @[Slice.scala 161:24]
  assign mshrAlloc_io_status_0_valid = abc_mshr_0_io_status_valid; // @[Slice.scala 168:30]
  assign mshrAlloc_io_status_0_bits_set = abc_mshr_0_io_status_bits_set; // @[Slice.scala 168:30]
  assign mshrAlloc_io_status_0_bits_nestB = abc_mshr_0_io_status_bits_nestB; // @[Slice.scala 168:30]
  assign mshrAlloc_io_status_0_bits_nestC = abc_mshr_0_io_status_bits_nestC; // @[Slice.scala 168:30]
  assign mshrAlloc_io_status_1_valid = abc_mshr_1_io_status_valid; // @[Slice.scala 168:30]
  assign mshrAlloc_io_status_1_bits_set = abc_mshr_1_io_status_bits_set; // @[Slice.scala 168:30]
  assign mshrAlloc_io_status_1_bits_nestB = abc_mshr_1_io_status_bits_nestB; // @[Slice.scala 168:30]
  assign mshrAlloc_io_status_1_bits_nestC = abc_mshr_1_io_status_bits_nestC; // @[Slice.scala 168:30]
  assign mshrAlloc_io_status_2_valid = abc_mshr_2_io_status_valid; // @[Slice.scala 168:30]
  assign mshrAlloc_io_status_2_bits_set = abc_mshr_2_io_status_bits_set; // @[Slice.scala 168:30]
  assign mshrAlloc_io_status_2_bits_nestB = abc_mshr_2_io_status_bits_nestB; // @[Slice.scala 168:30]
  assign mshrAlloc_io_status_2_bits_nestC = abc_mshr_2_io_status_bits_nestC; // @[Slice.scala 168:30]
  assign mshrAlloc_io_status_3_valid = abc_mshr_3_io_status_valid; // @[Slice.scala 168:30]
  assign mshrAlloc_io_status_3_bits_set = abc_mshr_3_io_status_bits_set; // @[Slice.scala 168:30]
  assign mshrAlloc_io_status_3_bits_nestB = abc_mshr_3_io_status_bits_nestB; // @[Slice.scala 168:30]
  assign mshrAlloc_io_status_3_bits_nestC = abc_mshr_3_io_status_bits_nestC; // @[Slice.scala 168:30]
  assign mshrAlloc_io_status_4_valid = abc_mshr_4_io_status_valid; // @[Slice.scala 168:30]
  assign mshrAlloc_io_status_4_bits_set = abc_mshr_4_io_status_bits_set; // @[Slice.scala 168:30]
  assign mshrAlloc_io_status_4_bits_nestB = abc_mshr_4_io_status_bits_nestB; // @[Slice.scala 168:30]
  assign mshrAlloc_io_status_4_bits_nestC = abc_mshr_4_io_status_bits_nestC; // @[Slice.scala 168:30]
  assign mshrAlloc_io_status_5_valid = abc_mshr_5_io_status_valid; // @[Slice.scala 168:30]
  assign mshrAlloc_io_status_5_bits_set = abc_mshr_5_io_status_bits_set; // @[Slice.scala 168:30]
  assign mshrAlloc_io_status_5_bits_nestB = abc_mshr_5_io_status_bits_nestB; // @[Slice.scala 168:30]
  assign mshrAlloc_io_status_5_bits_nestC = abc_mshr_5_io_status_bits_nestC; // @[Slice.scala 168:30]
  assign mshrAlloc_io_status_6_valid = abc_mshr_6_io_status_valid; // @[Slice.scala 168:30]
  assign mshrAlloc_io_status_6_bits_set = abc_mshr_6_io_status_bits_set; // @[Slice.scala 168:30]
  assign mshrAlloc_io_status_6_bits_nestB = abc_mshr_6_io_status_bits_nestB; // @[Slice.scala 168:30]
  assign mshrAlloc_io_status_6_bits_nestC = abc_mshr_6_io_status_bits_nestC; // @[Slice.scala 168:30]
  assign mshrAlloc_io_status_7_valid = abc_mshr_7_io_status_valid; // @[Slice.scala 168:30]
  assign mshrAlloc_io_status_7_bits_set = abc_mshr_7_io_status_bits_set; // @[Slice.scala 168:30]
  assign mshrAlloc_io_status_7_bits_nestB = abc_mshr_7_io_status_bits_nestB; // @[Slice.scala 168:30]
  assign mshrAlloc_io_status_7_bits_nestC = abc_mshr_7_io_status_bits_nestC; // @[Slice.scala 168:30]
  assign mshrAlloc_io_status_8_valid = abc_mshr_8_io_status_valid; // @[Slice.scala 168:30]
  assign mshrAlloc_io_status_8_bits_set = abc_mshr_8_io_status_bits_set; // @[Slice.scala 168:30]
  assign mshrAlloc_io_status_8_bits_nestB = abc_mshr_8_io_status_bits_nestB; // @[Slice.scala 168:30]
  assign mshrAlloc_io_status_8_bits_nestC = abc_mshr_8_io_status_bits_nestC; // @[Slice.scala 168:30]
  assign mshrAlloc_io_status_9_valid = abc_mshr_9_io_status_valid; // @[Slice.scala 168:30]
  assign mshrAlloc_io_status_9_bits_set = abc_mshr_9_io_status_bits_set; // @[Slice.scala 168:30]
  assign mshrAlloc_io_status_9_bits_nestB = abc_mshr_9_io_status_bits_nestB; // @[Slice.scala 168:30]
  assign mshrAlloc_io_status_9_bits_nestC = abc_mshr_9_io_status_bits_nestC; // @[Slice.scala 168:30]
  assign mshrAlloc_io_status_10_valid = abc_mshr_10_io_status_valid; // @[Slice.scala 168:30]
  assign mshrAlloc_io_status_10_bits_set = abc_mshr_10_io_status_bits_set; // @[Slice.scala 168:30]
  assign mshrAlloc_io_status_10_bits_nestB = abc_mshr_10_io_status_bits_nestB; // @[Slice.scala 168:30]
  assign mshrAlloc_io_status_10_bits_nestC = abc_mshr_10_io_status_bits_nestC; // @[Slice.scala 168:30]
  assign mshrAlloc_io_status_11_valid = abc_mshr_11_io_status_valid; // @[Slice.scala 168:30]
  assign mshrAlloc_io_status_11_bits_set = abc_mshr_11_io_status_bits_set; // @[Slice.scala 168:30]
  assign mshrAlloc_io_status_11_bits_nestB = abc_mshr_11_io_status_bits_nestB; // @[Slice.scala 168:30]
  assign mshrAlloc_io_status_11_bits_nestC = abc_mshr_11_io_status_bits_nestC; // @[Slice.scala 168:30]
  assign mshrAlloc_io_status_12_valid = abc_mshr_12_io_status_valid; // @[Slice.scala 168:30]
  assign mshrAlloc_io_status_12_bits_set = abc_mshr_12_io_status_bits_set; // @[Slice.scala 168:30]
  assign mshrAlloc_io_status_12_bits_nestB = abc_mshr_12_io_status_bits_nestB; // @[Slice.scala 168:30]
  assign mshrAlloc_io_status_12_bits_nestC = abc_mshr_12_io_status_bits_nestC; // @[Slice.scala 168:30]
  assign mshrAlloc_io_status_13_valid = abc_mshr_13_io_status_valid; // @[Slice.scala 168:30]
  assign mshrAlloc_io_status_13_bits_set = abc_mshr_13_io_status_bits_set; // @[Slice.scala 168:30]
  assign mshrAlloc_io_status_13_bits_nestB = abc_mshr_13_io_status_bits_nestB; // @[Slice.scala 168:30]
  assign mshrAlloc_io_status_13_bits_nestC = abc_mshr_13_io_status_bits_nestC; // @[Slice.scala 168:30]
  assign mshrAlloc_io_status_14_valid = bc_mshr_io_status_valid; // @[Slice.scala 168:30]
  assign mshrAlloc_io_status_14_bits_set = bc_mshr_io_status_bits_set; // @[Slice.scala 168:30]
  assign mshrAlloc_io_status_14_bits_nestC = bc_mshr_io_status_bits_nestC; // @[Slice.scala 168:30]
  assign mshrAlloc_io_status_15_valid = c_mshr_io_status_valid; // @[Slice.scala 168:30]
  assign mshrAlloc_io_status_15_bits_set = c_mshr_io_status_bits_set; // @[Slice.scala 168:30]
  assign mshrAlloc_io_dirRead_ready = directory_io_read_ready; // @[Slice.scala 376:21]
  assign a_req_buffer_clock = clock;
  assign a_req_buffer_reset = reset;
  assign a_req_buffer_io_in_valid = ~probeHelperOpt_io_full & sinkA_io_alloc_valid; // @[Slice.scala 389:26]
  assign a_req_buffer_io_in_bits_opcode = sinkA_io_alloc_bits_opcode; // @[Slice.scala 129:19 390:15]
  assign a_req_buffer_io_in_bits_param = sinkA_io_alloc_bits_param; // @[Slice.scala 129:19 390:15]
  assign a_req_buffer_io_in_bits_size = sinkA_io_alloc_bits_size; // @[Slice.scala 129:19 390:15]
  assign a_req_buffer_io_in_bits_source = sinkA_io_alloc_bits_source; // @[Slice.scala 129:19 390:15]
  assign a_req_buffer_io_in_bits_set = sinkA_io_alloc_bits_set; // @[Slice.scala 129:19 390:15]
  assign a_req_buffer_io_in_bits_tag = sinkA_io_alloc_bits_tag; // @[Slice.scala 129:19 390:15]
  assign a_req_buffer_io_in_bits_off = sinkA_io_alloc_bits_off; // @[Slice.scala 129:19 390:15]
  assign a_req_buffer_io_in_bits_mask = sinkA_io_alloc_bits_mask; // @[Slice.scala 129:19 390:15]
  assign a_req_buffer_io_in_bits_bufIdx = sinkA_io_alloc_bits_bufIdx; // @[Slice.scala 129:19 390:15]
  assign a_req_buffer_io_in_bits_preferCache = sinkA_io_alloc_bits_preferCache; // @[Slice.scala 129:19 390:15]
  assign a_req_buffer_io_out_ready = mshrAlloc_io_a_req_ready; // @[Slice.scala 150:22]
  assign a_req_buffer_io_mshr_status_0_valid = abc_mshr_0_io_status_valid; // @[Slice.scala 177:38]
  assign a_req_buffer_io_mshr_status_0_bits_set = abc_mshr_0_io_status_bits_set; // @[Slice.scala 177:38]
  assign a_req_buffer_io_mshr_status_0_bits_will_free = abc_mshr_0_io_status_bits_will_free; // @[Slice.scala 177:38]
  assign a_req_buffer_io_mshr_status_1_valid = abc_mshr_1_io_status_valid; // @[Slice.scala 177:38]
  assign a_req_buffer_io_mshr_status_1_bits_set = abc_mshr_1_io_status_bits_set; // @[Slice.scala 177:38]
  assign a_req_buffer_io_mshr_status_1_bits_will_free = abc_mshr_1_io_status_bits_will_free; // @[Slice.scala 177:38]
  assign a_req_buffer_io_mshr_status_2_valid = abc_mshr_2_io_status_valid; // @[Slice.scala 177:38]
  assign a_req_buffer_io_mshr_status_2_bits_set = abc_mshr_2_io_status_bits_set; // @[Slice.scala 177:38]
  assign a_req_buffer_io_mshr_status_2_bits_will_free = abc_mshr_2_io_status_bits_will_free; // @[Slice.scala 177:38]
  assign a_req_buffer_io_mshr_status_3_valid = abc_mshr_3_io_status_valid; // @[Slice.scala 177:38]
  assign a_req_buffer_io_mshr_status_3_bits_set = abc_mshr_3_io_status_bits_set; // @[Slice.scala 177:38]
  assign a_req_buffer_io_mshr_status_3_bits_will_free = abc_mshr_3_io_status_bits_will_free; // @[Slice.scala 177:38]
  assign a_req_buffer_io_mshr_status_4_valid = abc_mshr_4_io_status_valid; // @[Slice.scala 177:38]
  assign a_req_buffer_io_mshr_status_4_bits_set = abc_mshr_4_io_status_bits_set; // @[Slice.scala 177:38]
  assign a_req_buffer_io_mshr_status_4_bits_will_free = abc_mshr_4_io_status_bits_will_free; // @[Slice.scala 177:38]
  assign a_req_buffer_io_mshr_status_5_valid = abc_mshr_5_io_status_valid; // @[Slice.scala 177:38]
  assign a_req_buffer_io_mshr_status_5_bits_set = abc_mshr_5_io_status_bits_set; // @[Slice.scala 177:38]
  assign a_req_buffer_io_mshr_status_5_bits_will_free = abc_mshr_5_io_status_bits_will_free; // @[Slice.scala 177:38]
  assign a_req_buffer_io_mshr_status_6_valid = abc_mshr_6_io_status_valid; // @[Slice.scala 177:38]
  assign a_req_buffer_io_mshr_status_6_bits_set = abc_mshr_6_io_status_bits_set; // @[Slice.scala 177:38]
  assign a_req_buffer_io_mshr_status_6_bits_will_free = abc_mshr_6_io_status_bits_will_free; // @[Slice.scala 177:38]
  assign a_req_buffer_io_mshr_status_7_valid = abc_mshr_7_io_status_valid; // @[Slice.scala 177:38]
  assign a_req_buffer_io_mshr_status_7_bits_set = abc_mshr_7_io_status_bits_set; // @[Slice.scala 177:38]
  assign a_req_buffer_io_mshr_status_7_bits_will_free = abc_mshr_7_io_status_bits_will_free; // @[Slice.scala 177:38]
  assign a_req_buffer_io_mshr_status_8_valid = abc_mshr_8_io_status_valid; // @[Slice.scala 177:38]
  assign a_req_buffer_io_mshr_status_8_bits_set = abc_mshr_8_io_status_bits_set; // @[Slice.scala 177:38]
  assign a_req_buffer_io_mshr_status_8_bits_will_free = abc_mshr_8_io_status_bits_will_free; // @[Slice.scala 177:38]
  assign a_req_buffer_io_mshr_status_9_valid = abc_mshr_9_io_status_valid; // @[Slice.scala 177:38]
  assign a_req_buffer_io_mshr_status_9_bits_set = abc_mshr_9_io_status_bits_set; // @[Slice.scala 177:38]
  assign a_req_buffer_io_mshr_status_9_bits_will_free = abc_mshr_9_io_status_bits_will_free; // @[Slice.scala 177:38]
  assign a_req_buffer_io_mshr_status_10_valid = abc_mshr_10_io_status_valid; // @[Slice.scala 177:38]
  assign a_req_buffer_io_mshr_status_10_bits_set = abc_mshr_10_io_status_bits_set; // @[Slice.scala 177:38]
  assign a_req_buffer_io_mshr_status_10_bits_will_free = abc_mshr_10_io_status_bits_will_free; // @[Slice.scala 177:38]
  assign a_req_buffer_io_mshr_status_11_valid = abc_mshr_11_io_status_valid; // @[Slice.scala 177:38]
  assign a_req_buffer_io_mshr_status_11_bits_set = abc_mshr_11_io_status_bits_set; // @[Slice.scala 177:38]
  assign a_req_buffer_io_mshr_status_11_bits_will_free = abc_mshr_11_io_status_bits_will_free; // @[Slice.scala 177:38]
  assign a_req_buffer_io_mshr_status_12_valid = abc_mshr_12_io_status_valid; // @[Slice.scala 177:38]
  assign a_req_buffer_io_mshr_status_12_bits_set = abc_mshr_12_io_status_bits_set; // @[Slice.scala 177:38]
  assign a_req_buffer_io_mshr_status_12_bits_will_free = abc_mshr_12_io_status_bits_will_free; // @[Slice.scala 177:38]
  assign a_req_buffer_io_mshr_status_13_valid = abc_mshr_13_io_status_valid; // @[Slice.scala 177:38]
  assign a_req_buffer_io_mshr_status_13_bits_set = abc_mshr_13_io_status_bits_set; // @[Slice.scala 177:38]
  assign a_req_buffer_io_mshr_status_13_bits_will_free = abc_mshr_13_io_status_bits_will_free; // @[Slice.scala 177:38]
  assign probeHelperOpt_clock = clock;
  assign probeHelperOpt_reset = reset;
  assign probeHelperOpt_io_dirResult_valid = probeHelperOpt_io_dirResult_valid_REG; // @[Slice.scala 560:26]
  assign probeHelperOpt_io_dirResult_bits_clients_states_0_state = directory_io_result_bits_clients_states_0_state; // @[Slice.scala 559:25]
  assign probeHelperOpt_io_dirResult_bits_clients_states_0_hit = directory_io_result_bits_clients_states_0_hit; // @[Slice.scala 559:25]
  assign probeHelperOpt_io_dirResult_bits_clients_states_1_state = directory_io_result_bits_clients_states_1_state; // @[Slice.scala 559:25]
  assign probeHelperOpt_io_dirResult_bits_clients_states_1_hit = directory_io_result_bits_clients_states_1_hit; // @[Slice.scala 559:25]
  assign probeHelperOpt_io_dirResult_bits_clients_tag_match = directory_io_result_bits_clients_tag_match; // @[Slice.scala 559:25]
  assign probeHelperOpt_io_dirResult_bits_clients_tag = directory_io_result_bits_clients_tag; // @[Slice.scala 559:25]
  assign probeHelperOpt_io_dirResult_bits_sourceId = directory_io_result_bits_sourceId; // @[Slice.scala 559:25]
  assign probeHelperOpt_io_dirResult_bits_set = directory_io_result_bits_set; // @[Slice.scala 559:25]
  assign probeHelperOpt_io_dirResult_bits_replacerInfo_channel = directory_io_result_bits_replacerInfo_channel; // @[Slice.scala 559:25]
  assign probeHelperOpt_io_dirResult_bits_replacerInfo_opcode = directory_io_result_bits_replacerInfo_opcode; // @[Slice.scala 559:25]
  assign probeHelperOpt_io_probe_ready = b_arb_io_in_0_ready; // @[Slice.scala 137:20]
  assign b_arb_io_in_0_valid = probeHelperOpt_io_probe_valid; // @[Slice.scala 137:20]
  assign b_arb_io_in_0_bits_channel = probeHelperOpt_io_probe_bits_channel; // @[Slice.scala 137:20]
  assign b_arb_io_in_0_bits_opcode = probeHelperOpt_io_probe_bits_opcode; // @[Slice.scala 137:20]
  assign b_arb_io_in_0_bits_param = probeHelperOpt_io_probe_bits_param; // @[Slice.scala 137:20]
  assign b_arb_io_in_0_bits_size = probeHelperOpt_io_probe_bits_size; // @[Slice.scala 137:20]
  assign b_arb_io_in_0_bits_source = probeHelperOpt_io_probe_bits_source; // @[Slice.scala 137:20]
  assign b_arb_io_in_0_bits_set = probeHelperOpt_io_probe_bits_set; // @[Slice.scala 137:20]
  assign b_arb_io_in_0_bits_tag = probeHelperOpt_io_probe_bits_tag; // @[Slice.scala 137:20]
  assign b_arb_io_in_0_bits_off = probeHelperOpt_io_probe_bits_off; // @[Slice.scala 137:20]
  assign b_arb_io_in_0_bits_mask = probeHelperOpt_io_probe_bits_mask; // @[Slice.scala 137:20]
  assign b_arb_io_in_0_bits_bufIdx = probeHelperOpt_io_probe_bits_bufIdx; // @[Slice.scala 137:20]
  assign b_arb_io_in_0_bits_preferCache = probeHelperOpt_io_probe_bits_preferCache; // @[Slice.scala 137:20]
  assign b_arb_io_in_0_bits_dirty = probeHelperOpt_io_probe_bits_dirty; // @[Slice.scala 137:20]
  assign b_arb_io_in_0_bits_fromProbeHelper = probeHelperOpt_io_probe_bits_fromProbeHelper; // @[Slice.scala 137:20]
  assign b_arb_io_in_0_bits_fromCmoHelper = probeHelperOpt_io_probe_bits_fromCmoHelper; // @[Slice.scala 137:20]
  assign b_arb_io_in_0_bits_needProbeAckData = probeHelperOpt_io_probe_bits_needProbeAckData; // @[Slice.scala 137:20]
  assign b_arb_io_in_1_valid = sinkB_io_alloc_valid; // @[Slice.scala 138:20]
  assign b_arb_io_in_1_bits_opcode = sinkB_io_alloc_bits_opcode; // @[Slice.scala 138:20]
  assign b_arb_io_in_1_bits_param = sinkB_io_alloc_bits_param; // @[Slice.scala 138:20]
  assign b_arb_io_in_1_bits_size = sinkB_io_alloc_bits_size; // @[Slice.scala 138:20]
  assign b_arb_io_in_1_bits_source = sinkB_io_alloc_bits_source; // @[Slice.scala 138:20]
  assign b_arb_io_in_1_bits_set = sinkB_io_alloc_bits_set; // @[Slice.scala 138:20]
  assign b_arb_io_in_1_bits_tag = sinkB_io_alloc_bits_tag; // @[Slice.scala 138:20]
  assign b_arb_io_in_1_bits_off = sinkB_io_alloc_bits_off; // @[Slice.scala 138:20]
  assign b_arb_io_in_1_bits_mask = sinkB_io_alloc_bits_mask; // @[Slice.scala 138:20]
  assign b_arb_io_in_1_bits_needProbeAckData = sinkB_io_alloc_bits_needProbeAckData; // @[Slice.scala 138:20]
  assign b_arb_io_out_ready = mshrAlloc_io_breq_ready; // @[Slice.scala 139:24]
  assign directory_clock = clock;
  assign directory_reset = reset;
  assign directory_io_read_valid = mshrAlloc_io_dirRead_valid; // @[Slice.scala 376:21]
  assign directory_io_read_bits_idOH = mshrAlloc_io_dirRead_bits_idOH; // @[Slice.scala 376:21]
  assign directory_io_read_bits_tag = mshrAlloc_io_dirRead_bits_tag; // @[Slice.scala 376:21]
  assign directory_io_read_bits_set = mshrAlloc_io_dirRead_bits_set; // @[Slice.scala 376:21]
  assign directory_io_read_bits_replacerInfo_channel = mshrAlloc_io_dirRead_bits_replacerInfo_channel; // @[Slice.scala 376:21]
  assign directory_io_read_bits_replacerInfo_opcode = mshrAlloc_io_dirRead_bits_replacerInfo_opcode; // @[Slice.scala 376:21]
  assign directory_io_read_bits_source = mshrAlloc_io_dirRead_bits_source; // @[Slice.scala 376:21]
  assign directory_io_dirWReq_valid = pipeline_io_out_valid; // @[Pipeline.scala 41:9]
  assign directory_io_dirWReq_bits_set = pipeline_io_out_bits_set; // @[Pipeline.scala 41:9]
  assign directory_io_dirWReq_bits_way = pipeline_io_out_bits_way; // @[Pipeline.scala 41:9]
  assign directory_io_dirWReq_bits_data_dirty = pipeline_io_out_bits_data_dirty; // @[Pipeline.scala 41:9]
  assign directory_io_dirWReq_bits_data_state = pipeline_io_out_bits_data_state; // @[Pipeline.scala 41:9]
  assign directory_io_dirWReq_bits_data_clientStates_0 = pipeline_io_out_bits_data_clientStates_0; // @[Pipeline.scala 41:9]
  assign directory_io_dirWReq_bits_data_clientStates_1 = pipeline_io_out_bits_data_clientStates_1; // @[Pipeline.scala 41:9]
  assign directory_io_tagWReq_valid = pipeline_1_io_out_valid; // @[Pipeline.scala 41:9]
  assign directory_io_tagWReq_bits_set = pipeline_1_io_out_bits_set; // @[Pipeline.scala 41:9]
  assign directory_io_tagWReq_bits_way = pipeline_1_io_out_bits_way; // @[Pipeline.scala 41:9]
  assign directory_io_tagWReq_bits_tag = pipeline_1_io_out_bits_tag; // @[Pipeline.scala 41:9]
  assign directory_io_clientDirWReq_valid = pipeline_2_io_out_valid; // @[Pipeline.scala 41:9]
  assign directory_io_clientDirWReq_bits_set = pipeline_2_io_out_bits_set; // @[Pipeline.scala 41:9]
  assign directory_io_clientDirWReq_bits_way = pipeline_2_io_out_bits_way; // @[Pipeline.scala 41:9]
  assign directory_io_clientDirWReq_bits_data_0_state = pipeline_2_io_out_bits_data_0_state; // @[Pipeline.scala 41:9]
  assign directory_io_clientDirWReq_bits_data_1_state = pipeline_2_io_out_bits_data_1_state; // @[Pipeline.scala 41:9]
  assign directory_io_clientTagWreq_valid = pipeline_3_io_out_valid; // @[Pipeline.scala 41:9]
  assign directory_io_clientTagWreq_bits_set = pipeline_3_io_out_bits_set; // @[Pipeline.scala 41:9]
  assign directory_io_clientTagWreq_bits_way = pipeline_3_io_out_bits_way; // @[Pipeline.scala 41:9]
  assign directory_io_clientTagWreq_bits_tag = pipeline_3_io_out_bits_tag; // @[Pipeline.scala 41:9]
  assign pipeline_clock = clock;
  assign pipeline_reset = reset;
  assign pipeline_io_in_valid = arbiter_io_out_valid; // @[Slice.scala 409:10]
  assign pipeline_io_in_bits_set = arbiter_io_out_bits_set; // @[Slice.scala 409:10]
  assign pipeline_io_in_bits_way = arbiter_io_out_bits_way; // @[Slice.scala 409:10]
  assign pipeline_io_in_bits_data_dirty = arbiter_io_out_bits_data_dirty; // @[Slice.scala 409:10]
  assign pipeline_io_in_bits_data_state = arbiter_io_out_bits_data_state; // @[Slice.scala 409:10]
  assign pipeline_io_in_bits_data_clientStates_0 = arbiter_io_out_bits_data_clientStates_0; // @[Slice.scala 409:10]
  assign pipeline_io_in_bits_data_clientStates_1 = arbiter_io_out_bits_data_clientStates_1; // @[Slice.scala 409:10]
  assign arbiter_clock = clock;
  assign arbiter_reset = reset;
  assign arbiter_io_in_0_valid = abc_mshr_0_io_tasks_dir_write_valid; // @[Slice.scala 406:60]
  assign arbiter_io_in_0_bits_set = abc_mshr_0_io_tasks_dir_write_bits_set; // @[Slice.scala 406:60]
  assign arbiter_io_in_0_bits_way = abc_mshr_0_io_tasks_dir_write_bits_way; // @[Slice.scala 406:60]
  assign arbiter_io_in_0_bits_data_dirty = abc_mshr_0_io_tasks_dir_write_bits_data_dirty; // @[Slice.scala 406:60]
  assign arbiter_io_in_0_bits_data_state = abc_mshr_0_io_tasks_dir_write_bits_data_state; // @[Slice.scala 406:60]
  assign arbiter_io_in_0_bits_data_clientStates_0 = abc_mshr_0_io_tasks_dir_write_bits_data_clientStates_0; // @[Slice.scala 406:60]
  assign arbiter_io_in_0_bits_data_clientStates_1 = abc_mshr_0_io_tasks_dir_write_bits_data_clientStates_1; // @[Slice.scala 406:60]
  assign arbiter_io_in_1_valid = abc_mshr_1_io_tasks_dir_write_valid; // @[Slice.scala 406:60]
  assign arbiter_io_in_1_bits_set = abc_mshr_1_io_tasks_dir_write_bits_set; // @[Slice.scala 406:60]
  assign arbiter_io_in_1_bits_way = abc_mshr_1_io_tasks_dir_write_bits_way; // @[Slice.scala 406:60]
  assign arbiter_io_in_1_bits_data_dirty = abc_mshr_1_io_tasks_dir_write_bits_data_dirty; // @[Slice.scala 406:60]
  assign arbiter_io_in_1_bits_data_state = abc_mshr_1_io_tasks_dir_write_bits_data_state; // @[Slice.scala 406:60]
  assign arbiter_io_in_1_bits_data_clientStates_0 = abc_mshr_1_io_tasks_dir_write_bits_data_clientStates_0; // @[Slice.scala 406:60]
  assign arbiter_io_in_1_bits_data_clientStates_1 = abc_mshr_1_io_tasks_dir_write_bits_data_clientStates_1; // @[Slice.scala 406:60]
  assign arbiter_io_in_2_valid = abc_mshr_2_io_tasks_dir_write_valid; // @[Slice.scala 406:60]
  assign arbiter_io_in_2_bits_set = abc_mshr_2_io_tasks_dir_write_bits_set; // @[Slice.scala 406:60]
  assign arbiter_io_in_2_bits_way = abc_mshr_2_io_tasks_dir_write_bits_way; // @[Slice.scala 406:60]
  assign arbiter_io_in_2_bits_data_dirty = abc_mshr_2_io_tasks_dir_write_bits_data_dirty; // @[Slice.scala 406:60]
  assign arbiter_io_in_2_bits_data_state = abc_mshr_2_io_tasks_dir_write_bits_data_state; // @[Slice.scala 406:60]
  assign arbiter_io_in_2_bits_data_clientStates_0 = abc_mshr_2_io_tasks_dir_write_bits_data_clientStates_0; // @[Slice.scala 406:60]
  assign arbiter_io_in_2_bits_data_clientStates_1 = abc_mshr_2_io_tasks_dir_write_bits_data_clientStates_1; // @[Slice.scala 406:60]
  assign arbiter_io_in_3_valid = abc_mshr_3_io_tasks_dir_write_valid; // @[Slice.scala 406:60]
  assign arbiter_io_in_3_bits_set = abc_mshr_3_io_tasks_dir_write_bits_set; // @[Slice.scala 406:60]
  assign arbiter_io_in_3_bits_way = abc_mshr_3_io_tasks_dir_write_bits_way; // @[Slice.scala 406:60]
  assign arbiter_io_in_3_bits_data_dirty = abc_mshr_3_io_tasks_dir_write_bits_data_dirty; // @[Slice.scala 406:60]
  assign arbiter_io_in_3_bits_data_state = abc_mshr_3_io_tasks_dir_write_bits_data_state; // @[Slice.scala 406:60]
  assign arbiter_io_in_3_bits_data_clientStates_0 = abc_mshr_3_io_tasks_dir_write_bits_data_clientStates_0; // @[Slice.scala 406:60]
  assign arbiter_io_in_3_bits_data_clientStates_1 = abc_mshr_3_io_tasks_dir_write_bits_data_clientStates_1; // @[Slice.scala 406:60]
  assign arbiter_io_in_4_valid = abc_mshr_4_io_tasks_dir_write_valid; // @[Slice.scala 406:60]
  assign arbiter_io_in_4_bits_set = abc_mshr_4_io_tasks_dir_write_bits_set; // @[Slice.scala 406:60]
  assign arbiter_io_in_4_bits_way = abc_mshr_4_io_tasks_dir_write_bits_way; // @[Slice.scala 406:60]
  assign arbiter_io_in_4_bits_data_dirty = abc_mshr_4_io_tasks_dir_write_bits_data_dirty; // @[Slice.scala 406:60]
  assign arbiter_io_in_4_bits_data_state = abc_mshr_4_io_tasks_dir_write_bits_data_state; // @[Slice.scala 406:60]
  assign arbiter_io_in_4_bits_data_clientStates_0 = abc_mshr_4_io_tasks_dir_write_bits_data_clientStates_0; // @[Slice.scala 406:60]
  assign arbiter_io_in_4_bits_data_clientStates_1 = abc_mshr_4_io_tasks_dir_write_bits_data_clientStates_1; // @[Slice.scala 406:60]
  assign arbiter_io_in_5_valid = abc_mshr_5_io_tasks_dir_write_valid; // @[Slice.scala 406:60]
  assign arbiter_io_in_5_bits_set = abc_mshr_5_io_tasks_dir_write_bits_set; // @[Slice.scala 406:60]
  assign arbiter_io_in_5_bits_way = abc_mshr_5_io_tasks_dir_write_bits_way; // @[Slice.scala 406:60]
  assign arbiter_io_in_5_bits_data_dirty = abc_mshr_5_io_tasks_dir_write_bits_data_dirty; // @[Slice.scala 406:60]
  assign arbiter_io_in_5_bits_data_state = abc_mshr_5_io_tasks_dir_write_bits_data_state; // @[Slice.scala 406:60]
  assign arbiter_io_in_5_bits_data_clientStates_0 = abc_mshr_5_io_tasks_dir_write_bits_data_clientStates_0; // @[Slice.scala 406:60]
  assign arbiter_io_in_5_bits_data_clientStates_1 = abc_mshr_5_io_tasks_dir_write_bits_data_clientStates_1; // @[Slice.scala 406:60]
  assign arbiter_io_in_6_valid = abc_mshr_6_io_tasks_dir_write_valid; // @[Slice.scala 406:60]
  assign arbiter_io_in_6_bits_set = abc_mshr_6_io_tasks_dir_write_bits_set; // @[Slice.scala 406:60]
  assign arbiter_io_in_6_bits_way = abc_mshr_6_io_tasks_dir_write_bits_way; // @[Slice.scala 406:60]
  assign arbiter_io_in_6_bits_data_dirty = abc_mshr_6_io_tasks_dir_write_bits_data_dirty; // @[Slice.scala 406:60]
  assign arbiter_io_in_6_bits_data_state = abc_mshr_6_io_tasks_dir_write_bits_data_state; // @[Slice.scala 406:60]
  assign arbiter_io_in_6_bits_data_clientStates_0 = abc_mshr_6_io_tasks_dir_write_bits_data_clientStates_0; // @[Slice.scala 406:60]
  assign arbiter_io_in_6_bits_data_clientStates_1 = abc_mshr_6_io_tasks_dir_write_bits_data_clientStates_1; // @[Slice.scala 406:60]
  assign arbiter_io_in_7_valid = abc_mshr_7_io_tasks_dir_write_valid; // @[Slice.scala 406:60]
  assign arbiter_io_in_7_bits_set = abc_mshr_7_io_tasks_dir_write_bits_set; // @[Slice.scala 406:60]
  assign arbiter_io_in_7_bits_way = abc_mshr_7_io_tasks_dir_write_bits_way; // @[Slice.scala 406:60]
  assign arbiter_io_in_7_bits_data_dirty = abc_mshr_7_io_tasks_dir_write_bits_data_dirty; // @[Slice.scala 406:60]
  assign arbiter_io_in_7_bits_data_state = abc_mshr_7_io_tasks_dir_write_bits_data_state; // @[Slice.scala 406:60]
  assign arbiter_io_in_7_bits_data_clientStates_0 = abc_mshr_7_io_tasks_dir_write_bits_data_clientStates_0; // @[Slice.scala 406:60]
  assign arbiter_io_in_7_bits_data_clientStates_1 = abc_mshr_7_io_tasks_dir_write_bits_data_clientStates_1; // @[Slice.scala 406:60]
  assign arbiter_io_in_8_valid = abc_mshr_8_io_tasks_dir_write_valid; // @[Slice.scala 406:60]
  assign arbiter_io_in_8_bits_set = abc_mshr_8_io_tasks_dir_write_bits_set; // @[Slice.scala 406:60]
  assign arbiter_io_in_8_bits_way = abc_mshr_8_io_tasks_dir_write_bits_way; // @[Slice.scala 406:60]
  assign arbiter_io_in_8_bits_data_dirty = abc_mshr_8_io_tasks_dir_write_bits_data_dirty; // @[Slice.scala 406:60]
  assign arbiter_io_in_8_bits_data_state = abc_mshr_8_io_tasks_dir_write_bits_data_state; // @[Slice.scala 406:60]
  assign arbiter_io_in_8_bits_data_clientStates_0 = abc_mshr_8_io_tasks_dir_write_bits_data_clientStates_0; // @[Slice.scala 406:60]
  assign arbiter_io_in_8_bits_data_clientStates_1 = abc_mshr_8_io_tasks_dir_write_bits_data_clientStates_1; // @[Slice.scala 406:60]
  assign arbiter_io_in_9_valid = abc_mshr_9_io_tasks_dir_write_valid; // @[Slice.scala 406:60]
  assign arbiter_io_in_9_bits_set = abc_mshr_9_io_tasks_dir_write_bits_set; // @[Slice.scala 406:60]
  assign arbiter_io_in_9_bits_way = abc_mshr_9_io_tasks_dir_write_bits_way; // @[Slice.scala 406:60]
  assign arbiter_io_in_9_bits_data_dirty = abc_mshr_9_io_tasks_dir_write_bits_data_dirty; // @[Slice.scala 406:60]
  assign arbiter_io_in_9_bits_data_state = abc_mshr_9_io_tasks_dir_write_bits_data_state; // @[Slice.scala 406:60]
  assign arbiter_io_in_9_bits_data_clientStates_0 = abc_mshr_9_io_tasks_dir_write_bits_data_clientStates_0; // @[Slice.scala 406:60]
  assign arbiter_io_in_9_bits_data_clientStates_1 = abc_mshr_9_io_tasks_dir_write_bits_data_clientStates_1; // @[Slice.scala 406:60]
  assign arbiter_io_in_10_valid = abc_mshr_10_io_tasks_dir_write_valid; // @[Slice.scala 406:60]
  assign arbiter_io_in_10_bits_set = abc_mshr_10_io_tasks_dir_write_bits_set; // @[Slice.scala 406:60]
  assign arbiter_io_in_10_bits_way = abc_mshr_10_io_tasks_dir_write_bits_way; // @[Slice.scala 406:60]
  assign arbiter_io_in_10_bits_data_dirty = abc_mshr_10_io_tasks_dir_write_bits_data_dirty; // @[Slice.scala 406:60]
  assign arbiter_io_in_10_bits_data_state = abc_mshr_10_io_tasks_dir_write_bits_data_state; // @[Slice.scala 406:60]
  assign arbiter_io_in_10_bits_data_clientStates_0 = abc_mshr_10_io_tasks_dir_write_bits_data_clientStates_0; // @[Slice.scala 406:60]
  assign arbiter_io_in_10_bits_data_clientStates_1 = abc_mshr_10_io_tasks_dir_write_bits_data_clientStates_1; // @[Slice.scala 406:60]
  assign arbiter_io_in_11_valid = abc_mshr_11_io_tasks_dir_write_valid; // @[Slice.scala 406:60]
  assign arbiter_io_in_11_bits_set = abc_mshr_11_io_tasks_dir_write_bits_set; // @[Slice.scala 406:60]
  assign arbiter_io_in_11_bits_way = abc_mshr_11_io_tasks_dir_write_bits_way; // @[Slice.scala 406:60]
  assign arbiter_io_in_11_bits_data_dirty = abc_mshr_11_io_tasks_dir_write_bits_data_dirty; // @[Slice.scala 406:60]
  assign arbiter_io_in_11_bits_data_state = abc_mshr_11_io_tasks_dir_write_bits_data_state; // @[Slice.scala 406:60]
  assign arbiter_io_in_11_bits_data_clientStates_0 = abc_mshr_11_io_tasks_dir_write_bits_data_clientStates_0; // @[Slice.scala 406:60]
  assign arbiter_io_in_11_bits_data_clientStates_1 = abc_mshr_11_io_tasks_dir_write_bits_data_clientStates_1; // @[Slice.scala 406:60]
  assign arbiter_io_in_12_valid = abc_mshr_12_io_tasks_dir_write_valid; // @[Slice.scala 406:60]
  assign arbiter_io_in_12_bits_set = abc_mshr_12_io_tasks_dir_write_bits_set; // @[Slice.scala 406:60]
  assign arbiter_io_in_12_bits_way = abc_mshr_12_io_tasks_dir_write_bits_way; // @[Slice.scala 406:60]
  assign arbiter_io_in_12_bits_data_dirty = abc_mshr_12_io_tasks_dir_write_bits_data_dirty; // @[Slice.scala 406:60]
  assign arbiter_io_in_12_bits_data_state = abc_mshr_12_io_tasks_dir_write_bits_data_state; // @[Slice.scala 406:60]
  assign arbiter_io_in_12_bits_data_clientStates_0 = abc_mshr_12_io_tasks_dir_write_bits_data_clientStates_0; // @[Slice.scala 406:60]
  assign arbiter_io_in_12_bits_data_clientStates_1 = abc_mshr_12_io_tasks_dir_write_bits_data_clientStates_1; // @[Slice.scala 406:60]
  assign arbiter_io_in_13_valid = abc_mshr_13_io_tasks_dir_write_valid; // @[Slice.scala 406:60]
  assign arbiter_io_in_13_bits_set = abc_mshr_13_io_tasks_dir_write_bits_set; // @[Slice.scala 406:60]
  assign arbiter_io_in_13_bits_way = abc_mshr_13_io_tasks_dir_write_bits_way; // @[Slice.scala 406:60]
  assign arbiter_io_in_13_bits_data_dirty = abc_mshr_13_io_tasks_dir_write_bits_data_dirty; // @[Slice.scala 406:60]
  assign arbiter_io_in_13_bits_data_state = abc_mshr_13_io_tasks_dir_write_bits_data_state; // @[Slice.scala 406:60]
  assign arbiter_io_in_13_bits_data_clientStates_0 = abc_mshr_13_io_tasks_dir_write_bits_data_clientStates_0; // @[Slice.scala 406:60]
  assign arbiter_io_in_13_bits_data_clientStates_1 = abc_mshr_13_io_tasks_dir_write_bits_data_clientStates_1; // @[Slice.scala 406:60]
  assign arbiter_io_in_14_valid = _nestedWb_btoN_T & bc_mshr_io_tasks_dir_write_valid; // @[Slice.scala 389:26]
  assign arbiter_io_in_14_bits_set = bc_mshr_io_tasks_dir_write_bits_set; // @[Slice.scala 390:15]
  assign arbiter_io_in_14_bits_way = bc_mshr_io_tasks_dir_write_bits_way; // @[Slice.scala 390:15]
  assign arbiter_io_in_14_bits_data_dirty = bc_mshr_io_tasks_dir_write_bits_data_dirty; // @[Slice.scala 390:15]
  assign arbiter_io_in_14_bits_data_state = bc_mshr_io_tasks_dir_write_bits_data_state; // @[Slice.scala 390:15]
  assign arbiter_io_in_14_bits_data_clientStates_0 = bc_mshr_io_tasks_dir_write_bits_data_clientStates_0; // @[Slice.scala 390:15]
  assign arbiter_io_in_14_bits_data_clientStates_1 = bc_mshr_io_tasks_dir_write_bits_data_clientStates_1; // @[Slice.scala 390:15]
  assign arbiter_io_in_15_valid = c_mshr_io_tasks_dir_write_valid; // @[Slice.scala 408:24]
  assign arbiter_io_in_15_bits_set = c_mshr_io_tasks_dir_write_bits_set; // @[Slice.scala 408:24]
  assign arbiter_io_in_15_bits_way = c_mshr_io_tasks_dir_write_bits_way; // @[Slice.scala 408:24]
  assign arbiter_io_in_15_bits_data_dirty = c_mshr_io_tasks_dir_write_bits_data_dirty; // @[Slice.scala 408:24]
  assign arbiter_io_in_15_bits_data_state = c_mshr_io_tasks_dir_write_bits_data_state; // @[Slice.scala 408:24]
  assign arbiter_io_in_15_bits_data_clientStates_0 = c_mshr_io_tasks_dir_write_bits_data_clientStates_0; // @[Slice.scala 408:24]
  assign arbiter_io_in_15_bits_data_clientStates_1 = c_mshr_io_tasks_dir_write_bits_data_clientStates_1; // @[Slice.scala 408:24]
  assign sourceA_task_arb_clock = clock;
  assign sourceA_task_arb_reset = reset;
  assign sourceA_task_arb_io_in_0_valid = abc_mshr_0_io_tasks_source_a_valid; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_0_bits_tag = abc_mshr_0_io_tasks_source_a_bits_tag; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_0_bits_set = abc_mshr_0_io_tasks_source_a_bits_set; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_0_bits_off = abc_mshr_0_io_tasks_source_a_bits_off; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_0_bits_opcode = abc_mshr_0_io_tasks_source_a_bits_opcode; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_0_bits_param = abc_mshr_0_io_tasks_source_a_bits_param; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_0_bits_source = abc_mshr_0_io_tasks_source_a_bits_source; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_0_bits_bufIdx = abc_mshr_0_io_tasks_source_a_bits_bufIdx; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_0_bits_size = abc_mshr_0_io_tasks_source_a_bits_size; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_0_bits_putData = abc_mshr_0_io_tasks_source_a_bits_putData; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_1_valid = abc_mshr_1_io_tasks_source_a_valid; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_1_bits_tag = abc_mshr_1_io_tasks_source_a_bits_tag; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_1_bits_set = abc_mshr_1_io_tasks_source_a_bits_set; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_1_bits_off = abc_mshr_1_io_tasks_source_a_bits_off; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_1_bits_opcode = abc_mshr_1_io_tasks_source_a_bits_opcode; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_1_bits_param = abc_mshr_1_io_tasks_source_a_bits_param; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_1_bits_source = abc_mshr_1_io_tasks_source_a_bits_source; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_1_bits_bufIdx = abc_mshr_1_io_tasks_source_a_bits_bufIdx; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_1_bits_size = abc_mshr_1_io_tasks_source_a_bits_size; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_1_bits_putData = abc_mshr_1_io_tasks_source_a_bits_putData; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_2_valid = abc_mshr_2_io_tasks_source_a_valid; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_2_bits_tag = abc_mshr_2_io_tasks_source_a_bits_tag; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_2_bits_set = abc_mshr_2_io_tasks_source_a_bits_set; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_2_bits_off = abc_mshr_2_io_tasks_source_a_bits_off; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_2_bits_opcode = abc_mshr_2_io_tasks_source_a_bits_opcode; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_2_bits_param = abc_mshr_2_io_tasks_source_a_bits_param; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_2_bits_source = abc_mshr_2_io_tasks_source_a_bits_source; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_2_bits_bufIdx = abc_mshr_2_io_tasks_source_a_bits_bufIdx; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_2_bits_size = abc_mshr_2_io_tasks_source_a_bits_size; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_2_bits_putData = abc_mshr_2_io_tasks_source_a_bits_putData; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_3_valid = abc_mshr_3_io_tasks_source_a_valid; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_3_bits_tag = abc_mshr_3_io_tasks_source_a_bits_tag; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_3_bits_set = abc_mshr_3_io_tasks_source_a_bits_set; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_3_bits_off = abc_mshr_3_io_tasks_source_a_bits_off; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_3_bits_opcode = abc_mshr_3_io_tasks_source_a_bits_opcode; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_3_bits_param = abc_mshr_3_io_tasks_source_a_bits_param; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_3_bits_source = abc_mshr_3_io_tasks_source_a_bits_source; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_3_bits_bufIdx = abc_mshr_3_io_tasks_source_a_bits_bufIdx; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_3_bits_size = abc_mshr_3_io_tasks_source_a_bits_size; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_3_bits_putData = abc_mshr_3_io_tasks_source_a_bits_putData; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_4_valid = abc_mshr_4_io_tasks_source_a_valid; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_4_bits_tag = abc_mshr_4_io_tasks_source_a_bits_tag; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_4_bits_set = abc_mshr_4_io_tasks_source_a_bits_set; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_4_bits_off = abc_mshr_4_io_tasks_source_a_bits_off; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_4_bits_opcode = abc_mshr_4_io_tasks_source_a_bits_opcode; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_4_bits_param = abc_mshr_4_io_tasks_source_a_bits_param; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_4_bits_source = abc_mshr_4_io_tasks_source_a_bits_source; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_4_bits_bufIdx = abc_mshr_4_io_tasks_source_a_bits_bufIdx; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_4_bits_size = abc_mshr_4_io_tasks_source_a_bits_size; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_4_bits_putData = abc_mshr_4_io_tasks_source_a_bits_putData; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_5_valid = abc_mshr_5_io_tasks_source_a_valid; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_5_bits_tag = abc_mshr_5_io_tasks_source_a_bits_tag; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_5_bits_set = abc_mshr_5_io_tasks_source_a_bits_set; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_5_bits_off = abc_mshr_5_io_tasks_source_a_bits_off; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_5_bits_opcode = abc_mshr_5_io_tasks_source_a_bits_opcode; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_5_bits_param = abc_mshr_5_io_tasks_source_a_bits_param; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_5_bits_source = abc_mshr_5_io_tasks_source_a_bits_source; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_5_bits_bufIdx = abc_mshr_5_io_tasks_source_a_bits_bufIdx; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_5_bits_size = abc_mshr_5_io_tasks_source_a_bits_size; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_5_bits_putData = abc_mshr_5_io_tasks_source_a_bits_putData; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_6_valid = abc_mshr_6_io_tasks_source_a_valid; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_6_bits_tag = abc_mshr_6_io_tasks_source_a_bits_tag; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_6_bits_set = abc_mshr_6_io_tasks_source_a_bits_set; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_6_bits_off = abc_mshr_6_io_tasks_source_a_bits_off; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_6_bits_opcode = abc_mshr_6_io_tasks_source_a_bits_opcode; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_6_bits_param = abc_mshr_6_io_tasks_source_a_bits_param; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_6_bits_source = abc_mshr_6_io_tasks_source_a_bits_source; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_6_bits_bufIdx = abc_mshr_6_io_tasks_source_a_bits_bufIdx; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_6_bits_size = abc_mshr_6_io_tasks_source_a_bits_size; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_6_bits_putData = abc_mshr_6_io_tasks_source_a_bits_putData; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_7_valid = abc_mshr_7_io_tasks_source_a_valid; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_7_bits_tag = abc_mshr_7_io_tasks_source_a_bits_tag; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_7_bits_set = abc_mshr_7_io_tasks_source_a_bits_set; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_7_bits_off = abc_mshr_7_io_tasks_source_a_bits_off; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_7_bits_opcode = abc_mshr_7_io_tasks_source_a_bits_opcode; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_7_bits_param = abc_mshr_7_io_tasks_source_a_bits_param; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_7_bits_source = abc_mshr_7_io_tasks_source_a_bits_source; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_7_bits_bufIdx = abc_mshr_7_io_tasks_source_a_bits_bufIdx; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_7_bits_size = abc_mshr_7_io_tasks_source_a_bits_size; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_7_bits_putData = abc_mshr_7_io_tasks_source_a_bits_putData; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_8_valid = abc_mshr_8_io_tasks_source_a_valid; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_8_bits_tag = abc_mshr_8_io_tasks_source_a_bits_tag; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_8_bits_set = abc_mshr_8_io_tasks_source_a_bits_set; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_8_bits_off = abc_mshr_8_io_tasks_source_a_bits_off; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_8_bits_opcode = abc_mshr_8_io_tasks_source_a_bits_opcode; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_8_bits_param = abc_mshr_8_io_tasks_source_a_bits_param; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_8_bits_source = abc_mshr_8_io_tasks_source_a_bits_source; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_8_bits_bufIdx = abc_mshr_8_io_tasks_source_a_bits_bufIdx; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_8_bits_size = abc_mshr_8_io_tasks_source_a_bits_size; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_8_bits_putData = abc_mshr_8_io_tasks_source_a_bits_putData; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_9_valid = abc_mshr_9_io_tasks_source_a_valid; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_9_bits_tag = abc_mshr_9_io_tasks_source_a_bits_tag; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_9_bits_set = abc_mshr_9_io_tasks_source_a_bits_set; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_9_bits_off = abc_mshr_9_io_tasks_source_a_bits_off; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_9_bits_opcode = abc_mshr_9_io_tasks_source_a_bits_opcode; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_9_bits_param = abc_mshr_9_io_tasks_source_a_bits_param; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_9_bits_source = abc_mshr_9_io_tasks_source_a_bits_source; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_9_bits_bufIdx = abc_mshr_9_io_tasks_source_a_bits_bufIdx; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_9_bits_size = abc_mshr_9_io_tasks_source_a_bits_size; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_9_bits_putData = abc_mshr_9_io_tasks_source_a_bits_putData; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_10_valid = abc_mshr_10_io_tasks_source_a_valid; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_10_bits_tag = abc_mshr_10_io_tasks_source_a_bits_tag; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_10_bits_set = abc_mshr_10_io_tasks_source_a_bits_set; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_10_bits_off = abc_mshr_10_io_tasks_source_a_bits_off; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_10_bits_opcode = abc_mshr_10_io_tasks_source_a_bits_opcode; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_10_bits_param = abc_mshr_10_io_tasks_source_a_bits_param; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_10_bits_source = abc_mshr_10_io_tasks_source_a_bits_source; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_10_bits_bufIdx = abc_mshr_10_io_tasks_source_a_bits_bufIdx; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_10_bits_size = abc_mshr_10_io_tasks_source_a_bits_size; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_10_bits_putData = abc_mshr_10_io_tasks_source_a_bits_putData; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_11_valid = abc_mshr_11_io_tasks_source_a_valid; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_11_bits_tag = abc_mshr_11_io_tasks_source_a_bits_tag; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_11_bits_set = abc_mshr_11_io_tasks_source_a_bits_set; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_11_bits_off = abc_mshr_11_io_tasks_source_a_bits_off; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_11_bits_opcode = abc_mshr_11_io_tasks_source_a_bits_opcode; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_11_bits_param = abc_mshr_11_io_tasks_source_a_bits_param; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_11_bits_source = abc_mshr_11_io_tasks_source_a_bits_source; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_11_bits_bufIdx = abc_mshr_11_io_tasks_source_a_bits_bufIdx; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_11_bits_size = abc_mshr_11_io_tasks_source_a_bits_size; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_11_bits_putData = abc_mshr_11_io_tasks_source_a_bits_putData; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_12_valid = abc_mshr_12_io_tasks_source_a_valid; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_12_bits_tag = abc_mshr_12_io_tasks_source_a_bits_tag; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_12_bits_set = abc_mshr_12_io_tasks_source_a_bits_set; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_12_bits_off = abc_mshr_12_io_tasks_source_a_bits_off; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_12_bits_opcode = abc_mshr_12_io_tasks_source_a_bits_opcode; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_12_bits_param = abc_mshr_12_io_tasks_source_a_bits_param; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_12_bits_source = abc_mshr_12_io_tasks_source_a_bits_source; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_12_bits_bufIdx = abc_mshr_12_io_tasks_source_a_bits_bufIdx; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_12_bits_size = abc_mshr_12_io_tasks_source_a_bits_size; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_12_bits_putData = abc_mshr_12_io_tasks_source_a_bits_putData; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_13_valid = abc_mshr_13_io_tasks_source_a_valid; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_13_bits_tag = abc_mshr_13_io_tasks_source_a_bits_tag; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_13_bits_set = abc_mshr_13_io_tasks_source_a_bits_set; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_13_bits_off = abc_mshr_13_io_tasks_source_a_bits_off; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_13_bits_opcode = abc_mshr_13_io_tasks_source_a_bits_opcode; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_13_bits_param = abc_mshr_13_io_tasks_source_a_bits_param; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_13_bits_source = abc_mshr_13_io_tasks_source_a_bits_source; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_13_bits_bufIdx = abc_mshr_13_io_tasks_source_a_bits_bufIdx; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_13_bits_size = abc_mshr_13_io_tasks_source_a_bits_size; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_in_13_bits_putData = abc_mshr_13_io_tasks_source_a_bits_putData; // @[Slice.scala 472:13]
  assign sourceA_task_arb_io_out_ready = sourceA_io_task_ready & _ms_14_io_tasks_source_a_ready_T_1 & ~bc_real_valid; // @[Slice.scala 493:60]
  assign sourceB_task_arb_clock = clock;
  assign sourceB_task_arb_reset = reset;
  assign sourceB_task_arb_io_in_0_valid = abc_mshr_0_io_tasks_source_bvalid; // @[Slice.scala 472:13]
  assign sourceB_task_arb_io_in_0_bits_set = abc_mshr_0_io_tasks_source_bset; // @[Slice.scala 472:13]
  assign sourceB_task_arb_io_in_0_bits_tag = abc_mshr_0_io_tasks_source_btag; // @[Slice.scala 472:13]
  assign sourceB_task_arb_io_in_0_bits_param = abc_mshr_0_io_tasks_source_bparam; // @[Slice.scala 472:13]
  assign sourceB_task_arb_io_in_0_bits_clients = abc_mshr_0_io_tasks_source_bclients; // @[Slice.scala 472:13]
  assign sourceB_task_arb_io_in_0_bits_needData = abc_mshr_0_io_tasks_source_bneedData; // @[Slice.scala 472:13]
  assign sourceB_task_arb_io_in_1_valid = abc_mshr_1_io_tasks_source_bvalid; // @[Slice.scala 472:13]
  assign sourceB_task_arb_io_in_1_bits_set = abc_mshr_1_io_tasks_source_bset; // @[Slice.scala 472:13]
  assign sourceB_task_arb_io_in_1_bits_tag = abc_mshr_1_io_tasks_source_btag; // @[Slice.scala 472:13]
  assign sourceB_task_arb_io_in_1_bits_param = abc_mshr_1_io_tasks_source_bparam; // @[Slice.scala 472:13]
  assign sourceB_task_arb_io_in_1_bits_clients = abc_mshr_1_io_tasks_source_bclients; // @[Slice.scala 472:13]
  assign sourceB_task_arb_io_in_1_bits_needData = abc_mshr_1_io_tasks_source_bneedData; // @[Slice.scala 472:13]
  assign sourceB_task_arb_io_in_2_valid = abc_mshr_2_io_tasks_source_bvalid; // @[Slice.scala 472:13]
  assign sourceB_task_arb_io_in_2_bits_set = abc_mshr_2_io_tasks_source_bset; // @[Slice.scala 472:13]
  assign sourceB_task_arb_io_in_2_bits_tag = abc_mshr_2_io_tasks_source_btag; // @[Slice.scala 472:13]
  assign sourceB_task_arb_io_in_2_bits_param = abc_mshr_2_io_tasks_source_bparam; // @[Slice.scala 472:13]
  assign sourceB_task_arb_io_in_2_bits_clients = abc_mshr_2_io_tasks_source_bclients; // @[Slice.scala 472:13]
  assign sourceB_task_arb_io_in_2_bits_needData = abc_mshr_2_io_tasks_source_bneedData; // @[Slice.scala 472:13]
  assign sourceB_task_arb_io_in_3_valid = abc_mshr_3_io_tasks_source_bvalid; // @[Slice.scala 472:13]
  assign sourceB_task_arb_io_in_3_bits_set = abc_mshr_3_io_tasks_source_bset; // @[Slice.scala 472:13]
  assign sourceB_task_arb_io_in_3_bits_tag = abc_mshr_3_io_tasks_source_btag; // @[Slice.scala 472:13]
  assign sourceB_task_arb_io_in_3_bits_param = abc_mshr_3_io_tasks_source_bparam; // @[Slice.scala 472:13]
  assign sourceB_task_arb_io_in_3_bits_clients = abc_mshr_3_io_tasks_source_bclients; // @[Slice.scala 472:13]
  assign sourceB_task_arb_io_in_3_bits_needData = abc_mshr_3_io_tasks_source_bneedData; // @[Slice.scala 472:13]
  assign sourceB_task_arb_io_in_4_valid = abc_mshr_4_io_tasks_source_bvalid; // @[Slice.scala 472:13]
  assign sourceB_task_arb_io_in_4_bits_set = abc_mshr_4_io_tasks_source_bset; // @[Slice.scala 472:13]
  assign sourceB_task_arb_io_in_4_bits_tag = abc_mshr_4_io_tasks_source_btag; // @[Slice.scala 472:13]
  assign sourceB_task_arb_io_in_4_bits_param = abc_mshr_4_io_tasks_source_bparam; // @[Slice.scala 472:13]
  assign sourceB_task_arb_io_in_4_bits_clients = abc_mshr_4_io_tasks_source_bclients; // @[Slice.scala 472:13]
  assign sourceB_task_arb_io_in_4_bits_needData = abc_mshr_4_io_tasks_source_bneedData; // @[Slice.scala 472:13]
  assign sourceB_task_arb_io_in_5_valid = abc_mshr_5_io_tasks_source_bvalid; // @[Slice.scala 472:13]
  assign sourceB_task_arb_io_in_5_bits_set = abc_mshr_5_io_tasks_source_bset; // @[Slice.scala 472:13]
  assign sourceB_task_arb_io_in_5_bits_tag = abc_mshr_5_io_tasks_source_btag; // @[Slice.scala 472:13]
  assign sourceB_task_arb_io_in_5_bits_param = abc_mshr_5_io_tasks_source_bparam; // @[Slice.scala 472:13]
  assign sourceB_task_arb_io_in_5_bits_clients = abc_mshr_5_io_tasks_source_bclients; // @[Slice.scala 472:13]
  assign sourceB_task_arb_io_in_5_bits_needData = abc_mshr_5_io_tasks_source_bneedData; // @[Slice.scala 472:13]
  assign sourceB_task_arb_io_in_6_valid = abc_mshr_6_io_tasks_source_bvalid; // @[Slice.scala 472:13]
  assign sourceB_task_arb_io_in_6_bits_set = abc_mshr_6_io_tasks_source_bset; // @[Slice.scala 472:13]
  assign sourceB_task_arb_io_in_6_bits_tag = abc_mshr_6_io_tasks_source_btag; // @[Slice.scala 472:13]
  assign sourceB_task_arb_io_in_6_bits_param = abc_mshr_6_io_tasks_source_bparam; // @[Slice.scala 472:13]
  assign sourceB_task_arb_io_in_6_bits_clients = abc_mshr_6_io_tasks_source_bclients; // @[Slice.scala 472:13]
  assign sourceB_task_arb_io_in_6_bits_needData = abc_mshr_6_io_tasks_source_bneedData; // @[Slice.scala 472:13]
  assign sourceB_task_arb_io_in_7_valid = abc_mshr_7_io_tasks_source_bvalid; // @[Slice.scala 472:13]
  assign sourceB_task_arb_io_in_7_bits_set = abc_mshr_7_io_tasks_source_bset; // @[Slice.scala 472:13]
  assign sourceB_task_arb_io_in_7_bits_tag = abc_mshr_7_io_tasks_source_btag; // @[Slice.scala 472:13]
  assign sourceB_task_arb_io_in_7_bits_param = abc_mshr_7_io_tasks_source_bparam; // @[Slice.scala 472:13]
  assign sourceB_task_arb_io_in_7_bits_clients = abc_mshr_7_io_tasks_source_bclients; // @[Slice.scala 472:13]
  assign sourceB_task_arb_io_in_7_bits_needData = abc_mshr_7_io_tasks_source_bneedData; // @[Slice.scala 472:13]
  assign sourceB_task_arb_io_in_8_valid = abc_mshr_8_io_tasks_source_bvalid; // @[Slice.scala 472:13]
  assign sourceB_task_arb_io_in_8_bits_set = abc_mshr_8_io_tasks_source_bset; // @[Slice.scala 472:13]
  assign sourceB_task_arb_io_in_8_bits_tag = abc_mshr_8_io_tasks_source_btag; // @[Slice.scala 472:13]
  assign sourceB_task_arb_io_in_8_bits_param = abc_mshr_8_io_tasks_source_bparam; // @[Slice.scala 472:13]
  assign sourceB_task_arb_io_in_8_bits_clients = abc_mshr_8_io_tasks_source_bclients; // @[Slice.scala 472:13]
  assign sourceB_task_arb_io_in_8_bits_needData = abc_mshr_8_io_tasks_source_bneedData; // @[Slice.scala 472:13]
  assign sourceB_task_arb_io_in_9_valid = abc_mshr_9_io_tasks_source_bvalid; // @[Slice.scala 472:13]
  assign sourceB_task_arb_io_in_9_bits_set = abc_mshr_9_io_tasks_source_bset; // @[Slice.scala 472:13]
  assign sourceB_task_arb_io_in_9_bits_tag = abc_mshr_9_io_tasks_source_btag; // @[Slice.scala 472:13]
  assign sourceB_task_arb_io_in_9_bits_param = abc_mshr_9_io_tasks_source_bparam; // @[Slice.scala 472:13]
  assign sourceB_task_arb_io_in_9_bits_clients = abc_mshr_9_io_tasks_source_bclients; // @[Slice.scala 472:13]
  assign sourceB_task_arb_io_in_9_bits_needData = abc_mshr_9_io_tasks_source_bneedData; // @[Slice.scala 472:13]
  assign sourceB_task_arb_io_in_10_valid = abc_mshr_10_io_tasks_source_bvalid; // @[Slice.scala 472:13]
  assign sourceB_task_arb_io_in_10_bits_set = abc_mshr_10_io_tasks_source_bset; // @[Slice.scala 472:13]
  assign sourceB_task_arb_io_in_10_bits_tag = abc_mshr_10_io_tasks_source_btag; // @[Slice.scala 472:13]
  assign sourceB_task_arb_io_in_10_bits_param = abc_mshr_10_io_tasks_source_bparam; // @[Slice.scala 472:13]
  assign sourceB_task_arb_io_in_10_bits_clients = abc_mshr_10_io_tasks_source_bclients; // @[Slice.scala 472:13]
  assign sourceB_task_arb_io_in_10_bits_needData = abc_mshr_10_io_tasks_source_bneedData; // @[Slice.scala 472:13]
  assign sourceB_task_arb_io_in_11_valid = abc_mshr_11_io_tasks_source_bvalid; // @[Slice.scala 472:13]
  assign sourceB_task_arb_io_in_11_bits_set = abc_mshr_11_io_tasks_source_bset; // @[Slice.scala 472:13]
  assign sourceB_task_arb_io_in_11_bits_tag = abc_mshr_11_io_tasks_source_btag; // @[Slice.scala 472:13]
  assign sourceB_task_arb_io_in_11_bits_param = abc_mshr_11_io_tasks_source_bparam; // @[Slice.scala 472:13]
  assign sourceB_task_arb_io_in_11_bits_clients = abc_mshr_11_io_tasks_source_bclients; // @[Slice.scala 472:13]
  assign sourceB_task_arb_io_in_11_bits_needData = abc_mshr_11_io_tasks_source_bneedData; // @[Slice.scala 472:13]
  assign sourceB_task_arb_io_in_12_valid = abc_mshr_12_io_tasks_source_bvalid; // @[Slice.scala 472:13]
  assign sourceB_task_arb_io_in_12_bits_set = abc_mshr_12_io_tasks_source_bset; // @[Slice.scala 472:13]
  assign sourceB_task_arb_io_in_12_bits_tag = abc_mshr_12_io_tasks_source_btag; // @[Slice.scala 472:13]
  assign sourceB_task_arb_io_in_12_bits_param = abc_mshr_12_io_tasks_source_bparam; // @[Slice.scala 472:13]
  assign sourceB_task_arb_io_in_12_bits_clients = abc_mshr_12_io_tasks_source_bclients; // @[Slice.scala 472:13]
  assign sourceB_task_arb_io_in_12_bits_needData = abc_mshr_12_io_tasks_source_bneedData; // @[Slice.scala 472:13]
  assign sourceB_task_arb_io_in_13_valid = abc_mshr_13_io_tasks_source_bvalid; // @[Slice.scala 472:13]
  assign sourceB_task_arb_io_in_13_bits_set = abc_mshr_13_io_tasks_source_bset; // @[Slice.scala 472:13]
  assign sourceB_task_arb_io_in_13_bits_tag = abc_mshr_13_io_tasks_source_btag; // @[Slice.scala 472:13]
  assign sourceB_task_arb_io_in_13_bits_param = abc_mshr_13_io_tasks_source_bparam; // @[Slice.scala 472:13]
  assign sourceB_task_arb_io_in_13_bits_clients = abc_mshr_13_io_tasks_source_bclients; // @[Slice.scala 472:13]
  assign sourceB_task_arb_io_in_13_bits_needData = abc_mshr_13_io_tasks_source_bneedData; // @[Slice.scala 472:13]
  assign sourceB_task_arb_io_out_ready = sourceB_io_task_ready & _ms_14_io_tasks_source_bready_T_1 & ~bc_real_valid_1; // @[Slice.scala 493:60]
  assign sourceC_task_arb_clock = clock;
  assign sourceC_task_arb_reset = reset;
  assign sourceC_task_arb_io_in_0_valid = abc_mshr_0_io_tasks_source_c_valid; // @[Slice.scala 472:13]
  assign sourceC_task_arb_io_in_0_bits_opcode = abc_mshr_0_io_tasks_source_c_bits_opcode; // @[Slice.scala 472:13]
  assign sourceC_task_arb_io_in_0_bits_tag = abc_mshr_0_io_tasks_source_c_bits_tag; // @[Slice.scala 472:13]
  assign sourceC_task_arb_io_in_0_bits_set = abc_mshr_0_io_tasks_source_c_bits_set; // @[Slice.scala 472:13]
  assign sourceC_task_arb_io_in_0_bits_source = abc_mshr_0_io_tasks_source_c_bits_source; // @[Slice.scala 472:13]
  assign sourceC_task_arb_io_in_0_bits_way = abc_mshr_0_io_tasks_source_c_bits_way; // @[Slice.scala 472:13]
  assign sourceC_task_arb_io_in_1_valid = abc_mshr_1_io_tasks_source_c_valid; // @[Slice.scala 472:13]
  assign sourceC_task_arb_io_in_1_bits_opcode = abc_mshr_1_io_tasks_source_c_bits_opcode; // @[Slice.scala 472:13]
  assign sourceC_task_arb_io_in_1_bits_tag = abc_mshr_1_io_tasks_source_c_bits_tag; // @[Slice.scala 472:13]
  assign sourceC_task_arb_io_in_1_bits_set = abc_mshr_1_io_tasks_source_c_bits_set; // @[Slice.scala 472:13]
  assign sourceC_task_arb_io_in_1_bits_source = abc_mshr_1_io_tasks_source_c_bits_source; // @[Slice.scala 472:13]
  assign sourceC_task_arb_io_in_1_bits_way = abc_mshr_1_io_tasks_source_c_bits_way; // @[Slice.scala 472:13]
  assign sourceC_task_arb_io_in_2_valid = abc_mshr_2_io_tasks_source_c_valid; // @[Slice.scala 472:13]
  assign sourceC_task_arb_io_in_2_bits_opcode = abc_mshr_2_io_tasks_source_c_bits_opcode; // @[Slice.scala 472:13]
  assign sourceC_task_arb_io_in_2_bits_tag = abc_mshr_2_io_tasks_source_c_bits_tag; // @[Slice.scala 472:13]
  assign sourceC_task_arb_io_in_2_bits_set = abc_mshr_2_io_tasks_source_c_bits_set; // @[Slice.scala 472:13]
  assign sourceC_task_arb_io_in_2_bits_source = abc_mshr_2_io_tasks_source_c_bits_source; // @[Slice.scala 472:13]
  assign sourceC_task_arb_io_in_2_bits_way = abc_mshr_2_io_tasks_source_c_bits_way; // @[Slice.scala 472:13]
  assign sourceC_task_arb_io_in_3_valid = abc_mshr_3_io_tasks_source_c_valid; // @[Slice.scala 472:13]
  assign sourceC_task_arb_io_in_3_bits_opcode = abc_mshr_3_io_tasks_source_c_bits_opcode; // @[Slice.scala 472:13]
  assign sourceC_task_arb_io_in_3_bits_tag = abc_mshr_3_io_tasks_source_c_bits_tag; // @[Slice.scala 472:13]
  assign sourceC_task_arb_io_in_3_bits_set = abc_mshr_3_io_tasks_source_c_bits_set; // @[Slice.scala 472:13]
  assign sourceC_task_arb_io_in_3_bits_source = abc_mshr_3_io_tasks_source_c_bits_source; // @[Slice.scala 472:13]
  assign sourceC_task_arb_io_in_3_bits_way = abc_mshr_3_io_tasks_source_c_bits_way; // @[Slice.scala 472:13]
  assign sourceC_task_arb_io_in_4_valid = abc_mshr_4_io_tasks_source_c_valid; // @[Slice.scala 472:13]
  assign sourceC_task_arb_io_in_4_bits_opcode = abc_mshr_4_io_tasks_source_c_bits_opcode; // @[Slice.scala 472:13]
  assign sourceC_task_arb_io_in_4_bits_tag = abc_mshr_4_io_tasks_source_c_bits_tag; // @[Slice.scala 472:13]
  assign sourceC_task_arb_io_in_4_bits_set = abc_mshr_4_io_tasks_source_c_bits_set; // @[Slice.scala 472:13]
  assign sourceC_task_arb_io_in_4_bits_source = abc_mshr_4_io_tasks_source_c_bits_source; // @[Slice.scala 472:13]
  assign sourceC_task_arb_io_in_4_bits_way = abc_mshr_4_io_tasks_source_c_bits_way; // @[Slice.scala 472:13]
  assign sourceC_task_arb_io_in_5_valid = abc_mshr_5_io_tasks_source_c_valid; // @[Slice.scala 472:13]
  assign sourceC_task_arb_io_in_5_bits_opcode = abc_mshr_5_io_tasks_source_c_bits_opcode; // @[Slice.scala 472:13]
  assign sourceC_task_arb_io_in_5_bits_tag = abc_mshr_5_io_tasks_source_c_bits_tag; // @[Slice.scala 472:13]
  assign sourceC_task_arb_io_in_5_bits_set = abc_mshr_5_io_tasks_source_c_bits_set; // @[Slice.scala 472:13]
  assign sourceC_task_arb_io_in_5_bits_source = abc_mshr_5_io_tasks_source_c_bits_source; // @[Slice.scala 472:13]
  assign sourceC_task_arb_io_in_5_bits_way = abc_mshr_5_io_tasks_source_c_bits_way; // @[Slice.scala 472:13]
  assign sourceC_task_arb_io_in_6_valid = abc_mshr_6_io_tasks_source_c_valid; // @[Slice.scala 472:13]
  assign sourceC_task_arb_io_in_6_bits_opcode = abc_mshr_6_io_tasks_source_c_bits_opcode; // @[Slice.scala 472:13]
  assign sourceC_task_arb_io_in_6_bits_tag = abc_mshr_6_io_tasks_source_c_bits_tag; // @[Slice.scala 472:13]
  assign sourceC_task_arb_io_in_6_bits_set = abc_mshr_6_io_tasks_source_c_bits_set; // @[Slice.scala 472:13]
  assign sourceC_task_arb_io_in_6_bits_source = abc_mshr_6_io_tasks_source_c_bits_source; // @[Slice.scala 472:13]
  assign sourceC_task_arb_io_in_6_bits_way = abc_mshr_6_io_tasks_source_c_bits_way; // @[Slice.scala 472:13]
  assign sourceC_task_arb_io_in_7_valid = abc_mshr_7_io_tasks_source_c_valid; // @[Slice.scala 472:13]
  assign sourceC_task_arb_io_in_7_bits_opcode = abc_mshr_7_io_tasks_source_c_bits_opcode; // @[Slice.scala 472:13]
  assign sourceC_task_arb_io_in_7_bits_tag = abc_mshr_7_io_tasks_source_c_bits_tag; // @[Slice.scala 472:13]
  assign sourceC_task_arb_io_in_7_bits_set = abc_mshr_7_io_tasks_source_c_bits_set; // @[Slice.scala 472:13]
  assign sourceC_task_arb_io_in_7_bits_source = abc_mshr_7_io_tasks_source_c_bits_source; // @[Slice.scala 472:13]
  assign sourceC_task_arb_io_in_7_bits_way = abc_mshr_7_io_tasks_source_c_bits_way; // @[Slice.scala 472:13]
  assign sourceC_task_arb_io_in_8_valid = abc_mshr_8_io_tasks_source_c_valid; // @[Slice.scala 472:13]
  assign sourceC_task_arb_io_in_8_bits_opcode = abc_mshr_8_io_tasks_source_c_bits_opcode; // @[Slice.scala 472:13]
  assign sourceC_task_arb_io_in_8_bits_tag = abc_mshr_8_io_tasks_source_c_bits_tag; // @[Slice.scala 472:13]
  assign sourceC_task_arb_io_in_8_bits_set = abc_mshr_8_io_tasks_source_c_bits_set; // @[Slice.scala 472:13]
  assign sourceC_task_arb_io_in_8_bits_source = abc_mshr_8_io_tasks_source_c_bits_source; // @[Slice.scala 472:13]
  assign sourceC_task_arb_io_in_8_bits_way = abc_mshr_8_io_tasks_source_c_bits_way; // @[Slice.scala 472:13]
  assign sourceC_task_arb_io_in_9_valid = abc_mshr_9_io_tasks_source_c_valid; // @[Slice.scala 472:13]
  assign sourceC_task_arb_io_in_9_bits_opcode = abc_mshr_9_io_tasks_source_c_bits_opcode; // @[Slice.scala 472:13]
  assign sourceC_task_arb_io_in_9_bits_tag = abc_mshr_9_io_tasks_source_c_bits_tag; // @[Slice.scala 472:13]
  assign sourceC_task_arb_io_in_9_bits_set = abc_mshr_9_io_tasks_source_c_bits_set; // @[Slice.scala 472:13]
  assign sourceC_task_arb_io_in_9_bits_source = abc_mshr_9_io_tasks_source_c_bits_source; // @[Slice.scala 472:13]
  assign sourceC_task_arb_io_in_9_bits_way = abc_mshr_9_io_tasks_source_c_bits_way; // @[Slice.scala 472:13]
  assign sourceC_task_arb_io_in_10_valid = abc_mshr_10_io_tasks_source_c_valid; // @[Slice.scala 472:13]
  assign sourceC_task_arb_io_in_10_bits_opcode = abc_mshr_10_io_tasks_source_c_bits_opcode; // @[Slice.scala 472:13]
  assign sourceC_task_arb_io_in_10_bits_tag = abc_mshr_10_io_tasks_source_c_bits_tag; // @[Slice.scala 472:13]
  assign sourceC_task_arb_io_in_10_bits_set = abc_mshr_10_io_tasks_source_c_bits_set; // @[Slice.scala 472:13]
  assign sourceC_task_arb_io_in_10_bits_source = abc_mshr_10_io_tasks_source_c_bits_source; // @[Slice.scala 472:13]
  assign sourceC_task_arb_io_in_10_bits_way = abc_mshr_10_io_tasks_source_c_bits_way; // @[Slice.scala 472:13]
  assign sourceC_task_arb_io_in_11_valid = abc_mshr_11_io_tasks_source_c_valid; // @[Slice.scala 472:13]
  assign sourceC_task_arb_io_in_11_bits_opcode = abc_mshr_11_io_tasks_source_c_bits_opcode; // @[Slice.scala 472:13]
  assign sourceC_task_arb_io_in_11_bits_tag = abc_mshr_11_io_tasks_source_c_bits_tag; // @[Slice.scala 472:13]
  assign sourceC_task_arb_io_in_11_bits_set = abc_mshr_11_io_tasks_source_c_bits_set; // @[Slice.scala 472:13]
  assign sourceC_task_arb_io_in_11_bits_source = abc_mshr_11_io_tasks_source_c_bits_source; // @[Slice.scala 472:13]
  assign sourceC_task_arb_io_in_11_bits_way = abc_mshr_11_io_tasks_source_c_bits_way; // @[Slice.scala 472:13]
  assign sourceC_task_arb_io_in_12_valid = abc_mshr_12_io_tasks_source_c_valid; // @[Slice.scala 472:13]
  assign sourceC_task_arb_io_in_12_bits_opcode = abc_mshr_12_io_tasks_source_c_bits_opcode; // @[Slice.scala 472:13]
  assign sourceC_task_arb_io_in_12_bits_tag = abc_mshr_12_io_tasks_source_c_bits_tag; // @[Slice.scala 472:13]
  assign sourceC_task_arb_io_in_12_bits_set = abc_mshr_12_io_tasks_source_c_bits_set; // @[Slice.scala 472:13]
  assign sourceC_task_arb_io_in_12_bits_source = abc_mshr_12_io_tasks_source_c_bits_source; // @[Slice.scala 472:13]
  assign sourceC_task_arb_io_in_12_bits_way = abc_mshr_12_io_tasks_source_c_bits_way; // @[Slice.scala 472:13]
  assign sourceC_task_arb_io_in_13_valid = abc_mshr_13_io_tasks_source_c_valid; // @[Slice.scala 472:13]
  assign sourceC_task_arb_io_in_13_bits_opcode = abc_mshr_13_io_tasks_source_c_bits_opcode; // @[Slice.scala 472:13]
  assign sourceC_task_arb_io_in_13_bits_tag = abc_mshr_13_io_tasks_source_c_bits_tag; // @[Slice.scala 472:13]
  assign sourceC_task_arb_io_in_13_bits_set = abc_mshr_13_io_tasks_source_c_bits_set; // @[Slice.scala 472:13]
  assign sourceC_task_arb_io_in_13_bits_source = abc_mshr_13_io_tasks_source_c_bits_source; // @[Slice.scala 472:13]
  assign sourceC_task_arb_io_in_13_bits_way = abc_mshr_13_io_tasks_source_c_bits_way; // @[Slice.scala 472:13]
  assign sourceC_task_arb_io_out_ready = sourceC_io_task_ready & _ms_14_io_tasks_source_c_ready_T_1 & ~bc_real_valid_2; // @[Slice.scala 493:60]
  assign sourceD_task_arb_clock = clock;
  assign sourceD_task_arb_reset = reset;
  assign sourceD_task_arb_io_in_0_valid = abc_mshr_0_io_tasks_source_d_valid; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_0_bits_sourceId = abc_mshr_0_io_tasks_source_d_bits_sourceId; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_0_bits_set = abc_mshr_0_io_tasks_source_d_bits_set; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_0_bits_channel = abc_mshr_0_io_tasks_source_d_bits_channel; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_0_bits_opcode = abc_mshr_0_io_tasks_source_d_bits_opcode; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_0_bits_param = abc_mshr_0_io_tasks_source_d_bits_param; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_0_bits_size = abc_mshr_0_io_tasks_source_d_bits_size; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_0_bits_way = abc_mshr_0_io_tasks_source_d_bits_way; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_0_bits_off = abc_mshr_0_io_tasks_source_d_bits_off; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_0_bits_useBypass = abc_mshr_0_io_tasks_source_d_bits_useBypass; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_0_bits_bufIdx = abc_mshr_0_io_tasks_source_d_bits_bufIdx; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_0_bits_denied = abc_mshr_0_io_tasks_source_d_bits_denied; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_0_bits_sinkId = abc_mshr_0_io_tasks_source_d_bits_sinkId; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_0_bits_bypassPut = abc_mshr_0_io_tasks_source_d_bits_bypassPut; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_0_bits_dirty = abc_mshr_0_io_tasks_source_d_bits_dirty; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_1_valid = abc_mshr_1_io_tasks_source_d_valid; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_1_bits_sourceId = abc_mshr_1_io_tasks_source_d_bits_sourceId; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_1_bits_set = abc_mshr_1_io_tasks_source_d_bits_set; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_1_bits_channel = abc_mshr_1_io_tasks_source_d_bits_channel; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_1_bits_opcode = abc_mshr_1_io_tasks_source_d_bits_opcode; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_1_bits_param = abc_mshr_1_io_tasks_source_d_bits_param; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_1_bits_size = abc_mshr_1_io_tasks_source_d_bits_size; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_1_bits_way = abc_mshr_1_io_tasks_source_d_bits_way; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_1_bits_off = abc_mshr_1_io_tasks_source_d_bits_off; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_1_bits_useBypass = abc_mshr_1_io_tasks_source_d_bits_useBypass; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_1_bits_bufIdx = abc_mshr_1_io_tasks_source_d_bits_bufIdx; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_1_bits_denied = abc_mshr_1_io_tasks_source_d_bits_denied; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_1_bits_sinkId = abc_mshr_1_io_tasks_source_d_bits_sinkId; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_1_bits_bypassPut = abc_mshr_1_io_tasks_source_d_bits_bypassPut; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_1_bits_dirty = abc_mshr_1_io_tasks_source_d_bits_dirty; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_2_valid = abc_mshr_2_io_tasks_source_d_valid; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_2_bits_sourceId = abc_mshr_2_io_tasks_source_d_bits_sourceId; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_2_bits_set = abc_mshr_2_io_tasks_source_d_bits_set; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_2_bits_channel = abc_mshr_2_io_tasks_source_d_bits_channel; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_2_bits_opcode = abc_mshr_2_io_tasks_source_d_bits_opcode; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_2_bits_param = abc_mshr_2_io_tasks_source_d_bits_param; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_2_bits_size = abc_mshr_2_io_tasks_source_d_bits_size; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_2_bits_way = abc_mshr_2_io_tasks_source_d_bits_way; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_2_bits_off = abc_mshr_2_io_tasks_source_d_bits_off; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_2_bits_useBypass = abc_mshr_2_io_tasks_source_d_bits_useBypass; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_2_bits_bufIdx = abc_mshr_2_io_tasks_source_d_bits_bufIdx; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_2_bits_denied = abc_mshr_2_io_tasks_source_d_bits_denied; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_2_bits_sinkId = abc_mshr_2_io_tasks_source_d_bits_sinkId; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_2_bits_bypassPut = abc_mshr_2_io_tasks_source_d_bits_bypassPut; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_2_bits_dirty = abc_mshr_2_io_tasks_source_d_bits_dirty; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_3_valid = abc_mshr_3_io_tasks_source_d_valid; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_3_bits_sourceId = abc_mshr_3_io_tasks_source_d_bits_sourceId; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_3_bits_set = abc_mshr_3_io_tasks_source_d_bits_set; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_3_bits_channel = abc_mshr_3_io_tasks_source_d_bits_channel; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_3_bits_opcode = abc_mshr_3_io_tasks_source_d_bits_opcode; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_3_bits_param = abc_mshr_3_io_tasks_source_d_bits_param; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_3_bits_size = abc_mshr_3_io_tasks_source_d_bits_size; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_3_bits_way = abc_mshr_3_io_tasks_source_d_bits_way; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_3_bits_off = abc_mshr_3_io_tasks_source_d_bits_off; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_3_bits_useBypass = abc_mshr_3_io_tasks_source_d_bits_useBypass; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_3_bits_bufIdx = abc_mshr_3_io_tasks_source_d_bits_bufIdx; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_3_bits_denied = abc_mshr_3_io_tasks_source_d_bits_denied; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_3_bits_sinkId = abc_mshr_3_io_tasks_source_d_bits_sinkId; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_3_bits_bypassPut = abc_mshr_3_io_tasks_source_d_bits_bypassPut; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_3_bits_dirty = abc_mshr_3_io_tasks_source_d_bits_dirty; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_4_valid = abc_mshr_4_io_tasks_source_d_valid; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_4_bits_sourceId = abc_mshr_4_io_tasks_source_d_bits_sourceId; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_4_bits_set = abc_mshr_4_io_tasks_source_d_bits_set; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_4_bits_channel = abc_mshr_4_io_tasks_source_d_bits_channel; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_4_bits_opcode = abc_mshr_4_io_tasks_source_d_bits_opcode; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_4_bits_param = abc_mshr_4_io_tasks_source_d_bits_param; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_4_bits_size = abc_mshr_4_io_tasks_source_d_bits_size; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_4_bits_way = abc_mshr_4_io_tasks_source_d_bits_way; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_4_bits_off = abc_mshr_4_io_tasks_source_d_bits_off; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_4_bits_useBypass = abc_mshr_4_io_tasks_source_d_bits_useBypass; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_4_bits_bufIdx = abc_mshr_4_io_tasks_source_d_bits_bufIdx; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_4_bits_denied = abc_mshr_4_io_tasks_source_d_bits_denied; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_4_bits_sinkId = abc_mshr_4_io_tasks_source_d_bits_sinkId; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_4_bits_bypassPut = abc_mshr_4_io_tasks_source_d_bits_bypassPut; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_4_bits_dirty = abc_mshr_4_io_tasks_source_d_bits_dirty; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_5_valid = abc_mshr_5_io_tasks_source_d_valid; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_5_bits_sourceId = abc_mshr_5_io_tasks_source_d_bits_sourceId; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_5_bits_set = abc_mshr_5_io_tasks_source_d_bits_set; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_5_bits_channel = abc_mshr_5_io_tasks_source_d_bits_channel; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_5_bits_opcode = abc_mshr_5_io_tasks_source_d_bits_opcode; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_5_bits_param = abc_mshr_5_io_tasks_source_d_bits_param; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_5_bits_size = abc_mshr_5_io_tasks_source_d_bits_size; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_5_bits_way = abc_mshr_5_io_tasks_source_d_bits_way; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_5_bits_off = abc_mshr_5_io_tasks_source_d_bits_off; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_5_bits_useBypass = abc_mshr_5_io_tasks_source_d_bits_useBypass; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_5_bits_bufIdx = abc_mshr_5_io_tasks_source_d_bits_bufIdx; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_5_bits_denied = abc_mshr_5_io_tasks_source_d_bits_denied; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_5_bits_sinkId = abc_mshr_5_io_tasks_source_d_bits_sinkId; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_5_bits_bypassPut = abc_mshr_5_io_tasks_source_d_bits_bypassPut; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_5_bits_dirty = abc_mshr_5_io_tasks_source_d_bits_dirty; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_6_valid = abc_mshr_6_io_tasks_source_d_valid; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_6_bits_sourceId = abc_mshr_6_io_tasks_source_d_bits_sourceId; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_6_bits_set = abc_mshr_6_io_tasks_source_d_bits_set; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_6_bits_channel = abc_mshr_6_io_tasks_source_d_bits_channel; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_6_bits_opcode = abc_mshr_6_io_tasks_source_d_bits_opcode; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_6_bits_param = abc_mshr_6_io_tasks_source_d_bits_param; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_6_bits_size = abc_mshr_6_io_tasks_source_d_bits_size; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_6_bits_way = abc_mshr_6_io_tasks_source_d_bits_way; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_6_bits_off = abc_mshr_6_io_tasks_source_d_bits_off; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_6_bits_useBypass = abc_mshr_6_io_tasks_source_d_bits_useBypass; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_6_bits_bufIdx = abc_mshr_6_io_tasks_source_d_bits_bufIdx; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_6_bits_denied = abc_mshr_6_io_tasks_source_d_bits_denied; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_6_bits_sinkId = abc_mshr_6_io_tasks_source_d_bits_sinkId; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_6_bits_bypassPut = abc_mshr_6_io_tasks_source_d_bits_bypassPut; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_6_bits_dirty = abc_mshr_6_io_tasks_source_d_bits_dirty; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_7_valid = abc_mshr_7_io_tasks_source_d_valid; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_7_bits_sourceId = abc_mshr_7_io_tasks_source_d_bits_sourceId; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_7_bits_set = abc_mshr_7_io_tasks_source_d_bits_set; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_7_bits_channel = abc_mshr_7_io_tasks_source_d_bits_channel; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_7_bits_opcode = abc_mshr_7_io_tasks_source_d_bits_opcode; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_7_bits_param = abc_mshr_7_io_tasks_source_d_bits_param; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_7_bits_size = abc_mshr_7_io_tasks_source_d_bits_size; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_7_bits_way = abc_mshr_7_io_tasks_source_d_bits_way; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_7_bits_off = abc_mshr_7_io_tasks_source_d_bits_off; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_7_bits_useBypass = abc_mshr_7_io_tasks_source_d_bits_useBypass; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_7_bits_bufIdx = abc_mshr_7_io_tasks_source_d_bits_bufIdx; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_7_bits_denied = abc_mshr_7_io_tasks_source_d_bits_denied; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_7_bits_sinkId = abc_mshr_7_io_tasks_source_d_bits_sinkId; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_7_bits_bypassPut = abc_mshr_7_io_tasks_source_d_bits_bypassPut; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_7_bits_dirty = abc_mshr_7_io_tasks_source_d_bits_dirty; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_8_valid = abc_mshr_8_io_tasks_source_d_valid; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_8_bits_sourceId = abc_mshr_8_io_tasks_source_d_bits_sourceId; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_8_bits_set = abc_mshr_8_io_tasks_source_d_bits_set; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_8_bits_channel = abc_mshr_8_io_tasks_source_d_bits_channel; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_8_bits_opcode = abc_mshr_8_io_tasks_source_d_bits_opcode; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_8_bits_param = abc_mshr_8_io_tasks_source_d_bits_param; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_8_bits_size = abc_mshr_8_io_tasks_source_d_bits_size; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_8_bits_way = abc_mshr_8_io_tasks_source_d_bits_way; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_8_bits_off = abc_mshr_8_io_tasks_source_d_bits_off; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_8_bits_useBypass = abc_mshr_8_io_tasks_source_d_bits_useBypass; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_8_bits_bufIdx = abc_mshr_8_io_tasks_source_d_bits_bufIdx; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_8_bits_denied = abc_mshr_8_io_tasks_source_d_bits_denied; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_8_bits_sinkId = abc_mshr_8_io_tasks_source_d_bits_sinkId; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_8_bits_bypassPut = abc_mshr_8_io_tasks_source_d_bits_bypassPut; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_8_bits_dirty = abc_mshr_8_io_tasks_source_d_bits_dirty; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_9_valid = abc_mshr_9_io_tasks_source_d_valid; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_9_bits_sourceId = abc_mshr_9_io_tasks_source_d_bits_sourceId; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_9_bits_set = abc_mshr_9_io_tasks_source_d_bits_set; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_9_bits_channel = abc_mshr_9_io_tasks_source_d_bits_channel; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_9_bits_opcode = abc_mshr_9_io_tasks_source_d_bits_opcode; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_9_bits_param = abc_mshr_9_io_tasks_source_d_bits_param; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_9_bits_size = abc_mshr_9_io_tasks_source_d_bits_size; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_9_bits_way = abc_mshr_9_io_tasks_source_d_bits_way; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_9_bits_off = abc_mshr_9_io_tasks_source_d_bits_off; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_9_bits_useBypass = abc_mshr_9_io_tasks_source_d_bits_useBypass; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_9_bits_bufIdx = abc_mshr_9_io_tasks_source_d_bits_bufIdx; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_9_bits_denied = abc_mshr_9_io_tasks_source_d_bits_denied; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_9_bits_sinkId = abc_mshr_9_io_tasks_source_d_bits_sinkId; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_9_bits_bypassPut = abc_mshr_9_io_tasks_source_d_bits_bypassPut; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_9_bits_dirty = abc_mshr_9_io_tasks_source_d_bits_dirty; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_10_valid = abc_mshr_10_io_tasks_source_d_valid; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_10_bits_sourceId = abc_mshr_10_io_tasks_source_d_bits_sourceId; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_10_bits_set = abc_mshr_10_io_tasks_source_d_bits_set; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_10_bits_channel = abc_mshr_10_io_tasks_source_d_bits_channel; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_10_bits_opcode = abc_mshr_10_io_tasks_source_d_bits_opcode; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_10_bits_param = abc_mshr_10_io_tasks_source_d_bits_param; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_10_bits_size = abc_mshr_10_io_tasks_source_d_bits_size; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_10_bits_way = abc_mshr_10_io_tasks_source_d_bits_way; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_10_bits_off = abc_mshr_10_io_tasks_source_d_bits_off; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_10_bits_useBypass = abc_mshr_10_io_tasks_source_d_bits_useBypass; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_10_bits_bufIdx = abc_mshr_10_io_tasks_source_d_bits_bufIdx; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_10_bits_denied = abc_mshr_10_io_tasks_source_d_bits_denied; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_10_bits_sinkId = abc_mshr_10_io_tasks_source_d_bits_sinkId; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_10_bits_bypassPut = abc_mshr_10_io_tasks_source_d_bits_bypassPut; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_10_bits_dirty = abc_mshr_10_io_tasks_source_d_bits_dirty; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_11_valid = abc_mshr_11_io_tasks_source_d_valid; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_11_bits_sourceId = abc_mshr_11_io_tasks_source_d_bits_sourceId; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_11_bits_set = abc_mshr_11_io_tasks_source_d_bits_set; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_11_bits_channel = abc_mshr_11_io_tasks_source_d_bits_channel; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_11_bits_opcode = abc_mshr_11_io_tasks_source_d_bits_opcode; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_11_bits_param = abc_mshr_11_io_tasks_source_d_bits_param; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_11_bits_size = abc_mshr_11_io_tasks_source_d_bits_size; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_11_bits_way = abc_mshr_11_io_tasks_source_d_bits_way; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_11_bits_off = abc_mshr_11_io_tasks_source_d_bits_off; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_11_bits_useBypass = abc_mshr_11_io_tasks_source_d_bits_useBypass; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_11_bits_bufIdx = abc_mshr_11_io_tasks_source_d_bits_bufIdx; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_11_bits_denied = abc_mshr_11_io_tasks_source_d_bits_denied; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_11_bits_sinkId = abc_mshr_11_io_tasks_source_d_bits_sinkId; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_11_bits_bypassPut = abc_mshr_11_io_tasks_source_d_bits_bypassPut; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_11_bits_dirty = abc_mshr_11_io_tasks_source_d_bits_dirty; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_12_valid = abc_mshr_12_io_tasks_source_d_valid; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_12_bits_sourceId = abc_mshr_12_io_tasks_source_d_bits_sourceId; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_12_bits_set = abc_mshr_12_io_tasks_source_d_bits_set; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_12_bits_channel = abc_mshr_12_io_tasks_source_d_bits_channel; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_12_bits_opcode = abc_mshr_12_io_tasks_source_d_bits_opcode; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_12_bits_param = abc_mshr_12_io_tasks_source_d_bits_param; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_12_bits_size = abc_mshr_12_io_tasks_source_d_bits_size; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_12_bits_way = abc_mshr_12_io_tasks_source_d_bits_way; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_12_bits_off = abc_mshr_12_io_tasks_source_d_bits_off; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_12_bits_useBypass = abc_mshr_12_io_tasks_source_d_bits_useBypass; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_12_bits_bufIdx = abc_mshr_12_io_tasks_source_d_bits_bufIdx; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_12_bits_denied = abc_mshr_12_io_tasks_source_d_bits_denied; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_12_bits_sinkId = abc_mshr_12_io_tasks_source_d_bits_sinkId; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_12_bits_bypassPut = abc_mshr_12_io_tasks_source_d_bits_bypassPut; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_12_bits_dirty = abc_mshr_12_io_tasks_source_d_bits_dirty; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_13_valid = abc_mshr_13_io_tasks_source_d_valid; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_13_bits_sourceId = abc_mshr_13_io_tasks_source_d_bits_sourceId; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_13_bits_set = abc_mshr_13_io_tasks_source_d_bits_set; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_13_bits_channel = abc_mshr_13_io_tasks_source_d_bits_channel; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_13_bits_opcode = abc_mshr_13_io_tasks_source_d_bits_opcode; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_13_bits_param = abc_mshr_13_io_tasks_source_d_bits_param; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_13_bits_size = abc_mshr_13_io_tasks_source_d_bits_size; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_13_bits_way = abc_mshr_13_io_tasks_source_d_bits_way; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_13_bits_off = abc_mshr_13_io_tasks_source_d_bits_off; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_13_bits_useBypass = abc_mshr_13_io_tasks_source_d_bits_useBypass; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_13_bits_bufIdx = abc_mshr_13_io_tasks_source_d_bits_bufIdx; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_13_bits_denied = abc_mshr_13_io_tasks_source_d_bits_denied; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_13_bits_sinkId = abc_mshr_13_io_tasks_source_d_bits_sinkId; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_13_bits_bypassPut = abc_mshr_13_io_tasks_source_d_bits_bypassPut; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_in_13_bits_dirty = abc_mshr_13_io_tasks_source_d_bits_dirty; // @[Slice.scala 472:13]
  assign sourceD_task_arb_io_out_ready = sourceD_io_task_ready & _ms_14_io_tasks_source_d_ready_T_1 & ~bc_real_valid_3; // @[Slice.scala 493:60]
  assign sourceE_task_arb_clock = clock;
  assign sourceE_task_arb_reset = reset;
  assign sourceE_task_arb_io_in_0_valid = abc_mshr_0_io_tasks_source_e_valid; // @[Slice.scala 472:13]
  assign sourceE_task_arb_io_in_0_bits_sink = abc_mshr_0_io_tasks_source_e_bits_sink; // @[Slice.scala 472:13]
  assign sourceE_task_arb_io_in_1_valid = abc_mshr_1_io_tasks_source_e_valid; // @[Slice.scala 472:13]
  assign sourceE_task_arb_io_in_1_bits_sink = abc_mshr_1_io_tasks_source_e_bits_sink; // @[Slice.scala 472:13]
  assign sourceE_task_arb_io_in_2_valid = abc_mshr_2_io_tasks_source_e_valid; // @[Slice.scala 472:13]
  assign sourceE_task_arb_io_in_2_bits_sink = abc_mshr_2_io_tasks_source_e_bits_sink; // @[Slice.scala 472:13]
  assign sourceE_task_arb_io_in_3_valid = abc_mshr_3_io_tasks_source_e_valid; // @[Slice.scala 472:13]
  assign sourceE_task_arb_io_in_3_bits_sink = abc_mshr_3_io_tasks_source_e_bits_sink; // @[Slice.scala 472:13]
  assign sourceE_task_arb_io_in_4_valid = abc_mshr_4_io_tasks_source_e_valid; // @[Slice.scala 472:13]
  assign sourceE_task_arb_io_in_4_bits_sink = abc_mshr_4_io_tasks_source_e_bits_sink; // @[Slice.scala 472:13]
  assign sourceE_task_arb_io_in_5_valid = abc_mshr_5_io_tasks_source_e_valid; // @[Slice.scala 472:13]
  assign sourceE_task_arb_io_in_5_bits_sink = abc_mshr_5_io_tasks_source_e_bits_sink; // @[Slice.scala 472:13]
  assign sourceE_task_arb_io_in_6_valid = abc_mshr_6_io_tasks_source_e_valid; // @[Slice.scala 472:13]
  assign sourceE_task_arb_io_in_6_bits_sink = abc_mshr_6_io_tasks_source_e_bits_sink; // @[Slice.scala 472:13]
  assign sourceE_task_arb_io_in_7_valid = abc_mshr_7_io_tasks_source_e_valid; // @[Slice.scala 472:13]
  assign sourceE_task_arb_io_in_7_bits_sink = abc_mshr_7_io_tasks_source_e_bits_sink; // @[Slice.scala 472:13]
  assign sourceE_task_arb_io_in_8_valid = abc_mshr_8_io_tasks_source_e_valid; // @[Slice.scala 472:13]
  assign sourceE_task_arb_io_in_8_bits_sink = abc_mshr_8_io_tasks_source_e_bits_sink; // @[Slice.scala 472:13]
  assign sourceE_task_arb_io_in_9_valid = abc_mshr_9_io_tasks_source_e_valid; // @[Slice.scala 472:13]
  assign sourceE_task_arb_io_in_9_bits_sink = abc_mshr_9_io_tasks_source_e_bits_sink; // @[Slice.scala 472:13]
  assign sourceE_task_arb_io_in_10_valid = abc_mshr_10_io_tasks_source_e_valid; // @[Slice.scala 472:13]
  assign sourceE_task_arb_io_in_10_bits_sink = abc_mshr_10_io_tasks_source_e_bits_sink; // @[Slice.scala 472:13]
  assign sourceE_task_arb_io_in_11_valid = abc_mshr_11_io_tasks_source_e_valid; // @[Slice.scala 472:13]
  assign sourceE_task_arb_io_in_11_bits_sink = abc_mshr_11_io_tasks_source_e_bits_sink; // @[Slice.scala 472:13]
  assign sourceE_task_arb_io_in_12_valid = abc_mshr_12_io_tasks_source_e_valid; // @[Slice.scala 472:13]
  assign sourceE_task_arb_io_in_12_bits_sink = abc_mshr_12_io_tasks_source_e_bits_sink; // @[Slice.scala 472:13]
  assign sourceE_task_arb_io_in_13_valid = abc_mshr_13_io_tasks_source_e_valid; // @[Slice.scala 472:13]
  assign sourceE_task_arb_io_in_13_bits_sink = abc_mshr_13_io_tasks_source_e_bits_sink; // @[Slice.scala 472:13]
  assign sourceE_task_arb_io_out_ready = sourceE_io_task_ready & _ms_14_io_tasks_source_e_ready_T_1 & ~bc_real_valid_4; // @[Slice.scala 493:60]
  assign sinkC_task_arb_clock = clock;
  assign sinkC_task_arb_reset = reset;
  assign sinkC_task_arb_io_in_0_valid = abc_mshr_0_io_tasks_sink_c_valid; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_0_bits_set = abc_mshr_0_io_tasks_sink_c_bits_set; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_0_bits_tag = abc_mshr_0_io_tasks_sink_c_bits_tag; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_0_bits_way = abc_mshr_0_io_tasks_sink_c_bits_way; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_0_bits_bufIdx = abc_mshr_0_io_tasks_sink_c_bits_bufIdx; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_0_bits_opcode = abc_mshr_0_io_tasks_sink_c_bits_opcode; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_0_bits_source = abc_mshr_0_io_tasks_sink_c_bits_source; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_0_bits_save = abc_mshr_0_io_tasks_sink_c_bits_save; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_0_bits_drop = abc_mshr_0_io_tasks_sink_c_bits_drop; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_0_bits_release = abc_mshr_0_io_tasks_sink_c_bits_release; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_1_valid = abc_mshr_1_io_tasks_sink_c_valid; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_1_bits_set = abc_mshr_1_io_tasks_sink_c_bits_set; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_1_bits_tag = abc_mshr_1_io_tasks_sink_c_bits_tag; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_1_bits_way = abc_mshr_1_io_tasks_sink_c_bits_way; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_1_bits_bufIdx = abc_mshr_1_io_tasks_sink_c_bits_bufIdx; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_1_bits_opcode = abc_mshr_1_io_tasks_sink_c_bits_opcode; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_1_bits_source = abc_mshr_1_io_tasks_sink_c_bits_source; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_1_bits_save = abc_mshr_1_io_tasks_sink_c_bits_save; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_1_bits_drop = abc_mshr_1_io_tasks_sink_c_bits_drop; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_1_bits_release = abc_mshr_1_io_tasks_sink_c_bits_release; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_2_valid = abc_mshr_2_io_tasks_sink_c_valid; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_2_bits_set = abc_mshr_2_io_tasks_sink_c_bits_set; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_2_bits_tag = abc_mshr_2_io_tasks_sink_c_bits_tag; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_2_bits_way = abc_mshr_2_io_tasks_sink_c_bits_way; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_2_bits_bufIdx = abc_mshr_2_io_tasks_sink_c_bits_bufIdx; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_2_bits_opcode = abc_mshr_2_io_tasks_sink_c_bits_opcode; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_2_bits_source = abc_mshr_2_io_tasks_sink_c_bits_source; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_2_bits_save = abc_mshr_2_io_tasks_sink_c_bits_save; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_2_bits_drop = abc_mshr_2_io_tasks_sink_c_bits_drop; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_2_bits_release = abc_mshr_2_io_tasks_sink_c_bits_release; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_3_valid = abc_mshr_3_io_tasks_sink_c_valid; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_3_bits_set = abc_mshr_3_io_tasks_sink_c_bits_set; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_3_bits_tag = abc_mshr_3_io_tasks_sink_c_bits_tag; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_3_bits_way = abc_mshr_3_io_tasks_sink_c_bits_way; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_3_bits_bufIdx = abc_mshr_3_io_tasks_sink_c_bits_bufIdx; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_3_bits_opcode = abc_mshr_3_io_tasks_sink_c_bits_opcode; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_3_bits_source = abc_mshr_3_io_tasks_sink_c_bits_source; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_3_bits_save = abc_mshr_3_io_tasks_sink_c_bits_save; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_3_bits_drop = abc_mshr_3_io_tasks_sink_c_bits_drop; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_3_bits_release = abc_mshr_3_io_tasks_sink_c_bits_release; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_4_valid = abc_mshr_4_io_tasks_sink_c_valid; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_4_bits_set = abc_mshr_4_io_tasks_sink_c_bits_set; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_4_bits_tag = abc_mshr_4_io_tasks_sink_c_bits_tag; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_4_bits_way = abc_mshr_4_io_tasks_sink_c_bits_way; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_4_bits_bufIdx = abc_mshr_4_io_tasks_sink_c_bits_bufIdx; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_4_bits_opcode = abc_mshr_4_io_tasks_sink_c_bits_opcode; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_4_bits_source = abc_mshr_4_io_tasks_sink_c_bits_source; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_4_bits_save = abc_mshr_4_io_tasks_sink_c_bits_save; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_4_bits_drop = abc_mshr_4_io_tasks_sink_c_bits_drop; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_4_bits_release = abc_mshr_4_io_tasks_sink_c_bits_release; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_5_valid = abc_mshr_5_io_tasks_sink_c_valid; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_5_bits_set = abc_mshr_5_io_tasks_sink_c_bits_set; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_5_bits_tag = abc_mshr_5_io_tasks_sink_c_bits_tag; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_5_bits_way = abc_mshr_5_io_tasks_sink_c_bits_way; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_5_bits_bufIdx = abc_mshr_5_io_tasks_sink_c_bits_bufIdx; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_5_bits_opcode = abc_mshr_5_io_tasks_sink_c_bits_opcode; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_5_bits_source = abc_mshr_5_io_tasks_sink_c_bits_source; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_5_bits_save = abc_mshr_5_io_tasks_sink_c_bits_save; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_5_bits_drop = abc_mshr_5_io_tasks_sink_c_bits_drop; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_5_bits_release = abc_mshr_5_io_tasks_sink_c_bits_release; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_6_valid = abc_mshr_6_io_tasks_sink_c_valid; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_6_bits_set = abc_mshr_6_io_tasks_sink_c_bits_set; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_6_bits_tag = abc_mshr_6_io_tasks_sink_c_bits_tag; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_6_bits_way = abc_mshr_6_io_tasks_sink_c_bits_way; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_6_bits_bufIdx = abc_mshr_6_io_tasks_sink_c_bits_bufIdx; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_6_bits_opcode = abc_mshr_6_io_tasks_sink_c_bits_opcode; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_6_bits_source = abc_mshr_6_io_tasks_sink_c_bits_source; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_6_bits_save = abc_mshr_6_io_tasks_sink_c_bits_save; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_6_bits_drop = abc_mshr_6_io_tasks_sink_c_bits_drop; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_6_bits_release = abc_mshr_6_io_tasks_sink_c_bits_release; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_7_valid = abc_mshr_7_io_tasks_sink_c_valid; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_7_bits_set = abc_mshr_7_io_tasks_sink_c_bits_set; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_7_bits_tag = abc_mshr_7_io_tasks_sink_c_bits_tag; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_7_bits_way = abc_mshr_7_io_tasks_sink_c_bits_way; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_7_bits_bufIdx = abc_mshr_7_io_tasks_sink_c_bits_bufIdx; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_7_bits_opcode = abc_mshr_7_io_tasks_sink_c_bits_opcode; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_7_bits_source = abc_mshr_7_io_tasks_sink_c_bits_source; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_7_bits_save = abc_mshr_7_io_tasks_sink_c_bits_save; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_7_bits_drop = abc_mshr_7_io_tasks_sink_c_bits_drop; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_7_bits_release = abc_mshr_7_io_tasks_sink_c_bits_release; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_8_valid = abc_mshr_8_io_tasks_sink_c_valid; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_8_bits_set = abc_mshr_8_io_tasks_sink_c_bits_set; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_8_bits_tag = abc_mshr_8_io_tasks_sink_c_bits_tag; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_8_bits_way = abc_mshr_8_io_tasks_sink_c_bits_way; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_8_bits_bufIdx = abc_mshr_8_io_tasks_sink_c_bits_bufIdx; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_8_bits_opcode = abc_mshr_8_io_tasks_sink_c_bits_opcode; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_8_bits_source = abc_mshr_8_io_tasks_sink_c_bits_source; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_8_bits_save = abc_mshr_8_io_tasks_sink_c_bits_save; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_8_bits_drop = abc_mshr_8_io_tasks_sink_c_bits_drop; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_8_bits_release = abc_mshr_8_io_tasks_sink_c_bits_release; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_9_valid = abc_mshr_9_io_tasks_sink_c_valid; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_9_bits_set = abc_mshr_9_io_tasks_sink_c_bits_set; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_9_bits_tag = abc_mshr_9_io_tasks_sink_c_bits_tag; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_9_bits_way = abc_mshr_9_io_tasks_sink_c_bits_way; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_9_bits_bufIdx = abc_mshr_9_io_tasks_sink_c_bits_bufIdx; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_9_bits_opcode = abc_mshr_9_io_tasks_sink_c_bits_opcode; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_9_bits_source = abc_mshr_9_io_tasks_sink_c_bits_source; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_9_bits_save = abc_mshr_9_io_tasks_sink_c_bits_save; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_9_bits_drop = abc_mshr_9_io_tasks_sink_c_bits_drop; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_9_bits_release = abc_mshr_9_io_tasks_sink_c_bits_release; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_10_valid = abc_mshr_10_io_tasks_sink_c_valid; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_10_bits_set = abc_mshr_10_io_tasks_sink_c_bits_set; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_10_bits_tag = abc_mshr_10_io_tasks_sink_c_bits_tag; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_10_bits_way = abc_mshr_10_io_tasks_sink_c_bits_way; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_10_bits_bufIdx = abc_mshr_10_io_tasks_sink_c_bits_bufIdx; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_10_bits_opcode = abc_mshr_10_io_tasks_sink_c_bits_opcode; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_10_bits_source = abc_mshr_10_io_tasks_sink_c_bits_source; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_10_bits_save = abc_mshr_10_io_tasks_sink_c_bits_save; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_10_bits_drop = abc_mshr_10_io_tasks_sink_c_bits_drop; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_10_bits_release = abc_mshr_10_io_tasks_sink_c_bits_release; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_11_valid = abc_mshr_11_io_tasks_sink_c_valid; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_11_bits_set = abc_mshr_11_io_tasks_sink_c_bits_set; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_11_bits_tag = abc_mshr_11_io_tasks_sink_c_bits_tag; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_11_bits_way = abc_mshr_11_io_tasks_sink_c_bits_way; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_11_bits_bufIdx = abc_mshr_11_io_tasks_sink_c_bits_bufIdx; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_11_bits_opcode = abc_mshr_11_io_tasks_sink_c_bits_opcode; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_11_bits_source = abc_mshr_11_io_tasks_sink_c_bits_source; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_11_bits_save = abc_mshr_11_io_tasks_sink_c_bits_save; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_11_bits_drop = abc_mshr_11_io_tasks_sink_c_bits_drop; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_11_bits_release = abc_mshr_11_io_tasks_sink_c_bits_release; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_12_valid = abc_mshr_12_io_tasks_sink_c_valid; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_12_bits_set = abc_mshr_12_io_tasks_sink_c_bits_set; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_12_bits_tag = abc_mshr_12_io_tasks_sink_c_bits_tag; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_12_bits_way = abc_mshr_12_io_tasks_sink_c_bits_way; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_12_bits_bufIdx = abc_mshr_12_io_tasks_sink_c_bits_bufIdx; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_12_bits_opcode = abc_mshr_12_io_tasks_sink_c_bits_opcode; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_12_bits_source = abc_mshr_12_io_tasks_sink_c_bits_source; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_12_bits_save = abc_mshr_12_io_tasks_sink_c_bits_save; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_12_bits_drop = abc_mshr_12_io_tasks_sink_c_bits_drop; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_12_bits_release = abc_mshr_12_io_tasks_sink_c_bits_release; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_13_valid = abc_mshr_13_io_tasks_sink_c_valid; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_13_bits_set = abc_mshr_13_io_tasks_sink_c_bits_set; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_13_bits_tag = abc_mshr_13_io_tasks_sink_c_bits_tag; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_13_bits_way = abc_mshr_13_io_tasks_sink_c_bits_way; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_13_bits_bufIdx = abc_mshr_13_io_tasks_sink_c_bits_bufIdx; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_13_bits_opcode = abc_mshr_13_io_tasks_sink_c_bits_opcode; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_13_bits_source = abc_mshr_13_io_tasks_sink_c_bits_source; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_13_bits_save = abc_mshr_13_io_tasks_sink_c_bits_save; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_13_bits_drop = abc_mshr_13_io_tasks_sink_c_bits_drop; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_in_13_bits_release = abc_mshr_13_io_tasks_sink_c_bits_release; // @[Slice.scala 472:13]
  assign sinkC_task_arb_io_out_ready = sinkC_io_task_ready & _ms_14_io_tasks_sink_c_ready_T_1 & ~bc_real_valid_6; // @[Slice.scala 493:60]
  assign pipeline_1_clock = clock;
  assign pipeline_1_reset = reset;
  assign pipeline_1_io_in_valid = c_real_valid_7 | bc_real_valid_7 | tagWrite_task_arb_io_out_valid; // @[Slice.scala 489:52]
  assign pipeline_1_io_in_bits_set = c_real_valid_7 ? c_bits_latch_7_set : _pipeline_io_in_bits_T_set; // @[Slice.scala 490:24]
  assign pipeline_1_io_in_bits_way = c_real_valid_7 ? c_bits_latch_7_way : _pipeline_io_in_bits_T_way; // @[Slice.scala 490:24]
  assign pipeline_1_io_in_bits_tag = c_real_valid_7 ? c_bits_latch_7_tag : _pipeline_io_in_bits_T_tag; // @[Slice.scala 490:24]
  assign tagWrite_task_arb_clock = clock;
  assign tagWrite_task_arb_reset = reset;
  assign tagWrite_task_arb_io_in_0_valid = abc_mshr_0_io_tasks_tag_write_valid; // @[Slice.scala 472:13]
  assign tagWrite_task_arb_io_in_0_bits_set = abc_mshr_0_io_tasks_tag_write_bits_set; // @[Slice.scala 472:13]
  assign tagWrite_task_arb_io_in_0_bits_way = abc_mshr_0_io_tasks_tag_write_bits_way; // @[Slice.scala 472:13]
  assign tagWrite_task_arb_io_in_0_bits_tag = abc_mshr_0_io_tasks_tag_write_bits_tag; // @[Slice.scala 472:13]
  assign tagWrite_task_arb_io_in_1_valid = abc_mshr_1_io_tasks_tag_write_valid; // @[Slice.scala 472:13]
  assign tagWrite_task_arb_io_in_1_bits_set = abc_mshr_1_io_tasks_tag_write_bits_set; // @[Slice.scala 472:13]
  assign tagWrite_task_arb_io_in_1_bits_way = abc_mshr_1_io_tasks_tag_write_bits_way; // @[Slice.scala 472:13]
  assign tagWrite_task_arb_io_in_1_bits_tag = abc_mshr_1_io_tasks_tag_write_bits_tag; // @[Slice.scala 472:13]
  assign tagWrite_task_arb_io_in_2_valid = abc_mshr_2_io_tasks_tag_write_valid; // @[Slice.scala 472:13]
  assign tagWrite_task_arb_io_in_2_bits_set = abc_mshr_2_io_tasks_tag_write_bits_set; // @[Slice.scala 472:13]
  assign tagWrite_task_arb_io_in_2_bits_way = abc_mshr_2_io_tasks_tag_write_bits_way; // @[Slice.scala 472:13]
  assign tagWrite_task_arb_io_in_2_bits_tag = abc_mshr_2_io_tasks_tag_write_bits_tag; // @[Slice.scala 472:13]
  assign tagWrite_task_arb_io_in_3_valid = abc_mshr_3_io_tasks_tag_write_valid; // @[Slice.scala 472:13]
  assign tagWrite_task_arb_io_in_3_bits_set = abc_mshr_3_io_tasks_tag_write_bits_set; // @[Slice.scala 472:13]
  assign tagWrite_task_arb_io_in_3_bits_way = abc_mshr_3_io_tasks_tag_write_bits_way; // @[Slice.scala 472:13]
  assign tagWrite_task_arb_io_in_3_bits_tag = abc_mshr_3_io_tasks_tag_write_bits_tag; // @[Slice.scala 472:13]
  assign tagWrite_task_arb_io_in_4_valid = abc_mshr_4_io_tasks_tag_write_valid; // @[Slice.scala 472:13]
  assign tagWrite_task_arb_io_in_4_bits_set = abc_mshr_4_io_tasks_tag_write_bits_set; // @[Slice.scala 472:13]
  assign tagWrite_task_arb_io_in_4_bits_way = abc_mshr_4_io_tasks_tag_write_bits_way; // @[Slice.scala 472:13]
  assign tagWrite_task_arb_io_in_4_bits_tag = abc_mshr_4_io_tasks_tag_write_bits_tag; // @[Slice.scala 472:13]
  assign tagWrite_task_arb_io_in_5_valid = abc_mshr_5_io_tasks_tag_write_valid; // @[Slice.scala 472:13]
  assign tagWrite_task_arb_io_in_5_bits_set = abc_mshr_5_io_tasks_tag_write_bits_set; // @[Slice.scala 472:13]
  assign tagWrite_task_arb_io_in_5_bits_way = abc_mshr_5_io_tasks_tag_write_bits_way; // @[Slice.scala 472:13]
  assign tagWrite_task_arb_io_in_5_bits_tag = abc_mshr_5_io_tasks_tag_write_bits_tag; // @[Slice.scala 472:13]
  assign tagWrite_task_arb_io_in_6_valid = abc_mshr_6_io_tasks_tag_write_valid; // @[Slice.scala 472:13]
  assign tagWrite_task_arb_io_in_6_bits_set = abc_mshr_6_io_tasks_tag_write_bits_set; // @[Slice.scala 472:13]
  assign tagWrite_task_arb_io_in_6_bits_way = abc_mshr_6_io_tasks_tag_write_bits_way; // @[Slice.scala 472:13]
  assign tagWrite_task_arb_io_in_6_bits_tag = abc_mshr_6_io_tasks_tag_write_bits_tag; // @[Slice.scala 472:13]
  assign tagWrite_task_arb_io_in_7_valid = abc_mshr_7_io_tasks_tag_write_valid; // @[Slice.scala 472:13]
  assign tagWrite_task_arb_io_in_7_bits_set = abc_mshr_7_io_tasks_tag_write_bits_set; // @[Slice.scala 472:13]
  assign tagWrite_task_arb_io_in_7_bits_way = abc_mshr_7_io_tasks_tag_write_bits_way; // @[Slice.scala 472:13]
  assign tagWrite_task_arb_io_in_7_bits_tag = abc_mshr_7_io_tasks_tag_write_bits_tag; // @[Slice.scala 472:13]
  assign tagWrite_task_arb_io_in_8_valid = abc_mshr_8_io_tasks_tag_write_valid; // @[Slice.scala 472:13]
  assign tagWrite_task_arb_io_in_8_bits_set = abc_mshr_8_io_tasks_tag_write_bits_set; // @[Slice.scala 472:13]
  assign tagWrite_task_arb_io_in_8_bits_way = abc_mshr_8_io_tasks_tag_write_bits_way; // @[Slice.scala 472:13]
  assign tagWrite_task_arb_io_in_8_bits_tag = abc_mshr_8_io_tasks_tag_write_bits_tag; // @[Slice.scala 472:13]
  assign tagWrite_task_arb_io_in_9_valid = abc_mshr_9_io_tasks_tag_write_valid; // @[Slice.scala 472:13]
  assign tagWrite_task_arb_io_in_9_bits_set = abc_mshr_9_io_tasks_tag_write_bits_set; // @[Slice.scala 472:13]
  assign tagWrite_task_arb_io_in_9_bits_way = abc_mshr_9_io_tasks_tag_write_bits_way; // @[Slice.scala 472:13]
  assign tagWrite_task_arb_io_in_9_bits_tag = abc_mshr_9_io_tasks_tag_write_bits_tag; // @[Slice.scala 472:13]
  assign tagWrite_task_arb_io_in_10_valid = abc_mshr_10_io_tasks_tag_write_valid; // @[Slice.scala 472:13]
  assign tagWrite_task_arb_io_in_10_bits_set = abc_mshr_10_io_tasks_tag_write_bits_set; // @[Slice.scala 472:13]
  assign tagWrite_task_arb_io_in_10_bits_way = abc_mshr_10_io_tasks_tag_write_bits_way; // @[Slice.scala 472:13]
  assign tagWrite_task_arb_io_in_10_bits_tag = abc_mshr_10_io_tasks_tag_write_bits_tag; // @[Slice.scala 472:13]
  assign tagWrite_task_arb_io_in_11_valid = abc_mshr_11_io_tasks_tag_write_valid; // @[Slice.scala 472:13]
  assign tagWrite_task_arb_io_in_11_bits_set = abc_mshr_11_io_tasks_tag_write_bits_set; // @[Slice.scala 472:13]
  assign tagWrite_task_arb_io_in_11_bits_way = abc_mshr_11_io_tasks_tag_write_bits_way; // @[Slice.scala 472:13]
  assign tagWrite_task_arb_io_in_11_bits_tag = abc_mshr_11_io_tasks_tag_write_bits_tag; // @[Slice.scala 472:13]
  assign tagWrite_task_arb_io_in_12_valid = abc_mshr_12_io_tasks_tag_write_valid; // @[Slice.scala 472:13]
  assign tagWrite_task_arb_io_in_12_bits_set = abc_mshr_12_io_tasks_tag_write_bits_set; // @[Slice.scala 472:13]
  assign tagWrite_task_arb_io_in_12_bits_way = abc_mshr_12_io_tasks_tag_write_bits_way; // @[Slice.scala 472:13]
  assign tagWrite_task_arb_io_in_12_bits_tag = abc_mshr_12_io_tasks_tag_write_bits_tag; // @[Slice.scala 472:13]
  assign tagWrite_task_arb_io_in_13_valid = abc_mshr_13_io_tasks_tag_write_valid; // @[Slice.scala 472:13]
  assign tagWrite_task_arb_io_in_13_bits_set = abc_mshr_13_io_tasks_tag_write_bits_set; // @[Slice.scala 472:13]
  assign tagWrite_task_arb_io_in_13_bits_way = abc_mshr_13_io_tasks_tag_write_bits_way; // @[Slice.scala 472:13]
  assign tagWrite_task_arb_io_in_13_bits_tag = abc_mshr_13_io_tasks_tag_write_bits_tag; // @[Slice.scala 472:13]
  assign tagWrite_task_arb_io_out_ready = _ms_14_io_tasks_tag_write_ready_T_1 & ~bc_real_valid_7; // @[Slice.scala 493:60]
  assign pipeline_2_clock = clock;
  assign pipeline_2_reset = reset;
  assign pipeline_2_io_in_valid = arbiter_1_io_out_valid; // @[Slice.scala 409:10]
  assign pipeline_2_io_in_bits_set = arbiter_1_io_out_bits_set; // @[Slice.scala 409:10]
  assign pipeline_2_io_in_bits_way = arbiter_1_io_out_bits_way; // @[Slice.scala 409:10]
  assign pipeline_2_io_in_bits_data_0_state = arbiter_1_io_out_bits_data_0_state; // @[Slice.scala 409:10]
  assign pipeline_2_io_in_bits_data_1_state = arbiter_1_io_out_bits_data_1_state; // @[Slice.scala 409:10]
  assign arbiter_1_clock = clock;
  assign arbiter_1_reset = reset;
  assign arbiter_1_io_in_0_valid = abc_mshr_0_io_tasks_client_dir_write_valid; // @[Slice.scala 406:60]
  assign arbiter_1_io_in_0_bits_set = abc_mshr_0_io_tasks_client_dir_write_bits_set; // @[Slice.scala 406:60]
  assign arbiter_1_io_in_0_bits_way = abc_mshr_0_io_tasks_client_dir_write_bits_way; // @[Slice.scala 406:60]
  assign arbiter_1_io_in_0_bits_data_0_state = abc_mshr_0_io_tasks_client_dir_write_bits_data_0_state; // @[Slice.scala 406:60]
  assign arbiter_1_io_in_0_bits_data_1_state = abc_mshr_0_io_tasks_client_dir_write_bits_data_1_state; // @[Slice.scala 406:60]
  assign arbiter_1_io_in_1_valid = abc_mshr_1_io_tasks_client_dir_write_valid; // @[Slice.scala 406:60]
  assign arbiter_1_io_in_1_bits_set = abc_mshr_1_io_tasks_client_dir_write_bits_set; // @[Slice.scala 406:60]
  assign arbiter_1_io_in_1_bits_way = abc_mshr_1_io_tasks_client_dir_write_bits_way; // @[Slice.scala 406:60]
  assign arbiter_1_io_in_1_bits_data_0_state = abc_mshr_1_io_tasks_client_dir_write_bits_data_0_state; // @[Slice.scala 406:60]
  assign arbiter_1_io_in_1_bits_data_1_state = abc_mshr_1_io_tasks_client_dir_write_bits_data_1_state; // @[Slice.scala 406:60]
  assign arbiter_1_io_in_2_valid = abc_mshr_2_io_tasks_client_dir_write_valid; // @[Slice.scala 406:60]
  assign arbiter_1_io_in_2_bits_set = abc_mshr_2_io_tasks_client_dir_write_bits_set; // @[Slice.scala 406:60]
  assign arbiter_1_io_in_2_bits_way = abc_mshr_2_io_tasks_client_dir_write_bits_way; // @[Slice.scala 406:60]
  assign arbiter_1_io_in_2_bits_data_0_state = abc_mshr_2_io_tasks_client_dir_write_bits_data_0_state; // @[Slice.scala 406:60]
  assign arbiter_1_io_in_2_bits_data_1_state = abc_mshr_2_io_tasks_client_dir_write_bits_data_1_state; // @[Slice.scala 406:60]
  assign arbiter_1_io_in_3_valid = abc_mshr_3_io_tasks_client_dir_write_valid; // @[Slice.scala 406:60]
  assign arbiter_1_io_in_3_bits_set = abc_mshr_3_io_tasks_client_dir_write_bits_set; // @[Slice.scala 406:60]
  assign arbiter_1_io_in_3_bits_way = abc_mshr_3_io_tasks_client_dir_write_bits_way; // @[Slice.scala 406:60]
  assign arbiter_1_io_in_3_bits_data_0_state = abc_mshr_3_io_tasks_client_dir_write_bits_data_0_state; // @[Slice.scala 406:60]
  assign arbiter_1_io_in_3_bits_data_1_state = abc_mshr_3_io_tasks_client_dir_write_bits_data_1_state; // @[Slice.scala 406:60]
  assign arbiter_1_io_in_4_valid = abc_mshr_4_io_tasks_client_dir_write_valid; // @[Slice.scala 406:60]
  assign arbiter_1_io_in_4_bits_set = abc_mshr_4_io_tasks_client_dir_write_bits_set; // @[Slice.scala 406:60]
  assign arbiter_1_io_in_4_bits_way = abc_mshr_4_io_tasks_client_dir_write_bits_way; // @[Slice.scala 406:60]
  assign arbiter_1_io_in_4_bits_data_0_state = abc_mshr_4_io_tasks_client_dir_write_bits_data_0_state; // @[Slice.scala 406:60]
  assign arbiter_1_io_in_4_bits_data_1_state = abc_mshr_4_io_tasks_client_dir_write_bits_data_1_state; // @[Slice.scala 406:60]
  assign arbiter_1_io_in_5_valid = abc_mshr_5_io_tasks_client_dir_write_valid; // @[Slice.scala 406:60]
  assign arbiter_1_io_in_5_bits_set = abc_mshr_5_io_tasks_client_dir_write_bits_set; // @[Slice.scala 406:60]
  assign arbiter_1_io_in_5_bits_way = abc_mshr_5_io_tasks_client_dir_write_bits_way; // @[Slice.scala 406:60]
  assign arbiter_1_io_in_5_bits_data_0_state = abc_mshr_5_io_tasks_client_dir_write_bits_data_0_state; // @[Slice.scala 406:60]
  assign arbiter_1_io_in_5_bits_data_1_state = abc_mshr_5_io_tasks_client_dir_write_bits_data_1_state; // @[Slice.scala 406:60]
  assign arbiter_1_io_in_6_valid = abc_mshr_6_io_tasks_client_dir_write_valid; // @[Slice.scala 406:60]
  assign arbiter_1_io_in_6_bits_set = abc_mshr_6_io_tasks_client_dir_write_bits_set; // @[Slice.scala 406:60]
  assign arbiter_1_io_in_6_bits_way = abc_mshr_6_io_tasks_client_dir_write_bits_way; // @[Slice.scala 406:60]
  assign arbiter_1_io_in_6_bits_data_0_state = abc_mshr_6_io_tasks_client_dir_write_bits_data_0_state; // @[Slice.scala 406:60]
  assign arbiter_1_io_in_6_bits_data_1_state = abc_mshr_6_io_tasks_client_dir_write_bits_data_1_state; // @[Slice.scala 406:60]
  assign arbiter_1_io_in_7_valid = abc_mshr_7_io_tasks_client_dir_write_valid; // @[Slice.scala 406:60]
  assign arbiter_1_io_in_7_bits_set = abc_mshr_7_io_tasks_client_dir_write_bits_set; // @[Slice.scala 406:60]
  assign arbiter_1_io_in_7_bits_way = abc_mshr_7_io_tasks_client_dir_write_bits_way; // @[Slice.scala 406:60]
  assign arbiter_1_io_in_7_bits_data_0_state = abc_mshr_7_io_tasks_client_dir_write_bits_data_0_state; // @[Slice.scala 406:60]
  assign arbiter_1_io_in_7_bits_data_1_state = abc_mshr_7_io_tasks_client_dir_write_bits_data_1_state; // @[Slice.scala 406:60]
  assign arbiter_1_io_in_8_valid = abc_mshr_8_io_tasks_client_dir_write_valid; // @[Slice.scala 406:60]
  assign arbiter_1_io_in_8_bits_set = abc_mshr_8_io_tasks_client_dir_write_bits_set; // @[Slice.scala 406:60]
  assign arbiter_1_io_in_8_bits_way = abc_mshr_8_io_tasks_client_dir_write_bits_way; // @[Slice.scala 406:60]
  assign arbiter_1_io_in_8_bits_data_0_state = abc_mshr_8_io_tasks_client_dir_write_bits_data_0_state; // @[Slice.scala 406:60]
  assign arbiter_1_io_in_8_bits_data_1_state = abc_mshr_8_io_tasks_client_dir_write_bits_data_1_state; // @[Slice.scala 406:60]
  assign arbiter_1_io_in_9_valid = abc_mshr_9_io_tasks_client_dir_write_valid; // @[Slice.scala 406:60]
  assign arbiter_1_io_in_9_bits_set = abc_mshr_9_io_tasks_client_dir_write_bits_set; // @[Slice.scala 406:60]
  assign arbiter_1_io_in_9_bits_way = abc_mshr_9_io_tasks_client_dir_write_bits_way; // @[Slice.scala 406:60]
  assign arbiter_1_io_in_9_bits_data_0_state = abc_mshr_9_io_tasks_client_dir_write_bits_data_0_state; // @[Slice.scala 406:60]
  assign arbiter_1_io_in_9_bits_data_1_state = abc_mshr_9_io_tasks_client_dir_write_bits_data_1_state; // @[Slice.scala 406:60]
  assign arbiter_1_io_in_10_valid = abc_mshr_10_io_tasks_client_dir_write_valid; // @[Slice.scala 406:60]
  assign arbiter_1_io_in_10_bits_set = abc_mshr_10_io_tasks_client_dir_write_bits_set; // @[Slice.scala 406:60]
  assign arbiter_1_io_in_10_bits_way = abc_mshr_10_io_tasks_client_dir_write_bits_way; // @[Slice.scala 406:60]
  assign arbiter_1_io_in_10_bits_data_0_state = abc_mshr_10_io_tasks_client_dir_write_bits_data_0_state; // @[Slice.scala 406:60]
  assign arbiter_1_io_in_10_bits_data_1_state = abc_mshr_10_io_tasks_client_dir_write_bits_data_1_state; // @[Slice.scala 406:60]
  assign arbiter_1_io_in_11_valid = abc_mshr_11_io_tasks_client_dir_write_valid; // @[Slice.scala 406:60]
  assign arbiter_1_io_in_11_bits_set = abc_mshr_11_io_tasks_client_dir_write_bits_set; // @[Slice.scala 406:60]
  assign arbiter_1_io_in_11_bits_way = abc_mshr_11_io_tasks_client_dir_write_bits_way; // @[Slice.scala 406:60]
  assign arbiter_1_io_in_11_bits_data_0_state = abc_mshr_11_io_tasks_client_dir_write_bits_data_0_state; // @[Slice.scala 406:60]
  assign arbiter_1_io_in_11_bits_data_1_state = abc_mshr_11_io_tasks_client_dir_write_bits_data_1_state; // @[Slice.scala 406:60]
  assign arbiter_1_io_in_12_valid = abc_mshr_12_io_tasks_client_dir_write_valid; // @[Slice.scala 406:60]
  assign arbiter_1_io_in_12_bits_set = abc_mshr_12_io_tasks_client_dir_write_bits_set; // @[Slice.scala 406:60]
  assign arbiter_1_io_in_12_bits_way = abc_mshr_12_io_tasks_client_dir_write_bits_way; // @[Slice.scala 406:60]
  assign arbiter_1_io_in_12_bits_data_0_state = abc_mshr_12_io_tasks_client_dir_write_bits_data_0_state; // @[Slice.scala 406:60]
  assign arbiter_1_io_in_12_bits_data_1_state = abc_mshr_12_io_tasks_client_dir_write_bits_data_1_state; // @[Slice.scala 406:60]
  assign arbiter_1_io_in_13_valid = abc_mshr_13_io_tasks_client_dir_write_valid; // @[Slice.scala 406:60]
  assign arbiter_1_io_in_13_bits_set = abc_mshr_13_io_tasks_client_dir_write_bits_set; // @[Slice.scala 406:60]
  assign arbiter_1_io_in_13_bits_way = abc_mshr_13_io_tasks_client_dir_write_bits_way; // @[Slice.scala 406:60]
  assign arbiter_1_io_in_13_bits_data_0_state = abc_mshr_13_io_tasks_client_dir_write_bits_data_0_state; // @[Slice.scala 406:60]
  assign arbiter_1_io_in_13_bits_data_1_state = abc_mshr_13_io_tasks_client_dir_write_bits_data_1_state; // @[Slice.scala 406:60]
  assign arbiter_1_io_in_14_valid = _nestedWb_btoN_T & bc_mshr_io_tasks_client_dir_write_valid; // @[Slice.scala 389:26]
  assign arbiter_1_io_in_14_bits_set = bc_mshr_io_tasks_client_dir_write_bits_set; // @[Slice.scala 390:15]
  assign arbiter_1_io_in_14_bits_way = bc_mshr_io_tasks_client_dir_write_bits_way; // @[Slice.scala 390:15]
  assign arbiter_1_io_in_14_bits_data_0_state = bc_mshr_io_tasks_client_dir_write_bits_data_0_state; // @[Slice.scala 390:15]
  assign arbiter_1_io_in_14_bits_data_1_state = bc_mshr_io_tasks_client_dir_write_bits_data_1_state; // @[Slice.scala 390:15]
  assign arbiter_1_io_in_15_valid = c_mshr_io_tasks_client_dir_write_valid; // @[Slice.scala 408:24]
  assign arbiter_1_io_in_15_bits_set = c_mshr_io_tasks_client_dir_write_bits_set; // @[Slice.scala 408:24]
  assign arbiter_1_io_in_15_bits_way = c_mshr_io_tasks_client_dir_write_bits_way; // @[Slice.scala 408:24]
  assign arbiter_1_io_in_15_bits_data_0_state = c_mshr_io_tasks_client_dir_write_bits_data_0_state; // @[Slice.scala 408:24]
  assign arbiter_1_io_in_15_bits_data_1_state = c_mshr_io_tasks_client_dir_write_bits_data_1_state; // @[Slice.scala 408:24]
  assign pipeline_3_clock = clock;
  assign pipeline_3_reset = reset;
  assign pipeline_3_io_in_valid = c_real_valid_8 | bc_real_valid_8 | arbiter_2_io_out_valid; // @[Slice.scala 489:52]
  assign pipeline_3_io_in_bits_set = c_real_valid_8 ? c_bits_latch_8_set : _pipeline_io_in_bits_T_2_set; // @[Slice.scala 490:24]
  assign pipeline_3_io_in_bits_way = c_real_valid_8 ? c_bits_latch_8_way : _pipeline_io_in_bits_T_2_way; // @[Slice.scala 490:24]
  assign pipeline_3_io_in_bits_tag = c_real_valid_8 ? c_bits_latch_8_tag : _pipeline_io_in_bits_T_2_tag; // @[Slice.scala 490:24]
  assign arbiter_2_clock = clock;
  assign arbiter_2_reset = reset;
  assign arbiter_2_io_in_0_valid = abc_mshr_0_io_tasks_client_tag_write_valid; // @[Slice.scala 472:13]
  assign arbiter_2_io_in_0_bits_set = abc_mshr_0_io_tasks_client_tag_write_bits_set; // @[Slice.scala 472:13]
  assign arbiter_2_io_in_0_bits_way = abc_mshr_0_io_tasks_client_tag_write_bits_way; // @[Slice.scala 472:13]
  assign arbiter_2_io_in_0_bits_tag = abc_mshr_0_io_tasks_client_tag_write_bits_tag; // @[Slice.scala 472:13]
  assign arbiter_2_io_in_1_valid = abc_mshr_1_io_tasks_client_tag_write_valid; // @[Slice.scala 472:13]
  assign arbiter_2_io_in_1_bits_set = abc_mshr_1_io_tasks_client_tag_write_bits_set; // @[Slice.scala 472:13]
  assign arbiter_2_io_in_1_bits_way = abc_mshr_1_io_tasks_client_tag_write_bits_way; // @[Slice.scala 472:13]
  assign arbiter_2_io_in_1_bits_tag = abc_mshr_1_io_tasks_client_tag_write_bits_tag; // @[Slice.scala 472:13]
  assign arbiter_2_io_in_2_valid = abc_mshr_2_io_tasks_client_tag_write_valid; // @[Slice.scala 472:13]
  assign arbiter_2_io_in_2_bits_set = abc_mshr_2_io_tasks_client_tag_write_bits_set; // @[Slice.scala 472:13]
  assign arbiter_2_io_in_2_bits_way = abc_mshr_2_io_tasks_client_tag_write_bits_way; // @[Slice.scala 472:13]
  assign arbiter_2_io_in_2_bits_tag = abc_mshr_2_io_tasks_client_tag_write_bits_tag; // @[Slice.scala 472:13]
  assign arbiter_2_io_in_3_valid = abc_mshr_3_io_tasks_client_tag_write_valid; // @[Slice.scala 472:13]
  assign arbiter_2_io_in_3_bits_set = abc_mshr_3_io_tasks_client_tag_write_bits_set; // @[Slice.scala 472:13]
  assign arbiter_2_io_in_3_bits_way = abc_mshr_3_io_tasks_client_tag_write_bits_way; // @[Slice.scala 472:13]
  assign arbiter_2_io_in_3_bits_tag = abc_mshr_3_io_tasks_client_tag_write_bits_tag; // @[Slice.scala 472:13]
  assign arbiter_2_io_in_4_valid = abc_mshr_4_io_tasks_client_tag_write_valid; // @[Slice.scala 472:13]
  assign arbiter_2_io_in_4_bits_set = abc_mshr_4_io_tasks_client_tag_write_bits_set; // @[Slice.scala 472:13]
  assign arbiter_2_io_in_4_bits_way = abc_mshr_4_io_tasks_client_tag_write_bits_way; // @[Slice.scala 472:13]
  assign arbiter_2_io_in_4_bits_tag = abc_mshr_4_io_tasks_client_tag_write_bits_tag; // @[Slice.scala 472:13]
  assign arbiter_2_io_in_5_valid = abc_mshr_5_io_tasks_client_tag_write_valid; // @[Slice.scala 472:13]
  assign arbiter_2_io_in_5_bits_set = abc_mshr_5_io_tasks_client_tag_write_bits_set; // @[Slice.scala 472:13]
  assign arbiter_2_io_in_5_bits_way = abc_mshr_5_io_tasks_client_tag_write_bits_way; // @[Slice.scala 472:13]
  assign arbiter_2_io_in_5_bits_tag = abc_mshr_5_io_tasks_client_tag_write_bits_tag; // @[Slice.scala 472:13]
  assign arbiter_2_io_in_6_valid = abc_mshr_6_io_tasks_client_tag_write_valid; // @[Slice.scala 472:13]
  assign arbiter_2_io_in_6_bits_set = abc_mshr_6_io_tasks_client_tag_write_bits_set; // @[Slice.scala 472:13]
  assign arbiter_2_io_in_6_bits_way = abc_mshr_6_io_tasks_client_tag_write_bits_way; // @[Slice.scala 472:13]
  assign arbiter_2_io_in_6_bits_tag = abc_mshr_6_io_tasks_client_tag_write_bits_tag; // @[Slice.scala 472:13]
  assign arbiter_2_io_in_7_valid = abc_mshr_7_io_tasks_client_tag_write_valid; // @[Slice.scala 472:13]
  assign arbiter_2_io_in_7_bits_set = abc_mshr_7_io_tasks_client_tag_write_bits_set; // @[Slice.scala 472:13]
  assign arbiter_2_io_in_7_bits_way = abc_mshr_7_io_tasks_client_tag_write_bits_way; // @[Slice.scala 472:13]
  assign arbiter_2_io_in_7_bits_tag = abc_mshr_7_io_tasks_client_tag_write_bits_tag; // @[Slice.scala 472:13]
  assign arbiter_2_io_in_8_valid = abc_mshr_8_io_tasks_client_tag_write_valid; // @[Slice.scala 472:13]
  assign arbiter_2_io_in_8_bits_set = abc_mshr_8_io_tasks_client_tag_write_bits_set; // @[Slice.scala 472:13]
  assign arbiter_2_io_in_8_bits_way = abc_mshr_8_io_tasks_client_tag_write_bits_way; // @[Slice.scala 472:13]
  assign arbiter_2_io_in_8_bits_tag = abc_mshr_8_io_tasks_client_tag_write_bits_tag; // @[Slice.scala 472:13]
  assign arbiter_2_io_in_9_valid = abc_mshr_9_io_tasks_client_tag_write_valid; // @[Slice.scala 472:13]
  assign arbiter_2_io_in_9_bits_set = abc_mshr_9_io_tasks_client_tag_write_bits_set; // @[Slice.scala 472:13]
  assign arbiter_2_io_in_9_bits_way = abc_mshr_9_io_tasks_client_tag_write_bits_way; // @[Slice.scala 472:13]
  assign arbiter_2_io_in_9_bits_tag = abc_mshr_9_io_tasks_client_tag_write_bits_tag; // @[Slice.scala 472:13]
  assign arbiter_2_io_in_10_valid = abc_mshr_10_io_tasks_client_tag_write_valid; // @[Slice.scala 472:13]
  assign arbiter_2_io_in_10_bits_set = abc_mshr_10_io_tasks_client_tag_write_bits_set; // @[Slice.scala 472:13]
  assign arbiter_2_io_in_10_bits_way = abc_mshr_10_io_tasks_client_tag_write_bits_way; // @[Slice.scala 472:13]
  assign arbiter_2_io_in_10_bits_tag = abc_mshr_10_io_tasks_client_tag_write_bits_tag; // @[Slice.scala 472:13]
  assign arbiter_2_io_in_11_valid = abc_mshr_11_io_tasks_client_tag_write_valid; // @[Slice.scala 472:13]
  assign arbiter_2_io_in_11_bits_set = abc_mshr_11_io_tasks_client_tag_write_bits_set; // @[Slice.scala 472:13]
  assign arbiter_2_io_in_11_bits_way = abc_mshr_11_io_tasks_client_tag_write_bits_way; // @[Slice.scala 472:13]
  assign arbiter_2_io_in_11_bits_tag = abc_mshr_11_io_tasks_client_tag_write_bits_tag; // @[Slice.scala 472:13]
  assign arbiter_2_io_in_12_valid = abc_mshr_12_io_tasks_client_tag_write_valid; // @[Slice.scala 472:13]
  assign arbiter_2_io_in_12_bits_set = abc_mshr_12_io_tasks_client_tag_write_bits_set; // @[Slice.scala 472:13]
  assign arbiter_2_io_in_12_bits_way = abc_mshr_12_io_tasks_client_tag_write_bits_way; // @[Slice.scala 472:13]
  assign arbiter_2_io_in_12_bits_tag = abc_mshr_12_io_tasks_client_tag_write_bits_tag; // @[Slice.scala 472:13]
  assign arbiter_2_io_in_13_valid = abc_mshr_13_io_tasks_client_tag_write_valid; // @[Slice.scala 472:13]
  assign arbiter_2_io_in_13_bits_set = abc_mshr_13_io_tasks_client_tag_write_bits_set; // @[Slice.scala 472:13]
  assign arbiter_2_io_in_13_bits_way = abc_mshr_13_io_tasks_client_tag_write_bits_way; // @[Slice.scala 472:13]
  assign arbiter_2_io_in_13_bits_tag = abc_mshr_13_io_tasks_client_tag_write_bits_tag; // @[Slice.scala 472:13]
  assign arbiter_2_io_out_ready = _ms_14_io_tasks_client_tag_write_ready_T_1 & ~bc_real_valid_8; // @[Slice.scala 493:60]
  always @(posedge clock) begin
    if (bc_mshr_io_tasks_source_a_valid) begin // @[Reg.scala 17:18]
      bc_bits_latch_tag <= bc_mshr_io_tasks_source_a_bits_tag; // @[Reg.scala 17:22]
    end
    if (bc_mshr_io_tasks_source_a_valid) begin // @[Reg.scala 17:18]
      bc_bits_latch_set <= bc_mshr_io_tasks_source_a_bits_set; // @[Reg.scala 17:22]
    end
    if (bc_mshr_io_tasks_source_a_valid) begin // @[Reg.scala 17:18]
      bc_bits_latch_off <= bc_mshr_io_tasks_source_a_bits_off; // @[Reg.scala 17:22]
    end
    if (bc_mshr_io_tasks_source_a_valid) begin // @[Reg.scala 17:18]
      bc_bits_latch_opcode <= bc_mshr_io_tasks_source_a_bits_opcode; // @[Reg.scala 17:22]
    end
    if (bc_mshr_io_tasks_source_a_valid) begin // @[Reg.scala 17:18]
      bc_bits_latch_param <= bc_mshr_io_tasks_source_a_bits_param; // @[Reg.scala 17:22]
    end
    if (bc_mshr_io_tasks_source_a_valid) begin // @[Reg.scala 17:18]
      bc_bits_latch_source <= bc_mshr_io_tasks_source_a_bits_source; // @[Reg.scala 17:22]
    end
    if (bc_mshr_io_tasks_source_a_valid) begin // @[Reg.scala 17:18]
      bc_bits_latch_bufIdx <= bc_mshr_io_tasks_source_a_bits_bufIdx; // @[Reg.scala 17:22]
    end
    if (bc_mshr_io_tasks_source_a_valid) begin // @[Reg.scala 17:18]
      bc_bits_latch_size <= bc_mshr_io_tasks_source_a_bits_size; // @[Reg.scala 17:22]
    end
    if (bc_mshr_io_tasks_source_a_valid) begin // @[Reg.scala 17:18]
      bc_bits_latch_putData <= bc_mshr_io_tasks_source_a_bits_putData; // @[Reg.scala 17:22]
    end
    bc_valid_latch <= bc_mshr_io_tasks_source_a_valid; // @[Slice.scala 484:37]
    if (c_mshr_io_tasks_source_a_valid) begin // @[Reg.scala 17:18]
      c_bits_latch_tag <= c_mshr_io_tasks_source_a_bits_tag; // @[Reg.scala 17:22]
    end
    if (c_mshr_io_tasks_source_a_valid) begin // @[Reg.scala 17:18]
      c_bits_latch_set <= c_mshr_io_tasks_source_a_bits_set; // @[Reg.scala 17:22]
    end
    if (c_mshr_io_tasks_source_a_valid) begin // @[Reg.scala 17:18]
      c_bits_latch_off <= c_mshr_io_tasks_source_a_bits_off; // @[Reg.scala 17:22]
    end
    if (c_mshr_io_tasks_source_a_valid) begin // @[Reg.scala 17:18]
      c_bits_latch_opcode <= c_mshr_io_tasks_source_a_bits_opcode; // @[Reg.scala 17:22]
    end
    if (c_mshr_io_tasks_source_a_valid) begin // @[Reg.scala 17:18]
      c_bits_latch_param <= c_mshr_io_tasks_source_a_bits_param; // @[Reg.scala 17:22]
    end
    if (c_mshr_io_tasks_source_a_valid) begin // @[Reg.scala 17:18]
      c_bits_latch_source <= c_mshr_io_tasks_source_a_bits_source; // @[Reg.scala 17:22]
    end
    if (c_mshr_io_tasks_source_a_valid) begin // @[Reg.scala 17:18]
      c_bits_latch_bufIdx <= c_mshr_io_tasks_source_a_bits_bufIdx; // @[Reg.scala 17:22]
    end
    if (c_mshr_io_tasks_source_a_valid) begin // @[Reg.scala 17:18]
      c_bits_latch_size <= c_mshr_io_tasks_source_a_bits_size; // @[Reg.scala 17:22]
    end
    if (c_mshr_io_tasks_source_a_valid) begin // @[Reg.scala 17:18]
      c_bits_latch_putData <= c_mshr_io_tasks_source_a_bits_putData; // @[Reg.scala 17:22]
    end
    c_valid_latch <= c_mshr_io_tasks_source_a_valid; // @[Slice.scala 486:36]
    if (bc_mshr_io_tasks_source_bvalid) begin // @[Reg.scala 17:18]
      bc_bits_latch_1_set <= bc_mshr_io_tasks_source_bset; // @[Reg.scala 17:22]
    end
    if (bc_mshr_io_tasks_source_bvalid) begin // @[Reg.scala 17:18]
      bc_bits_latch_1_tag <= bc_mshr_io_tasks_source_btag; // @[Reg.scala 17:22]
    end
    if (bc_mshr_io_tasks_source_bvalid) begin // @[Reg.scala 17:18]
      bc_bits_latch_1_param <= bc_mshr_io_tasks_source_bparam; // @[Reg.scala 17:22]
    end
    if (bc_mshr_io_tasks_source_bvalid) begin // @[Reg.scala 17:18]
      bc_bits_latch_1_clients <= bc_mshr_io_tasks_source_bclients; // @[Reg.scala 17:22]
    end
    if (bc_mshr_io_tasks_source_bvalid) begin // @[Reg.scala 17:18]
      bc_bits_latch_1_needData <= bc_mshr_io_tasks_source_bneedData; // @[Reg.scala 17:22]
    end
    bc_valid_latch_1 <= bc_mshr_io_tasks_source_bvalid; // @[Slice.scala 484:37]
    if (c_mshr_io_tasks_source_bvalid) begin // @[Reg.scala 17:18]
      c_bits_latch_1_set <= c_mshr_io_tasks_source_bset; // @[Reg.scala 17:22]
    end
    if (c_mshr_io_tasks_source_bvalid) begin // @[Reg.scala 17:18]
      c_bits_latch_1_tag <= c_mshr_io_tasks_source_btag; // @[Reg.scala 17:22]
    end
    if (c_mshr_io_tasks_source_bvalid) begin // @[Reg.scala 17:18]
      c_bits_latch_1_param <= c_mshr_io_tasks_source_bparam; // @[Reg.scala 17:22]
    end
    if (c_mshr_io_tasks_source_bvalid) begin // @[Reg.scala 17:18]
      c_bits_latch_1_clients <= c_mshr_io_tasks_source_bclients; // @[Reg.scala 17:22]
    end
    if (c_mshr_io_tasks_source_bvalid) begin // @[Reg.scala 17:18]
      c_bits_latch_1_needData <= c_mshr_io_tasks_source_bneedData; // @[Reg.scala 17:22]
    end
    c_valid_latch_1 <= c_mshr_io_tasks_source_bvalid; // @[Slice.scala 486:36]
    if (bc_mshr_io_tasks_source_c_valid) begin // @[Reg.scala 17:18]
      bc_bits_latch_2_opcode <= bc_mshr_io_tasks_source_c_bits_opcode; // @[Reg.scala 17:22]
    end
    if (bc_mshr_io_tasks_source_c_valid) begin // @[Reg.scala 17:18]
      bc_bits_latch_2_tag <= bc_mshr_io_tasks_source_c_bits_tag; // @[Reg.scala 17:22]
    end
    if (bc_mshr_io_tasks_source_c_valid) begin // @[Reg.scala 17:18]
      bc_bits_latch_2_set <= bc_mshr_io_tasks_source_c_bits_set; // @[Reg.scala 17:22]
    end
    if (bc_mshr_io_tasks_source_c_valid) begin // @[Reg.scala 17:18]
      bc_bits_latch_2_source <= bc_mshr_io_tasks_source_c_bits_source; // @[Reg.scala 17:22]
    end
    if (bc_mshr_io_tasks_source_c_valid) begin // @[Reg.scala 17:18]
      bc_bits_latch_2_way <= bc_mshr_io_tasks_source_c_bits_way; // @[Reg.scala 17:22]
    end
    bc_valid_latch_2 <= bc_mshr_io_tasks_source_c_valid; // @[Slice.scala 484:37]
    if (c_mshr_io_tasks_source_c_valid) begin // @[Reg.scala 17:18]
      c_bits_latch_2_opcode <= c_mshr_io_tasks_source_c_bits_opcode; // @[Reg.scala 17:22]
    end
    if (c_mshr_io_tasks_source_c_valid) begin // @[Reg.scala 17:18]
      c_bits_latch_2_tag <= c_mshr_io_tasks_source_c_bits_tag; // @[Reg.scala 17:22]
    end
    if (c_mshr_io_tasks_source_c_valid) begin // @[Reg.scala 17:18]
      c_bits_latch_2_set <= c_mshr_io_tasks_source_c_bits_set; // @[Reg.scala 17:22]
    end
    if (c_mshr_io_tasks_source_c_valid) begin // @[Reg.scala 17:18]
      c_bits_latch_2_source <= c_mshr_io_tasks_source_c_bits_source; // @[Reg.scala 17:22]
    end
    if (c_mshr_io_tasks_source_c_valid) begin // @[Reg.scala 17:18]
      c_bits_latch_2_way <= c_mshr_io_tasks_source_c_bits_way; // @[Reg.scala 17:22]
    end
    c_valid_latch_2 <= c_mshr_io_tasks_source_c_valid; // @[Slice.scala 486:36]
    if (bc_mshr_io_tasks_source_d_valid) begin // @[Reg.scala 17:18]
      bc_bits_latch_3_sourceId <= bc_mshr_io_tasks_source_d_bits_sourceId; // @[Reg.scala 17:22]
    end
    if (bc_mshr_io_tasks_source_d_valid) begin // @[Reg.scala 17:18]
      bc_bits_latch_3_set <= bc_mshr_io_tasks_source_d_bits_set; // @[Reg.scala 17:22]
    end
    if (bc_mshr_io_tasks_source_d_valid) begin // @[Reg.scala 17:18]
      bc_bits_latch_3_channel <= bc_mshr_io_tasks_source_d_bits_channel; // @[Reg.scala 17:22]
    end
    if (bc_mshr_io_tasks_source_d_valid) begin // @[Reg.scala 17:18]
      bc_bits_latch_3_opcode <= bc_mshr_io_tasks_source_d_bits_opcode; // @[Reg.scala 17:22]
    end
    if (bc_mshr_io_tasks_source_d_valid) begin // @[Reg.scala 17:18]
      bc_bits_latch_3_param <= bc_mshr_io_tasks_source_d_bits_param; // @[Reg.scala 17:22]
    end
    if (bc_mshr_io_tasks_source_d_valid) begin // @[Reg.scala 17:18]
      bc_bits_latch_3_size <= bc_mshr_io_tasks_source_d_bits_size; // @[Reg.scala 17:22]
    end
    if (bc_mshr_io_tasks_source_d_valid) begin // @[Reg.scala 17:18]
      bc_bits_latch_3_way <= bc_mshr_io_tasks_source_d_bits_way; // @[Reg.scala 17:22]
    end
    if (bc_mshr_io_tasks_source_d_valid) begin // @[Reg.scala 17:18]
      bc_bits_latch_3_off <= bc_mshr_io_tasks_source_d_bits_off; // @[Reg.scala 17:22]
    end
    if (bc_mshr_io_tasks_source_d_valid) begin // @[Reg.scala 17:18]
      bc_bits_latch_3_useBypass <= bc_mshr_io_tasks_source_d_bits_useBypass; // @[Reg.scala 17:22]
    end
    if (bc_mshr_io_tasks_source_d_valid) begin // @[Reg.scala 17:18]
      bc_bits_latch_3_bufIdx <= bc_mshr_io_tasks_source_d_bits_bufIdx; // @[Reg.scala 17:22]
    end
    if (bc_mshr_io_tasks_source_d_valid) begin // @[Reg.scala 17:18]
      bc_bits_latch_3_denied <= bc_mshr_io_tasks_source_d_bits_denied; // @[Reg.scala 17:22]
    end
    if (bc_mshr_io_tasks_source_d_valid) begin // @[Reg.scala 17:18]
      bc_bits_latch_3_sinkId <= bc_mshr_io_tasks_source_d_bits_sinkId; // @[Reg.scala 17:22]
    end
    if (bc_mshr_io_tasks_source_d_valid) begin // @[Reg.scala 17:18]
      bc_bits_latch_3_bypassPut <= bc_mshr_io_tasks_source_d_bits_bypassPut; // @[Reg.scala 17:22]
    end
    if (bc_mshr_io_tasks_source_d_valid) begin // @[Reg.scala 17:18]
      bc_bits_latch_3_dirty <= bc_mshr_io_tasks_source_d_bits_dirty; // @[Reg.scala 17:22]
    end
    bc_valid_latch_3 <= bc_mshr_io_tasks_source_d_valid; // @[Slice.scala 484:37]
    if (c_mshr_io_tasks_source_d_valid) begin // @[Reg.scala 17:18]
      c_bits_latch_3_sourceId <= c_mshr_io_tasks_source_d_bits_sourceId; // @[Reg.scala 17:22]
    end
    if (c_mshr_io_tasks_source_d_valid) begin // @[Reg.scala 17:18]
      c_bits_latch_3_set <= c_mshr_io_tasks_source_d_bits_set; // @[Reg.scala 17:22]
    end
    if (c_mshr_io_tasks_source_d_valid) begin // @[Reg.scala 17:18]
      c_bits_latch_3_channel <= c_mshr_io_tasks_source_d_bits_channel; // @[Reg.scala 17:22]
    end
    if (c_mshr_io_tasks_source_d_valid) begin // @[Reg.scala 17:18]
      c_bits_latch_3_opcode <= c_mshr_io_tasks_source_d_bits_opcode; // @[Reg.scala 17:22]
    end
    if (c_mshr_io_tasks_source_d_valid) begin // @[Reg.scala 17:18]
      c_bits_latch_3_param <= c_mshr_io_tasks_source_d_bits_param; // @[Reg.scala 17:22]
    end
    if (c_mshr_io_tasks_source_d_valid) begin // @[Reg.scala 17:18]
      c_bits_latch_3_size <= c_mshr_io_tasks_source_d_bits_size; // @[Reg.scala 17:22]
    end
    if (c_mshr_io_tasks_source_d_valid) begin // @[Reg.scala 17:18]
      c_bits_latch_3_way <= c_mshr_io_tasks_source_d_bits_way; // @[Reg.scala 17:22]
    end
    if (c_mshr_io_tasks_source_d_valid) begin // @[Reg.scala 17:18]
      c_bits_latch_3_off <= c_mshr_io_tasks_source_d_bits_off; // @[Reg.scala 17:22]
    end
    if (c_mshr_io_tasks_source_d_valid) begin // @[Reg.scala 17:18]
      c_bits_latch_3_useBypass <= c_mshr_io_tasks_source_d_bits_useBypass; // @[Reg.scala 17:22]
    end
    if (c_mshr_io_tasks_source_d_valid) begin // @[Reg.scala 17:18]
      c_bits_latch_3_bufIdx <= c_mshr_io_tasks_source_d_bits_bufIdx; // @[Reg.scala 17:22]
    end
    if (c_mshr_io_tasks_source_d_valid) begin // @[Reg.scala 17:18]
      c_bits_latch_3_denied <= c_mshr_io_tasks_source_d_bits_denied; // @[Reg.scala 17:22]
    end
    if (c_mshr_io_tasks_source_d_valid) begin // @[Reg.scala 17:18]
      c_bits_latch_3_sinkId <= c_mshr_io_tasks_source_d_bits_sinkId; // @[Reg.scala 17:22]
    end
    if (c_mshr_io_tasks_source_d_valid) begin // @[Reg.scala 17:18]
      c_bits_latch_3_bypassPut <= c_mshr_io_tasks_source_d_bits_bypassPut; // @[Reg.scala 17:22]
    end
    if (c_mshr_io_tasks_source_d_valid) begin // @[Reg.scala 17:18]
      c_bits_latch_3_dirty <= c_mshr_io_tasks_source_d_bits_dirty; // @[Reg.scala 17:22]
    end
    c_valid_latch_3 <= c_mshr_io_tasks_source_d_valid; // @[Slice.scala 486:36]
    if (bc_mshr_io_tasks_source_e_valid) begin // @[Reg.scala 17:18]
      bc_bits_latch_4_sink <= bc_mshr_io_tasks_source_e_bits_sink; // @[Reg.scala 17:22]
    end
    bc_valid_latch_4 <= bc_mshr_io_tasks_source_e_valid; // @[Slice.scala 484:37]
    if (c_mshr_io_tasks_source_e_valid) begin // @[Reg.scala 17:18]
      c_bits_latch_4_sink <= c_mshr_io_tasks_source_e_bits_sink; // @[Reg.scala 17:22]
    end
    c_valid_latch_4 <= c_mshr_io_tasks_source_e_valid; // @[Slice.scala 486:36]
    if (bc_mshr_io_tasks_sink_c_valid) begin // @[Reg.scala 17:18]
      bc_bits_latch_6_set <= bc_mshr_io_tasks_sink_c_bits_set; // @[Reg.scala 17:22]
    end
    if (bc_mshr_io_tasks_sink_c_valid) begin // @[Reg.scala 17:18]
      bc_bits_latch_6_tag <= bc_mshr_io_tasks_sink_c_bits_tag; // @[Reg.scala 17:22]
    end
    if (bc_mshr_io_tasks_sink_c_valid) begin // @[Reg.scala 17:18]
      bc_bits_latch_6_way <= bc_mshr_io_tasks_sink_c_bits_way; // @[Reg.scala 17:22]
    end
    if (bc_mshr_io_tasks_sink_c_valid) begin // @[Reg.scala 17:18]
      bc_bits_latch_6_bufIdx <= bc_mshr_io_tasks_sink_c_bits_bufIdx; // @[Reg.scala 17:22]
    end
    if (bc_mshr_io_tasks_sink_c_valid) begin // @[Reg.scala 17:18]
      bc_bits_latch_6_opcode <= bc_mshr_io_tasks_sink_c_bits_opcode; // @[Reg.scala 17:22]
    end
    if (bc_mshr_io_tasks_sink_c_valid) begin // @[Reg.scala 17:18]
      bc_bits_latch_6_source <= bc_mshr_io_tasks_sink_c_bits_source; // @[Reg.scala 17:22]
    end
    if (bc_mshr_io_tasks_sink_c_valid) begin // @[Reg.scala 17:18]
      bc_bits_latch_6_save <= bc_mshr_io_tasks_sink_c_bits_save; // @[Reg.scala 17:22]
    end
    if (bc_mshr_io_tasks_sink_c_valid) begin // @[Reg.scala 17:18]
      bc_bits_latch_6_drop <= bc_mshr_io_tasks_sink_c_bits_drop; // @[Reg.scala 17:22]
    end
    if (bc_mshr_io_tasks_sink_c_valid) begin // @[Reg.scala 17:18]
      bc_bits_latch_6_release <= bc_mshr_io_tasks_sink_c_bits_release; // @[Reg.scala 17:22]
    end
    bc_valid_latch_6 <= bc_mshr_io_tasks_sink_c_valid; // @[Slice.scala 484:37]
    if (c_mshr_io_tasks_sink_c_valid) begin // @[Reg.scala 17:18]
      c_bits_latch_6_set <= c_mshr_io_tasks_sink_c_bits_set; // @[Reg.scala 17:22]
    end
    if (c_mshr_io_tasks_sink_c_valid) begin // @[Reg.scala 17:18]
      c_bits_latch_6_tag <= c_mshr_io_tasks_sink_c_bits_tag; // @[Reg.scala 17:22]
    end
    if (c_mshr_io_tasks_sink_c_valid) begin // @[Reg.scala 17:18]
      c_bits_latch_6_way <= c_mshr_io_tasks_sink_c_bits_way; // @[Reg.scala 17:22]
    end
    if (c_mshr_io_tasks_sink_c_valid) begin // @[Reg.scala 17:18]
      c_bits_latch_6_bufIdx <= c_mshr_io_tasks_sink_c_bits_bufIdx; // @[Reg.scala 17:22]
    end
    if (c_mshr_io_tasks_sink_c_valid) begin // @[Reg.scala 17:18]
      c_bits_latch_6_opcode <= c_mshr_io_tasks_sink_c_bits_opcode; // @[Reg.scala 17:22]
    end
    if (c_mshr_io_tasks_sink_c_valid) begin // @[Reg.scala 17:18]
      c_bits_latch_6_source <= c_mshr_io_tasks_sink_c_bits_source; // @[Reg.scala 17:22]
    end
    if (c_mshr_io_tasks_sink_c_valid) begin // @[Reg.scala 17:18]
      c_bits_latch_6_save <= c_mshr_io_tasks_sink_c_bits_save; // @[Reg.scala 17:22]
    end
    if (c_mshr_io_tasks_sink_c_valid) begin // @[Reg.scala 17:18]
      c_bits_latch_6_drop <= c_mshr_io_tasks_sink_c_bits_drop; // @[Reg.scala 17:22]
    end
    if (c_mshr_io_tasks_sink_c_valid) begin // @[Reg.scala 17:18]
      c_bits_latch_6_release <= c_mshr_io_tasks_sink_c_bits_release; // @[Reg.scala 17:22]
    end
    c_valid_latch_6 <= c_mshr_io_tasks_sink_c_valid; // @[Slice.scala 486:36]
    if (bc_mshr_io_tasks_tag_write_valid) begin // @[Reg.scala 17:18]
      bc_bits_latch_7_set <= bc_mshr_io_tasks_tag_write_bits_set; // @[Reg.scala 17:22]
    end
    if (bc_mshr_io_tasks_tag_write_valid) begin // @[Reg.scala 17:18]
      bc_bits_latch_7_way <= bc_mshr_io_tasks_tag_write_bits_way; // @[Reg.scala 17:22]
    end
    if (bc_mshr_io_tasks_tag_write_valid) begin // @[Reg.scala 17:18]
      bc_bits_latch_7_tag <= bc_mshr_io_tasks_tag_write_bits_tag; // @[Reg.scala 17:22]
    end
    bc_valid_latch_7 <= bc_mshr_io_tasks_tag_write_valid; // @[Slice.scala 484:37]
    if (c_mshr_io_tasks_tag_write_valid) begin // @[Reg.scala 17:18]
      c_bits_latch_7_set <= c_mshr_io_tasks_tag_write_bits_set; // @[Reg.scala 17:22]
    end
    if (c_mshr_io_tasks_tag_write_valid) begin // @[Reg.scala 17:18]
      c_bits_latch_7_way <= c_mshr_io_tasks_tag_write_bits_way; // @[Reg.scala 17:22]
    end
    if (c_mshr_io_tasks_tag_write_valid) begin // @[Reg.scala 17:18]
      c_bits_latch_7_tag <= c_mshr_io_tasks_tag_write_bits_tag; // @[Reg.scala 17:22]
    end
    c_valid_latch_7 <= c_mshr_io_tasks_tag_write_valid; // @[Slice.scala 486:36]
    if (bc_mshr_io_tasks_client_tag_write_valid) begin // @[Reg.scala 17:18]
      bc_bits_latch_8_set <= bc_mshr_io_tasks_client_tag_write_bits_set; // @[Reg.scala 17:22]
    end
    if (bc_mshr_io_tasks_client_tag_write_valid) begin // @[Reg.scala 17:18]
      bc_bits_latch_8_way <= bc_mshr_io_tasks_client_tag_write_bits_way; // @[Reg.scala 17:22]
    end
    if (bc_mshr_io_tasks_client_tag_write_valid) begin // @[Reg.scala 17:18]
      bc_bits_latch_8_tag <= bc_mshr_io_tasks_client_tag_write_bits_tag; // @[Reg.scala 17:22]
    end
    bc_valid_latch_8 <= bc_mshr_io_tasks_client_tag_write_valid; // @[Slice.scala 484:37]
    if (c_mshr_io_tasks_client_tag_write_valid) begin // @[Reg.scala 17:18]
      c_bits_latch_8_set <= c_mshr_io_tasks_client_tag_write_bits_set; // @[Reg.scala 17:22]
    end
    if (c_mshr_io_tasks_client_tag_write_valid) begin // @[Reg.scala 17:18]
      c_bits_latch_8_way <= c_mshr_io_tasks_client_tag_write_bits_way; // @[Reg.scala 17:22]
    end
    if (c_mshr_io_tasks_client_tag_write_valid) begin // @[Reg.scala 17:18]
      c_bits_latch_8_tag <= c_mshr_io_tasks_client_tag_write_bits_tag; // @[Reg.scala 17:22]
    end
    c_valid_latch_8 <= c_mshr_io_tasks_client_tag_write_valid; // @[Slice.scala 486:36]
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Arbiter.scala 113:23]
      beatsLeft <= 1'h0;
    end else if (latch) begin
      beatsLeft <= initBeats;
    end else begin
      beatsLeft <= beatsLeft - _beatsLeft_T_2;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Arbiter.scala 118:30]
      state_0 <= 1'h0;
    end else if (idle) begin
      state_0 <= earlyWinner_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Arbiter.scala 118:30]
      state_1 <= 1'h0;
    end else if (idle) begin
      state_1 <= earlyWinner_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Slice.scala 188:36]
      bc_mask_latch_0 <= 1'h0; // @[Slice.scala 189:19]
    end else if (mshrAlloc_io_bc_mask_valid) begin // @[Slice.scala 186:30]
      bc_mask_latch_0 <= mshrAlloc_io_bc_mask_bits_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Slice.scala 188:36]
      bc_mask_latch_1 <= 1'h0; // @[Slice.scala 189:19]
    end else if (mshrAlloc_io_bc_mask_valid) begin // @[Slice.scala 186:30]
      bc_mask_latch_1 <= mshrAlloc_io_bc_mask_bits_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Slice.scala 188:36]
      bc_mask_latch_2 <= 1'h0; // @[Slice.scala 189:19]
    end else if (mshrAlloc_io_bc_mask_valid) begin // @[Slice.scala 186:30]
      bc_mask_latch_2 <= mshrAlloc_io_bc_mask_bits_2;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Slice.scala 188:36]
      bc_mask_latch_3 <= 1'h0; // @[Slice.scala 189:19]
    end else if (mshrAlloc_io_bc_mask_valid) begin // @[Slice.scala 186:30]
      bc_mask_latch_3 <= mshrAlloc_io_bc_mask_bits_3;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Slice.scala 188:36]
      bc_mask_latch_4 <= 1'h0; // @[Slice.scala 189:19]
    end else if (mshrAlloc_io_bc_mask_valid) begin // @[Slice.scala 186:30]
      bc_mask_latch_4 <= mshrAlloc_io_bc_mask_bits_4;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Slice.scala 188:36]
      bc_mask_latch_5 <= 1'h0; // @[Slice.scala 189:19]
    end else if (mshrAlloc_io_bc_mask_valid) begin // @[Slice.scala 186:30]
      bc_mask_latch_5 <= mshrAlloc_io_bc_mask_bits_5;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Slice.scala 188:36]
      bc_mask_latch_6 <= 1'h0; // @[Slice.scala 189:19]
    end else if (mshrAlloc_io_bc_mask_valid) begin // @[Slice.scala 186:30]
      bc_mask_latch_6 <= mshrAlloc_io_bc_mask_bits_6;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Slice.scala 188:36]
      bc_mask_latch_7 <= 1'h0; // @[Slice.scala 189:19]
    end else if (mshrAlloc_io_bc_mask_valid) begin // @[Slice.scala 186:30]
      bc_mask_latch_7 <= mshrAlloc_io_bc_mask_bits_7;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Slice.scala 188:36]
      bc_mask_latch_8 <= 1'h0; // @[Slice.scala 189:19]
    end else if (mshrAlloc_io_bc_mask_valid) begin // @[Slice.scala 186:30]
      bc_mask_latch_8 <= mshrAlloc_io_bc_mask_bits_8;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Slice.scala 188:36]
      bc_mask_latch_9 <= 1'h0; // @[Slice.scala 189:19]
    end else if (mshrAlloc_io_bc_mask_valid) begin // @[Slice.scala 186:30]
      bc_mask_latch_9 <= mshrAlloc_io_bc_mask_bits_9;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Slice.scala 188:36]
      bc_mask_latch_10 <= 1'h0; // @[Slice.scala 189:19]
    end else if (mshrAlloc_io_bc_mask_valid) begin // @[Slice.scala 186:30]
      bc_mask_latch_10 <= mshrAlloc_io_bc_mask_bits_10;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Slice.scala 188:36]
      bc_mask_latch_11 <= 1'h0; // @[Slice.scala 189:19]
    end else if (mshrAlloc_io_bc_mask_valid) begin // @[Slice.scala 186:30]
      bc_mask_latch_11 <= mshrAlloc_io_bc_mask_bits_11;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Slice.scala 188:36]
      bc_mask_latch_12 <= 1'h0; // @[Slice.scala 189:19]
    end else if (mshrAlloc_io_bc_mask_valid) begin // @[Slice.scala 186:30]
      bc_mask_latch_12 <= mshrAlloc_io_bc_mask_bits_12;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Slice.scala 188:36]
      bc_mask_latch_13 <= 1'h0; // @[Slice.scala 189:19]
    end else if (mshrAlloc_io_bc_mask_valid) begin // @[Slice.scala 186:30]
      bc_mask_latch_13 <= mshrAlloc_io_bc_mask_bits_13;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Slice.scala 191:35]
      c_mask_latch_0 <= 1'h0; // @[Slice.scala 192:18]
    end else if (mshrAlloc_io_c_mask_valid) begin // @[Slice.scala 187:29]
      c_mask_latch_0 <= mshrAlloc_io_c_mask_bits_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Slice.scala 191:35]
      c_mask_latch_1 <= 1'h0; // @[Slice.scala 192:18]
    end else if (mshrAlloc_io_c_mask_valid) begin // @[Slice.scala 187:29]
      c_mask_latch_1 <= mshrAlloc_io_c_mask_bits_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Slice.scala 191:35]
      c_mask_latch_2 <= 1'h0; // @[Slice.scala 192:18]
    end else if (mshrAlloc_io_c_mask_valid) begin // @[Slice.scala 187:29]
      c_mask_latch_2 <= mshrAlloc_io_c_mask_bits_2;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Slice.scala 191:35]
      c_mask_latch_3 <= 1'h0; // @[Slice.scala 192:18]
    end else if (mshrAlloc_io_c_mask_valid) begin // @[Slice.scala 187:29]
      c_mask_latch_3 <= mshrAlloc_io_c_mask_bits_3;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Slice.scala 191:35]
      c_mask_latch_4 <= 1'h0; // @[Slice.scala 192:18]
    end else if (mshrAlloc_io_c_mask_valid) begin // @[Slice.scala 187:29]
      c_mask_latch_4 <= mshrAlloc_io_c_mask_bits_4;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Slice.scala 191:35]
      c_mask_latch_5 <= 1'h0; // @[Slice.scala 192:18]
    end else if (mshrAlloc_io_c_mask_valid) begin // @[Slice.scala 187:29]
      c_mask_latch_5 <= mshrAlloc_io_c_mask_bits_5;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Slice.scala 191:35]
      c_mask_latch_6 <= 1'h0; // @[Slice.scala 192:18]
    end else if (mshrAlloc_io_c_mask_valid) begin // @[Slice.scala 187:29]
      c_mask_latch_6 <= mshrAlloc_io_c_mask_bits_6;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Slice.scala 191:35]
      c_mask_latch_7 <= 1'h0; // @[Slice.scala 192:18]
    end else if (mshrAlloc_io_c_mask_valid) begin // @[Slice.scala 187:29]
      c_mask_latch_7 <= mshrAlloc_io_c_mask_bits_7;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Slice.scala 191:35]
      c_mask_latch_8 <= 1'h0; // @[Slice.scala 192:18]
    end else if (mshrAlloc_io_c_mask_valid) begin // @[Slice.scala 187:29]
      c_mask_latch_8 <= mshrAlloc_io_c_mask_bits_8;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Slice.scala 191:35]
      c_mask_latch_9 <= 1'h0; // @[Slice.scala 192:18]
    end else if (mshrAlloc_io_c_mask_valid) begin // @[Slice.scala 187:29]
      c_mask_latch_9 <= mshrAlloc_io_c_mask_bits_9;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Slice.scala 191:35]
      c_mask_latch_10 <= 1'h0; // @[Slice.scala 192:18]
    end else if (mshrAlloc_io_c_mask_valid) begin // @[Slice.scala 187:29]
      c_mask_latch_10 <= mshrAlloc_io_c_mask_bits_10;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Slice.scala 191:35]
      c_mask_latch_11 <= 1'h0; // @[Slice.scala 192:18]
    end else if (mshrAlloc_io_c_mask_valid) begin // @[Slice.scala 187:29]
      c_mask_latch_11 <= mshrAlloc_io_c_mask_bits_11;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Slice.scala 191:35]
      c_mask_latch_12 <= 1'h0; // @[Slice.scala 192:18]
    end else if (mshrAlloc_io_c_mask_valid) begin // @[Slice.scala 187:29]
      c_mask_latch_12 <= mshrAlloc_io_c_mask_bits_12;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Slice.scala 191:35]
      c_mask_latch_13 <= 1'h0; // @[Slice.scala 192:18]
    end else if (mshrAlloc_io_c_mask_valid) begin // @[Slice.scala 187:29]
      c_mask_latch_13 <= mshrAlloc_io_c_mask_bits_13;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Slice.scala 191:35]
      c_mask_latch_14 <= 1'h0; // @[Slice.scala 192:18]
    end else if (mshrAlloc_io_c_mask_valid) begin // @[Slice.scala 187:29]
      c_mask_latch_14 <= mshrAlloc_io_c_mask_bits_14;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Slice.scala 554:74]
      ms_0_io_dirResult_valid_REG <= 1'h0;
    end else begin
      ms_0_io_dirResult_valid_REG <= ~is_ctrl_dir_res & directory_io_result_valid & directory_io_result_bits_idOH[0];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Slice.scala 554:74]
      ms_1_io_dirResult_valid_REG <= 1'h0;
    end else begin
      ms_1_io_dirResult_valid_REG <= ~is_ctrl_dir_res & directory_io_result_valid & directory_io_result_bits_idOH[1];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Slice.scala 554:74]
      ms_2_io_dirResult_valid_REG <= 1'h0;
    end else begin
      ms_2_io_dirResult_valid_REG <= ~is_ctrl_dir_res & directory_io_result_valid & directory_io_result_bits_idOH[2];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Slice.scala 554:74]
      ms_3_io_dirResult_valid_REG <= 1'h0;
    end else begin
      ms_3_io_dirResult_valid_REG <= ~is_ctrl_dir_res & directory_io_result_valid & directory_io_result_bits_idOH[3];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Slice.scala 554:74]
      ms_4_io_dirResult_valid_REG <= 1'h0;
    end else begin
      ms_4_io_dirResult_valid_REG <= ~is_ctrl_dir_res & directory_io_result_valid & directory_io_result_bits_idOH[4];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Slice.scala 554:74]
      ms_5_io_dirResult_valid_REG <= 1'h0;
    end else begin
      ms_5_io_dirResult_valid_REG <= ~is_ctrl_dir_res & directory_io_result_valid & directory_io_result_bits_idOH[5];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Slice.scala 554:74]
      ms_6_io_dirResult_valid_REG <= 1'h0;
    end else begin
      ms_6_io_dirResult_valid_REG <= ~is_ctrl_dir_res & directory_io_result_valid & directory_io_result_bits_idOH[6];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Slice.scala 554:74]
      ms_7_io_dirResult_valid_REG <= 1'h0;
    end else begin
      ms_7_io_dirResult_valid_REG <= ~is_ctrl_dir_res & directory_io_result_valid & directory_io_result_bits_idOH[7];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Slice.scala 554:74]
      ms_8_io_dirResult_valid_REG <= 1'h0;
    end else begin
      ms_8_io_dirResult_valid_REG <= ~is_ctrl_dir_res & directory_io_result_valid & directory_io_result_bits_idOH[8];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Slice.scala 554:74]
      ms_9_io_dirResult_valid_REG <= 1'h0;
    end else begin
      ms_9_io_dirResult_valid_REG <= ~is_ctrl_dir_res & directory_io_result_valid & directory_io_result_bits_idOH[9];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Slice.scala 554:74]
      ms_10_io_dirResult_valid_REG <= 1'h0;
    end else begin
      ms_10_io_dirResult_valid_REG <= ~is_ctrl_dir_res & directory_io_result_valid & directory_io_result_bits_idOH[10];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Slice.scala 554:74]
      ms_11_io_dirResult_valid_REG <= 1'h0;
    end else begin
      ms_11_io_dirResult_valid_REG <= ~is_ctrl_dir_res & directory_io_result_valid & directory_io_result_bits_idOH[11];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Slice.scala 554:74]
      ms_12_io_dirResult_valid_REG <= 1'h0;
    end else begin
      ms_12_io_dirResult_valid_REG <= ~is_ctrl_dir_res & directory_io_result_valid & directory_io_result_bits_idOH[12];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Slice.scala 554:74]
      ms_13_io_dirResult_valid_REG <= 1'h0;
    end else begin
      ms_13_io_dirResult_valid_REG <= ~is_ctrl_dir_res & directory_io_result_valid & directory_io_result_bits_idOH[13];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Slice.scala 554:74]
      ms_14_io_dirResult_valid_REG <= 1'h0;
    end else begin
      ms_14_io_dirResult_valid_REG <= ~is_ctrl_dir_res & directory_io_result_valid & directory_io_result_bits_idOH[14];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Slice.scala 554:74]
      ms_15_io_dirResult_valid_REG <= 1'h0;
    end else begin
      ms_15_io_dirResult_valid_REG <= ~is_ctrl_dir_res & directory_io_result_valid & directory_io_result_bits_idOH[15];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Slice.scala 560:36]
      probeHelperOpt_io_dirResult_valid_REG <= 1'h0; // @[Slice.scala 560:36]
    end else begin
      probeHelperOpt_io_dirResult_valid_REG <= directory_io_result_valid; // @[Slice.scala 560:36]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  beatsLeft = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  state_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  state_1 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  bc_mask_latch_0 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  bc_mask_latch_1 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  bc_mask_latch_2 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  bc_mask_latch_3 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  bc_mask_latch_4 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  bc_mask_latch_5 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  bc_mask_latch_6 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  bc_mask_latch_7 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  bc_mask_latch_8 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  bc_mask_latch_9 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  bc_mask_latch_10 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  bc_mask_latch_11 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  bc_mask_latch_12 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  bc_mask_latch_13 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  c_mask_latch_0 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  c_mask_latch_1 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  c_mask_latch_2 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  c_mask_latch_3 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  c_mask_latch_4 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  c_mask_latch_5 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  c_mask_latch_6 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  c_mask_latch_7 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  c_mask_latch_8 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  c_mask_latch_9 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  c_mask_latch_10 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  c_mask_latch_11 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  c_mask_latch_12 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  c_mask_latch_13 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  c_mask_latch_14 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  bc_bits_latch_tag = _RAND_32[19:0];
  _RAND_33 = {1{`RANDOM}};
  bc_bits_latch_set = _RAND_33[9:0];
  _RAND_34 = {1{`RANDOM}};
  bc_bits_latch_off = _RAND_34[5:0];
  _RAND_35 = {1{`RANDOM}};
  bc_bits_latch_opcode = _RAND_35[2:0];
  _RAND_36 = {1{`RANDOM}};
  bc_bits_latch_param = _RAND_36[2:0];
  _RAND_37 = {1{`RANDOM}};
  bc_bits_latch_source = _RAND_37[3:0];
  _RAND_38 = {1{`RANDOM}};
  bc_bits_latch_bufIdx = _RAND_38[2:0];
  _RAND_39 = {1{`RANDOM}};
  bc_bits_latch_size = _RAND_39[2:0];
  _RAND_40 = {1{`RANDOM}};
  bc_bits_latch_putData = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  bc_valid_latch = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  c_bits_latch_tag = _RAND_42[19:0];
  _RAND_43 = {1{`RANDOM}};
  c_bits_latch_set = _RAND_43[9:0];
  _RAND_44 = {1{`RANDOM}};
  c_bits_latch_off = _RAND_44[5:0];
  _RAND_45 = {1{`RANDOM}};
  c_bits_latch_opcode = _RAND_45[2:0];
  _RAND_46 = {1{`RANDOM}};
  c_bits_latch_param = _RAND_46[2:0];
  _RAND_47 = {1{`RANDOM}};
  c_bits_latch_source = _RAND_47[3:0];
  _RAND_48 = {1{`RANDOM}};
  c_bits_latch_bufIdx = _RAND_48[2:0];
  _RAND_49 = {1{`RANDOM}};
  c_bits_latch_size = _RAND_49[2:0];
  _RAND_50 = {1{`RANDOM}};
  c_bits_latch_putData = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  c_valid_latch = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  bc_bits_latch_1_set = _RAND_52[9:0];
  _RAND_53 = {1{`RANDOM}};
  bc_bits_latch_1_tag = _RAND_53[19:0];
  _RAND_54 = {1{`RANDOM}};
  bc_bits_latch_1_param = _RAND_54[2:0];
  _RAND_55 = {1{`RANDOM}};
  bc_bits_latch_1_clients = _RAND_55[1:0];
  _RAND_56 = {1{`RANDOM}};
  bc_bits_latch_1_needData = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  bc_valid_latch_1 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  c_bits_latch_1_set = _RAND_58[9:0];
  _RAND_59 = {1{`RANDOM}};
  c_bits_latch_1_tag = _RAND_59[19:0];
  _RAND_60 = {1{`RANDOM}};
  c_bits_latch_1_param = _RAND_60[2:0];
  _RAND_61 = {1{`RANDOM}};
  c_bits_latch_1_clients = _RAND_61[1:0];
  _RAND_62 = {1{`RANDOM}};
  c_bits_latch_1_needData = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  c_valid_latch_1 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  bc_bits_latch_2_opcode = _RAND_64[2:0];
  _RAND_65 = {1{`RANDOM}};
  bc_bits_latch_2_tag = _RAND_65[19:0];
  _RAND_66 = {1{`RANDOM}};
  bc_bits_latch_2_set = _RAND_66[9:0];
  _RAND_67 = {1{`RANDOM}};
  bc_bits_latch_2_source = _RAND_67[3:0];
  _RAND_68 = {1{`RANDOM}};
  bc_bits_latch_2_way = _RAND_68[2:0];
  _RAND_69 = {1{`RANDOM}};
  bc_valid_latch_2 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  c_bits_latch_2_opcode = _RAND_70[2:0];
  _RAND_71 = {1{`RANDOM}};
  c_bits_latch_2_tag = _RAND_71[19:0];
  _RAND_72 = {1{`RANDOM}};
  c_bits_latch_2_set = _RAND_72[9:0];
  _RAND_73 = {1{`RANDOM}};
  c_bits_latch_2_source = _RAND_73[3:0];
  _RAND_74 = {1{`RANDOM}};
  c_bits_latch_2_way = _RAND_74[2:0];
  _RAND_75 = {1{`RANDOM}};
  c_valid_latch_2 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  bc_bits_latch_3_sourceId = _RAND_76[5:0];
  _RAND_77 = {1{`RANDOM}};
  bc_bits_latch_3_set = _RAND_77[9:0];
  _RAND_78 = {1{`RANDOM}};
  bc_bits_latch_3_channel = _RAND_78[2:0];
  _RAND_79 = {1{`RANDOM}};
  bc_bits_latch_3_opcode = _RAND_79[2:0];
  _RAND_80 = {1{`RANDOM}};
  bc_bits_latch_3_param = _RAND_80[2:0];
  _RAND_81 = {1{`RANDOM}};
  bc_bits_latch_3_size = _RAND_81[2:0];
  _RAND_82 = {1{`RANDOM}};
  bc_bits_latch_3_way = _RAND_82[2:0];
  _RAND_83 = {1{`RANDOM}};
  bc_bits_latch_3_off = _RAND_83[5:0];
  _RAND_84 = {1{`RANDOM}};
  bc_bits_latch_3_useBypass = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  bc_bits_latch_3_bufIdx = _RAND_85[2:0];
  _RAND_86 = {1{`RANDOM}};
  bc_bits_latch_3_denied = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  bc_bits_latch_3_sinkId = _RAND_87[3:0];
  _RAND_88 = {1{`RANDOM}};
  bc_bits_latch_3_bypassPut = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  bc_bits_latch_3_dirty = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  bc_valid_latch_3 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  c_bits_latch_3_sourceId = _RAND_91[5:0];
  _RAND_92 = {1{`RANDOM}};
  c_bits_latch_3_set = _RAND_92[9:0];
  _RAND_93 = {1{`RANDOM}};
  c_bits_latch_3_channel = _RAND_93[2:0];
  _RAND_94 = {1{`RANDOM}};
  c_bits_latch_3_opcode = _RAND_94[2:0];
  _RAND_95 = {1{`RANDOM}};
  c_bits_latch_3_param = _RAND_95[2:0];
  _RAND_96 = {1{`RANDOM}};
  c_bits_latch_3_size = _RAND_96[2:0];
  _RAND_97 = {1{`RANDOM}};
  c_bits_latch_3_way = _RAND_97[2:0];
  _RAND_98 = {1{`RANDOM}};
  c_bits_latch_3_off = _RAND_98[5:0];
  _RAND_99 = {1{`RANDOM}};
  c_bits_latch_3_useBypass = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  c_bits_latch_3_bufIdx = _RAND_100[2:0];
  _RAND_101 = {1{`RANDOM}};
  c_bits_latch_3_denied = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  c_bits_latch_3_sinkId = _RAND_102[3:0];
  _RAND_103 = {1{`RANDOM}};
  c_bits_latch_3_bypassPut = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  c_bits_latch_3_dirty = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  c_valid_latch_3 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  bc_bits_latch_4_sink = _RAND_106[2:0];
  _RAND_107 = {1{`RANDOM}};
  bc_valid_latch_4 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  c_bits_latch_4_sink = _RAND_108[2:0];
  _RAND_109 = {1{`RANDOM}};
  c_valid_latch_4 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  bc_bits_latch_6_set = _RAND_110[9:0];
  _RAND_111 = {1{`RANDOM}};
  bc_bits_latch_6_tag = _RAND_111[19:0];
  _RAND_112 = {1{`RANDOM}};
  bc_bits_latch_6_way = _RAND_112[2:0];
  _RAND_113 = {1{`RANDOM}};
  bc_bits_latch_6_bufIdx = _RAND_113[2:0];
  _RAND_114 = {1{`RANDOM}};
  bc_bits_latch_6_opcode = _RAND_114[2:0];
  _RAND_115 = {1{`RANDOM}};
  bc_bits_latch_6_source = _RAND_115[3:0];
  _RAND_116 = {1{`RANDOM}};
  bc_bits_latch_6_save = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  bc_bits_latch_6_drop = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  bc_bits_latch_6_release = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  bc_valid_latch_6 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  c_bits_latch_6_set = _RAND_120[9:0];
  _RAND_121 = {1{`RANDOM}};
  c_bits_latch_6_tag = _RAND_121[19:0];
  _RAND_122 = {1{`RANDOM}};
  c_bits_latch_6_way = _RAND_122[2:0];
  _RAND_123 = {1{`RANDOM}};
  c_bits_latch_6_bufIdx = _RAND_123[2:0];
  _RAND_124 = {1{`RANDOM}};
  c_bits_latch_6_opcode = _RAND_124[2:0];
  _RAND_125 = {1{`RANDOM}};
  c_bits_latch_6_source = _RAND_125[3:0];
  _RAND_126 = {1{`RANDOM}};
  c_bits_latch_6_save = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  c_bits_latch_6_drop = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  c_bits_latch_6_release = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  c_valid_latch_6 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  bc_bits_latch_7_set = _RAND_130[9:0];
  _RAND_131 = {1{`RANDOM}};
  bc_bits_latch_7_way = _RAND_131[2:0];
  _RAND_132 = {1{`RANDOM}};
  bc_bits_latch_7_tag = _RAND_132[19:0];
  _RAND_133 = {1{`RANDOM}};
  bc_valid_latch_7 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  c_bits_latch_7_set = _RAND_134[9:0];
  _RAND_135 = {1{`RANDOM}};
  c_bits_latch_7_way = _RAND_135[2:0];
  _RAND_136 = {1{`RANDOM}};
  c_bits_latch_7_tag = _RAND_136[19:0];
  _RAND_137 = {1{`RANDOM}};
  c_valid_latch_7 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  bc_bits_latch_8_set = _RAND_138[6:0];
  _RAND_139 = {1{`RANDOM}};
  bc_bits_latch_8_way = _RAND_139[3:0];
  _RAND_140 = {1{`RANDOM}};
  bc_bits_latch_8_tag = _RAND_140[22:0];
  _RAND_141 = {1{`RANDOM}};
  bc_valid_latch_8 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  c_bits_latch_8_set = _RAND_142[6:0];
  _RAND_143 = {1{`RANDOM}};
  c_bits_latch_8_way = _RAND_143[3:0];
  _RAND_144 = {1{`RANDOM}};
  c_bits_latch_8_tag = _RAND_144[22:0];
  _RAND_145 = {1{`RANDOM}};
  c_valid_latch_8 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  ms_0_io_dirResult_valid_REG = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  ms_1_io_dirResult_valid_REG = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  ms_2_io_dirResult_valid_REG = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  ms_3_io_dirResult_valid_REG = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  ms_4_io_dirResult_valid_REG = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  ms_5_io_dirResult_valid_REG = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  ms_6_io_dirResult_valid_REG = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  ms_7_io_dirResult_valid_REG = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  ms_8_io_dirResult_valid_REG = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  ms_9_io_dirResult_valid_REG = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  ms_10_io_dirResult_valid_REG = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  ms_11_io_dirResult_valid_REG = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  ms_12_io_dirResult_valid_REG = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  ms_13_io_dirResult_valid_REG = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  ms_14_io_dirResult_valid_REG = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  ms_15_io_dirResult_valid_REG = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  probeHelperOpt_io_dirResult_valid_REG = _RAND_162[0:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    beatsLeft = 1'h0;
  end
  if (reset) begin
    state_0 = 1'h0;
  end
  if (reset) begin
    state_1 = 1'h0;
  end
  if (reset) begin
    bc_mask_latch_0 = 1'h0;
  end
  if (reset) begin
    bc_mask_latch_1 = 1'h0;
  end
  if (reset) begin
    bc_mask_latch_2 = 1'h0;
  end
  if (reset) begin
    bc_mask_latch_3 = 1'h0;
  end
  if (reset) begin
    bc_mask_latch_4 = 1'h0;
  end
  if (reset) begin
    bc_mask_latch_5 = 1'h0;
  end
  if (reset) begin
    bc_mask_latch_6 = 1'h0;
  end
  if (reset) begin
    bc_mask_latch_7 = 1'h0;
  end
  if (reset) begin
    bc_mask_latch_8 = 1'h0;
  end
  if (reset) begin
    bc_mask_latch_9 = 1'h0;
  end
  if (reset) begin
    bc_mask_latch_10 = 1'h0;
  end
  if (reset) begin
    bc_mask_latch_11 = 1'h0;
  end
  if (reset) begin
    bc_mask_latch_12 = 1'h0;
  end
  if (reset) begin
    bc_mask_latch_13 = 1'h0;
  end
  if (reset) begin
    c_mask_latch_0 = 1'h0;
  end
  if (reset) begin
    c_mask_latch_1 = 1'h0;
  end
  if (reset) begin
    c_mask_latch_2 = 1'h0;
  end
  if (reset) begin
    c_mask_latch_3 = 1'h0;
  end
  if (reset) begin
    c_mask_latch_4 = 1'h0;
  end
  if (reset) begin
    c_mask_latch_5 = 1'h0;
  end
  if (reset) begin
    c_mask_latch_6 = 1'h0;
  end
  if (reset) begin
    c_mask_latch_7 = 1'h0;
  end
  if (reset) begin
    c_mask_latch_8 = 1'h0;
  end
  if (reset) begin
    c_mask_latch_9 = 1'h0;
  end
  if (reset) begin
    c_mask_latch_10 = 1'h0;
  end
  if (reset) begin
    c_mask_latch_11 = 1'h0;
  end
  if (reset) begin
    c_mask_latch_12 = 1'h0;
  end
  if (reset) begin
    c_mask_latch_13 = 1'h0;
  end
  if (reset) begin
    c_mask_latch_14 = 1'h0;
  end
  if (reset) begin
    ms_0_io_dirResult_valid_REG = 1'h0;
  end
  if (reset) begin
    ms_1_io_dirResult_valid_REG = 1'h0;
  end
  if (reset) begin
    ms_2_io_dirResult_valid_REG = 1'h0;
  end
  if (reset) begin
    ms_3_io_dirResult_valid_REG = 1'h0;
  end
  if (reset) begin
    ms_4_io_dirResult_valid_REG = 1'h0;
  end
  if (reset) begin
    ms_5_io_dirResult_valid_REG = 1'h0;
  end
  if (reset) begin
    ms_6_io_dirResult_valid_REG = 1'h0;
  end
  if (reset) begin
    ms_7_io_dirResult_valid_REG = 1'h0;
  end
  if (reset) begin
    ms_8_io_dirResult_valid_REG = 1'h0;
  end
  if (reset) begin
    ms_9_io_dirResult_valid_REG = 1'h0;
  end
  if (reset) begin
    ms_10_io_dirResult_valid_REG = 1'h0;
  end
  if (reset) begin
    ms_11_io_dirResult_valid_REG = 1'h0;
  end
  if (reset) begin
    ms_12_io_dirResult_valid_REG = 1'h0;
  end
  if (reset) begin
    ms_13_io_dirResult_valid_REG = 1'h0;
  end
  if (reset) begin
    ms_14_io_dirResult_valid_REG = 1'h0;
  end
  if (reset) begin
    ms_15_io_dirResult_valid_REG = 1'h0;
  end
  if (reset) begin
    probeHelperOpt_io_dirResult_valid_REG = 1'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule

