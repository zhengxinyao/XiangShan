module RVCExpander(
  input  [31:0] io_in,
  output [31:0] io_out_bits
);
  wire [6:0] io_out_s_opc = |io_in[12:5] ? 7'h13 : 7'h1f; // @[RVC.scala 53:20]
  wire [29:0] _io_out_s_T_7 = {io_in[10:7],io_in[12:11],io_in[5],io_in[6],2'h0,5'h2,3'h0,2'h1,io_in[4:2],io_out_s_opc}; // @[Cat.scala 31:58]
  wire [7:0] _io_out_s_T_15 = {io_in[6:5],io_in[12:10],3'h0}; // @[Cat.scala 31:58]
  wire [27:0] _io_out_s_T_20 = {io_in[6:5],io_in[12:10],3'h0,2'h1,io_in[9:7],3'h3,2'h1,io_in[4:2],7'h7}; // @[Cat.scala 31:58]
  wire [6:0] _io_out_s_T_31 = {io_in[5],io_in[12:10],io_in[6],2'h0}; // @[Cat.scala 31:58]
  wire [26:0] _io_out_s_T_36 = {io_in[5],io_in[12:10],io_in[6],2'h0,2'h1,io_in[9:7],3'h2,2'h1,io_in[4:2],7'h3}; // @[Cat.scala 31:58]
  wire [27:0] _io_out_s_T_51 = {io_in[6:5],io_in[12:10],3'h0,2'h1,io_in[9:7],3'h3,2'h1,io_in[4:2],7'h3}; // @[Cat.scala 31:58]
  wire [26:0] _io_out_s_T_73 = {_io_out_s_T_31[6:5],2'h1,io_in[4:2],2'h1,io_in[9:7],3'h2,_io_out_s_T_31[4:0],7'h3f}; // @[Cat.scala 31:58]
  wire [27:0] _io_out_s_T_93 = {_io_out_s_T_15[7:5],2'h1,io_in[4:2],2'h1,io_in[9:7],3'h3,_io_out_s_T_15[4:0],7'h27}; // @[Cat.scala 31:58]
  wire [26:0] _io_out_s_T_115 = {_io_out_s_T_31[6:5],2'h1,io_in[4:2],2'h1,io_in[9:7],3'h2,_io_out_s_T_31[4:0],7'h23}; // @[Cat.scala 31:58]
  wire [27:0] _io_out_s_T_135 = {_io_out_s_T_15[7:5],2'h1,io_in[4:2],2'h1,io_in[9:7],3'h3,_io_out_s_T_15[4:0],7'h23}; // @[Cat.scala 31:58]
  wire [6:0] _io_out_s_T_145 = io_in[12] ? 7'h7f : 7'h0; // @[Bitwise.scala 74:12]
  wire [11:0] _io_out_s_T_147 = {_io_out_s_T_145,io_in[6:2]}; // @[Cat.scala 31:58]
  wire [31:0] io_out_s_8_bits = {_io_out_s_T_145,io_in[6:2],io_in[11:7],3'h0,io_in[11:7],7'h13}; // @[Cat.scala 31:58]
  wire  _io_out_s_opc_T_3 = |io_in[11:7]; // @[RVC.scala 77:24]
  wire [6:0] io_out_s_opc_1 = |io_in[11:7] ? 7'h1b : 7'h1f; // @[RVC.scala 77:20]
  wire [31:0] io_out_s_9_bits = {_io_out_s_T_145,io_in[6:2],io_in[11:7],3'h0,io_in[11:7],io_out_s_opc_1}; // @[Cat.scala 31:58]
  wire [31:0] io_out_s_10_bits = {_io_out_s_T_145,io_in[6:2],5'h0,3'h0,io_in[11:7],7'h13}; // @[Cat.scala 31:58]
  wire  _io_out_s_opc_T_9 = |_io_out_s_T_147; // @[RVC.scala 90:29]
  wire [6:0] io_out_s_opc_2 = |_io_out_s_T_147 ? 7'h37 : 7'h3f; // @[RVC.scala 90:20]
  wire [14:0] _io_out_s_me_T_2 = io_in[12] ? 15'h7fff : 15'h0; // @[Bitwise.scala 74:12]
  wire [31:0] _io_out_s_me_T_4 = {_io_out_s_me_T_2,io_in[6:2],12'h0}; // @[Cat.scala 31:58]
  wire [31:0] io_out_s_me_bits = {_io_out_s_me_T_4[31:12],io_in[11:7],io_out_s_opc_2}; // @[Cat.scala 31:58]
  wire [6:0] io_out_s_opc_3 = _io_out_s_opc_T_9 ? 7'h13 : 7'h1f; // @[RVC.scala 86:20]
  wire [2:0] _io_out_s_T_187 = io_in[12] ? 3'h7 : 3'h0; // @[Bitwise.scala 74:12]
  wire [31:0] io_out_s_res_bits = {_io_out_s_T_187,io_in[4:3],io_in[5],io_in[2],io_in[6],4'h0,io_in[11:7],3'h0,io_in[11:
    7],io_out_s_opc_3}; // @[Cat.scala 31:58]
  wire [31:0] io_out_s_11_bits = io_in[11:7] == 5'h0 | io_in[11:7] == 5'h2 ? io_out_s_res_bits : io_out_s_me_bits; // @[RVC.scala 92:10]
  wire [25:0] _io_out_s_T_208 = {io_in[12],io_in[6:2],2'h1,io_in[9:7],3'h5,2'h1,io_in[9:7],7'h13}; // @[Cat.scala 31:58]
  wire [30:0] _GEN_0 = {{5'd0}, _io_out_s_T_208}; // @[RVC.scala 99:23]
  wire [30:0] _io_out_s_T_217 = _GEN_0 | 31'h40000000; // @[RVC.scala 99:23]
  wire [31:0] _io_out_s_T_227 = {_io_out_s_T_145,io_in[6:2],2'h1,io_in[9:7],3'h7,2'h1,io_in[9:7],7'h13}; // @[Cat.scala 31:58]
  wire [2:0] _io_out_s_funct_T_2 = {io_in[12],io_in[6:5]}; // @[Cat.scala 31:58]
  wire [2:0] _io_out_s_funct_T_4 = _io_out_s_funct_T_2 == 3'h1 ? 3'h4 : 3'h0; // @[package.scala 32:76]
  wire [2:0] _io_out_s_funct_T_6 = _io_out_s_funct_T_2 == 3'h2 ? 3'h6 : _io_out_s_funct_T_4; // @[package.scala 32:76]
  wire [2:0] _io_out_s_funct_T_8 = _io_out_s_funct_T_2 == 3'h3 ? 3'h7 : _io_out_s_funct_T_6; // @[package.scala 32:76]
  wire [2:0] _io_out_s_funct_T_10 = _io_out_s_funct_T_2 == 3'h4 ? 3'h0 : _io_out_s_funct_T_8; // @[package.scala 32:76]
  wire [2:0] _io_out_s_funct_T_12 = _io_out_s_funct_T_2 == 3'h5 ? 3'h0 : _io_out_s_funct_T_10; // @[package.scala 32:76]
  wire [2:0] _io_out_s_funct_T_14 = _io_out_s_funct_T_2 == 3'h6 ? 3'h2 : _io_out_s_funct_T_12; // @[package.scala 32:76]
  wire [2:0] io_out_s_funct = _io_out_s_funct_T_2 == 3'h7 ? 3'h3 : _io_out_s_funct_T_14; // @[package.scala 32:76]
  wire [30:0] io_out_s_sub = io_in[6:5] == 2'h0 ? 31'h40000000 : 31'h0; // @[RVC.scala 103:22]
  wire [6:0] io_out_s_opc_4 = io_in[12] ? 7'h3b : 7'h33; // @[RVC.scala 104:22]
  wire [24:0] _io_out_s_T_234 = {2'h1,io_in[4:2],2'h1,io_in[9:7],io_out_s_funct,2'h1,io_in[9:7],io_out_s_opc_4}; // @[Cat.scala 31:58]
  wire [30:0] _GEN_1 = {{6'd0}, _io_out_s_T_234}; // @[RVC.scala 105:43]
  wire [30:0] _io_out_s_T_235 = _GEN_1 | io_out_s_sub; // @[RVC.scala 105:43]
  wire [30:0] _io_out_s_T_238 = io_in[11:10] == 2'h1 ? _io_out_s_T_217 : {{5'd0}, _io_out_s_T_208}; // @[package.scala 32:76]
  wire [31:0] _io_out_s_T_240 = io_in[11:10] == 2'h2 ? _io_out_s_T_227 : {{1'd0}, _io_out_s_T_238}; // @[package.scala 32:76]
  wire [31:0] io_out_s_12_bits = io_in[11:10] == 2'h3 ? {{1'd0}, _io_out_s_T_235} : _io_out_s_T_240; // @[package.scala 32:76]
  wire [9:0] _io_out_s_T_252 = io_in[12] ? 10'h3ff : 10'h0; // @[Bitwise.scala 74:12]
  wire [20:0] _io_out_s_T_260 = {_io_out_s_T_252,io_in[8],io_in[10:9],io_in[6],io_in[7],io_in[2],io_in[11],io_in[5:3],1'h0
    }; // @[Cat.scala 31:58]
  wire [31:0] io_out_s_13_bits = {_io_out_s_T_260[20],_io_out_s_T_260[10:1],_io_out_s_T_260[11],_io_out_s_T_260[19:12],5'h0
    ,7'h6f}; // @[Cat.scala 31:58]
  wire [4:0] _io_out_s_T_306 = io_in[12] ? 5'h1f : 5'h0; // @[Bitwise.scala 74:12]
  wire [12:0] _io_out_s_T_311 = {_io_out_s_T_306,io_in[6:5],io_in[2],io_in[11:10],io_in[4:3],1'h0}; // @[Cat.scala 31:58]
  wire [31:0] io_out_s_14_bits = {_io_out_s_T_311[12],_io_out_s_T_311[10:5],5'h0,2'h1,io_in[9:7],3'h0,_io_out_s_T_311[4:
    1],_io_out_s_T_311[11],7'h63}; // @[Cat.scala 31:58]
  wire [31:0] io_out_s_15_bits = {_io_out_s_T_311[12],_io_out_s_T_311[10:5],5'h0,2'h1,io_in[9:7],3'h1,_io_out_s_T_311[4:
    1],_io_out_s_T_311[11],7'h63}; // @[Cat.scala 31:58]
  wire [6:0] io_out_s_load_opc = _io_out_s_opc_T_3 ? 7'h3 : 7'h1f; // @[RVC.scala 113:23]
  wire [25:0] _io_out_s_T_395 = {io_in[12],io_in[6:2],io_in[11:7],3'h1,io_in[11:7],7'h13}; // @[Cat.scala 31:58]
  wire [28:0] _io_out_s_T_405 = {io_in[4:2],io_in[12],io_in[6:5],3'h0,5'h2,3'h3,io_in[11:7],7'h7}; // @[Cat.scala 31:58]
  wire [27:0] _io_out_s_T_414 = {io_in[3:2],io_in[12],io_in[6:4],2'h0,5'h2,3'h2,io_in[11:7],io_out_s_load_opc}; // @[Cat.scala 31:58]
  wire [28:0] _io_out_s_T_423 = {io_in[4:2],io_in[12],io_in[6:5],3'h0,5'h2,3'h3,io_in[11:7],io_out_s_load_opc}; // @[Cat.scala 31:58]
  wire [19:0] _io_out_s_mv_T_2 = {io_in[6:2],3'h0,io_in[11:7],7'h13}; // @[Cat.scala 31:58]
  wire [24:0] _io_out_s_add_T_3 = {io_in[6:2],io_in[11:7],3'h0,io_in[11:7],7'h33}; // @[Cat.scala 31:58]
  wire [24:0] io_out_s_jr = {io_in[6:2],io_in[11:7],3'h0,12'h67}; // @[Cat.scala 31:58]
  wire [24:0] io_out_s_reserved = {io_out_s_jr[24:7],7'h1f}; // @[Cat.scala 31:58]
  wire [24:0] _io_out_s_jr_reserved_T_2 = _io_out_s_opc_T_3 ? io_out_s_jr : io_out_s_reserved; // @[RVC.scala 134:33]
  wire  _io_out_s_jr_mv_T_1 = |io_in[6:2]; // @[RVC.scala 135:27]
  wire [31:0] io_out_s_mv_bits = {{12'd0}, _io_out_s_mv_T_2}; // @[RVC.scala 21:19 22:14]
  wire [31:0] io_out_s_jr_reserved_bits = {{7'd0}, _io_out_s_jr_reserved_T_2}; // @[RVC.scala 21:19 22:14]
  wire [31:0] io_out_s_jr_mv_bits = |io_in[6:2] ? io_out_s_mv_bits : io_out_s_jr_reserved_bits; // @[RVC.scala 135:22]
  wire [24:0] io_out_s_jalr = {io_in[6:2],io_in[11:7],3'h0,12'he7}; // @[Cat.scala 31:58]
  wire [24:0] _io_out_s_ebreak_T_1 = {io_out_s_jr[24:7],7'h73}; // @[Cat.scala 31:58]
  wire [24:0] io_out_s_ebreak = _io_out_s_ebreak_T_1 | 25'h100000; // @[RVC.scala 137:46]
  wire [24:0] _io_out_s_jalr_ebreak_T_2 = _io_out_s_opc_T_3 ? io_out_s_jalr : io_out_s_ebreak; // @[RVC.scala 138:33]
  wire [31:0] io_out_s_add_bits = {{7'd0}, _io_out_s_add_T_3}; // @[RVC.scala 21:19 22:14]
  wire [31:0] io_out_s_jalr_ebreak_bits = {{7'd0}, _io_out_s_jalr_ebreak_T_2}; // @[RVC.scala 21:19 22:14]
  wire [31:0] io_out_s_jalr_add_bits = _io_out_s_jr_mv_T_1 ? io_out_s_add_bits : io_out_s_jalr_ebreak_bits; // @[RVC.scala 139:25]
  wire [31:0] io_out_s_20_bits = io_in[12] ? io_out_s_jalr_add_bits : io_out_s_jr_mv_bits; // @[RVC.scala 140:10]
  wire [8:0] _io_out_s_T_430 = {io_in[9:7],io_in[12:10],3'h0}; // @[Cat.scala 31:58]
  wire [28:0] _io_out_s_T_437 = {_io_out_s_T_430[8:5],io_in[6:2],5'h2,3'h3,_io_out_s_T_430[4:0],7'h27}; // @[Cat.scala 31:58]
  wire [7:0] _io_out_s_T_443 = {io_in[8:7],io_in[12:9],2'h0}; // @[Cat.scala 31:58]
  wire [27:0] _io_out_s_T_450 = {_io_out_s_T_443[7:5],io_in[6:2],5'h2,3'h2,_io_out_s_T_443[4:0],7'h23}; // @[Cat.scala 31:58]
  wire [28:0] _io_out_s_T_463 = {_io_out_s_T_430[8:5],io_in[6:2],5'h2,3'h3,_io_out_s_T_430[4:0],7'h23}; // @[Cat.scala 31:58]
  wire [4:0] _io_out_T_2 = {io_in[1:0],io_in[15:13]}; // @[Cat.scala 31:58]
  wire [31:0] io_out_s_1_bits = {{4'd0}, _io_out_s_T_20}; // @[RVC.scala 21:19 22:14]
  wire [31:0] io_out_s_0_bits = {{2'd0}, _io_out_s_T_7}; // @[RVC.scala 21:19 22:14]
  wire [31:0] _io_out_T_4_bits = _io_out_T_2 == 5'h1 ? io_out_s_1_bits : io_out_s_0_bits; // @[package.scala 32:76]
  wire [31:0] io_out_s_2_bits = {{5'd0}, _io_out_s_T_36}; // @[RVC.scala 21:19 22:14]
  wire [31:0] _io_out_T_6_bits = _io_out_T_2 == 5'h2 ? io_out_s_2_bits : _io_out_T_4_bits; // @[package.scala 32:76]
  wire [31:0] io_out_s_3_bits = {{4'd0}, _io_out_s_T_51}; // @[RVC.scala 21:19 22:14]
  wire [31:0] _io_out_T_8_bits = _io_out_T_2 == 5'h3 ? io_out_s_3_bits : _io_out_T_6_bits; // @[package.scala 32:76]
  wire [31:0] io_out_s_4_bits = {{5'd0}, _io_out_s_T_73}; // @[RVC.scala 21:19 22:14]
  wire [31:0] _io_out_T_10_bits = _io_out_T_2 == 5'h4 ? io_out_s_4_bits : _io_out_T_8_bits; // @[package.scala 32:76]
  wire [31:0] io_out_s_5_bits = {{4'd0}, _io_out_s_T_93}; // @[RVC.scala 21:19 22:14]
  wire [31:0] _io_out_T_12_bits = _io_out_T_2 == 5'h5 ? io_out_s_5_bits : _io_out_T_10_bits; // @[package.scala 32:76]
  wire [31:0] io_out_s_6_bits = {{5'd0}, _io_out_s_T_115}; // @[RVC.scala 21:19 22:14]
  wire [31:0] _io_out_T_14_bits = _io_out_T_2 == 5'h6 ? io_out_s_6_bits : _io_out_T_12_bits; // @[package.scala 32:76]
  wire [31:0] io_out_s_7_bits = {{4'd0}, _io_out_s_T_135}; // @[RVC.scala 21:19 22:14]
  wire [31:0] _io_out_T_16_bits = _io_out_T_2 == 5'h7 ? io_out_s_7_bits : _io_out_T_14_bits; // @[package.scala 32:76]
  wire [31:0] _io_out_T_18_bits = _io_out_T_2 == 5'h8 ? io_out_s_8_bits : _io_out_T_16_bits; // @[package.scala 32:76]
  wire [31:0] _io_out_T_20_bits = _io_out_T_2 == 5'h9 ? io_out_s_9_bits : _io_out_T_18_bits; // @[package.scala 32:76]
  wire [31:0] _io_out_T_22_bits = _io_out_T_2 == 5'ha ? io_out_s_10_bits : _io_out_T_20_bits; // @[package.scala 32:76]
  wire [31:0] _io_out_T_24_bits = _io_out_T_2 == 5'hb ? io_out_s_11_bits : _io_out_T_22_bits; // @[package.scala 32:76]
  wire [31:0] _io_out_T_26_bits = _io_out_T_2 == 5'hc ? io_out_s_12_bits : _io_out_T_24_bits; // @[package.scala 32:76]
  wire [31:0] _io_out_T_28_bits = _io_out_T_2 == 5'hd ? io_out_s_13_bits : _io_out_T_26_bits; // @[package.scala 32:76]
  wire [31:0] _io_out_T_30_bits = _io_out_T_2 == 5'he ? io_out_s_14_bits : _io_out_T_28_bits; // @[package.scala 32:76]
  wire [31:0] _io_out_T_32_bits = _io_out_T_2 == 5'hf ? io_out_s_15_bits : _io_out_T_30_bits; // @[package.scala 32:76]
  wire [31:0] io_out_s_16_bits = {{6'd0}, _io_out_s_T_395}; // @[RVC.scala 21:19 22:14]
  wire [31:0] _io_out_T_34_bits = _io_out_T_2 == 5'h10 ? io_out_s_16_bits : _io_out_T_32_bits; // @[package.scala 32:76]
  wire [31:0] io_out_s_17_bits = {{3'd0}, _io_out_s_T_405}; // @[RVC.scala 21:19 22:14]
  wire [31:0] _io_out_T_36_bits = _io_out_T_2 == 5'h11 ? io_out_s_17_bits : _io_out_T_34_bits; // @[package.scala 32:76]
  wire [31:0] io_out_s_18_bits = {{4'd0}, _io_out_s_T_414}; // @[RVC.scala 21:19 22:14]
  wire [31:0] _io_out_T_38_bits = _io_out_T_2 == 5'h12 ? io_out_s_18_bits : _io_out_T_36_bits; // @[package.scala 32:76]
  wire [31:0] io_out_s_19_bits = {{3'd0}, _io_out_s_T_423}; // @[RVC.scala 21:19 22:14]
  wire [31:0] _io_out_T_40_bits = _io_out_T_2 == 5'h13 ? io_out_s_19_bits : _io_out_T_38_bits; // @[package.scala 32:76]
  wire [31:0] _io_out_T_42_bits = _io_out_T_2 == 5'h14 ? io_out_s_20_bits : _io_out_T_40_bits; // @[package.scala 32:76]
  wire [31:0] io_out_s_21_bits = {{3'd0}, _io_out_s_T_437}; // @[RVC.scala 21:19 22:14]
  wire [31:0] _io_out_T_44_bits = _io_out_T_2 == 5'h15 ? io_out_s_21_bits : _io_out_T_42_bits; // @[package.scala 32:76]
  wire [31:0] io_out_s_22_bits = {{4'd0}, _io_out_s_T_450}; // @[RVC.scala 21:19 22:14]
  wire [31:0] _io_out_T_46_bits = _io_out_T_2 == 5'h16 ? io_out_s_22_bits : _io_out_T_44_bits; // @[package.scala 32:76]
  wire [31:0] io_out_s_23_bits = {{3'd0}, _io_out_s_T_463}; // @[RVC.scala 21:19 22:14]
  wire [31:0] _io_out_T_48_bits = _io_out_T_2 == 5'h17 ? io_out_s_23_bits : _io_out_T_46_bits; // @[package.scala 32:76]
  wire [31:0] _io_out_T_50_bits = _io_out_T_2 == 5'h18 ? io_in : _io_out_T_48_bits; // @[package.scala 32:76]
  wire [31:0] _io_out_T_52_bits = _io_out_T_2 == 5'h19 ? io_in : _io_out_T_50_bits; // @[package.scala 32:76]
  wire [31:0] _io_out_T_54_bits = _io_out_T_2 == 5'h1a ? io_in : _io_out_T_52_bits; // @[package.scala 32:76]
  wire [31:0] _io_out_T_56_bits = _io_out_T_2 == 5'h1b ? io_in : _io_out_T_54_bits; // @[package.scala 32:76]
  wire [31:0] _io_out_T_58_bits = _io_out_T_2 == 5'h1c ? io_in : _io_out_T_56_bits; // @[package.scala 32:76]
  wire [31:0] _io_out_T_60_bits = _io_out_T_2 == 5'h1d ? io_in : _io_out_T_58_bits; // @[package.scala 32:76]
  wire [31:0] _io_out_T_62_bits = _io_out_T_2 == 5'h1e ? io_in : _io_out_T_60_bits; // @[package.scala 32:76]
  assign io_out_bits = _io_out_T_2 == 5'h1f ? io_in : _io_out_T_62_bits; // @[package.scala 32:76]
endmodule

