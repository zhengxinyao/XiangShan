module DelayN_66(
  input  [1:0] io_in,
  output [1:0] io_out
);
  assign io_out = io_in; // @[Hold.scala 92:10]
endmodule

