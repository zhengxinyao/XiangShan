module MemBlock(
  input          clock,
  input          reset,
  input          auto_uncache_client_out_a_ready,
  output         auto_uncache_client_out_a_valid,
  output [2:0]   auto_uncache_client_out_a_bits_opcode,
  output [2:0]   auto_uncache_client_out_a_bits_size,
  output [1:0]   auto_uncache_client_out_a_bits_source,
  output [35:0]  auto_uncache_client_out_a_bits_address,
  output [7:0]   auto_uncache_client_out_a_bits_mask,
  output [63:0]  auto_uncache_client_out_a_bits_data,
  output         auto_uncache_client_out_d_ready,
  input          auto_uncache_client_out_d_valid,
  input  [2:0]   auto_uncache_client_out_d_bits_opcode,
  input  [63:0]  auto_uncache_client_out_d_bits_data,
  input          auto_dcache_client_out_a_ready,
  output         auto_dcache_client_out_a_valid,
  output [2:0]   auto_dcache_client_out_a_bits_opcode,
  output [2:0]   auto_dcache_client_out_a_bits_param,
  output [2:0]   auto_dcache_client_out_a_bits_size,
  output [3:0]   auto_dcache_client_out_a_bits_source,
  output [35:0]  auto_dcache_client_out_a_bits_address,
  output [31:0]  auto_dcache_client_out_a_bits_mask,
  output         auto_dcache_client_out_bready,
  input          auto_dcache_client_out_bvalid,
  input  [1:0]   auto_dcache_client_out_bparam,
  input  [35:0]  auto_dcache_client_out_baddress,
  input  [255:0] auto_dcache_client_out_bdata,
  input          auto_dcache_client_out_c_ready,
  output         auto_dcache_client_out_c_valid,
  output [2:0]   auto_dcache_client_out_c_bits_opcode,
  output [2:0]   auto_dcache_client_out_c_bits_param,
  output [2:0]   auto_dcache_client_out_c_bits_size,
  output [3:0]   auto_dcache_client_out_c_bits_source,
  output [35:0]  auto_dcache_client_out_c_bits_address,
  output         auto_dcache_client_out_c_bits_echo_blockisdirty,
  output [255:0] auto_dcache_client_out_c_bits_data,
  output         auto_dcache_client_out_d_ready,
  input          auto_dcache_client_out_d_valid,
  input  [2:0]   auto_dcache_client_out_d_bits_opcode,
  input  [1:0]   auto_dcache_client_out_d_bits_param,
  input  [2:0]   auto_dcache_client_out_d_bits_size,
  input  [3:0]   auto_dcache_client_out_d_bits_source,
  input  [3:0]   auto_dcache_client_out_d_bits_sink,
  input          auto_dcache_client_out_d_bits_denied,
  input          auto_dcache_client_out_d_bits_echo_blockisdirty,
  input  [255:0] auto_dcache_client_out_d_bits_data,
  input          auto_dcache_client_out_d_bits_corrupt,
  input          auto_dcache_client_out_e_ready,
  output         auto_dcache_client_out_e_valid,
  output [3:0]   auto_dcache_client_out_e_bits_sink,
  input  [7:0]   io_hartId,
  input          io_redirect_valid,
  input          io_redirect_bits_robIdx_flag,
  input  [4:0]   io_redirect_bits_robIdx_value,
  input          io_redirect_bits_level,
  output         io_issue_0_ready,
  input          io_issue_0_valid,
  input  [9:0]   io_issue_0_bits_uop_cf_foldpc,
  input          io_issue_0_bits_uop_cf_trigger_backendEn_1,
  input          io_issue_0_bits_uop_cf_waitForRobIdx_flag,
  input  [4:0]   io_issue_0_bits_uop_cf_waitForRobIdx_value,
  input          io_issue_0_bits_uop_cf_loadWaitBit,
  input          io_issue_0_bits_uop_cf_loadWaitStrict,
  input          io_issue_0_bits_uop_cf_ftqPtr_flag,
  input  [2:0]   io_issue_0_bits_uop_cf_ftqPtr_value,
  input  [2:0]   io_issue_0_bits_uop_cf_ftqOffset,
  input  [3:0]   io_issue_0_bits_uop_ctrl_fuType,
  input  [6:0]   io_issue_0_bits_uop_ctrl_fuOpType,
  input          io_issue_0_bits_uop_ctrl_rfWen,
  input          io_issue_0_bits_uop_ctrl_fpWen,
  input  [19:0]  io_issue_0_bits_uop_ctrl_imm,
  input  [5:0]   io_issue_0_bits_uop_pdest,
  input          io_issue_0_bits_uop_robIdx_flag,
  input  [4:0]   io_issue_0_bits_uop_robIdx_value,
  input          io_issue_0_bits_uop_lqIdx_flag,
  input  [3:0]   io_issue_0_bits_uop_lqIdx_value,
  input          io_issue_0_bits_uop_sqIdx_flag,
  input  [3:0]   io_issue_0_bits_uop_sqIdx_value,
  input  [63:0]  io_issue_0_bits_src_0,
  output         io_issue_1_ready,
  input          io_issue_1_valid,
  input  [9:0]   io_issue_1_bits_uop_cf_foldpc,
  input          io_issue_1_bits_uop_cf_trigger_backendEn_1,
  input          io_issue_1_bits_uop_cf_waitForRobIdx_flag,
  input  [4:0]   io_issue_1_bits_uop_cf_waitForRobIdx_value,
  input          io_issue_1_bits_uop_cf_loadWaitBit,
  input          io_issue_1_bits_uop_cf_loadWaitStrict,
  input          io_issue_1_bits_uop_cf_ftqPtr_flag,
  input  [2:0]   io_issue_1_bits_uop_cf_ftqPtr_value,
  input  [2:0]   io_issue_1_bits_uop_cf_ftqOffset,
  input  [3:0]   io_issue_1_bits_uop_ctrl_fuType,
  input  [6:0]   io_issue_1_bits_uop_ctrl_fuOpType,
  input          io_issue_1_bits_uop_ctrl_rfWen,
  input          io_issue_1_bits_uop_ctrl_fpWen,
  input  [19:0]  io_issue_1_bits_uop_ctrl_imm,
  input  [5:0]   io_issue_1_bits_uop_pdest,
  input          io_issue_1_bits_uop_robIdx_flag,
  input  [4:0]   io_issue_1_bits_uop_robIdx_value,
  input          io_issue_1_bits_uop_lqIdx_flag,
  input  [3:0]   io_issue_1_bits_uop_lqIdx_value,
  input          io_issue_1_bits_uop_sqIdx_flag,
  input  [3:0]   io_issue_1_bits_uop_sqIdx_value,
  input  [63:0]  io_issue_1_bits_src_0,
  output         io_issue_2_ready,
  input          io_issue_2_valid,
  input          io_issue_2_bits_uop_cf_trigger_backendEn_0,
  input          io_issue_2_bits_uop_cf_trigger_backendEn_1,
  input          io_issue_2_bits_uop_cf_storeSetHit,
  input  [4:0]   io_issue_2_bits_uop_cf_ssid,
  input  [2:0]   io_issue_2_bits_uop_cf_ftqPtr_value,
  input  [2:0]   io_issue_2_bits_uop_cf_ftqOffset,
  input  [3:0]   io_issue_2_bits_uop_ctrl_fuType,
  input  [6:0]   io_issue_2_bits_uop_ctrl_fuOpType,
  input          io_issue_2_bits_uop_ctrl_rfWen,
  input          io_issue_2_bits_uop_ctrl_fpWen,
  input  [19:0]  io_issue_2_bits_uop_ctrl_imm,
  input  [5:0]   io_issue_2_bits_uop_pdest,
  input          io_issue_2_bits_uop_robIdx_flag,
  input  [4:0]   io_issue_2_bits_uop_robIdx_value,
  input          io_issue_2_bits_uop_sqIdx_flag,
  input  [3:0]   io_issue_2_bits_uop_sqIdx_value,
  input  [63:0]  io_issue_2_bits_src_0,
  output         io_issue_3_ready,
  input          io_issue_3_valid,
  input          io_issue_3_bits_uop_cf_trigger_backendEn_0,
  input          io_issue_3_bits_uop_cf_trigger_backendEn_1,
  input          io_issue_3_bits_uop_cf_storeSetHit,
  input  [4:0]   io_issue_3_bits_uop_cf_ssid,
  input  [2:0]   io_issue_3_bits_uop_cf_ftqPtr_value,
  input  [2:0]   io_issue_3_bits_uop_cf_ftqOffset,
  input  [3:0]   io_issue_3_bits_uop_ctrl_fuType,
  input  [6:0]   io_issue_3_bits_uop_ctrl_fuOpType,
  input          io_issue_3_bits_uop_ctrl_rfWen,
  input          io_issue_3_bits_uop_ctrl_fpWen,
  input  [19:0]  io_issue_3_bits_uop_ctrl_imm,
  input  [5:0]   io_issue_3_bits_uop_pdest,
  input          io_issue_3_bits_uop_robIdx_flag,
  input  [4:0]   io_issue_3_bits_uop_robIdx_value,
  input          io_issue_3_bits_uop_sqIdx_flag,
  input  [3:0]   io_issue_3_bits_uop_sqIdx_value,
  input  [63:0]  io_issue_3_bits_src_0,
  output         io_issue_4_ready,
  input          io_issue_4_valid,
  input  [3:0]   io_issue_4_bits_uop_ctrl_fuType,
  input  [6:0]   io_issue_4_bits_uop_ctrl_fuOpType,
  input          io_issue_4_bits_uop_robIdx_flag,
  input  [4:0]   io_issue_4_bits_uop_robIdx_value,
  input          io_issue_4_bits_uop_sqIdx_flag,
  input  [3:0]   io_issue_4_bits_uop_sqIdx_value,
  input  [63:0]  io_issue_4_bits_src_0,
  output         io_issue_5_ready,
  input          io_issue_5_valid,
  input  [3:0]   io_issue_5_bits_uop_ctrl_fuType,
  input  [6:0]   io_issue_5_bits_uop_ctrl_fuOpType,
  input          io_issue_5_bits_uop_robIdx_flag,
  input  [4:0]   io_issue_5_bits_uop_robIdx_value,
  input          io_issue_5_bits_uop_sqIdx_flag,
  input  [3:0]   io_issue_5_bits_uop_sqIdx_value,
  input  [63:0]  io_issue_5_bits_src_0,
  input  [1:0]   io_loadFastMatch_0,
  input  [1:0]   io_loadFastMatch_1,
  input  [11:0]  io_loadFastImm_0,
  input  [11:0]  io_loadFastImm_1,
  output         io_rsfeedback_0_feedbackSlow_valid,
  output [3:0]   io_rsfeedback_0_feedbackSlow_bits_rsIdx,
  output         io_rsfeedback_0_feedbackSlow_bits_hit,
  input  [3:0]   io_rsfeedback_0_rsIdx,
  output         io_rsfeedback_1_feedbackSlow_valid,
  output [3:0]   io_rsfeedback_1_feedbackSlow_bits_rsIdx,
  output         io_rsfeedback_1_feedbackSlow_bits_hit,
  input  [3:0]   io_rsfeedback_1_rsIdx,
  input          io_writeback_0_ready,
  output         io_writeback_0_valid,
  output         io_writeback_0_bits_uop_cf_exceptionVec_4,
  output         io_writeback_0_bits_uop_cf_exceptionVec_5,
  output         io_writeback_0_bits_uop_cf_exceptionVec_13,
  output         io_writeback_0_bits_uop_cf_trigger_backendEn_1,
  output         io_writeback_0_bits_uop_cf_trigger_backendHit_0,
  output         io_writeback_0_bits_uop_cf_trigger_backendHit_1,
  output         io_writeback_0_bits_uop_cf_trigger_backendHit_2,
  output         io_writeback_0_bits_uop_cf_trigger_backendHit_3,
  output         io_writeback_0_bits_uop_cf_trigger_backendHit_4,
  output         io_writeback_0_bits_uop_cf_trigger_backendHit_5,
  output         io_writeback_0_bits_uop_ctrl_rfWen,
  output         io_writeback_0_bits_uop_ctrl_fpWen,
  output         io_writeback_0_bits_uop_ctrl_flushPipe,
  output         io_writeback_0_bits_uop_ctrl_replayInst,
  output [5:0]   io_writeback_0_bits_uop_pdest,
  output         io_writeback_0_bits_uop_robIdx_flag,
  output [4:0]   io_writeback_0_bits_uop_robIdx_value,
  output [63:0]  io_writeback_0_bits_data,
  output         io_writeback_0_bits_debug_isMMIO,
  input          io_writeback_1_ready,
  output         io_writeback_1_valid,
  output         io_writeback_1_bits_uop_cf_exceptionVec_4,
  output         io_writeback_1_bits_uop_cf_exceptionVec_5,
  output         io_writeback_1_bits_uop_cf_exceptionVec_13,
  output         io_writeback_1_bits_uop_cf_trigger_backendEn_1,
  output         io_writeback_1_bits_uop_cf_trigger_backendHit_0,
  output         io_writeback_1_bits_uop_cf_trigger_backendHit_1,
  output         io_writeback_1_bits_uop_cf_trigger_backendHit_2,
  output         io_writeback_1_bits_uop_cf_trigger_backendHit_3,
  output         io_writeback_1_bits_uop_cf_trigger_backendHit_4,
  output         io_writeback_1_bits_uop_cf_trigger_backendHit_5,
  output         io_writeback_1_bits_uop_ctrl_rfWen,
  output         io_writeback_1_bits_uop_ctrl_fpWen,
  output         io_writeback_1_bits_uop_ctrl_flushPipe,
  output         io_writeback_1_bits_uop_ctrl_replayInst,
  output [5:0]   io_writeback_1_bits_uop_pdest,
  output         io_writeback_1_bits_uop_robIdx_flag,
  output [4:0]   io_writeback_1_bits_uop_robIdx_value,
  output [63:0]  io_writeback_1_bits_data,
  output         io_writeback_1_bits_debug_isMMIO,
  input          io_writeback_2_ready,
  output         io_writeback_2_valid,
  output         io_writeback_2_bits_uop_cf_exceptionVec_4,
  output         io_writeback_2_bits_uop_cf_exceptionVec_5,
  output         io_writeback_2_bits_uop_cf_exceptionVec_6,
  output         io_writeback_2_bits_uop_cf_exceptionVec_7,
  output         io_writeback_2_bits_uop_cf_exceptionVec_13,
  output         io_writeback_2_bits_uop_cf_exceptionVec_15,
  output         io_writeback_2_bits_uop_cf_trigger_backendEn_0,
  output         io_writeback_2_bits_uop_cf_trigger_backendHit_0,
  output         io_writeback_2_bits_uop_cf_trigger_backendHit_1,
  output         io_writeback_2_bits_uop_cf_trigger_backendHit_2,
  output         io_writeback_2_bits_uop_cf_trigger_backendHit_3,
  output         io_writeback_2_bits_uop_cf_trigger_backendHit_4,
  output         io_writeback_2_bits_uop_cf_trigger_backendHit_5,
  output         io_writeback_2_bits_uop_robIdx_flag,
  output [4:0]   io_writeback_2_bits_uop_robIdx_value,
  output         io_writeback_2_bits_debug_isMMIO,
  output [38:0]  io_writeback_2_bits_debug_vaddr,
  input          io_writeback_3_ready,
  output         io_writeback_3_valid,
  output         io_writeback_3_bits_uop_cf_exceptionVec_6,
  output         io_writeback_3_bits_uop_cf_exceptionVec_7,
  output         io_writeback_3_bits_uop_cf_exceptionVec_15,
  output         io_writeback_3_bits_uop_cf_trigger_backendEn_0,
  output         io_writeback_3_bits_uop_cf_trigger_backendHit_0,
  output         io_writeback_3_bits_uop_cf_trigger_backendHit_1,
  output         io_writeback_3_bits_uop_cf_trigger_backendHit_4,
  output         io_writeback_3_bits_uop_robIdx_flag,
  output [4:0]   io_writeback_3_bits_uop_robIdx_value,
  output         io_writeback_3_bits_debug_isMMIO,
  output [38:0]  io_writeback_3_bits_debug_vaddr,
  output         io_writeback_4_valid,
  output         io_writeback_4_bits_uop_robIdx_flag,
  output [4:0]   io_writeback_4_bits_uop_robIdx_value,
  output         io_writeback_5_valid,
  output         io_writeback_5_bits_uop_robIdx_flag,
  output [4:0]   io_writeback_5_bits_uop_robIdx_value,
  output         io_stIn_0_valid,
  output         io_stIn_0_bits_uop_cf_storeSetHit,
  output [4:0]   io_stIn_0_bits_uop_cf_ssid,
  output [4:0]   io_stIn_0_bits_uop_robIdx_value,
  output         io_stIn_1_valid,
  output         io_stIn_1_bits_uop_cf_storeSetHit,
  output [4:0]   io_stIn_1_bits_uop_cf_ssid,
  output [4:0]   io_stIn_1_bits_uop_robIdx_value,
  output         io_memoryViolation_valid,
  output         io_memoryViolation_bits_robIdx_flag,
  output [4:0]   io_memoryViolation_bits_robIdx_value,
  output         io_memoryViolation_bits_ftqIdx_flag,
  output [2:0]   io_memoryViolation_bits_ftqIdx_value,
  output [2:0]   io_memoryViolation_bits_ftqOffset,
  output [2:0]   io_memoryViolation_bits_stFtqIdx_value,
  output [2:0]   io_memoryViolation_bits_stFtqOffset,
  output         io_ptw_req_0_valid,
  output [26:0]  io_ptw_req_0_bits_vpn,
  output         io_ptw_req_1_valid,
  output [26:0]  io_ptw_req_1_bits_vpn,
  output         io_ptw_req_2_valid,
  output [26:0]  io_ptw_req_2_bits_vpn,
  output         io_ptw_req_3_valid,
  output [26:0]  io_ptw_req_3_bits_vpn,
  input          io_ptw_resp_valid,
  input  [26:0]  io_ptw_resp_bits_data_entry_tag,
  input  [15:0]  io_ptw_resp_bits_data_entry_asid,
  input  [23:0]  io_ptw_resp_bits_data_entry_ppn,
  input          io_ptw_resp_bits_data_entry_perm_d,
  input          io_ptw_resp_bits_data_entry_perm_a,
  input          io_ptw_resp_bits_data_entry_perm_g,
  input          io_ptw_resp_bits_data_entry_perm_u,
  input          io_ptw_resp_bits_data_entry_perm_x,
  input          io_ptw_resp_bits_data_entry_perm_w,
  input          io_ptw_resp_bits_data_entry_perm_r,
  input  [1:0]   io_ptw_resp_bits_data_entry_level,
  input          io_ptw_resp_bits_data_pf,
  input          io_ptw_resp_bits_data_af,
  input          io_ptw_resp_bits_vector_0,
  input          io_ptw_resp_bits_vector_1,
  input          io_ptw_resp_bits_vector_2,
  input          io_ptw_resp_bits_vector_3,
  input          io_ptw_resp_bits_vector_4,
  input          io_sfence_valid,
  input          io_sfence_bits_rs1,
  input          io_sfence_bits_rs2,
  input  [38:0]  io_sfence_bits_addr,
  input  [15:0]  io_sfence_bits_asid,
  input  [3:0]   io_tlbCsr_satp_mode,
  input  [15:0]  io_tlbCsr_satp_asid,
  input          io_tlbCsr_satp_changed,
  input          io_tlbCsr_priv_mxr,
  input          io_tlbCsr_priv_sum,
  input  [1:0]   io_tlbCsr_priv_dmode,
  input          io_fenceToSbuffer_flushSb,
  output         io_fenceToSbuffer_sbIsEmpty,
  input  [1:0]   io_enqLsq_needAlloc_0,
  input  [1:0]   io_enqLsq_needAlloc_1,
  input  [1:0]   io_enqLsq_needAlloc_2,
  input  [1:0]   io_enqLsq_needAlloc_3,
  input          io_enqLsq_req_0_valid,
  input          io_enqLsq_req_0_bits_cf_trigger_backendEn_0,
  input          io_enqLsq_req_0_bits_cf_trigger_backendEn_1,
  input  [6:0]   io_enqLsq_req_0_bits_ctrl_fuOpType,
  input          io_enqLsq_req_0_bits_ctrl_rfWen,
  input          io_enqLsq_req_0_bits_ctrl_fpWen,
  input          io_enqLsq_req_0_bits_ctrl_flushPipe,
  input          io_enqLsq_req_0_bits_ctrl_replayInst,
  input  [5:0]   io_enqLsq_req_0_bits_pdest,
  input          io_enqLsq_req_0_bits_robIdx_flag,
  input  [4:0]   io_enqLsq_req_0_bits_robIdx_value,
  input  [3:0]   io_enqLsq_req_0_bits_lqIdx_value,
  input  [3:0]   io_enqLsq_req_0_bits_sqIdx_value,
  input          io_enqLsq_req_1_valid,
  input          io_enqLsq_req_1_bits_cf_trigger_backendEn_0,
  input          io_enqLsq_req_1_bits_cf_trigger_backendEn_1,
  input  [6:0]   io_enqLsq_req_1_bits_ctrl_fuOpType,
  input          io_enqLsq_req_1_bits_ctrl_rfWen,
  input          io_enqLsq_req_1_bits_ctrl_fpWen,
  input          io_enqLsq_req_1_bits_ctrl_flushPipe,
  input          io_enqLsq_req_1_bits_ctrl_replayInst,
  input  [5:0]   io_enqLsq_req_1_bits_pdest,
  input          io_enqLsq_req_1_bits_robIdx_flag,
  input  [4:0]   io_enqLsq_req_1_bits_robIdx_value,
  input  [3:0]   io_enqLsq_req_1_bits_lqIdx_value,
  input  [3:0]   io_enqLsq_req_1_bits_sqIdx_value,
  input          io_enqLsq_req_2_valid,
  input          io_enqLsq_req_2_bits_cf_trigger_backendEn_0,
  input          io_enqLsq_req_2_bits_cf_trigger_backendEn_1,
  input  [6:0]   io_enqLsq_req_2_bits_ctrl_fuOpType,
  input          io_enqLsq_req_2_bits_ctrl_rfWen,
  input          io_enqLsq_req_2_bits_ctrl_fpWen,
  input          io_enqLsq_req_2_bits_ctrl_flushPipe,
  input          io_enqLsq_req_2_bits_ctrl_replayInst,
  input  [5:0]   io_enqLsq_req_2_bits_pdest,
  input          io_enqLsq_req_2_bits_robIdx_flag,
  input  [4:0]   io_enqLsq_req_2_bits_robIdx_value,
  input  [3:0]   io_enqLsq_req_2_bits_lqIdx_value,
  input  [3:0]   io_enqLsq_req_2_bits_sqIdx_value,
  input          io_enqLsq_req_3_valid,
  input          io_enqLsq_req_3_bits_cf_trigger_backendEn_0,
  input          io_enqLsq_req_3_bits_cf_trigger_backendEn_1,
  input  [6:0]   io_enqLsq_req_3_bits_ctrl_fuOpType,
  input          io_enqLsq_req_3_bits_ctrl_rfWen,
  input          io_enqLsq_req_3_bits_ctrl_fpWen,
  input          io_enqLsq_req_3_bits_ctrl_flushPipe,
  input          io_enqLsq_req_3_bits_ctrl_replayInst,
  input  [5:0]   io_enqLsq_req_3_bits_pdest,
  input          io_enqLsq_req_3_bits_robIdx_flag,
  input  [4:0]   io_enqLsq_req_3_bits_robIdx_value,
  input  [3:0]   io_enqLsq_req_3_bits_lqIdx_value,
  input  [3:0]   io_enqLsq_req_3_bits_sqIdx_value,
  input          io_lsqio_exceptionAddr_isStore,
  output [38:0]  io_lsqio_exceptionAddr_vaddr,
  input  [1:0]   io_lsqio_rob_scommit,
  input          io_lsqio_rob_pendingld,
  input          io_lsqio_rob_pendingst,
  input          io_lsqio_rob_commit,
  output         io_lsqio_rob_isMMIO_0,
  output         io_lsqio_rob_isMMIO_1,
  output [4:0]   io_lsqio_rob_uop_0_robIdx_value,
  output [4:0]   io_lsqio_rob_uop_1_robIdx_value,
  input          io_csrCtrl_icache_parity_enable,
  input          io_csrCtrl_lvpred_disable,
  input          io_csrCtrl_no_spec_load,
  input          io_csrCtrl_storeset_wait_store,
  input  [4:0]   io_csrCtrl_lvpred_timeout,
  input          io_csrCtrl_bp_ctrl_ubtb_enable,
  input          io_csrCtrl_bp_ctrl_btb_enable,
  input          io_csrCtrl_bp_ctrl_tage_enable,
  input          io_csrCtrl_bp_ctrl_sc_enable,
  input          io_csrCtrl_bp_ctrl_ras_enable,
  input  [3:0]   io_csrCtrl_sbuffer_threshold,
  input          io_csrCtrl_ldld_vio_check_enable,
  input          io_csrCtrl_cache_error_enable,
  input          io_csrCtrl_uncache_write_outstanding_enable,
  input          io_csrCtrl_fusion_enable,
  input          io_csrCtrl_wfi_enable,
  input          io_csrCtrl_svinval_enable,
  input          io_csrCtrl_distribute_csr_wvalid,
  input  [11:0]  io_csrCtrl_distribute_csr_waddr,
  input  [63:0]  io_csrCtrl_distribute_csr_wdata,
  input          io_csrCtrl_singlestep,
  input          io_csrCtrl_frontend_trigger_t_valid,
  input  [1:0]   io_csrCtrl_frontend_trigger_t_bits_addr,
  input  [1:0]   io_csrCtrl_frontend_trigger_t_bits_tdata_matchType,
  input          io_csrCtrl_frontend_trigger_t_bits_tdata_select,
  input          io_csrCtrl_frontend_trigger_t_bits_tdata_timing,
  input          io_csrCtrl_frontend_trigger_t_bits_tdata_chain,
  input  [63:0]  io_csrCtrl_frontend_trigger_t_bits_tdata_tdata2,
  input          io_csrCtrl_mem_trigger_t_valid,
  input  [2:0]   io_csrCtrl_mem_trigger_t_bits_addr,
  input  [1:0]   io_csrCtrl_mem_trigger_t_bits_tdata_matchType,
  input          io_csrCtrl_mem_trigger_t_bits_tdata_select,
  input          io_csrCtrl_mem_trigger_t_bits_tdata_chain,
  input  [63:0]  io_csrCtrl_mem_trigger_t_bits_tdata_tdata2,
  input          io_csrCtrl_trigger_enable_0,
  input          io_csrCtrl_trigger_enable_1,
  input          io_csrCtrl_trigger_enable_2,
  input          io_csrCtrl_trigger_enable_3,
  input          io_csrCtrl_trigger_enable_4,
  input          io_csrCtrl_trigger_enable_5,
  input          io_csrCtrl_trigger_enable_6,
  input          io_csrCtrl_trigger_enable_7,
  input          io_csrCtrl_trigger_enable_8,
  input          io_csrCtrl_trigger_enable_9,
  output         io_csrUpdate_wvalid,
  output [11:0]  io_csrUpdate_waddr,
  output [63:0]  io_csrUpdate_wdata,
  output [35:0]  io_error_paddr,
  output         io_error_report_to_beu,
  input  [5:0]   io_perfEventsPTW_0_value,
  input  [5:0]   io_perfEventsPTW_1_value,
  input  [5:0]   io_perfEventsPTW_2_value,
  input  [5:0]   io_perfEventsPTW_3_value,
  input  [5:0]   io_perfEventsPTW_4_value,
  input  [5:0]   io_perfEventsPTW_5_value,
  input  [5:0]   io_perfEventsPTW_6_value,
  input  [5:0]   io_perfEventsPTW_7_value,
  input  [5:0]   io_perfEventsPTW_8_value,
  input  [5:0]   io_perfEventsPTW_9_value,
  input  [5:0]   io_perfEventsPTW_10_value,
  input  [5:0]   io_perfEventsPTW_11_value,
  input  [5:0]   io_perfEventsPTW_12_value,
  input  [5:0]   io_perfEventsPTW_13_value,
  input  [5:0]   io_perfEventsPTW_14_value,
  input  [5:0]   io_perfEventsPTW_15_value,
  input  [5:0]   io_perfEventsPTW_16_value,
  input  [5:0]   io_perfEventsPTW_17_value,
  input  [5:0]   io_perfEventsPTW_18_value,
  output [4:0]   io_lqCancelCnt,
  output [3:0]   io_sqCancelCnt,
  output [1:0]   io_sqDeq,
  output [1:0]   io_lqDeq,
  output [5:0]   io_perf_0_value,
  output [5:0]   io_perf_1_value,
  output [5:0]   io_perf_2_value,
  output [5:0]   io_perf_3_value,
  output [5:0]   io_perf_4_value,
  output [5:0]   io_perf_5_value,
  output [5:0]   io_perf_6_value,
  output [5:0]   io_perf_7_value
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [63:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [63:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [63:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [63:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [63:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [63:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [63:0] _RAND_84;
  reg [63:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
`endif // RANDOMIZE_REG_INIT
  wire  dcache_clock; // @[MemBlock.scala 47:26]
  wire  dcache_reset; // @[MemBlock.scala 47:26]
  wire  dcache_auto_client_out_a_ready; // @[MemBlock.scala 47:26]
  wire  dcache_auto_client_out_a_valid; // @[MemBlock.scala 47:26]
  wire [2:0] dcache_auto_client_out_a_bits_opcode; // @[MemBlock.scala 47:26]
  wire [2:0] dcache_auto_client_out_a_bits_param; // @[MemBlock.scala 47:26]
  wire [2:0] dcache_auto_client_out_a_bits_size; // @[MemBlock.scala 47:26]
  wire [3:0] dcache_auto_client_out_a_bits_source; // @[MemBlock.scala 47:26]
  wire [35:0] dcache_auto_client_out_a_bits_address; // @[MemBlock.scala 47:26]
  wire [31:0] dcache_auto_client_out_a_bits_mask; // @[MemBlock.scala 47:26]
  wire  dcache_auto_client_out_bready; // @[MemBlock.scala 47:26]
  wire  dcache_auto_client_out_bvalid; // @[MemBlock.scala 47:26]
  wire [1:0] dcache_auto_client_out_bparam; // @[MemBlock.scala 47:26]
  wire [35:0] dcache_auto_client_out_baddress; // @[MemBlock.scala 47:26]
  wire [255:0] dcache_auto_client_out_bdata; // @[MemBlock.scala 47:26]
  wire  dcache_auto_client_out_c_ready; // @[MemBlock.scala 47:26]
  wire  dcache_auto_client_out_c_valid; // @[MemBlock.scala 47:26]
  wire [2:0] dcache_auto_client_out_c_bits_opcode; // @[MemBlock.scala 47:26]
  wire [2:0] dcache_auto_client_out_c_bits_param; // @[MemBlock.scala 47:26]
  wire [2:0] dcache_auto_client_out_c_bits_size; // @[MemBlock.scala 47:26]
  wire [3:0] dcache_auto_client_out_c_bits_source; // @[MemBlock.scala 47:26]
  wire [35:0] dcache_auto_client_out_c_bits_address; // @[MemBlock.scala 47:26]
  wire  dcache_auto_client_out_c_bits_echo_blockisdirty; // @[MemBlock.scala 47:26]
  wire [255:0] dcache_auto_client_out_c_bits_data; // @[MemBlock.scala 47:26]
  wire  dcache_auto_client_out_d_ready; // @[MemBlock.scala 47:26]
  wire  dcache_auto_client_out_d_valid; // @[MemBlock.scala 47:26]
  wire [2:0] dcache_auto_client_out_d_bits_opcode; // @[MemBlock.scala 47:26]
  wire [1:0] dcache_auto_client_out_d_bits_param; // @[MemBlock.scala 47:26]
  wire [2:0] dcache_auto_client_out_d_bits_size; // @[MemBlock.scala 47:26]
  wire [3:0] dcache_auto_client_out_d_bits_source; // @[MemBlock.scala 47:26]
  wire [3:0] dcache_auto_client_out_d_bits_sink; // @[MemBlock.scala 47:26]
  wire  dcache_auto_client_out_d_bits_denied; // @[MemBlock.scala 47:26]
  wire  dcache_auto_client_out_d_bits_echo_blockisdirty; // @[MemBlock.scala 47:26]
  wire [255:0] dcache_auto_client_out_d_bits_data; // @[MemBlock.scala 47:26]
  wire  dcache_auto_client_out_d_bits_corrupt; // @[MemBlock.scala 47:26]
  wire  dcache_auto_client_out_e_ready; // @[MemBlock.scala 47:26]
  wire  dcache_auto_client_out_e_valid; // @[MemBlock.scala 47:26]
  wire [3:0] dcache_auto_client_out_e_bits_sink; // @[MemBlock.scala 47:26]
  wire  dcache_io_lsu_load_0_req_ready; // @[MemBlock.scala 47:26]
  wire  dcache_io_lsu_load_0_req_valid; // @[MemBlock.scala 47:26]
  wire [4:0] dcache_io_lsu_load_0_req_bits_cmd; // @[MemBlock.scala 47:26]
  wire [35:0] dcache_io_lsu_load_0_req_bits_addr; // @[MemBlock.scala 47:26]
  wire [3:0] dcache_io_lsu_load_0_req_bits_instrtype; // @[MemBlock.scala 47:26]
  wire [7:0] dcache_io_lsu_load_0_req_bits_replayCarry_real_way_en; // @[MemBlock.scala 47:26]
  wire  dcache_io_lsu_load_0_req_bits_replayCarry_valid; // @[MemBlock.scala 47:26]
  wire [127:0] dcache_io_lsu_load_0_resp_bits_data_delayed; // @[MemBlock.scala 47:26]
  wire  dcache_io_lsu_load_0_resp_bits_miss; // @[MemBlock.scala 47:26]
  wire  dcache_io_lsu_load_0_resp_bits_replay; // @[MemBlock.scala 47:26]
  wire [7:0] dcache_io_lsu_load_0_resp_bits_replayCarry_real_way_en; // @[MemBlock.scala 47:26]
  wire  dcache_io_lsu_load_0_resp_bits_replayCarry_valid; // @[MemBlock.scala 47:26]
  wire  dcache_io_lsu_load_0_resp_bits_tag_error; // @[MemBlock.scala 47:26]
  wire [1:0] dcache_io_lsu_load_0_resp_bits_mshr_id; // @[MemBlock.scala 47:26]
  wire  dcache_io_lsu_load_0_resp_bits_error_delayed; // @[MemBlock.scala 47:26]
  wire  dcache_io_lsu_load_0_s1_kill; // @[MemBlock.scala 47:26]
  wire  dcache_io_lsu_load_0_s2_kill; // @[MemBlock.scala 47:26]
  wire [35:0] dcache_io_lsu_load_0_s1_paddr_dup_lsu; // @[MemBlock.scala 47:26]
  wire [35:0] dcache_io_lsu_load_0_s1_paddr_dup_dcache; // @[MemBlock.scala 47:26]
  wire  dcache_io_lsu_load_0_s1_bank_conflict; // @[MemBlock.scala 47:26]
  wire  dcache_io_lsu_load_1_req_ready; // @[MemBlock.scala 47:26]
  wire  dcache_io_lsu_load_1_req_valid; // @[MemBlock.scala 47:26]
  wire [4:0] dcache_io_lsu_load_1_req_bits_cmd; // @[MemBlock.scala 47:26]
  wire [35:0] dcache_io_lsu_load_1_req_bits_addr; // @[MemBlock.scala 47:26]
  wire [3:0] dcache_io_lsu_load_1_req_bits_instrtype; // @[MemBlock.scala 47:26]
  wire [7:0] dcache_io_lsu_load_1_req_bits_replayCarry_real_way_en; // @[MemBlock.scala 47:26]
  wire  dcache_io_lsu_load_1_req_bits_replayCarry_valid; // @[MemBlock.scala 47:26]
  wire [127:0] dcache_io_lsu_load_1_resp_bits_data_delayed; // @[MemBlock.scala 47:26]
  wire  dcache_io_lsu_load_1_resp_bits_miss; // @[MemBlock.scala 47:26]
  wire  dcache_io_lsu_load_1_resp_bits_replay; // @[MemBlock.scala 47:26]
  wire [7:0] dcache_io_lsu_load_1_resp_bits_replayCarry_real_way_en; // @[MemBlock.scala 47:26]
  wire  dcache_io_lsu_load_1_resp_bits_replayCarry_valid; // @[MemBlock.scala 47:26]
  wire  dcache_io_lsu_load_1_resp_bits_tag_error; // @[MemBlock.scala 47:26]
  wire [1:0] dcache_io_lsu_load_1_resp_bits_mshr_id; // @[MemBlock.scala 47:26]
  wire  dcache_io_lsu_load_1_resp_bits_error_delayed; // @[MemBlock.scala 47:26]
  wire  dcache_io_lsu_load_1_s1_kill; // @[MemBlock.scala 47:26]
  wire  dcache_io_lsu_load_1_s2_kill; // @[MemBlock.scala 47:26]
  wire [35:0] dcache_io_lsu_load_1_s1_paddr_dup_lsu; // @[MemBlock.scala 47:26]
  wire [35:0] dcache_io_lsu_load_1_s1_paddr_dup_dcache; // @[MemBlock.scala 47:26]
  wire  dcache_io_lsu_load_1_s1_bank_conflict; // @[MemBlock.scala 47:26]
  wire  dcache_io_lsu_lsq_valid; // @[MemBlock.scala 47:26]
  wire [1:0] dcache_io_lsu_lsq_bits_id; // @[MemBlock.scala 47:26]
  wire  dcache_io_lsu_store_req_ready; // @[MemBlock.scala 47:26]
  wire  dcache_io_lsu_store_req_valid; // @[MemBlock.scala 47:26]
  wire [38:0] dcache_io_lsu_store_req_bits_vaddr; // @[MemBlock.scala 47:26]
  wire [35:0] dcache_io_lsu_store_req_bits_addr; // @[MemBlock.scala 47:26]
  wire [511:0] dcache_io_lsu_store_req_bits_data; // @[MemBlock.scala 47:26]
  wire [63:0] dcache_io_lsu_store_req_bits_mask; // @[MemBlock.scala 47:26]
  wire [3:0] dcache_io_lsu_store_req_bits_id; // @[MemBlock.scala 47:26]
  wire  dcache_io_lsu_store_main_pipe_hit_resp_valid; // @[MemBlock.scala 47:26]
  wire [3:0] dcache_io_lsu_store_main_pipe_hit_resp_bits_id; // @[MemBlock.scala 47:26]
  wire  dcache_io_lsu_store_refill_hit_resp_valid; // @[MemBlock.scala 47:26]
  wire [3:0] dcache_io_lsu_store_refill_hit_resp_bits_id; // @[MemBlock.scala 47:26]
  wire  dcache_io_lsu_store_replay_resp_valid; // @[MemBlock.scala 47:26]
  wire [3:0] dcache_io_lsu_store_replay_resp_bits_id; // @[MemBlock.scala 47:26]
  wire  dcache_io_lsu_atomics_req_ready; // @[MemBlock.scala 47:26]
  wire  dcache_io_lsu_atomics_req_valid; // @[MemBlock.scala 47:26]
  wire [4:0] dcache_io_lsu_atomics_req_bits_cmd; // @[MemBlock.scala 47:26]
  wire [38:0] dcache_io_lsu_atomics_req_bits_vaddr; // @[MemBlock.scala 47:26]
  wire [35:0] dcache_io_lsu_atomics_req_bits_addr; // @[MemBlock.scala 47:26]
  wire [2:0] dcache_io_lsu_atomics_req_bits_word_idx; // @[MemBlock.scala 47:26]
  wire [63:0] dcache_io_lsu_atomics_req_bits_amo_data; // @[MemBlock.scala 47:26]
  wire [7:0] dcache_io_lsu_atomics_req_bits_amo_mask; // @[MemBlock.scala 47:26]
  wire  dcache_io_lsu_atomics_resp_valid; // @[MemBlock.scala 47:26]
  wire [63:0] dcache_io_lsu_atomics_resp_bits_data; // @[MemBlock.scala 47:26]
  wire  dcache_io_lsu_atomics_resp_bits_miss; // @[MemBlock.scala 47:26]
  wire  dcache_io_lsu_atomics_resp_bits_replay; // @[MemBlock.scala 47:26]
  wire  dcache_io_lsu_atomics_resp_bits_error; // @[MemBlock.scala 47:26]
  wire [3:0] dcache_io_lsu_atomics_resp_bits_id; // @[MemBlock.scala 47:26]
  wire  dcache_io_lsu_atomics_block_lr; // @[MemBlock.scala 47:26]
  wire  dcache_io_lsu_release_valid; // @[MemBlock.scala 47:26]
  wire [35:0] dcache_io_lsu_release_bits_paddr; // @[MemBlock.scala 47:26]
  wire  dcache_io_lsu_forward_D_0_valid; // @[MemBlock.scala 47:26]
  wire [255:0] dcache_io_lsu_forward_D_0_data; // @[MemBlock.scala 47:26]
  wire [1:0] dcache_io_lsu_forward_D_0_mshrid; // @[MemBlock.scala 47:26]
  wire  dcache_io_lsu_forward_D_0_last; // @[MemBlock.scala 47:26]
  wire  dcache_io_lsu_forward_D_1_valid; // @[MemBlock.scala 47:26]
  wire [255:0] dcache_io_lsu_forward_D_1_data; // @[MemBlock.scala 47:26]
  wire [1:0] dcache_io_lsu_forward_D_1_mshrid; // @[MemBlock.scala 47:26]
  wire  dcache_io_lsu_forward_D_1_last; // @[MemBlock.scala 47:26]
  wire  dcache_io_lsu_forward_mshr_0_valid; // @[MemBlock.scala 47:26]
  wire [1:0] dcache_io_lsu_forward_mshr_0_mshrid; // @[MemBlock.scala 47:26]
  wire [35:0] dcache_io_lsu_forward_mshr_0_paddr; // @[MemBlock.scala 47:26]
  wire  dcache_io_lsu_forward_mshr_0_forward_mshr; // @[MemBlock.scala 47:26]
  wire [7:0] dcache_io_lsu_forward_mshr_0_forwardData_0; // @[MemBlock.scala 47:26]
  wire [7:0] dcache_io_lsu_forward_mshr_0_forwardData_1; // @[MemBlock.scala 47:26]
  wire [7:0] dcache_io_lsu_forward_mshr_0_forwardData_2; // @[MemBlock.scala 47:26]
  wire [7:0] dcache_io_lsu_forward_mshr_0_forwardData_3; // @[MemBlock.scala 47:26]
  wire [7:0] dcache_io_lsu_forward_mshr_0_forwardData_4; // @[MemBlock.scala 47:26]
  wire [7:0] dcache_io_lsu_forward_mshr_0_forwardData_5; // @[MemBlock.scala 47:26]
  wire [7:0] dcache_io_lsu_forward_mshr_0_forwardData_6; // @[MemBlock.scala 47:26]
  wire [7:0] dcache_io_lsu_forward_mshr_0_forwardData_7; // @[MemBlock.scala 47:26]
  wire [7:0] dcache_io_lsu_forward_mshr_0_forwardData_8; // @[MemBlock.scala 47:26]
  wire [7:0] dcache_io_lsu_forward_mshr_0_forwardData_9; // @[MemBlock.scala 47:26]
  wire [7:0] dcache_io_lsu_forward_mshr_0_forwardData_10; // @[MemBlock.scala 47:26]
  wire [7:0] dcache_io_lsu_forward_mshr_0_forwardData_11; // @[MemBlock.scala 47:26]
  wire [7:0] dcache_io_lsu_forward_mshr_0_forwardData_12; // @[MemBlock.scala 47:26]
  wire [7:0] dcache_io_lsu_forward_mshr_0_forwardData_13; // @[MemBlock.scala 47:26]
  wire [7:0] dcache_io_lsu_forward_mshr_0_forwardData_14; // @[MemBlock.scala 47:26]
  wire [7:0] dcache_io_lsu_forward_mshr_0_forwardData_15; // @[MemBlock.scala 47:26]
  wire  dcache_io_lsu_forward_mshr_0_forward_result_valid; // @[MemBlock.scala 47:26]
  wire  dcache_io_lsu_forward_mshr_1_valid; // @[MemBlock.scala 47:26]
  wire [1:0] dcache_io_lsu_forward_mshr_1_mshrid; // @[MemBlock.scala 47:26]
  wire [35:0] dcache_io_lsu_forward_mshr_1_paddr; // @[MemBlock.scala 47:26]
  wire  dcache_io_lsu_forward_mshr_1_forward_mshr; // @[MemBlock.scala 47:26]
  wire [7:0] dcache_io_lsu_forward_mshr_1_forwardData_0; // @[MemBlock.scala 47:26]
  wire [7:0] dcache_io_lsu_forward_mshr_1_forwardData_1; // @[MemBlock.scala 47:26]
  wire [7:0] dcache_io_lsu_forward_mshr_1_forwardData_2; // @[MemBlock.scala 47:26]
  wire [7:0] dcache_io_lsu_forward_mshr_1_forwardData_3; // @[MemBlock.scala 47:26]
  wire [7:0] dcache_io_lsu_forward_mshr_1_forwardData_4; // @[MemBlock.scala 47:26]
  wire [7:0] dcache_io_lsu_forward_mshr_1_forwardData_5; // @[MemBlock.scala 47:26]
  wire [7:0] dcache_io_lsu_forward_mshr_1_forwardData_6; // @[MemBlock.scala 47:26]
  wire [7:0] dcache_io_lsu_forward_mshr_1_forwardData_7; // @[MemBlock.scala 47:26]
  wire [7:0] dcache_io_lsu_forward_mshr_1_forwardData_8; // @[MemBlock.scala 47:26]
  wire [7:0] dcache_io_lsu_forward_mshr_1_forwardData_9; // @[MemBlock.scala 47:26]
  wire [7:0] dcache_io_lsu_forward_mshr_1_forwardData_10; // @[MemBlock.scala 47:26]
  wire [7:0] dcache_io_lsu_forward_mshr_1_forwardData_11; // @[MemBlock.scala 47:26]
  wire [7:0] dcache_io_lsu_forward_mshr_1_forwardData_12; // @[MemBlock.scala 47:26]
  wire [7:0] dcache_io_lsu_forward_mshr_1_forwardData_13; // @[MemBlock.scala 47:26]
  wire [7:0] dcache_io_lsu_forward_mshr_1_forwardData_14; // @[MemBlock.scala 47:26]
  wire [7:0] dcache_io_lsu_forward_mshr_1_forwardData_15; // @[MemBlock.scala 47:26]
  wire  dcache_io_lsu_forward_mshr_1_forward_result_valid; // @[MemBlock.scala 47:26]
  wire  dcache_io_csr_distribute_csr_wvalid; // @[MemBlock.scala 47:26]
  wire [11:0] dcache_io_csr_distribute_csr_waddr; // @[MemBlock.scala 47:26]
  wire [63:0] dcache_io_csr_distribute_csr_wdata; // @[MemBlock.scala 47:26]
  wire  dcache_io_csr_update_wvalid; // @[MemBlock.scala 47:26]
  wire [11:0] dcache_io_csr_update_waddr; // @[MemBlock.scala 47:26]
  wire [63:0] dcache_io_csr_update_wdata; // @[MemBlock.scala 47:26]
  wire [35:0] dcache_io_error_paddr; // @[MemBlock.scala 47:26]
  wire  dcache_io_error_report_to_beu; // @[MemBlock.scala 47:26]
  wire [5:0] dcache_io_perf_0_value; // @[MemBlock.scala 47:26]
  wire [5:0] dcache_io_perf_1_value; // @[MemBlock.scala 47:26]
  wire [5:0] dcache_io_perf_2_value; // @[MemBlock.scala 47:26]
  wire [5:0] dcache_io_perf_3_value; // @[MemBlock.scala 47:26]
  wire [5:0] dcache_io_perf_4_value; // @[MemBlock.scala 47:26]
  wire [5:0] dcache_io_perf_5_value; // @[MemBlock.scala 47:26]
  wire [5:0] dcache_io_perf_6_value; // @[MemBlock.scala 47:26]
  wire [5:0] dcache_io_perf_7_value; // @[MemBlock.scala 47:26]
  wire [5:0] dcache_io_perf_8_value; // @[MemBlock.scala 47:26]
  wire [5:0] dcache_io_perf_9_value; // @[MemBlock.scala 47:26]
  wire [5:0] dcache_io_perf_10_value; // @[MemBlock.scala 47:26]
  wire [5:0] dcache_io_perf_11_value; // @[MemBlock.scala 47:26]
  wire [5:0] dcache_io_perf_12_value; // @[MemBlock.scala 47:26]
  wire [5:0] dcache_io_perf_13_value; // @[MemBlock.scala 47:26]
  wire [5:0] dcache_io_perf_14_value; // @[MemBlock.scala 47:26]
  wire [5:0] dcache_io_perf_15_value; // @[MemBlock.scala 47:26]
  wire [5:0] dcache_io_perf_16_value; // @[MemBlock.scala 47:26]
  wire [5:0] dcache_io_perf_17_value; // @[MemBlock.scala 47:26]
  wire [5:0] dcache_io_perf_18_value; // @[MemBlock.scala 47:26]
  wire [5:0] dcache_io_perf_19_value; // @[MemBlock.scala 47:26]
  wire [5:0] dcache_io_perf_20_value; // @[MemBlock.scala 47:26]
  wire [5:0] dcache_io_perf_21_value; // @[MemBlock.scala 47:26]
  wire [5:0] dcache_io_perf_22_value; // @[MemBlock.scala 47:26]
  wire [5:0] dcache_io_perf_23_value; // @[MemBlock.scala 47:26]
  wire [5:0] dcache_io_perf_24_value; // @[MemBlock.scala 47:26]
  wire [5:0] dcache_io_perf_25_value; // @[MemBlock.scala 47:26]
  wire [5:0] dcache_io_perf_26_value; // @[MemBlock.scala 47:26]
  wire  uncache_clock; // @[MemBlock.scala 48:27]
  wire  uncache_reset; // @[MemBlock.scala 48:27]
  wire  uncache_auto_client_out_a_ready; // @[MemBlock.scala 48:27]
  wire  uncache_auto_client_out_a_valid; // @[MemBlock.scala 48:27]
  wire [2:0] uncache_auto_client_out_a_bits_opcode; // @[MemBlock.scala 48:27]
  wire [2:0] uncache_auto_client_out_a_bits_size; // @[MemBlock.scala 48:27]
  wire [1:0] uncache_auto_client_out_a_bits_source; // @[MemBlock.scala 48:27]
  wire [35:0] uncache_auto_client_out_a_bits_address; // @[MemBlock.scala 48:27]
  wire [7:0] uncache_auto_client_out_a_bits_mask; // @[MemBlock.scala 48:27]
  wire [63:0] uncache_auto_client_out_a_bits_data; // @[MemBlock.scala 48:27]
  wire  uncache_auto_client_out_d_ready; // @[MemBlock.scala 48:27]
  wire  uncache_auto_client_out_d_valid; // @[MemBlock.scala 48:27]
  wire [2:0] uncache_auto_client_out_d_bits_opcode; // @[MemBlock.scala 48:27]
  wire [63:0] uncache_auto_client_out_d_bits_data; // @[MemBlock.scala 48:27]
  wire [7:0] uncache_io_hartId; // @[MemBlock.scala 48:27]
  wire  uncache_io_enableOutstanding; // @[MemBlock.scala 48:27]
  wire  uncache_io_flush_empty; // @[MemBlock.scala 48:27]
  wire  uncache_io_lsq_req_ready; // @[MemBlock.scala 48:27]
  wire  uncache_io_lsq_req_valid; // @[MemBlock.scala 48:27]
  wire [4:0] uncache_io_lsq_req_bits_cmd; // @[MemBlock.scala 48:27]
  wire [35:0] uncache_io_lsq_req_bits_addr; // @[MemBlock.scala 48:27]
  wire [63:0] uncache_io_lsq_req_bits_data; // @[MemBlock.scala 48:27]
  wire [7:0] uncache_io_lsq_req_bits_mask; // @[MemBlock.scala 48:27]
  wire  uncache_io_lsq_req_bits_atomic; // @[MemBlock.scala 48:27]
  wire  uncache_io_lsq_resp_valid; // @[MemBlock.scala 48:27]
  wire [63:0] uncache_io_lsq_resp_bits_data; // @[MemBlock.scala 48:27]
  wire  csrCtrl_delay_clock; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_in_icache_parity_enable; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_in_lvpred_disable; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_in_no_spec_load; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_in_storeset_wait_store; // @[Hold.scala 97:23]
  wire [4:0] csrCtrl_delay_io_in_lvpred_timeout; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_in_bp_ctrl_ubtb_enable; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_in_bp_ctrl_btb_enable; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_in_bp_ctrl_tage_enable; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_in_bp_ctrl_sc_enable; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_in_bp_ctrl_ras_enable; // @[Hold.scala 97:23]
  wire [3:0] csrCtrl_delay_io_in_sbuffer_threshold; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_in_ldld_vio_check_enable; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_in_cache_error_enable; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_in_uncache_write_outstanding_enable; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_in_fusion_enable; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_in_wfi_enable; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_in_svinval_enable; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_in_distribute_csr_wvalid; // @[Hold.scala 97:23]
  wire [11:0] csrCtrl_delay_io_in_distribute_csr_waddr; // @[Hold.scala 97:23]
  wire [63:0] csrCtrl_delay_io_in_distribute_csr_wdata; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_in_singlestep; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_in_frontend_trigger_t_valid; // @[Hold.scala 97:23]
  wire [1:0] csrCtrl_delay_io_in_frontend_trigger_t_bits_addr; // @[Hold.scala 97:23]
  wire [1:0] csrCtrl_delay_io_in_frontend_trigger_t_bits_tdata_matchType; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_in_frontend_trigger_t_bits_tdata_select; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_in_frontend_trigger_t_bits_tdata_timing; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_in_frontend_trigger_t_bits_tdata_chain; // @[Hold.scala 97:23]
  wire [63:0] csrCtrl_delay_io_in_frontend_trigger_t_bits_tdata_tdata2; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_in_mem_trigger_t_valid; // @[Hold.scala 97:23]
  wire [2:0] csrCtrl_delay_io_in_mem_trigger_t_bits_addr; // @[Hold.scala 97:23]
  wire [1:0] csrCtrl_delay_io_in_mem_trigger_t_bits_tdata_matchType; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_in_mem_trigger_t_bits_tdata_select; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_in_mem_trigger_t_bits_tdata_chain; // @[Hold.scala 97:23]
  wire [63:0] csrCtrl_delay_io_in_mem_trigger_t_bits_tdata_tdata2; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_in_trigger_enable_0; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_in_trigger_enable_1; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_in_trigger_enable_2; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_in_trigger_enable_3; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_in_trigger_enable_4; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_in_trigger_enable_5; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_in_trigger_enable_6; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_in_trigger_enable_7; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_in_trigger_enable_8; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_in_trigger_enable_9; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_out_icache_parity_enable; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_out_lvpred_disable; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_out_no_spec_load; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_out_storeset_wait_store; // @[Hold.scala 97:23]
  wire [4:0] csrCtrl_delay_io_out_lvpred_timeout; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_out_bp_ctrl_ubtb_enable; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_out_bp_ctrl_btb_enable; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_out_bp_ctrl_tage_enable; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_out_bp_ctrl_sc_enable; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_out_bp_ctrl_ras_enable; // @[Hold.scala 97:23]
  wire [3:0] csrCtrl_delay_io_out_sbuffer_threshold; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_out_ldld_vio_check_enable; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_out_cache_error_enable; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_out_uncache_write_outstanding_enable; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_out_fusion_enable; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_out_wfi_enable; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_out_svinval_enable; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_out_distribute_csr_wvalid; // @[Hold.scala 97:23]
  wire [11:0] csrCtrl_delay_io_out_distribute_csr_waddr; // @[Hold.scala 97:23]
  wire [63:0] csrCtrl_delay_io_out_distribute_csr_wdata; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_out_singlestep; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_out_frontend_trigger_t_valid; // @[Hold.scala 97:23]
  wire [1:0] csrCtrl_delay_io_out_frontend_trigger_t_bits_addr; // @[Hold.scala 97:23]
  wire [1:0] csrCtrl_delay_io_out_frontend_trigger_t_bits_tdata_matchType; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_out_frontend_trigger_t_bits_tdata_select; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_out_frontend_trigger_t_bits_tdata_timing; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_out_frontend_trigger_t_bits_tdata_chain; // @[Hold.scala 97:23]
  wire [63:0] csrCtrl_delay_io_out_frontend_trigger_t_bits_tdata_tdata2; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_out_mem_trigger_t_valid; // @[Hold.scala 97:23]
  wire [2:0] csrCtrl_delay_io_out_mem_trigger_t_bits_addr; // @[Hold.scala 97:23]
  wire [1:0] csrCtrl_delay_io_out_mem_trigger_t_bits_tdata_matchType; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_out_mem_trigger_t_bits_tdata_select; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_out_mem_trigger_t_bits_tdata_chain; // @[Hold.scala 97:23]
  wire [63:0] csrCtrl_delay_io_out_mem_trigger_t_bits_tdata_tdata2; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_out_trigger_enable_0; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_out_trigger_enable_1; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_out_trigger_enable_2; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_out_trigger_enable_3; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_out_trigger_enable_4; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_out_trigger_enable_5; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_out_trigger_enable_6; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_out_trigger_enable_7; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_out_trigger_enable_8; // @[Hold.scala 97:23]
  wire  csrCtrl_delay_io_out_trigger_enable_9; // @[Hold.scala 97:23]
  wire  LoadUnit_0_clock; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_reset; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_loadIn_ready; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_loadIn_valid; // @[MemBlock.scala 139:56]
  wire [9:0] LoadUnit_0_io_loadIn_bits_uop_cf_foldpc; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_loadIn_bits_uop_cf_trigger_backendEn_1; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_loadIn_bits_uop_cf_waitForRobIdx_flag; // @[MemBlock.scala 139:56]
  wire [4:0] LoadUnit_0_io_loadIn_bits_uop_cf_waitForRobIdx_value; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_loadIn_bits_uop_cf_loadWaitBit; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_loadIn_bits_uop_cf_loadWaitStrict; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_loadIn_bits_uop_cf_ftqPtr_flag; // @[MemBlock.scala 139:56]
  wire [2:0] LoadUnit_0_io_loadIn_bits_uop_cf_ftqPtr_value; // @[MemBlock.scala 139:56]
  wire [2:0] LoadUnit_0_io_loadIn_bits_uop_cf_ftqOffset; // @[MemBlock.scala 139:56]
  wire [3:0] LoadUnit_0_io_loadIn_bits_uop_ctrl_fuType; // @[MemBlock.scala 139:56]
  wire [6:0] LoadUnit_0_io_loadIn_bits_uop_ctrl_fuOpType; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_loadIn_bits_uop_ctrl_rfWen; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_loadIn_bits_uop_ctrl_fpWen; // @[MemBlock.scala 139:56]
  wire [19:0] LoadUnit_0_io_loadIn_bits_uop_ctrl_imm; // @[MemBlock.scala 139:56]
  wire [5:0] LoadUnit_0_io_loadIn_bits_uop_pdest; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_loadIn_bits_uop_robIdx_flag; // @[MemBlock.scala 139:56]
  wire [4:0] LoadUnit_0_io_loadIn_bits_uop_robIdx_value; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_loadIn_bits_uop_lqIdx_flag; // @[MemBlock.scala 139:56]
  wire [3:0] LoadUnit_0_io_loadIn_bits_uop_lqIdx_value; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_loadIn_bits_uop_sqIdx_flag; // @[MemBlock.scala 139:56]
  wire [3:0] LoadUnit_0_io_loadIn_bits_uop_sqIdx_value; // @[MemBlock.scala 139:56]
  wire [63:0] LoadUnit_0_io_loadIn_bits_src_0; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_VecloadIn_ready; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_VecloadIn_valid; // @[MemBlock.scala 139:56]
  wire [38:0] LoadUnit_0_io_VecloadIn_bits_vaddr; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_loadOut_valid; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_loadOut_bits_uop_cf_exceptionVec_4; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_loadOut_bits_uop_cf_exceptionVec_5; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_loadOut_bits_uop_cf_exceptionVec_13; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_loadOut_bits_uop_cf_trigger_backendEn_1; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_loadOut_bits_uop_cf_trigger_backendHit_0; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_loadOut_bits_uop_cf_trigger_backendHit_1; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_loadOut_bits_uop_cf_trigger_backendHit_4; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_loadOut_bits_uop_ctrl_rfWen; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_loadOut_bits_uop_ctrl_fpWen; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_loadOut_bits_uop_ctrl_flushPipe; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_loadOut_bits_uop_ctrl_replayInst; // @[MemBlock.scala 139:56]
  wire [5:0] LoadUnit_0_io_loadOut_bits_uop_pdest; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_loadOut_bits_uop_robIdx_flag; // @[MemBlock.scala 139:56]
  wire [4:0] LoadUnit_0_io_loadOut_bits_uop_robIdx_value; // @[MemBlock.scala 139:56]
  wire [63:0] LoadUnit_0_io_loadOut_bits_data; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_loadOut_bits_debug_isMMIO; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_redirect_valid; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_redirect_bits_robIdx_flag; // @[MemBlock.scala 139:56]
  wire [4:0] LoadUnit_0_io_redirect_bits_robIdx_value; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_redirect_bits_level; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_dcache_req_ready; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_dcache_req_valid; // @[MemBlock.scala 139:56]
  wire [4:0] LoadUnit_0_io_dcache_req_bits_cmd; // @[MemBlock.scala 139:56]
  wire [35:0] LoadUnit_0_io_dcache_req_bits_addr; // @[MemBlock.scala 139:56]
  wire [3:0] LoadUnit_0_io_dcache_req_bits_instrtype; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_0_io_dcache_req_bits_replayCarry_real_way_en; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_dcache_req_bits_replayCarry_valid; // @[MemBlock.scala 139:56]
  wire [127:0] LoadUnit_0_io_dcache_resp_bits_data_delayed; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_dcache_resp_bits_miss; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_dcache_resp_bits_replay; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_0_io_dcache_resp_bits_replayCarry_real_way_en; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_dcache_resp_bits_replayCarry_valid; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_dcache_resp_bits_tag_error; // @[MemBlock.scala 139:56]
  wire [1:0] LoadUnit_0_io_dcache_resp_bits_mshr_id; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_dcache_resp_bits_error_delayed; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_dcache_s1_kill; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_dcache_s2_kill; // @[MemBlock.scala 139:56]
  wire [35:0] LoadUnit_0_io_dcache_s1_paddr_dup_lsu; // @[MemBlock.scala 139:56]
  wire [35:0] LoadUnit_0_io_dcache_s1_paddr_dup_dcache; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_dcache_s1_bank_conflict; // @[MemBlock.scala 139:56]
  wire [38:0] LoadUnit_0_io_sbuffer_vaddr; // @[MemBlock.scala 139:56]
  wire [35:0] LoadUnit_0_io_sbuffer_paddr; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_sbuffer_valid; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_sbuffer_forwardMask_0; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_sbuffer_forwardMask_1; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_sbuffer_forwardMask_2; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_sbuffer_forwardMask_3; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_sbuffer_forwardMask_4; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_sbuffer_forwardMask_5; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_sbuffer_forwardMask_6; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_sbuffer_forwardMask_7; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_sbuffer_forwardMask_8; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_sbuffer_forwardMask_9; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_sbuffer_forwardMask_10; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_sbuffer_forwardMask_11; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_sbuffer_forwardMask_12; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_sbuffer_forwardMask_13; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_sbuffer_forwardMask_14; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_sbuffer_forwardMask_15; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_0_io_sbuffer_forwardData_0; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_0_io_sbuffer_forwardData_1; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_0_io_sbuffer_forwardData_2; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_0_io_sbuffer_forwardData_3; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_0_io_sbuffer_forwardData_4; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_0_io_sbuffer_forwardData_5; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_0_io_sbuffer_forwardData_6; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_0_io_sbuffer_forwardData_7; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_0_io_sbuffer_forwardData_8; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_0_io_sbuffer_forwardData_9; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_0_io_sbuffer_forwardData_10; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_0_io_sbuffer_forwardData_11; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_0_io_sbuffer_forwardData_12; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_0_io_sbuffer_forwardData_13; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_0_io_sbuffer_forwardData_14; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_0_io_sbuffer_forwardData_15; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_sbuffer_matchInvalid; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_loadIn_valid; // @[MemBlock.scala 139:56]
  wire [9:0] LoadUnit_0_io_lsq_loadIn_bits_uop_cf_foldpc; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_loadIn_bits_uop_cf_exceptionVec_4; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_loadIn_bits_uop_cf_exceptionVec_5; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_loadIn_bits_uop_cf_exceptionVec_13; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_loadIn_bits_uop_cf_trigger_backendEn_1; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_loadIn_bits_uop_cf_trigger_backendHit_0; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_loadIn_bits_uop_cf_trigger_backendHit_1; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_loadIn_bits_uop_cf_trigger_backendHit_4; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_loadIn_bits_uop_cf_waitForRobIdx_flag; // @[MemBlock.scala 139:56]
  wire [4:0] LoadUnit_0_io_lsq_loadIn_bits_uop_cf_waitForRobIdx_value; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_loadIn_bits_uop_cf_loadWaitBit; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_loadIn_bits_uop_cf_loadWaitStrict; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_loadIn_bits_uop_cf_ftqPtr_flag; // @[MemBlock.scala 139:56]
  wire [2:0] LoadUnit_0_io_lsq_loadIn_bits_uop_cf_ftqPtr_value; // @[MemBlock.scala 139:56]
  wire [2:0] LoadUnit_0_io_lsq_loadIn_bits_uop_cf_ftqOffset; // @[MemBlock.scala 139:56]
  wire [3:0] LoadUnit_0_io_lsq_loadIn_bits_uop_ctrl_fuType; // @[MemBlock.scala 139:56]
  wire [6:0] LoadUnit_0_io_lsq_loadIn_bits_uop_ctrl_fuOpType; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_loadIn_bits_uop_ctrl_rfWen; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_loadIn_bits_uop_ctrl_fpWen; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_loadIn_bits_uop_ctrl_replayInst; // @[MemBlock.scala 139:56]
  wire [5:0] LoadUnit_0_io_lsq_loadIn_bits_uop_pdest; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_loadIn_bits_uop_robIdx_flag; // @[MemBlock.scala 139:56]
  wire [4:0] LoadUnit_0_io_lsq_loadIn_bits_uop_robIdx_value; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_loadIn_bits_uop_lqIdx_flag; // @[MemBlock.scala 139:56]
  wire [3:0] LoadUnit_0_io_lsq_loadIn_bits_uop_lqIdx_value; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_loadIn_bits_uop_sqIdx_flag; // @[MemBlock.scala 139:56]
  wire [3:0] LoadUnit_0_io_lsq_loadIn_bits_uop_sqIdx_value; // @[MemBlock.scala 139:56]
  wire [38:0] LoadUnit_0_io_lsq_loadIn_bits_vaddr; // @[MemBlock.scala 139:56]
  wire [35:0] LoadUnit_0_io_lsq_loadIn_bits_paddr; // @[MemBlock.scala 139:56]
  wire [15:0] LoadUnit_0_io_lsq_loadIn_bits_mask; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_loadIn_bits_miss; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_loadIn_bits_tlbMiss; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_loadIn_bits_mmio; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_loadIn_bits_rarAllocated; // @[MemBlock.scala 139:56]
  wire [3:0] LoadUnit_0_io_lsq_loadIn_bits_rarIndex; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_loadIn_bits_rawAllocated; // @[MemBlock.scala 139:56]
  wire [2:0] LoadUnit_0_io_lsq_loadIn_bits_rawIndex; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_loadIn_bits_canAccept; // @[MemBlock.scala 139:56]
  wire [1:0] LoadUnit_0_io_lsq_loadIn_bits_replayInfo_missMSHRId; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_loadIn_bits_replayInfo_canForwardFullData; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_loadIn_bits_replayInfo_dataInvalidSqIdx_flag; // @[MemBlock.scala 139:56]
  wire [3:0] LoadUnit_0_io_lsq_loadIn_bits_replayInfo_dataInvalidSqIdx_value; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_loadIn_bits_replayInfo_addrInvalidSqIdx_flag; // @[MemBlock.scala 139:56]
  wire [3:0] LoadUnit_0_io_lsq_loadIn_bits_replayInfo_addrInvalidSqIdx_value; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_0_io_lsq_loadIn_bits_replayInfo_replayCarry_real_way_en; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_loadIn_bits_replayInfo_replayCarry_valid; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_loadIn_bits_replayInfo_dataInLastBeat; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_loadIn_bits_replayInfo_cause_0; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_loadIn_bits_replayInfo_cause_1; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_loadIn_bits_replayInfo_cause_2; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_loadIn_bits_replayInfo_cause_3; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_loadIn_bits_replayInfo_cause_4; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_loadIn_bits_replayInfo_cause_5; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_loadIn_bits_replayInfo_cause_6; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_loadIn_bits_replayInfo_cause_7; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_loadIn_bits_lqDataWenDup_1; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_loadIn_bits_lqDataWenDup_2; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_loadIn_bits_lqDataWenDup_3; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_loadIn_bits_lqDataWenDup_5; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_loadOut_ready; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_loadOut_valid; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_loadOut_bits_uop_cf_exceptionVec_4; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_loadOut_bits_uop_cf_exceptionVec_5; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_loadOut_bits_uop_cf_exceptionVec_13; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_loadOut_bits_uop_cf_trigger_backendEn_1; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_loadOut_bits_uop_cf_trigger_backendHit_0; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_loadOut_bits_uop_cf_trigger_backendHit_1; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_loadOut_bits_uop_cf_trigger_backendHit_4; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_loadOut_bits_uop_ctrl_rfWen; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_loadOut_bits_uop_ctrl_fpWen; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_loadOut_bits_uop_ctrl_flushPipe; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_loadOut_bits_uop_ctrl_replayInst; // @[MemBlock.scala 139:56]
  wire [5:0] LoadUnit_0_io_lsq_loadOut_bits_uop_pdest; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_loadOut_bits_uop_robIdx_flag; // @[MemBlock.scala 139:56]
  wire [4:0] LoadUnit_0_io_lsq_loadOut_bits_uop_robIdx_value; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_loadOut_bits_debug_isMMIO; // @[MemBlock.scala 139:56]
  wire [63:0] LoadUnit_0_io_lsq_ldRawData_lqData; // @[MemBlock.scala 139:56]
  wire [6:0] LoadUnit_0_io_lsq_ldRawData_uop_ctrl_fuOpType; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_ldRawData_uop_ctrl_fpWen; // @[MemBlock.scala 139:56]
  wire [2:0] LoadUnit_0_io_lsq_ldRawData_addrOffset; // @[MemBlock.scala 139:56]
  wire [38:0] LoadUnit_0_io_lsq_forward_vaddr; // @[MemBlock.scala 139:56]
  wire [35:0] LoadUnit_0_io_lsq_forward_paddr; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_forward_uop_cf_waitForRobIdx_flag; // @[MemBlock.scala 139:56]
  wire [4:0] LoadUnit_0_io_lsq_forward_uop_cf_waitForRobIdx_value; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_forward_uop_sqIdx_flag; // @[MemBlock.scala 139:56]
  wire [3:0] LoadUnit_0_io_lsq_forward_uop_sqIdx_value; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_forward_valid; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_forward_forwardMask_0; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_forward_forwardMask_1; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_forward_forwardMask_2; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_forward_forwardMask_3; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_forward_forwardMask_4; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_forward_forwardMask_5; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_forward_forwardMask_6; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_forward_forwardMask_7; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_forward_forwardMask_8; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_forward_forwardMask_9; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_forward_forwardMask_10; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_forward_forwardMask_11; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_forward_forwardMask_12; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_forward_forwardMask_13; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_forward_forwardMask_14; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_forward_forwardMask_15; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_0_io_lsq_forward_forwardData_0; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_0_io_lsq_forward_forwardData_1; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_0_io_lsq_forward_forwardData_2; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_0_io_lsq_forward_forwardData_3; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_0_io_lsq_forward_forwardData_4; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_0_io_lsq_forward_forwardData_5; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_0_io_lsq_forward_forwardData_6; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_0_io_lsq_forward_forwardData_7; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_0_io_lsq_forward_forwardData_8; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_0_io_lsq_forward_forwardData_9; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_0_io_lsq_forward_forwardData_10; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_0_io_lsq_forward_forwardData_11; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_0_io_lsq_forward_forwardData_12; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_0_io_lsq_forward_forwardData_13; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_0_io_lsq_forward_forwardData_14; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_0_io_lsq_forward_forwardData_15; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_forward_sqIdx_flag; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_forward_dataInvalid; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_forward_matchInvalid; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_forward_schedWait; // @[MemBlock.scala 139:56]
  wire [11:0] LoadUnit_0_io_lsq_forward_sqIdxMask; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_forward_dataInvalidSqIdx_flag; // @[MemBlock.scala 139:56]
  wire [3:0] LoadUnit_0_io_lsq_forward_dataInvalidSqIdx_value; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_forward_addrInvalidSqIdx_flag; // @[MemBlock.scala 139:56]
  wire [3:0] LoadUnit_0_io_lsq_forward_addrInvalidSqIdx_value; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_storeLoadViolationQuery_req_valid; // @[MemBlock.scala 139:56]
  wire [9:0] LoadUnit_0_io_lsq_storeLoadViolationQuery_req_bits_uop_cf_foldpc; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_storeLoadViolationQuery_req_bits_uop_cf_ftqPtr_flag; // @[MemBlock.scala 139:56]
  wire [2:0] LoadUnit_0_io_lsq_storeLoadViolationQuery_req_bits_uop_cf_ftqPtr_value; // @[MemBlock.scala 139:56]
  wire [2:0] LoadUnit_0_io_lsq_storeLoadViolationQuery_req_bits_uop_cf_ftqOffset; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_storeLoadViolationQuery_req_bits_uop_robIdx_flag; // @[MemBlock.scala 139:56]
  wire [4:0] LoadUnit_0_io_lsq_storeLoadViolationQuery_req_bits_uop_robIdx_value; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_storeLoadViolationQuery_req_bits_uop_sqIdx_flag; // @[MemBlock.scala 139:56]
  wire [3:0] LoadUnit_0_io_lsq_storeLoadViolationQuery_req_bits_uop_sqIdx_value; // @[MemBlock.scala 139:56]
  wire [2:0] LoadUnit_0_io_lsq_storeLoadViolationQuery_req_bits_index; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_storeLoadViolationQuery_req_bits_allocated; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_storeLoadViolationQuery_req_bits_datavalid; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_0_io_lsq_storeLoadViolationQuery_req_bits_mask; // @[MemBlock.scala 139:56]
  wire [35:0] LoadUnit_0_io_lsq_storeLoadViolationQuery_req_bits_paddr; // @[MemBlock.scala 139:56]
  wire [2:0] LoadUnit_0_io_lsq_storeLoadViolationQuery_resp_bits_index; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_storeLoadViolationQuery_resp_bits_canAccept; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_storeLoadViolationQuery_resp_bits_allocated; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_loadLoadViolationQuery_req_valid; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_loadLoadViolationQuery_req_bits_uop_robIdx_flag; // @[MemBlock.scala 139:56]
  wire [4:0] LoadUnit_0_io_lsq_loadLoadViolationQuery_req_bits_uop_robIdx_value; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_loadLoadViolationQuery_req_bits_uop_lqIdx_flag; // @[MemBlock.scala 139:56]
  wire [3:0] LoadUnit_0_io_lsq_loadLoadViolationQuery_req_bits_uop_lqIdx_value; // @[MemBlock.scala 139:56]
  wire [3:0] LoadUnit_0_io_lsq_loadLoadViolationQuery_req_bits_index; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_loadLoadViolationQuery_req_bits_allocated; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_loadLoadViolationQuery_req_bits_datavalid; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_loadLoadViolationQuery_req_bits_miss; // @[MemBlock.scala 139:56]
  wire [35:0] LoadUnit_0_io_lsq_loadLoadViolationQuery_req_bits_paddr; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_loadLoadViolationQuery_resp_valid; // @[MemBlock.scala 139:56]
  wire [3:0] LoadUnit_0_io_lsq_loadLoadViolationQuery_resp_bits_index; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_loadLoadViolationQuery_resp_bits_canAccept; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_loadLoadViolationQuery_resp_bits_allocated; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_loadLoadViolationQuery_resp_bits_replayFromFetch; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_trigger_hitLoadAddrTriggerHitVec_0; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_trigger_hitLoadAddrTriggerHitVec_1; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_trigger_hitLoadAddrTriggerHitVec_2; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_trigger_lqLoadAddrTriggerHitVec_0; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_trigger_lqLoadAddrTriggerHitVec_1; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lsq_trigger_lqLoadAddrTriggerHitVec_2; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_tlDchannel_valid; // @[MemBlock.scala 139:56]
  wire [255:0] LoadUnit_0_io_tlDchannel_data; // @[MemBlock.scala 139:56]
  wire [1:0] LoadUnit_0_io_tlDchannel_mshrid; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_tlDchannel_last; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_forward_mshr_valid; // @[MemBlock.scala 139:56]
  wire [1:0] LoadUnit_0_io_forward_mshr_mshrid; // @[MemBlock.scala 139:56]
  wire [35:0] LoadUnit_0_io_forward_mshr_paddr; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_forward_mshr_forward_mshr; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_0_io_forward_mshr_forwardData_0; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_0_io_forward_mshr_forwardData_1; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_0_io_forward_mshr_forwardData_2; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_0_io_forward_mshr_forwardData_3; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_0_io_forward_mshr_forwardData_4; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_0_io_forward_mshr_forwardData_5; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_0_io_forward_mshr_forwardData_6; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_0_io_forward_mshr_forwardData_7; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_0_io_forward_mshr_forwardData_8; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_0_io_forward_mshr_forwardData_9; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_0_io_forward_mshr_forwardData_10; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_0_io_forward_mshr_forwardData_11; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_0_io_forward_mshr_forwardData_12; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_0_io_forward_mshr_forwardData_13; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_0_io_forward_mshr_forwardData_14; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_0_io_forward_mshr_forwardData_15; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_forward_mshr_forward_result_valid; // @[MemBlock.scala 139:56]
  wire [63:0] LoadUnit_0_io_trigger_0_tdata2; // @[MemBlock.scala 139:56]
  wire [1:0] LoadUnit_0_io_trigger_0_matchType; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_trigger_0_tEnable; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_trigger_0_addrHit; // @[MemBlock.scala 139:56]
  wire [63:0] LoadUnit_0_io_trigger_1_tdata2; // @[MemBlock.scala 139:56]
  wire [1:0] LoadUnit_0_io_trigger_1_matchType; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_trigger_1_tEnable; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_trigger_1_addrHit; // @[MemBlock.scala 139:56]
  wire [63:0] LoadUnit_0_io_trigger_2_tdata2; // @[MemBlock.scala 139:56]
  wire [1:0] LoadUnit_0_io_trigger_2_matchType; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_trigger_2_tEnable; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_trigger_2_addrHit; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_tlb_req_valid; // @[MemBlock.scala 139:56]
  wire [38:0] LoadUnit_0_io_tlb_req_bits_vaddr; // @[MemBlock.scala 139:56]
  wire [2:0] LoadUnit_0_io_tlb_req_bits_cmd; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_tlb_req_bits_no_translate; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_tlb_req_kill; // @[MemBlock.scala 139:56]
  wire [35:0] LoadUnit_0_io_tlb_resp_bits_paddr_0; // @[MemBlock.scala 139:56]
  wire [35:0] LoadUnit_0_io_tlb_resp_bits_paddr_1; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_tlb_resp_bits_miss; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_tlb_resp_bits_excp_0_pf_ld; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_tlb_resp_bits_excp_0_af_ld; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_tlb_resp_bits_static_pm_valid; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_tlb_resp_bits_static_pm_bits; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_pmp_ld; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_pmp_mmio; // @[MemBlock.scala 139:56]
  wire [63:0] LoadUnit_0_io_fastpathOut_data; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_fastpathOut_valid; // @[MemBlock.scala 139:56]
  wire [63:0] LoadUnit_0_io_fastpathIn_data; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_fastpathIn_valid; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_loadFastMatch; // @[MemBlock.scala 139:56]
  wire [11:0] LoadUnit_0_io_loadFastImm; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_csrCtrl_ldld_vio_check_enable; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_csrCtrl_cache_error_enable; // @[MemBlock.scala 139:56]
  wire [9:0] LoadUnit_0_io_correctTableQuery_req_addr; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_correctTableQuery_resp_strict; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_correctTableUpdate_valid; // @[MemBlock.scala 139:56]
  wire [9:0] LoadUnit_0_io_correctTableUpdate_bits_addr; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_correctTableUpdate_bits_strict; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_correctTableUpdate_bits_violation; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_reExecuteQuery_0_valid; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_reExecuteQuery_0_bits_robIdx_flag; // @[MemBlock.scala 139:56]
  wire [4:0] LoadUnit_0_io_reExecuteQuery_0_bits_robIdx_value; // @[MemBlock.scala 139:56]
  wire [35:0] LoadUnit_0_io_reExecuteQuery_0_bits_paddr; // @[MemBlock.scala 139:56]
  wire [15:0] LoadUnit_0_io_reExecuteQuery_0_bits_mask; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_reExecuteQuery_1_valid; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_reExecuteQuery_1_bits_robIdx_flag; // @[MemBlock.scala 139:56]
  wire [4:0] LoadUnit_0_io_reExecuteQuery_1_bits_robIdx_value; // @[MemBlock.scala 139:56]
  wire [35:0] LoadUnit_0_io_reExecuteQuery_1_bits_paddr; // @[MemBlock.scala 139:56]
  wire [15:0] LoadUnit_0_io_reExecuteQuery_1_bits_mask; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_replay_ready; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_replay_valid; // @[MemBlock.scala 139:56]
  wire [9:0] LoadUnit_0_io_replay_bits_uop_cf_foldpc; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_replay_bits_uop_cf_trigger_backendEn_1; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_replay_bits_uop_cf_trigger_backendHit_0; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_replay_bits_uop_cf_trigger_backendHit_1; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_replay_bits_uop_cf_trigger_backendHit_4; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_replay_bits_uop_cf_waitForRobIdx_flag; // @[MemBlock.scala 139:56]
  wire [4:0] LoadUnit_0_io_replay_bits_uop_cf_waitForRobIdx_value; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_replay_bits_uop_cf_loadWaitBit; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_replay_bits_uop_cf_loadWaitStrict; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_replay_bits_uop_cf_ftqPtr_flag; // @[MemBlock.scala 139:56]
  wire [2:0] LoadUnit_0_io_replay_bits_uop_cf_ftqPtr_value; // @[MemBlock.scala 139:56]
  wire [2:0] LoadUnit_0_io_replay_bits_uop_cf_ftqOffset; // @[MemBlock.scala 139:56]
  wire [3:0] LoadUnit_0_io_replay_bits_uop_ctrl_fuType; // @[MemBlock.scala 139:56]
  wire [6:0] LoadUnit_0_io_replay_bits_uop_ctrl_fuOpType; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_replay_bits_uop_ctrl_rfWen; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_replay_bits_uop_ctrl_fpWen; // @[MemBlock.scala 139:56]
  wire [5:0] LoadUnit_0_io_replay_bits_uop_pdest; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_replay_bits_uop_robIdx_flag; // @[MemBlock.scala 139:56]
  wire [4:0] LoadUnit_0_io_replay_bits_uop_robIdx_value; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_replay_bits_uop_lqIdx_flag; // @[MemBlock.scala 139:56]
  wire [3:0] LoadUnit_0_io_replay_bits_uop_lqIdx_value; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_replay_bits_uop_sqIdx_flag; // @[MemBlock.scala 139:56]
  wire [3:0] LoadUnit_0_io_replay_bits_uop_sqIdx_value; // @[MemBlock.scala 139:56]
  wire [38:0] LoadUnit_0_io_replay_bits_vaddr; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_replay_bits_isFirstIssue; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_0_io_replay_bits_replayCarry_real_way_en; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_replay_bits_replayCarry_valid; // @[MemBlock.scala 139:56]
  wire [1:0] LoadUnit_0_io_replay_bits_mshrid; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_replay_bits_forward_tlDchannel; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_replay_bits_rarAllocated; // @[MemBlock.scala 139:56]
  wire [3:0] LoadUnit_0_io_replay_bits_rarIndex; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_replay_bits_rawAllocated; // @[MemBlock.scala 139:56]
  wire [2:0] LoadUnit_0_io_replay_bits_rawIndex; // @[MemBlock.scala 139:56]
  wire  LoadUnit_0_io_lqReplayFull; // @[MemBlock.scala 139:56]
  wire [5:0] LoadUnit_0_io_perf_0_value; // @[MemBlock.scala 139:56]
  wire [5:0] LoadUnit_0_io_perf_1_value; // @[MemBlock.scala 139:56]
  wire [5:0] LoadUnit_0_io_perf_2_value; // @[MemBlock.scala 139:56]
  wire [5:0] LoadUnit_0_io_perf_3_value; // @[MemBlock.scala 139:56]
  wire [5:0] LoadUnit_0_io_perf_4_value; // @[MemBlock.scala 139:56]
  wire [5:0] LoadUnit_0_io_perf_5_value; // @[MemBlock.scala 139:56]
  wire [5:0] LoadUnit_0_io_perf_6_value; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_clock; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_reset; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_loadIn_ready; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_loadIn_valid; // @[MemBlock.scala 139:56]
  wire [9:0] LoadUnit_1_io_loadIn_bits_uop_cf_foldpc; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_loadIn_bits_uop_cf_trigger_backendEn_1; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_loadIn_bits_uop_cf_waitForRobIdx_flag; // @[MemBlock.scala 139:56]
  wire [4:0] LoadUnit_1_io_loadIn_bits_uop_cf_waitForRobIdx_value; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_loadIn_bits_uop_cf_loadWaitBit; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_loadIn_bits_uop_cf_loadWaitStrict; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_loadIn_bits_uop_cf_ftqPtr_flag; // @[MemBlock.scala 139:56]
  wire [2:0] LoadUnit_1_io_loadIn_bits_uop_cf_ftqPtr_value; // @[MemBlock.scala 139:56]
  wire [2:0] LoadUnit_1_io_loadIn_bits_uop_cf_ftqOffset; // @[MemBlock.scala 139:56]
  wire [3:0] LoadUnit_1_io_loadIn_bits_uop_ctrl_fuType; // @[MemBlock.scala 139:56]
  wire [6:0] LoadUnit_1_io_loadIn_bits_uop_ctrl_fuOpType; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_loadIn_bits_uop_ctrl_rfWen; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_loadIn_bits_uop_ctrl_fpWen; // @[MemBlock.scala 139:56]
  wire [19:0] LoadUnit_1_io_loadIn_bits_uop_ctrl_imm; // @[MemBlock.scala 139:56]
  wire [5:0] LoadUnit_1_io_loadIn_bits_uop_pdest; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_loadIn_bits_uop_robIdx_flag; // @[MemBlock.scala 139:56]
  wire [4:0] LoadUnit_1_io_loadIn_bits_uop_robIdx_value; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_loadIn_bits_uop_lqIdx_flag; // @[MemBlock.scala 139:56]
  wire [3:0] LoadUnit_1_io_loadIn_bits_uop_lqIdx_value; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_loadIn_bits_uop_sqIdx_flag; // @[MemBlock.scala 139:56]
  wire [3:0] LoadUnit_1_io_loadIn_bits_uop_sqIdx_value; // @[MemBlock.scala 139:56]
  wire [63:0] LoadUnit_1_io_loadIn_bits_src_0; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_VecloadIn_ready; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_VecloadIn_valid; // @[MemBlock.scala 139:56]
  wire [38:0] LoadUnit_1_io_VecloadIn_bits_vaddr; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_loadOut_valid; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_loadOut_bits_uop_cf_exceptionVec_4; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_loadOut_bits_uop_cf_exceptionVec_5; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_loadOut_bits_uop_cf_exceptionVec_13; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_loadOut_bits_uop_cf_trigger_backendEn_1; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_loadOut_bits_uop_cf_trigger_backendHit_0; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_loadOut_bits_uop_cf_trigger_backendHit_1; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_loadOut_bits_uop_cf_trigger_backendHit_4; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_loadOut_bits_uop_ctrl_rfWen; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_loadOut_bits_uop_ctrl_fpWen; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_loadOut_bits_uop_ctrl_flushPipe; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_loadOut_bits_uop_ctrl_replayInst; // @[MemBlock.scala 139:56]
  wire [5:0] LoadUnit_1_io_loadOut_bits_uop_pdest; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_loadOut_bits_uop_robIdx_flag; // @[MemBlock.scala 139:56]
  wire [4:0] LoadUnit_1_io_loadOut_bits_uop_robIdx_value; // @[MemBlock.scala 139:56]
  wire [63:0] LoadUnit_1_io_loadOut_bits_data; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_loadOut_bits_debug_isMMIO; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_redirect_valid; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_redirect_bits_robIdx_flag; // @[MemBlock.scala 139:56]
  wire [4:0] LoadUnit_1_io_redirect_bits_robIdx_value; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_redirect_bits_level; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_dcache_req_ready; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_dcache_req_valid; // @[MemBlock.scala 139:56]
  wire [4:0] LoadUnit_1_io_dcache_req_bits_cmd; // @[MemBlock.scala 139:56]
  wire [35:0] LoadUnit_1_io_dcache_req_bits_addr; // @[MemBlock.scala 139:56]
  wire [3:0] LoadUnit_1_io_dcache_req_bits_instrtype; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_1_io_dcache_req_bits_replayCarry_real_way_en; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_dcache_req_bits_replayCarry_valid; // @[MemBlock.scala 139:56]
  wire [127:0] LoadUnit_1_io_dcache_resp_bits_data_delayed; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_dcache_resp_bits_miss; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_dcache_resp_bits_replay; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_1_io_dcache_resp_bits_replayCarry_real_way_en; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_dcache_resp_bits_replayCarry_valid; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_dcache_resp_bits_tag_error; // @[MemBlock.scala 139:56]
  wire [1:0] LoadUnit_1_io_dcache_resp_bits_mshr_id; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_dcache_resp_bits_error_delayed; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_dcache_s1_kill; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_dcache_s2_kill; // @[MemBlock.scala 139:56]
  wire [35:0] LoadUnit_1_io_dcache_s1_paddr_dup_lsu; // @[MemBlock.scala 139:56]
  wire [35:0] LoadUnit_1_io_dcache_s1_paddr_dup_dcache; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_dcache_s1_bank_conflict; // @[MemBlock.scala 139:56]
  wire [38:0] LoadUnit_1_io_sbuffer_vaddr; // @[MemBlock.scala 139:56]
  wire [35:0] LoadUnit_1_io_sbuffer_paddr; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_sbuffer_valid; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_sbuffer_forwardMask_0; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_sbuffer_forwardMask_1; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_sbuffer_forwardMask_2; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_sbuffer_forwardMask_3; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_sbuffer_forwardMask_4; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_sbuffer_forwardMask_5; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_sbuffer_forwardMask_6; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_sbuffer_forwardMask_7; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_sbuffer_forwardMask_8; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_sbuffer_forwardMask_9; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_sbuffer_forwardMask_10; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_sbuffer_forwardMask_11; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_sbuffer_forwardMask_12; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_sbuffer_forwardMask_13; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_sbuffer_forwardMask_14; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_sbuffer_forwardMask_15; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_1_io_sbuffer_forwardData_0; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_1_io_sbuffer_forwardData_1; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_1_io_sbuffer_forwardData_2; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_1_io_sbuffer_forwardData_3; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_1_io_sbuffer_forwardData_4; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_1_io_sbuffer_forwardData_5; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_1_io_sbuffer_forwardData_6; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_1_io_sbuffer_forwardData_7; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_1_io_sbuffer_forwardData_8; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_1_io_sbuffer_forwardData_9; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_1_io_sbuffer_forwardData_10; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_1_io_sbuffer_forwardData_11; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_1_io_sbuffer_forwardData_12; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_1_io_sbuffer_forwardData_13; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_1_io_sbuffer_forwardData_14; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_1_io_sbuffer_forwardData_15; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_sbuffer_matchInvalid; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_loadIn_valid; // @[MemBlock.scala 139:56]
  wire [9:0] LoadUnit_1_io_lsq_loadIn_bits_uop_cf_foldpc; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_loadIn_bits_uop_cf_exceptionVec_4; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_loadIn_bits_uop_cf_exceptionVec_5; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_loadIn_bits_uop_cf_exceptionVec_13; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_loadIn_bits_uop_cf_trigger_backendEn_1; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_loadIn_bits_uop_cf_trigger_backendHit_0; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_loadIn_bits_uop_cf_trigger_backendHit_1; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_loadIn_bits_uop_cf_trigger_backendHit_4; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_loadIn_bits_uop_cf_waitForRobIdx_flag; // @[MemBlock.scala 139:56]
  wire [4:0] LoadUnit_1_io_lsq_loadIn_bits_uop_cf_waitForRobIdx_value; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_loadIn_bits_uop_cf_loadWaitBit; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_loadIn_bits_uop_cf_loadWaitStrict; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_loadIn_bits_uop_cf_ftqPtr_flag; // @[MemBlock.scala 139:56]
  wire [2:0] LoadUnit_1_io_lsq_loadIn_bits_uop_cf_ftqPtr_value; // @[MemBlock.scala 139:56]
  wire [2:0] LoadUnit_1_io_lsq_loadIn_bits_uop_cf_ftqOffset; // @[MemBlock.scala 139:56]
  wire [3:0] LoadUnit_1_io_lsq_loadIn_bits_uop_ctrl_fuType; // @[MemBlock.scala 139:56]
  wire [6:0] LoadUnit_1_io_lsq_loadIn_bits_uop_ctrl_fuOpType; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_loadIn_bits_uop_ctrl_rfWen; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_loadIn_bits_uop_ctrl_fpWen; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_loadIn_bits_uop_ctrl_replayInst; // @[MemBlock.scala 139:56]
  wire [5:0] LoadUnit_1_io_lsq_loadIn_bits_uop_pdest; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_loadIn_bits_uop_robIdx_flag; // @[MemBlock.scala 139:56]
  wire [4:0] LoadUnit_1_io_lsq_loadIn_bits_uop_robIdx_value; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_loadIn_bits_uop_lqIdx_flag; // @[MemBlock.scala 139:56]
  wire [3:0] LoadUnit_1_io_lsq_loadIn_bits_uop_lqIdx_value; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_loadIn_bits_uop_sqIdx_flag; // @[MemBlock.scala 139:56]
  wire [3:0] LoadUnit_1_io_lsq_loadIn_bits_uop_sqIdx_value; // @[MemBlock.scala 139:56]
  wire [38:0] LoadUnit_1_io_lsq_loadIn_bits_vaddr; // @[MemBlock.scala 139:56]
  wire [35:0] LoadUnit_1_io_lsq_loadIn_bits_paddr; // @[MemBlock.scala 139:56]
  wire [15:0] LoadUnit_1_io_lsq_loadIn_bits_mask; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_loadIn_bits_miss; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_loadIn_bits_tlbMiss; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_loadIn_bits_mmio; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_loadIn_bits_rarAllocated; // @[MemBlock.scala 139:56]
  wire [3:0] LoadUnit_1_io_lsq_loadIn_bits_rarIndex; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_loadIn_bits_rawAllocated; // @[MemBlock.scala 139:56]
  wire [2:0] LoadUnit_1_io_lsq_loadIn_bits_rawIndex; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_loadIn_bits_canAccept; // @[MemBlock.scala 139:56]
  wire [1:0] LoadUnit_1_io_lsq_loadIn_bits_replayInfo_missMSHRId; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_loadIn_bits_replayInfo_canForwardFullData; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_loadIn_bits_replayInfo_dataInvalidSqIdx_flag; // @[MemBlock.scala 139:56]
  wire [3:0] LoadUnit_1_io_lsq_loadIn_bits_replayInfo_dataInvalidSqIdx_value; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_loadIn_bits_replayInfo_addrInvalidSqIdx_flag; // @[MemBlock.scala 139:56]
  wire [3:0] LoadUnit_1_io_lsq_loadIn_bits_replayInfo_addrInvalidSqIdx_value; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_1_io_lsq_loadIn_bits_replayInfo_replayCarry_real_way_en; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_loadIn_bits_replayInfo_replayCarry_valid; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_loadIn_bits_replayInfo_dataInLastBeat; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_loadIn_bits_replayInfo_cause_0; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_loadIn_bits_replayInfo_cause_1; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_loadIn_bits_replayInfo_cause_2; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_loadIn_bits_replayInfo_cause_3; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_loadIn_bits_replayInfo_cause_4; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_loadIn_bits_replayInfo_cause_5; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_loadIn_bits_replayInfo_cause_6; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_loadIn_bits_replayInfo_cause_7; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_loadIn_bits_lqDataWenDup_1; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_loadIn_bits_lqDataWenDup_2; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_loadIn_bits_lqDataWenDup_3; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_loadIn_bits_lqDataWenDup_5; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_loadOut_ready; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_loadOut_valid; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_loadOut_bits_uop_cf_exceptionVec_4; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_loadOut_bits_uop_cf_exceptionVec_5; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_loadOut_bits_uop_cf_exceptionVec_13; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_loadOut_bits_uop_cf_trigger_backendEn_1; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_loadOut_bits_uop_cf_trigger_backendHit_0; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_loadOut_bits_uop_cf_trigger_backendHit_1; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_loadOut_bits_uop_cf_trigger_backendHit_4; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_loadOut_bits_uop_ctrl_rfWen; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_loadOut_bits_uop_ctrl_fpWen; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_loadOut_bits_uop_ctrl_flushPipe; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_loadOut_bits_uop_ctrl_replayInst; // @[MemBlock.scala 139:56]
  wire [5:0] LoadUnit_1_io_lsq_loadOut_bits_uop_pdest; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_loadOut_bits_uop_robIdx_flag; // @[MemBlock.scala 139:56]
  wire [4:0] LoadUnit_1_io_lsq_loadOut_bits_uop_robIdx_value; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_loadOut_bits_debug_isMMIO; // @[MemBlock.scala 139:56]
  wire [63:0] LoadUnit_1_io_lsq_ldRawData_lqData; // @[MemBlock.scala 139:56]
  wire [6:0] LoadUnit_1_io_lsq_ldRawData_uop_ctrl_fuOpType; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_ldRawData_uop_ctrl_fpWen; // @[MemBlock.scala 139:56]
  wire [2:0] LoadUnit_1_io_lsq_ldRawData_addrOffset; // @[MemBlock.scala 139:56]
  wire [38:0] LoadUnit_1_io_lsq_forward_vaddr; // @[MemBlock.scala 139:56]
  wire [35:0] LoadUnit_1_io_lsq_forward_paddr; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_forward_uop_cf_waitForRobIdx_flag; // @[MemBlock.scala 139:56]
  wire [4:0] LoadUnit_1_io_lsq_forward_uop_cf_waitForRobIdx_value; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_forward_uop_sqIdx_flag; // @[MemBlock.scala 139:56]
  wire [3:0] LoadUnit_1_io_lsq_forward_uop_sqIdx_value; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_forward_valid; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_forward_forwardMask_0; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_forward_forwardMask_1; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_forward_forwardMask_2; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_forward_forwardMask_3; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_forward_forwardMask_4; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_forward_forwardMask_5; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_forward_forwardMask_6; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_forward_forwardMask_7; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_forward_forwardMask_8; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_forward_forwardMask_9; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_forward_forwardMask_10; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_forward_forwardMask_11; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_forward_forwardMask_12; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_forward_forwardMask_13; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_forward_forwardMask_14; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_forward_forwardMask_15; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_1_io_lsq_forward_forwardData_0; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_1_io_lsq_forward_forwardData_1; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_1_io_lsq_forward_forwardData_2; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_1_io_lsq_forward_forwardData_3; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_1_io_lsq_forward_forwardData_4; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_1_io_lsq_forward_forwardData_5; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_1_io_lsq_forward_forwardData_6; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_1_io_lsq_forward_forwardData_7; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_1_io_lsq_forward_forwardData_8; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_1_io_lsq_forward_forwardData_9; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_1_io_lsq_forward_forwardData_10; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_1_io_lsq_forward_forwardData_11; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_1_io_lsq_forward_forwardData_12; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_1_io_lsq_forward_forwardData_13; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_1_io_lsq_forward_forwardData_14; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_1_io_lsq_forward_forwardData_15; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_forward_sqIdx_flag; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_forward_dataInvalid; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_forward_matchInvalid; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_forward_schedWait; // @[MemBlock.scala 139:56]
  wire [11:0] LoadUnit_1_io_lsq_forward_sqIdxMask; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_forward_dataInvalidSqIdx_flag; // @[MemBlock.scala 139:56]
  wire [3:0] LoadUnit_1_io_lsq_forward_dataInvalidSqIdx_value; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_forward_addrInvalidSqIdx_flag; // @[MemBlock.scala 139:56]
  wire [3:0] LoadUnit_1_io_lsq_forward_addrInvalidSqIdx_value; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_storeLoadViolationQuery_req_valid; // @[MemBlock.scala 139:56]
  wire [9:0] LoadUnit_1_io_lsq_storeLoadViolationQuery_req_bits_uop_cf_foldpc; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_storeLoadViolationQuery_req_bits_uop_cf_ftqPtr_flag; // @[MemBlock.scala 139:56]
  wire [2:0] LoadUnit_1_io_lsq_storeLoadViolationQuery_req_bits_uop_cf_ftqPtr_value; // @[MemBlock.scala 139:56]
  wire [2:0] LoadUnit_1_io_lsq_storeLoadViolationQuery_req_bits_uop_cf_ftqOffset; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_storeLoadViolationQuery_req_bits_uop_robIdx_flag; // @[MemBlock.scala 139:56]
  wire [4:0] LoadUnit_1_io_lsq_storeLoadViolationQuery_req_bits_uop_robIdx_value; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_storeLoadViolationQuery_req_bits_uop_sqIdx_flag; // @[MemBlock.scala 139:56]
  wire [3:0] LoadUnit_1_io_lsq_storeLoadViolationQuery_req_bits_uop_sqIdx_value; // @[MemBlock.scala 139:56]
  wire [2:0] LoadUnit_1_io_lsq_storeLoadViolationQuery_req_bits_index; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_storeLoadViolationQuery_req_bits_allocated; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_storeLoadViolationQuery_req_bits_datavalid; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_1_io_lsq_storeLoadViolationQuery_req_bits_mask; // @[MemBlock.scala 139:56]
  wire [35:0] LoadUnit_1_io_lsq_storeLoadViolationQuery_req_bits_paddr; // @[MemBlock.scala 139:56]
  wire [2:0] LoadUnit_1_io_lsq_storeLoadViolationQuery_resp_bits_index; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_storeLoadViolationQuery_resp_bits_canAccept; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_storeLoadViolationQuery_resp_bits_allocated; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_loadLoadViolationQuery_req_valid; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_loadLoadViolationQuery_req_bits_uop_robIdx_flag; // @[MemBlock.scala 139:56]
  wire [4:0] LoadUnit_1_io_lsq_loadLoadViolationQuery_req_bits_uop_robIdx_value; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_loadLoadViolationQuery_req_bits_uop_lqIdx_flag; // @[MemBlock.scala 139:56]
  wire [3:0] LoadUnit_1_io_lsq_loadLoadViolationQuery_req_bits_uop_lqIdx_value; // @[MemBlock.scala 139:56]
  wire [3:0] LoadUnit_1_io_lsq_loadLoadViolationQuery_req_bits_index; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_loadLoadViolationQuery_req_bits_allocated; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_loadLoadViolationQuery_req_bits_datavalid; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_loadLoadViolationQuery_req_bits_miss; // @[MemBlock.scala 139:56]
  wire [35:0] LoadUnit_1_io_lsq_loadLoadViolationQuery_req_bits_paddr; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_loadLoadViolationQuery_resp_valid; // @[MemBlock.scala 139:56]
  wire [3:0] LoadUnit_1_io_lsq_loadLoadViolationQuery_resp_bits_index; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_loadLoadViolationQuery_resp_bits_canAccept; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_loadLoadViolationQuery_resp_bits_allocated; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_loadLoadViolationQuery_resp_bits_replayFromFetch; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_trigger_hitLoadAddrTriggerHitVec_0; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_trigger_hitLoadAddrTriggerHitVec_1; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_trigger_hitLoadAddrTriggerHitVec_2; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_trigger_lqLoadAddrTriggerHitVec_0; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_trigger_lqLoadAddrTriggerHitVec_1; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lsq_trigger_lqLoadAddrTriggerHitVec_2; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_tlDchannel_valid; // @[MemBlock.scala 139:56]
  wire [255:0] LoadUnit_1_io_tlDchannel_data; // @[MemBlock.scala 139:56]
  wire [1:0] LoadUnit_1_io_tlDchannel_mshrid; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_tlDchannel_last; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_forward_mshr_valid; // @[MemBlock.scala 139:56]
  wire [1:0] LoadUnit_1_io_forward_mshr_mshrid; // @[MemBlock.scala 139:56]
  wire [35:0] LoadUnit_1_io_forward_mshr_paddr; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_forward_mshr_forward_mshr; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_1_io_forward_mshr_forwardData_0; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_1_io_forward_mshr_forwardData_1; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_1_io_forward_mshr_forwardData_2; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_1_io_forward_mshr_forwardData_3; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_1_io_forward_mshr_forwardData_4; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_1_io_forward_mshr_forwardData_5; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_1_io_forward_mshr_forwardData_6; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_1_io_forward_mshr_forwardData_7; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_1_io_forward_mshr_forwardData_8; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_1_io_forward_mshr_forwardData_9; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_1_io_forward_mshr_forwardData_10; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_1_io_forward_mshr_forwardData_11; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_1_io_forward_mshr_forwardData_12; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_1_io_forward_mshr_forwardData_13; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_1_io_forward_mshr_forwardData_14; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_1_io_forward_mshr_forwardData_15; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_forward_mshr_forward_result_valid; // @[MemBlock.scala 139:56]
  wire [63:0] LoadUnit_1_io_trigger_0_tdata2; // @[MemBlock.scala 139:56]
  wire [1:0] LoadUnit_1_io_trigger_0_matchType; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_trigger_0_tEnable; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_trigger_0_addrHit; // @[MemBlock.scala 139:56]
  wire [63:0] LoadUnit_1_io_trigger_1_tdata2; // @[MemBlock.scala 139:56]
  wire [1:0] LoadUnit_1_io_trigger_1_matchType; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_trigger_1_tEnable; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_trigger_1_addrHit; // @[MemBlock.scala 139:56]
  wire [63:0] LoadUnit_1_io_trigger_2_tdata2; // @[MemBlock.scala 139:56]
  wire [1:0] LoadUnit_1_io_trigger_2_matchType; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_trigger_2_tEnable; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_trigger_2_addrHit; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_tlb_req_valid; // @[MemBlock.scala 139:56]
  wire [38:0] LoadUnit_1_io_tlb_req_bits_vaddr; // @[MemBlock.scala 139:56]
  wire [2:0] LoadUnit_1_io_tlb_req_bits_cmd; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_tlb_req_bits_no_translate; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_tlb_req_kill; // @[MemBlock.scala 139:56]
  wire [35:0] LoadUnit_1_io_tlb_resp_bits_paddr_0; // @[MemBlock.scala 139:56]
  wire [35:0] LoadUnit_1_io_tlb_resp_bits_paddr_1; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_tlb_resp_bits_miss; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_tlb_resp_bits_excp_0_pf_ld; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_tlb_resp_bits_excp_0_af_ld; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_tlb_resp_bits_static_pm_valid; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_tlb_resp_bits_static_pm_bits; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_pmp_ld; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_pmp_mmio; // @[MemBlock.scala 139:56]
  wire [63:0] LoadUnit_1_io_fastpathOut_data; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_fastpathOut_valid; // @[MemBlock.scala 139:56]
  wire [63:0] LoadUnit_1_io_fastpathIn_data; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_fastpathIn_valid; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_loadFastMatch; // @[MemBlock.scala 139:56]
  wire [11:0] LoadUnit_1_io_loadFastImm; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_csrCtrl_ldld_vio_check_enable; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_csrCtrl_cache_error_enable; // @[MemBlock.scala 139:56]
  wire [9:0] LoadUnit_1_io_correctTableQuery_req_addr; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_correctTableQuery_resp_strict; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_correctTableUpdate_valid; // @[MemBlock.scala 139:56]
  wire [9:0] LoadUnit_1_io_correctTableUpdate_bits_addr; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_correctTableUpdate_bits_strict; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_correctTableUpdate_bits_violation; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_reExecuteQuery_0_valid; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_reExecuteQuery_0_bits_robIdx_flag; // @[MemBlock.scala 139:56]
  wire [4:0] LoadUnit_1_io_reExecuteQuery_0_bits_robIdx_value; // @[MemBlock.scala 139:56]
  wire [35:0] LoadUnit_1_io_reExecuteQuery_0_bits_paddr; // @[MemBlock.scala 139:56]
  wire [15:0] LoadUnit_1_io_reExecuteQuery_0_bits_mask; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_reExecuteQuery_1_valid; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_reExecuteQuery_1_bits_robIdx_flag; // @[MemBlock.scala 139:56]
  wire [4:0] LoadUnit_1_io_reExecuteQuery_1_bits_robIdx_value; // @[MemBlock.scala 139:56]
  wire [35:0] LoadUnit_1_io_reExecuteQuery_1_bits_paddr; // @[MemBlock.scala 139:56]
  wire [15:0] LoadUnit_1_io_reExecuteQuery_1_bits_mask; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_replay_ready; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_replay_valid; // @[MemBlock.scala 139:56]
  wire [9:0] LoadUnit_1_io_replay_bits_uop_cf_foldpc; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_replay_bits_uop_cf_trigger_backendEn_1; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_replay_bits_uop_cf_trigger_backendHit_0; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_replay_bits_uop_cf_trigger_backendHit_1; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_replay_bits_uop_cf_trigger_backendHit_4; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_replay_bits_uop_cf_waitForRobIdx_flag; // @[MemBlock.scala 139:56]
  wire [4:0] LoadUnit_1_io_replay_bits_uop_cf_waitForRobIdx_value; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_replay_bits_uop_cf_loadWaitBit; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_replay_bits_uop_cf_loadWaitStrict; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_replay_bits_uop_cf_ftqPtr_flag; // @[MemBlock.scala 139:56]
  wire [2:0] LoadUnit_1_io_replay_bits_uop_cf_ftqPtr_value; // @[MemBlock.scala 139:56]
  wire [2:0] LoadUnit_1_io_replay_bits_uop_cf_ftqOffset; // @[MemBlock.scala 139:56]
  wire [3:0] LoadUnit_1_io_replay_bits_uop_ctrl_fuType; // @[MemBlock.scala 139:56]
  wire [6:0] LoadUnit_1_io_replay_bits_uop_ctrl_fuOpType; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_replay_bits_uop_ctrl_rfWen; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_replay_bits_uop_ctrl_fpWen; // @[MemBlock.scala 139:56]
  wire [5:0] LoadUnit_1_io_replay_bits_uop_pdest; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_replay_bits_uop_robIdx_flag; // @[MemBlock.scala 139:56]
  wire [4:0] LoadUnit_1_io_replay_bits_uop_robIdx_value; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_replay_bits_uop_lqIdx_flag; // @[MemBlock.scala 139:56]
  wire [3:0] LoadUnit_1_io_replay_bits_uop_lqIdx_value; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_replay_bits_uop_sqIdx_flag; // @[MemBlock.scala 139:56]
  wire [3:0] LoadUnit_1_io_replay_bits_uop_sqIdx_value; // @[MemBlock.scala 139:56]
  wire [38:0] LoadUnit_1_io_replay_bits_vaddr; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_replay_bits_isFirstIssue; // @[MemBlock.scala 139:56]
  wire [7:0] LoadUnit_1_io_replay_bits_replayCarry_real_way_en; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_replay_bits_replayCarry_valid; // @[MemBlock.scala 139:56]
  wire [1:0] LoadUnit_1_io_replay_bits_mshrid; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_replay_bits_forward_tlDchannel; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_replay_bits_rarAllocated; // @[MemBlock.scala 139:56]
  wire [3:0] LoadUnit_1_io_replay_bits_rarIndex; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_replay_bits_rawAllocated; // @[MemBlock.scala 139:56]
  wire [2:0] LoadUnit_1_io_replay_bits_rawIndex; // @[MemBlock.scala 139:56]
  wire  LoadUnit_1_io_lqReplayFull; // @[MemBlock.scala 139:56]
  wire [5:0] LoadUnit_1_io_perf_0_value; // @[MemBlock.scala 139:56]
  wire [5:0] LoadUnit_1_io_perf_1_value; // @[MemBlock.scala 139:56]
  wire [5:0] LoadUnit_1_io_perf_2_value; // @[MemBlock.scala 139:56]
  wire [5:0] LoadUnit_1_io_perf_3_value; // @[MemBlock.scala 139:56]
  wire [5:0] LoadUnit_1_io_perf_4_value; // @[MemBlock.scala 139:56]
  wire [5:0] LoadUnit_1_io_perf_5_value; // @[MemBlock.scala 139:56]
  wire [5:0] LoadUnit_1_io_perf_6_value; // @[MemBlock.scala 139:56]
  wire  StoreUnit_0_clock; // @[MemBlock.scala 140:57]
  wire  StoreUnit_0_reset; // @[MemBlock.scala 140:57]
  wire  StoreUnit_0_io_stin_valid; // @[MemBlock.scala 140:57]
  wire  StoreUnit_0_io_stin_bits_uop_cf_trigger_backendEn_0; // @[MemBlock.scala 140:57]
  wire  StoreUnit_0_io_stin_bits_uop_cf_storeSetHit; // @[MemBlock.scala 140:57]
  wire [4:0] StoreUnit_0_io_stin_bits_uop_cf_ssid; // @[MemBlock.scala 140:57]
  wire [2:0] StoreUnit_0_io_stin_bits_uop_cf_ftqPtr_value; // @[MemBlock.scala 140:57]
  wire [2:0] StoreUnit_0_io_stin_bits_uop_cf_ftqOffset; // @[MemBlock.scala 140:57]
  wire [6:0] StoreUnit_0_io_stin_bits_uop_ctrl_fuOpType; // @[MemBlock.scala 140:57]
  wire [19:0] StoreUnit_0_io_stin_bits_uop_ctrl_imm; // @[MemBlock.scala 140:57]
  wire  StoreUnit_0_io_stin_bits_uop_robIdx_flag; // @[MemBlock.scala 140:57]
  wire [4:0] StoreUnit_0_io_stin_bits_uop_robIdx_value; // @[MemBlock.scala 140:57]
  wire  StoreUnit_0_io_stin_bits_uop_sqIdx_flag; // @[MemBlock.scala 140:57]
  wire [3:0] StoreUnit_0_io_stin_bits_uop_sqIdx_value; // @[MemBlock.scala 140:57]
  wire [63:0] StoreUnit_0_io_stin_bits_src_0; // @[MemBlock.scala 140:57]
  wire  StoreUnit_0_io_redirect_valid; // @[MemBlock.scala 140:57]
  wire  StoreUnit_0_io_redirect_bits_robIdx_flag; // @[MemBlock.scala 140:57]
  wire [4:0] StoreUnit_0_io_redirect_bits_robIdx_value; // @[MemBlock.scala 140:57]
  wire  StoreUnit_0_io_redirect_bits_level; // @[MemBlock.scala 140:57]
  wire  StoreUnit_0_io_feedbackSlow_valid; // @[MemBlock.scala 140:57]
  wire [3:0] StoreUnit_0_io_feedbackSlow_bits_rsIdx; // @[MemBlock.scala 140:57]
  wire  StoreUnit_0_io_feedbackSlow_bits_hit; // @[MemBlock.scala 140:57]
  wire  StoreUnit_0_io_tlb_req_valid; // @[MemBlock.scala 140:57]
  wire [38:0] StoreUnit_0_io_tlb_req_bits_vaddr; // @[MemBlock.scala 140:57]
  wire [35:0] StoreUnit_0_io_tlb_resp_bits_paddr_0; // @[MemBlock.scala 140:57]
  wire  StoreUnit_0_io_tlb_resp_bits_miss; // @[MemBlock.scala 140:57]
  wire  StoreUnit_0_io_tlb_resp_bits_excp_0_pf_st; // @[MemBlock.scala 140:57]
  wire  StoreUnit_0_io_tlb_resp_bits_excp_0_af_st; // @[MemBlock.scala 140:57]
  wire  StoreUnit_0_io_tlb_resp_bits_static_pm_valid; // @[MemBlock.scala 140:57]
  wire  StoreUnit_0_io_tlb_resp_bits_static_pm_bits; // @[MemBlock.scala 140:57]
  wire  StoreUnit_0_io_pmp_st; // @[MemBlock.scala 140:57]
  wire  StoreUnit_0_io_pmp_mmio; // @[MemBlock.scala 140:57]
  wire  StoreUnit_0_io_pmp_atomic; // @[MemBlock.scala 140:57]
  wire [3:0] StoreUnit_0_io_rsIdx; // @[MemBlock.scala 140:57]
  wire  StoreUnit_0_io_lsq_valid; // @[MemBlock.scala 140:57]
  wire [2:0] StoreUnit_0_io_lsq_bits_uop_cf_ftqPtr_value; // @[MemBlock.scala 140:57]
  wire [2:0] StoreUnit_0_io_lsq_bits_uop_cf_ftqOffset; // @[MemBlock.scala 140:57]
  wire [6:0] StoreUnit_0_io_lsq_bits_uop_ctrl_fuOpType; // @[MemBlock.scala 140:57]
  wire  StoreUnit_0_io_lsq_bits_uop_robIdx_flag; // @[MemBlock.scala 140:57]
  wire [4:0] StoreUnit_0_io_lsq_bits_uop_robIdx_value; // @[MemBlock.scala 140:57]
  wire  StoreUnit_0_io_lsq_bits_uop_sqIdx_flag; // @[MemBlock.scala 140:57]
  wire [3:0] StoreUnit_0_io_lsq_bits_uop_sqIdx_value; // @[MemBlock.scala 140:57]
  wire [38:0] StoreUnit_0_io_lsq_bits_vaddr; // @[MemBlock.scala 140:57]
  wire [35:0] StoreUnit_0_io_lsq_bits_paddr; // @[MemBlock.scala 140:57]
  wire [15:0] StoreUnit_0_io_lsq_bits_mask; // @[MemBlock.scala 140:57]
  wire  StoreUnit_0_io_lsq_bits_wlineflag; // @[MemBlock.scala 140:57]
  wire  StoreUnit_0_io_lsq_bits_miss; // @[MemBlock.scala 140:57]
  wire  StoreUnit_0_io_lsq_replenish_mmio; // @[MemBlock.scala 140:57]
  wire  StoreUnit_0_io_lsq_replenish_atomic; // @[MemBlock.scala 140:57]
  wire  StoreUnit_0_io_stout_valid; // @[MemBlock.scala 140:57]
  wire  StoreUnit_0_io_stout_bits_uop_cf_exceptionVec_6; // @[MemBlock.scala 140:57]
  wire  StoreUnit_0_io_stout_bits_uop_cf_exceptionVec_7; // @[MemBlock.scala 140:57]
  wire  StoreUnit_0_io_stout_bits_uop_cf_exceptionVec_15; // @[MemBlock.scala 140:57]
  wire  StoreUnit_0_io_stout_bits_uop_cf_trigger_backendEn_0; // @[MemBlock.scala 140:57]
  wire  StoreUnit_0_io_stout_bits_uop_robIdx_flag; // @[MemBlock.scala 140:57]
  wire [4:0] StoreUnit_0_io_stout_bits_uop_robIdx_value; // @[MemBlock.scala 140:57]
  wire  StoreUnit_0_io_stout_bits_debug_isMMIO; // @[MemBlock.scala 140:57]
  wire [38:0] StoreUnit_0_io_stout_bits_debug_vaddr; // @[MemBlock.scala 140:57]
  wire  StoreUnit_0_io_storeMaskOut_valid; // @[MemBlock.scala 140:57]
  wire [3:0] StoreUnit_0_io_storeMaskOut_bits_sqIdx_value; // @[MemBlock.scala 140:57]
  wire [15:0] StoreUnit_0_io_storeMaskOut_bits_mask; // @[MemBlock.scala 140:57]
  wire  StoreUnit_0_io_reExecuteQuery_valid; // @[MemBlock.scala 140:57]
  wire  StoreUnit_0_io_reExecuteQuery_bits_robIdx_flag; // @[MemBlock.scala 140:57]
  wire [4:0] StoreUnit_0_io_reExecuteQuery_bits_robIdx_value; // @[MemBlock.scala 140:57]
  wire [35:0] StoreUnit_0_io_reExecuteQuery_bits_paddr; // @[MemBlock.scala 140:57]
  wire [15:0] StoreUnit_0_io_reExecuteQuery_bits_mask; // @[MemBlock.scala 140:57]
  wire  StoreUnit_0_io_issue_valid; // @[MemBlock.scala 140:57]
  wire  StoreUnit_0_io_issue_bits_uop_cf_storeSetHit; // @[MemBlock.scala 140:57]
  wire [4:0] StoreUnit_0_io_issue_bits_uop_cf_ssid; // @[MemBlock.scala 140:57]
  wire [4:0] StoreUnit_0_io_issue_bits_uop_robIdx_value; // @[MemBlock.scala 140:57]
  wire  StoreUnit_1_clock; // @[MemBlock.scala 140:57]
  wire  StoreUnit_1_reset; // @[MemBlock.scala 140:57]
  wire  StoreUnit_1_io_stin_valid; // @[MemBlock.scala 140:57]
  wire  StoreUnit_1_io_stin_bits_uop_cf_trigger_backendEn_0; // @[MemBlock.scala 140:57]
  wire  StoreUnit_1_io_stin_bits_uop_cf_storeSetHit; // @[MemBlock.scala 140:57]
  wire [4:0] StoreUnit_1_io_stin_bits_uop_cf_ssid; // @[MemBlock.scala 140:57]
  wire [2:0] StoreUnit_1_io_stin_bits_uop_cf_ftqPtr_value; // @[MemBlock.scala 140:57]
  wire [2:0] StoreUnit_1_io_stin_bits_uop_cf_ftqOffset; // @[MemBlock.scala 140:57]
  wire [6:0] StoreUnit_1_io_stin_bits_uop_ctrl_fuOpType; // @[MemBlock.scala 140:57]
  wire [19:0] StoreUnit_1_io_stin_bits_uop_ctrl_imm; // @[MemBlock.scala 140:57]
  wire  StoreUnit_1_io_stin_bits_uop_robIdx_flag; // @[MemBlock.scala 140:57]
  wire [4:0] StoreUnit_1_io_stin_bits_uop_robIdx_value; // @[MemBlock.scala 140:57]
  wire  StoreUnit_1_io_stin_bits_uop_sqIdx_flag; // @[MemBlock.scala 140:57]
  wire [3:0] StoreUnit_1_io_stin_bits_uop_sqIdx_value; // @[MemBlock.scala 140:57]
  wire [63:0] StoreUnit_1_io_stin_bits_src_0; // @[MemBlock.scala 140:57]
  wire  StoreUnit_1_io_redirect_valid; // @[MemBlock.scala 140:57]
  wire  StoreUnit_1_io_redirect_bits_robIdx_flag; // @[MemBlock.scala 140:57]
  wire [4:0] StoreUnit_1_io_redirect_bits_robIdx_value; // @[MemBlock.scala 140:57]
  wire  StoreUnit_1_io_redirect_bits_level; // @[MemBlock.scala 140:57]
  wire  StoreUnit_1_io_feedbackSlow_valid; // @[MemBlock.scala 140:57]
  wire [3:0] StoreUnit_1_io_feedbackSlow_bits_rsIdx; // @[MemBlock.scala 140:57]
  wire  StoreUnit_1_io_feedbackSlow_bits_hit; // @[MemBlock.scala 140:57]
  wire  StoreUnit_1_io_tlb_req_valid; // @[MemBlock.scala 140:57]
  wire [38:0] StoreUnit_1_io_tlb_req_bits_vaddr; // @[MemBlock.scala 140:57]
  wire [35:0] StoreUnit_1_io_tlb_resp_bits_paddr_0; // @[MemBlock.scala 140:57]
  wire  StoreUnit_1_io_tlb_resp_bits_miss; // @[MemBlock.scala 140:57]
  wire  StoreUnit_1_io_tlb_resp_bits_excp_0_pf_st; // @[MemBlock.scala 140:57]
  wire  StoreUnit_1_io_tlb_resp_bits_excp_0_af_st; // @[MemBlock.scala 140:57]
  wire  StoreUnit_1_io_tlb_resp_bits_static_pm_valid; // @[MemBlock.scala 140:57]
  wire  StoreUnit_1_io_tlb_resp_bits_static_pm_bits; // @[MemBlock.scala 140:57]
  wire  StoreUnit_1_io_pmp_st; // @[MemBlock.scala 140:57]
  wire  StoreUnit_1_io_pmp_mmio; // @[MemBlock.scala 140:57]
  wire  StoreUnit_1_io_pmp_atomic; // @[MemBlock.scala 140:57]
  wire [3:0] StoreUnit_1_io_rsIdx; // @[MemBlock.scala 140:57]
  wire  StoreUnit_1_io_lsq_valid; // @[MemBlock.scala 140:57]
  wire [2:0] StoreUnit_1_io_lsq_bits_uop_cf_ftqPtr_value; // @[MemBlock.scala 140:57]
  wire [2:0] StoreUnit_1_io_lsq_bits_uop_cf_ftqOffset; // @[MemBlock.scala 140:57]
  wire [6:0] StoreUnit_1_io_lsq_bits_uop_ctrl_fuOpType; // @[MemBlock.scala 140:57]
  wire  StoreUnit_1_io_lsq_bits_uop_robIdx_flag; // @[MemBlock.scala 140:57]
  wire [4:0] StoreUnit_1_io_lsq_bits_uop_robIdx_value; // @[MemBlock.scala 140:57]
  wire  StoreUnit_1_io_lsq_bits_uop_sqIdx_flag; // @[MemBlock.scala 140:57]
  wire [3:0] StoreUnit_1_io_lsq_bits_uop_sqIdx_value; // @[MemBlock.scala 140:57]
  wire [38:0] StoreUnit_1_io_lsq_bits_vaddr; // @[MemBlock.scala 140:57]
  wire [35:0] StoreUnit_1_io_lsq_bits_paddr; // @[MemBlock.scala 140:57]
  wire [15:0] StoreUnit_1_io_lsq_bits_mask; // @[MemBlock.scala 140:57]
  wire  StoreUnit_1_io_lsq_bits_wlineflag; // @[MemBlock.scala 140:57]
  wire  StoreUnit_1_io_lsq_bits_miss; // @[MemBlock.scala 140:57]
  wire  StoreUnit_1_io_lsq_replenish_mmio; // @[MemBlock.scala 140:57]
  wire  StoreUnit_1_io_lsq_replenish_atomic; // @[MemBlock.scala 140:57]
  wire  StoreUnit_1_io_stout_valid; // @[MemBlock.scala 140:57]
  wire  StoreUnit_1_io_stout_bits_uop_cf_exceptionVec_6; // @[MemBlock.scala 140:57]
  wire  StoreUnit_1_io_stout_bits_uop_cf_exceptionVec_7; // @[MemBlock.scala 140:57]
  wire  StoreUnit_1_io_stout_bits_uop_cf_exceptionVec_15; // @[MemBlock.scala 140:57]
  wire  StoreUnit_1_io_stout_bits_uop_cf_trigger_backendEn_0; // @[MemBlock.scala 140:57]
  wire  StoreUnit_1_io_stout_bits_uop_robIdx_flag; // @[MemBlock.scala 140:57]
  wire [4:0] StoreUnit_1_io_stout_bits_uop_robIdx_value; // @[MemBlock.scala 140:57]
  wire  StoreUnit_1_io_stout_bits_debug_isMMIO; // @[MemBlock.scala 140:57]
  wire [38:0] StoreUnit_1_io_stout_bits_debug_vaddr; // @[MemBlock.scala 140:57]
  wire  StoreUnit_1_io_storeMaskOut_valid; // @[MemBlock.scala 140:57]
  wire [3:0] StoreUnit_1_io_storeMaskOut_bits_sqIdx_value; // @[MemBlock.scala 140:57]
  wire [15:0] StoreUnit_1_io_storeMaskOut_bits_mask; // @[MemBlock.scala 140:57]
  wire  StoreUnit_1_io_reExecuteQuery_valid; // @[MemBlock.scala 140:57]
  wire  StoreUnit_1_io_reExecuteQuery_bits_robIdx_flag; // @[MemBlock.scala 140:57]
  wire [4:0] StoreUnit_1_io_reExecuteQuery_bits_robIdx_value; // @[MemBlock.scala 140:57]
  wire [35:0] StoreUnit_1_io_reExecuteQuery_bits_paddr; // @[MemBlock.scala 140:57]
  wire [15:0] StoreUnit_1_io_reExecuteQuery_bits_mask; // @[MemBlock.scala 140:57]
  wire  StoreUnit_1_io_issue_valid; // @[MemBlock.scala 140:57]
  wire  StoreUnit_1_io_issue_bits_uop_cf_storeSetHit; // @[MemBlock.scala 140:57]
  wire [4:0] StoreUnit_1_io_issue_bits_uop_cf_ssid; // @[MemBlock.scala 140:57]
  wire [4:0] StoreUnit_1_io_issue_bits_uop_robIdx_value; // @[MemBlock.scala 140:57]
  wire  stdExeUnits_0_io_fromInt_ready; // @[MemBlock.scala 141:58]
  wire  stdExeUnits_0_io_fromInt_valid; // @[MemBlock.scala 141:58]
  wire [3:0] stdExeUnits_0_io_fromInt_bits_uop_ctrl_fuType; // @[MemBlock.scala 141:58]
  wire [6:0] stdExeUnits_0_io_fromInt_bits_uop_ctrl_fuOpType; // @[MemBlock.scala 141:58]
  wire  stdExeUnits_0_io_fromInt_bits_uop_robIdx_flag; // @[MemBlock.scala 141:58]
  wire [4:0] stdExeUnits_0_io_fromInt_bits_uop_robIdx_value; // @[MemBlock.scala 141:58]
  wire  stdExeUnits_0_io_fromInt_bits_uop_sqIdx_flag; // @[MemBlock.scala 141:58]
  wire [3:0] stdExeUnits_0_io_fromInt_bits_uop_sqIdx_value; // @[MemBlock.scala 141:58]
  wire [63:0] stdExeUnits_0_io_fromInt_bits_src_0; // @[MemBlock.scala 141:58]
  wire  stdExeUnits_0_io_out_valid; // @[MemBlock.scala 141:58]
  wire [3:0] stdExeUnits_0_io_out_bits_uop_ctrl_fuType; // @[MemBlock.scala 141:58]
  wire [6:0] stdExeUnits_0_io_out_bits_uop_ctrl_fuOpType; // @[MemBlock.scala 141:58]
  wire  stdExeUnits_0_io_out_bits_uop_robIdx_flag; // @[MemBlock.scala 141:58]
  wire [4:0] stdExeUnits_0_io_out_bits_uop_robIdx_value; // @[MemBlock.scala 141:58]
  wire  stdExeUnits_0_io_out_bits_uop_sqIdx_flag; // @[MemBlock.scala 141:58]
  wire [3:0] stdExeUnits_0_io_out_bits_uop_sqIdx_value; // @[MemBlock.scala 141:58]
  wire [63:0] stdExeUnits_0_io_out_bits_data; // @[MemBlock.scala 141:58]
  wire  stdExeUnits_1_io_fromInt_ready; // @[MemBlock.scala 141:58]
  wire  stdExeUnits_1_io_fromInt_valid; // @[MemBlock.scala 141:58]
  wire [3:0] stdExeUnits_1_io_fromInt_bits_uop_ctrl_fuType; // @[MemBlock.scala 141:58]
  wire [6:0] stdExeUnits_1_io_fromInt_bits_uop_ctrl_fuOpType; // @[MemBlock.scala 141:58]
  wire  stdExeUnits_1_io_fromInt_bits_uop_robIdx_flag; // @[MemBlock.scala 141:58]
  wire [4:0] stdExeUnits_1_io_fromInt_bits_uop_robIdx_value; // @[MemBlock.scala 141:58]
  wire  stdExeUnits_1_io_fromInt_bits_uop_sqIdx_flag; // @[MemBlock.scala 141:58]
  wire [3:0] stdExeUnits_1_io_fromInt_bits_uop_sqIdx_value; // @[MemBlock.scala 141:58]
  wire [63:0] stdExeUnits_1_io_fromInt_bits_src_0; // @[MemBlock.scala 141:58]
  wire  stdExeUnits_1_io_out_valid; // @[MemBlock.scala 141:58]
  wire [3:0] stdExeUnits_1_io_out_bits_uop_ctrl_fuType; // @[MemBlock.scala 141:58]
  wire [6:0] stdExeUnits_1_io_out_bits_uop_ctrl_fuOpType; // @[MemBlock.scala 141:58]
  wire  stdExeUnits_1_io_out_bits_uop_robIdx_flag; // @[MemBlock.scala 141:58]
  wire [4:0] stdExeUnits_1_io_out_bits_uop_robIdx_value; // @[MemBlock.scala 141:58]
  wire  stdExeUnits_1_io_out_bits_uop_sqIdx_flag; // @[MemBlock.scala 141:58]
  wire [3:0] stdExeUnits_1_io_out_bits_uop_sqIdx_value; // @[MemBlock.scala 141:58]
  wire [63:0] stdExeUnits_1_io_out_bits_data; // @[MemBlock.scala 141:58]
  wire  correctTable_clock; // @[MemBlock.scala 144:28]
  wire [9:0] correctTable_io_issue_0_req_addr; // @[MemBlock.scala 144:28]
  wire  correctTable_io_issue_0_resp_strict; // @[MemBlock.scala 144:28]
  wire [9:0] correctTable_io_issue_1_req_addr; // @[MemBlock.scala 144:28]
  wire  correctTable_io_issue_1_resp_strict; // @[MemBlock.scala 144:28]
  wire  correctTable_io_update_0_valid; // @[MemBlock.scala 144:28]
  wire [9:0] correctTable_io_update_0_bits_addr; // @[MemBlock.scala 144:28]
  wire  correctTable_io_update_0_bits_strict; // @[MemBlock.scala 144:28]
  wire  correctTable_io_update_0_bits_violation; // @[MemBlock.scala 144:28]
  wire  correctTable_io_update_1_valid; // @[MemBlock.scala 144:28]
  wire [9:0] correctTable_io_update_1_bits_addr; // @[MemBlock.scala 144:28]
  wire  correctTable_io_update_1_bits_strict; // @[MemBlock.scala 144:28]
  wire  correctTable_io_update_1_bits_violation; // @[MemBlock.scala 144:28]
  wire  correctTable_io_update_2_valid; // @[MemBlock.scala 144:28]
  wire [9:0] correctTable_io_update_2_bits_addr; // @[MemBlock.scala 144:28]
  wire  atomicsUnit_clock; // @[MemBlock.scala 174:27]
  wire  atomicsUnit_reset; // @[MemBlock.scala 174:27]
  wire [7:0] atomicsUnit_io_hartId; // @[MemBlock.scala 174:27]
  wire  atomicsUnit_io_in_ready; // @[MemBlock.scala 174:27]
  wire  atomicsUnit_io_in_valid; // @[MemBlock.scala 174:27]
  wire  atomicsUnit_io_in_bits_uop_cf_trigger_backendEn_0; // @[MemBlock.scala 174:27]
  wire  atomicsUnit_io_in_bits_uop_cf_trigger_backendEn_1; // @[MemBlock.scala 174:27]
  wire [6:0] atomicsUnit_io_in_bits_uop_ctrl_fuOpType; // @[MemBlock.scala 174:27]
  wire  atomicsUnit_io_in_bits_uop_ctrl_rfWen; // @[MemBlock.scala 174:27]
  wire  atomicsUnit_io_in_bits_uop_ctrl_fpWen; // @[MemBlock.scala 174:27]
  wire [5:0] atomicsUnit_io_in_bits_uop_pdest; // @[MemBlock.scala 174:27]
  wire  atomicsUnit_io_in_bits_uop_robIdx_flag; // @[MemBlock.scala 174:27]
  wire [4:0] atomicsUnit_io_in_bits_uop_robIdx_value; // @[MemBlock.scala 174:27]
  wire [63:0] atomicsUnit_io_in_bits_src_0; // @[MemBlock.scala 174:27]
  wire  atomicsUnit_io_storeDataIn_valid; // @[MemBlock.scala 174:27]
  wire [63:0] atomicsUnit_io_storeDataIn_bits_data; // @[MemBlock.scala 174:27]
  wire  atomicsUnit_io_out_valid; // @[MemBlock.scala 174:27]
  wire  atomicsUnit_io_out_bits_uop_cf_exceptionVec_4; // @[MemBlock.scala 174:27]
  wire  atomicsUnit_io_out_bits_uop_cf_exceptionVec_5; // @[MemBlock.scala 174:27]
  wire  atomicsUnit_io_out_bits_uop_cf_exceptionVec_6; // @[MemBlock.scala 174:27]
  wire  atomicsUnit_io_out_bits_uop_cf_exceptionVec_7; // @[MemBlock.scala 174:27]
  wire  atomicsUnit_io_out_bits_uop_cf_exceptionVec_13; // @[MemBlock.scala 174:27]
  wire  atomicsUnit_io_out_bits_uop_cf_exceptionVec_15; // @[MemBlock.scala 174:27]
  wire  atomicsUnit_io_out_bits_uop_cf_trigger_backendEn_0; // @[MemBlock.scala 174:27]
  wire  atomicsUnit_io_out_bits_uop_cf_trigger_backendEn_1; // @[MemBlock.scala 174:27]
  wire  atomicsUnit_io_out_bits_uop_cf_trigger_backendHit_0; // @[MemBlock.scala 174:27]
  wire  atomicsUnit_io_out_bits_uop_cf_trigger_backendHit_1; // @[MemBlock.scala 174:27]
  wire  atomicsUnit_io_out_bits_uop_cf_trigger_backendHit_2; // @[MemBlock.scala 174:27]
  wire  atomicsUnit_io_out_bits_uop_cf_trigger_backendHit_3; // @[MemBlock.scala 174:27]
  wire  atomicsUnit_io_out_bits_uop_cf_trigger_backendHit_4; // @[MemBlock.scala 174:27]
  wire  atomicsUnit_io_out_bits_uop_cf_trigger_backendHit_5; // @[MemBlock.scala 174:27]
  wire [6:0] atomicsUnit_io_out_bits_uop_ctrl_fuOpType; // @[MemBlock.scala 174:27]
  wire  atomicsUnit_io_out_bits_uop_ctrl_rfWen; // @[MemBlock.scala 174:27]
  wire  atomicsUnit_io_out_bits_uop_ctrl_fpWen; // @[MemBlock.scala 174:27]
  wire [5:0] atomicsUnit_io_out_bits_uop_pdest; // @[MemBlock.scala 174:27]
  wire  atomicsUnit_io_out_bits_uop_robIdx_flag; // @[MemBlock.scala 174:27]
  wire [4:0] atomicsUnit_io_out_bits_uop_robIdx_value; // @[MemBlock.scala 174:27]
  wire [63:0] atomicsUnit_io_out_bits_data; // @[MemBlock.scala 174:27]
  wire  atomicsUnit_io_out_bits_debug_isMMIO; // @[MemBlock.scala 174:27]
  wire  atomicsUnit_io_dcache_req_ready; // @[MemBlock.scala 174:27]
  wire  atomicsUnit_io_dcache_req_valid; // @[MemBlock.scala 174:27]
  wire [4:0] atomicsUnit_io_dcache_req_bits_cmd; // @[MemBlock.scala 174:27]
  wire [38:0] atomicsUnit_io_dcache_req_bits_vaddr; // @[MemBlock.scala 174:27]
  wire [35:0] atomicsUnit_io_dcache_req_bits_addr; // @[MemBlock.scala 174:27]
  wire [2:0] atomicsUnit_io_dcache_req_bits_word_idx; // @[MemBlock.scala 174:27]
  wire [63:0] atomicsUnit_io_dcache_req_bits_amo_data; // @[MemBlock.scala 174:27]
  wire [7:0] atomicsUnit_io_dcache_req_bits_amo_mask; // @[MemBlock.scala 174:27]
  wire  atomicsUnit_io_dcache_resp_valid; // @[MemBlock.scala 174:27]
  wire [63:0] atomicsUnit_io_dcache_resp_bits_data; // @[MemBlock.scala 174:27]
  wire  atomicsUnit_io_dcache_resp_bits_miss; // @[MemBlock.scala 174:27]
  wire  atomicsUnit_io_dcache_resp_bits_replay; // @[MemBlock.scala 174:27]
  wire  atomicsUnit_io_dcache_resp_bits_error; // @[MemBlock.scala 174:27]
  wire [3:0] atomicsUnit_io_dcache_resp_bits_id; // @[MemBlock.scala 174:27]
  wire  atomicsUnit_io_dcache_block_lr; // @[MemBlock.scala 174:27]
  wire  atomicsUnit_io_dtlb_req_valid; // @[MemBlock.scala 174:27]
  wire [38:0] atomicsUnit_io_dtlb_req_bits_vaddr; // @[MemBlock.scala 174:27]
  wire [2:0] atomicsUnit_io_dtlb_req_bits_cmd; // @[MemBlock.scala 174:27]
  wire  atomicsUnit_io_dtlb_resp_ready; // @[MemBlock.scala 174:27]
  wire  atomicsUnit_io_dtlb_resp_valid; // @[MemBlock.scala 174:27]
  wire [35:0] atomicsUnit_io_dtlb_resp_bits_paddr_0; // @[MemBlock.scala 174:27]
  wire  atomicsUnit_io_dtlb_resp_bits_miss; // @[MemBlock.scala 174:27]
  wire  atomicsUnit_io_dtlb_resp_bits_excp_0_pf_ld; // @[MemBlock.scala 174:27]
  wire  atomicsUnit_io_dtlb_resp_bits_excp_0_pf_st; // @[MemBlock.scala 174:27]
  wire  atomicsUnit_io_dtlb_resp_bits_excp_0_af_ld; // @[MemBlock.scala 174:27]
  wire  atomicsUnit_io_dtlb_resp_bits_excp_0_af_st; // @[MemBlock.scala 174:27]
  wire  atomicsUnit_io_dtlb_resp_bits_static_pm_valid; // @[MemBlock.scala 174:27]
  wire  atomicsUnit_io_dtlb_resp_bits_static_pm_bits; // @[MemBlock.scala 174:27]
  wire  atomicsUnit_io_pmpResp_ld; // @[MemBlock.scala 174:27]
  wire  atomicsUnit_io_pmpResp_st; // @[MemBlock.scala 174:27]
  wire  atomicsUnit_io_pmpResp_mmio; // @[MemBlock.scala 174:27]
  wire [3:0] atomicsUnit_io_rsIdx; // @[MemBlock.scala 174:27]
  wire  atomicsUnit_io_flush_sbuffer_valid; // @[MemBlock.scala 174:27]
  wire  atomicsUnit_io_flush_sbuffer_empty; // @[MemBlock.scala 174:27]
  wire  atomicsUnit_io_feedbackSlow_valid; // @[MemBlock.scala 174:27]
  wire [3:0] atomicsUnit_io_feedbackSlow_bits_rsIdx; // @[MemBlock.scala 174:27]
  wire  atomicsUnit_io_redirect_valid; // @[MemBlock.scala 174:27]
  wire  atomicsUnit_io_exceptionAddr_valid; // @[MemBlock.scala 174:27]
  wire [38:0] atomicsUnit_io_exceptionAddr_bits; // @[MemBlock.scala 174:27]
  wire  atomicsUnit_io_csrCtrl_cache_error_enable; // @[MemBlock.scala 174:27]
  wire  atomicsUnit_io_csrCtrl_mem_trigger_t_valid; // @[MemBlock.scala 174:27]
  wire [2:0] atomicsUnit_io_csrCtrl_mem_trigger_t_bits_addr; // @[MemBlock.scala 174:27]
  wire [1:0] atomicsUnit_io_csrCtrl_mem_trigger_t_bits_tdata_matchType; // @[MemBlock.scala 174:27]
  wire  atomicsUnit_io_csrCtrl_mem_trigger_t_bits_tdata_select; // @[MemBlock.scala 174:27]
  wire  atomicsUnit_io_csrCtrl_mem_trigger_t_bits_tdata_chain; // @[MemBlock.scala 174:27]
  wire [63:0] atomicsUnit_io_csrCtrl_mem_trigger_t_bits_tdata_tdata2; // @[MemBlock.scala 174:27]
  wire  atomicsUnit_io_csrCtrl_trigger_enable_2; // @[MemBlock.scala 174:27]
  wire  atomicsUnit_io_csrCtrl_trigger_enable_3; // @[MemBlock.scala 174:27]
  wire  atomicsUnit_io_csrCtrl_trigger_enable_4; // @[MemBlock.scala 174:27]
  wire  atomicsUnit_io_csrCtrl_trigger_enable_5; // @[MemBlock.scala 174:27]
  wire  atomicsUnit_io_csrCtrl_trigger_enable_7; // @[MemBlock.scala 174:27]
  wire  atomicsUnit_io_csrCtrl_trigger_enable_9; // @[MemBlock.scala 174:27]
  wire  vlflowqueue_clock; // @[MemBlock.scala 226:27]
  wire  vlflowqueue_reset; // @[MemBlock.scala 226:27]
  wire  vlflowqueue_io_loadRegIn_0_valid; // @[MemBlock.scala 226:27]
  wire [4:0] vlflowqueue_io_loadRegIn_0_bits_uop_robIdx_value; // @[MemBlock.scala 226:27]
  wire [38:0] vlflowqueue_io_loadRegIn_0_bits_baseaddr; // @[MemBlock.scala 226:27]
  wire  vlflowqueue_io_loadRegIn_1_valid; // @[MemBlock.scala 226:27]
  wire [4:0] vlflowqueue_io_loadRegIn_1_bits_uop_robIdx_value; // @[MemBlock.scala 226:27]
  wire [38:0] vlflowqueue_io_loadRegIn_1_bits_baseaddr; // @[MemBlock.scala 226:27]
  wire  vlflowqueue_io_loadPipeOut_0_ready; // @[MemBlock.scala 226:27]
  wire  vlflowqueue_io_loadPipeOut_0_valid; // @[MemBlock.scala 226:27]
  wire [38:0] vlflowqueue_io_loadPipeOut_0_bits_vaddr; // @[MemBlock.scala 226:27]
  wire  vlflowqueue_io_loadPipeOut_1_ready; // @[MemBlock.scala 226:27]
  wire  vlflowqueue_io_loadPipeOut_1_valid; // @[MemBlock.scala 226:27]
  wire [38:0] vlflowqueue_io_loadPipeOut_1_bits_vaddr; // @[MemBlock.scala 226:27]
  wire  vlExcSignal_clock; // @[MemBlock.scala 228:27]
  wire  vlExcSignal_reset; // @[MemBlock.scala 228:27]
  wire  vlExcSignal_io_vecloadRegIn_0_valid; // @[MemBlock.scala 228:27]
  wire [4:0] vlExcSignal_io_vecloadRegIn_0_bits_uop_robIdx_value; // @[MemBlock.scala 228:27]
  wire [38:0] vlExcSignal_io_vecloadRegIn_0_bits_baseaddr; // @[MemBlock.scala 228:27]
  wire  vlExcSignal_io_vecloadRegIn_1_valid; // @[MemBlock.scala 228:27]
  wire [4:0] vlExcSignal_io_vecloadRegIn_1_bits_uop_robIdx_value; // @[MemBlock.scala 228:27]
  wire [38:0] vlExcSignal_io_vecloadRegIn_1_bits_baseaddr; // @[MemBlock.scala 228:27]
  wire  lsq_clock; // @[MemBlock.scala 231:23]
  wire  lsq_reset; // @[MemBlock.scala 231:23]
  wire  lsq_io_brqRedirect_valid; // @[MemBlock.scala 231:23]
  wire  lsq_io_brqRedirect_bits_robIdx_flag; // @[MemBlock.scala 231:23]
  wire [4:0] lsq_io_brqRedirect_bits_robIdx_value; // @[MemBlock.scala 231:23]
  wire  lsq_io_brqRedirect_bits_level; // @[MemBlock.scala 231:23]
  wire [1:0] lsq_io_enq_needAlloc_0; // @[MemBlock.scala 231:23]
  wire [1:0] lsq_io_enq_needAlloc_1; // @[MemBlock.scala 231:23]
  wire [1:0] lsq_io_enq_needAlloc_2; // @[MemBlock.scala 231:23]
  wire [1:0] lsq_io_enq_needAlloc_3; // @[MemBlock.scala 231:23]
  wire  lsq_io_enq_req_0_valid; // @[MemBlock.scala 231:23]
  wire  lsq_io_enq_req_0_bits_cf_trigger_backendEn_0; // @[MemBlock.scala 231:23]
  wire  lsq_io_enq_req_0_bits_cf_trigger_backendEn_1; // @[MemBlock.scala 231:23]
  wire [6:0] lsq_io_enq_req_0_bits_ctrl_fuOpType; // @[MemBlock.scala 231:23]
  wire  lsq_io_enq_req_0_bits_ctrl_rfWen; // @[MemBlock.scala 231:23]
  wire  lsq_io_enq_req_0_bits_ctrl_fpWen; // @[MemBlock.scala 231:23]
  wire  lsq_io_enq_req_0_bits_ctrl_flushPipe; // @[MemBlock.scala 231:23]
  wire  lsq_io_enq_req_0_bits_ctrl_replayInst; // @[MemBlock.scala 231:23]
  wire [5:0] lsq_io_enq_req_0_bits_pdest; // @[MemBlock.scala 231:23]
  wire  lsq_io_enq_req_0_bits_robIdx_flag; // @[MemBlock.scala 231:23]
  wire [4:0] lsq_io_enq_req_0_bits_robIdx_value; // @[MemBlock.scala 231:23]
  wire [3:0] lsq_io_enq_req_0_bits_lqIdx_value; // @[MemBlock.scala 231:23]
  wire [3:0] lsq_io_enq_req_0_bits_sqIdx_value; // @[MemBlock.scala 231:23]
  wire  lsq_io_enq_req_1_valid; // @[MemBlock.scala 231:23]
  wire  lsq_io_enq_req_1_bits_cf_trigger_backendEn_0; // @[MemBlock.scala 231:23]
  wire  lsq_io_enq_req_1_bits_cf_trigger_backendEn_1; // @[MemBlock.scala 231:23]
  wire [6:0] lsq_io_enq_req_1_bits_ctrl_fuOpType; // @[MemBlock.scala 231:23]
  wire  lsq_io_enq_req_1_bits_ctrl_rfWen; // @[MemBlock.scala 231:23]
  wire  lsq_io_enq_req_1_bits_ctrl_fpWen; // @[MemBlock.scala 231:23]
  wire  lsq_io_enq_req_1_bits_ctrl_flushPipe; // @[MemBlock.scala 231:23]
  wire  lsq_io_enq_req_1_bits_ctrl_replayInst; // @[MemBlock.scala 231:23]
  wire [5:0] lsq_io_enq_req_1_bits_pdest; // @[MemBlock.scala 231:23]
  wire  lsq_io_enq_req_1_bits_robIdx_flag; // @[MemBlock.scala 231:23]
  wire [4:0] lsq_io_enq_req_1_bits_robIdx_value; // @[MemBlock.scala 231:23]
  wire [3:0] lsq_io_enq_req_1_bits_lqIdx_value; // @[MemBlock.scala 231:23]
  wire [3:0] lsq_io_enq_req_1_bits_sqIdx_value; // @[MemBlock.scala 231:23]
  wire  lsq_io_enq_req_2_valid; // @[MemBlock.scala 231:23]
  wire  lsq_io_enq_req_2_bits_cf_trigger_backendEn_0; // @[MemBlock.scala 231:23]
  wire  lsq_io_enq_req_2_bits_cf_trigger_backendEn_1; // @[MemBlock.scala 231:23]
  wire [6:0] lsq_io_enq_req_2_bits_ctrl_fuOpType; // @[MemBlock.scala 231:23]
  wire  lsq_io_enq_req_2_bits_ctrl_rfWen; // @[MemBlock.scala 231:23]
  wire  lsq_io_enq_req_2_bits_ctrl_fpWen; // @[MemBlock.scala 231:23]
  wire  lsq_io_enq_req_2_bits_ctrl_flushPipe; // @[MemBlock.scala 231:23]
  wire  lsq_io_enq_req_2_bits_ctrl_replayInst; // @[MemBlock.scala 231:23]
  wire [5:0] lsq_io_enq_req_2_bits_pdest; // @[MemBlock.scala 231:23]
  wire  lsq_io_enq_req_2_bits_robIdx_flag; // @[MemBlock.scala 231:23]
  wire [4:0] lsq_io_enq_req_2_bits_robIdx_value; // @[MemBlock.scala 231:23]
  wire [3:0] lsq_io_enq_req_2_bits_lqIdx_value; // @[MemBlock.scala 231:23]
  wire [3:0] lsq_io_enq_req_2_bits_sqIdx_value; // @[MemBlock.scala 231:23]
  wire  lsq_io_enq_req_3_valid; // @[MemBlock.scala 231:23]
  wire  lsq_io_enq_req_3_bits_cf_trigger_backendEn_0; // @[MemBlock.scala 231:23]
  wire  lsq_io_enq_req_3_bits_cf_trigger_backendEn_1; // @[MemBlock.scala 231:23]
  wire [6:0] lsq_io_enq_req_3_bits_ctrl_fuOpType; // @[MemBlock.scala 231:23]
  wire  lsq_io_enq_req_3_bits_ctrl_rfWen; // @[MemBlock.scala 231:23]
  wire  lsq_io_enq_req_3_bits_ctrl_fpWen; // @[MemBlock.scala 231:23]
  wire  lsq_io_enq_req_3_bits_ctrl_flushPipe; // @[MemBlock.scala 231:23]
  wire  lsq_io_enq_req_3_bits_ctrl_replayInst; // @[MemBlock.scala 231:23]
  wire [5:0] lsq_io_enq_req_3_bits_pdest; // @[MemBlock.scala 231:23]
  wire  lsq_io_enq_req_3_bits_robIdx_flag; // @[MemBlock.scala 231:23]
  wire [4:0] lsq_io_enq_req_3_bits_robIdx_value; // @[MemBlock.scala 231:23]
  wire [3:0] lsq_io_enq_req_3_bits_lqIdx_value; // @[MemBlock.scala 231:23]
  wire [3:0] lsq_io_enq_req_3_bits_sqIdx_value; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s2_storeLoadViolationQuery_0_req_valid; // @[MemBlock.scala 231:23]
  wire [9:0] lsq_io_ldu_s2_storeLoadViolationQuery_0_req_bits_uop_cf_foldpc; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s2_storeLoadViolationQuery_0_req_bits_uop_cf_ftqPtr_flag; // @[MemBlock.scala 231:23]
  wire [2:0] lsq_io_ldu_s2_storeLoadViolationQuery_0_req_bits_uop_cf_ftqPtr_value; // @[MemBlock.scala 231:23]
  wire [2:0] lsq_io_ldu_s2_storeLoadViolationQuery_0_req_bits_uop_cf_ftqOffset; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s2_storeLoadViolationQuery_0_req_bits_uop_robIdx_flag; // @[MemBlock.scala 231:23]
  wire [4:0] lsq_io_ldu_s2_storeLoadViolationQuery_0_req_bits_uop_robIdx_value; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s2_storeLoadViolationQuery_0_req_bits_uop_sqIdx_flag; // @[MemBlock.scala 231:23]
  wire [3:0] lsq_io_ldu_s2_storeLoadViolationQuery_0_req_bits_uop_sqIdx_value; // @[MemBlock.scala 231:23]
  wire [2:0] lsq_io_ldu_s2_storeLoadViolationQuery_0_req_bits_index; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s2_storeLoadViolationQuery_0_req_bits_allocated; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s2_storeLoadViolationQuery_0_req_bits_datavalid; // @[MemBlock.scala 231:23]
  wire [7:0] lsq_io_ldu_s2_storeLoadViolationQuery_0_req_bits_mask; // @[MemBlock.scala 231:23]
  wire [35:0] lsq_io_ldu_s2_storeLoadViolationQuery_0_req_bits_paddr; // @[MemBlock.scala 231:23]
  wire [2:0] lsq_io_ldu_s2_storeLoadViolationQuery_0_resp_bits_index; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s2_storeLoadViolationQuery_0_resp_bits_canAccept; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s2_storeLoadViolationQuery_0_resp_bits_allocated; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s2_storeLoadViolationQuery_1_req_valid; // @[MemBlock.scala 231:23]
  wire [9:0] lsq_io_ldu_s2_storeLoadViolationQuery_1_req_bits_uop_cf_foldpc; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s2_storeLoadViolationQuery_1_req_bits_uop_cf_ftqPtr_flag; // @[MemBlock.scala 231:23]
  wire [2:0] lsq_io_ldu_s2_storeLoadViolationQuery_1_req_bits_uop_cf_ftqPtr_value; // @[MemBlock.scala 231:23]
  wire [2:0] lsq_io_ldu_s2_storeLoadViolationQuery_1_req_bits_uop_cf_ftqOffset; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s2_storeLoadViolationQuery_1_req_bits_uop_robIdx_flag; // @[MemBlock.scala 231:23]
  wire [4:0] lsq_io_ldu_s2_storeLoadViolationQuery_1_req_bits_uop_robIdx_value; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s2_storeLoadViolationQuery_1_req_bits_uop_sqIdx_flag; // @[MemBlock.scala 231:23]
  wire [3:0] lsq_io_ldu_s2_storeLoadViolationQuery_1_req_bits_uop_sqIdx_value; // @[MemBlock.scala 231:23]
  wire [2:0] lsq_io_ldu_s2_storeLoadViolationQuery_1_req_bits_index; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s2_storeLoadViolationQuery_1_req_bits_allocated; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s2_storeLoadViolationQuery_1_req_bits_datavalid; // @[MemBlock.scala 231:23]
  wire [7:0] lsq_io_ldu_s2_storeLoadViolationQuery_1_req_bits_mask; // @[MemBlock.scala 231:23]
  wire [35:0] lsq_io_ldu_s2_storeLoadViolationQuery_1_req_bits_paddr; // @[MemBlock.scala 231:23]
  wire [2:0] lsq_io_ldu_s2_storeLoadViolationQuery_1_resp_bits_index; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s2_storeLoadViolationQuery_1_resp_bits_canAccept; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s2_storeLoadViolationQuery_1_resp_bits_allocated; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s2_loadLoadViolationQuery_0_req_valid; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s2_loadLoadViolationQuery_0_req_bits_uop_robIdx_flag; // @[MemBlock.scala 231:23]
  wire [4:0] lsq_io_ldu_s2_loadLoadViolationQuery_0_req_bits_uop_robIdx_value; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s2_loadLoadViolationQuery_0_req_bits_uop_lqIdx_flag; // @[MemBlock.scala 231:23]
  wire [3:0] lsq_io_ldu_s2_loadLoadViolationQuery_0_req_bits_uop_lqIdx_value; // @[MemBlock.scala 231:23]
  wire [3:0] lsq_io_ldu_s2_loadLoadViolationQuery_0_req_bits_index; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s2_loadLoadViolationQuery_0_req_bits_allocated; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s2_loadLoadViolationQuery_0_req_bits_datavalid; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s2_loadLoadViolationQuery_0_req_bits_miss; // @[MemBlock.scala 231:23]
  wire [35:0] lsq_io_ldu_s2_loadLoadViolationQuery_0_req_bits_paddr; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s2_loadLoadViolationQuery_0_resp_valid; // @[MemBlock.scala 231:23]
  wire [3:0] lsq_io_ldu_s2_loadLoadViolationQuery_0_resp_bits_index; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s2_loadLoadViolationQuery_0_resp_bits_canAccept; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s2_loadLoadViolationQuery_0_resp_bits_allocated; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s2_loadLoadViolationQuery_0_resp_bits_replayFromFetch; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s2_loadLoadViolationQuery_1_req_valid; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s2_loadLoadViolationQuery_1_req_bits_uop_robIdx_flag; // @[MemBlock.scala 231:23]
  wire [4:0] lsq_io_ldu_s2_loadLoadViolationQuery_1_req_bits_uop_robIdx_value; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s2_loadLoadViolationQuery_1_req_bits_uop_lqIdx_flag; // @[MemBlock.scala 231:23]
  wire [3:0] lsq_io_ldu_s2_loadLoadViolationQuery_1_req_bits_uop_lqIdx_value; // @[MemBlock.scala 231:23]
  wire [3:0] lsq_io_ldu_s2_loadLoadViolationQuery_1_req_bits_index; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s2_loadLoadViolationQuery_1_req_bits_allocated; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s2_loadLoadViolationQuery_1_req_bits_datavalid; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s2_loadLoadViolationQuery_1_req_bits_miss; // @[MemBlock.scala 231:23]
  wire [35:0] lsq_io_ldu_s2_loadLoadViolationQuery_1_req_bits_paddr; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s2_loadLoadViolationQuery_1_resp_valid; // @[MemBlock.scala 231:23]
  wire [3:0] lsq_io_ldu_s2_loadLoadViolationQuery_1_resp_bits_index; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s2_loadLoadViolationQuery_1_resp_bits_canAccept; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s2_loadLoadViolationQuery_1_resp_bits_allocated; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s2_loadLoadViolationQuery_1_resp_bits_replayFromFetch; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s3_loadIn_0_valid; // @[MemBlock.scala 231:23]
  wire [9:0] lsq_io_ldu_s3_loadIn_0_bits_uop_cf_foldpc; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s3_loadIn_0_bits_uop_cf_exceptionVec_4; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s3_loadIn_0_bits_uop_cf_exceptionVec_5; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s3_loadIn_0_bits_uop_cf_exceptionVec_13; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s3_loadIn_0_bits_uop_cf_trigger_backendEn_1; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s3_loadIn_0_bits_uop_cf_trigger_backendHit_0; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s3_loadIn_0_bits_uop_cf_trigger_backendHit_1; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s3_loadIn_0_bits_uop_cf_trigger_backendHit_4; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s3_loadIn_0_bits_uop_cf_waitForRobIdx_flag; // @[MemBlock.scala 231:23]
  wire [4:0] lsq_io_ldu_s3_loadIn_0_bits_uop_cf_waitForRobIdx_value; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s3_loadIn_0_bits_uop_cf_loadWaitBit; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s3_loadIn_0_bits_uop_cf_loadWaitStrict; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s3_loadIn_0_bits_uop_cf_ftqPtr_flag; // @[MemBlock.scala 231:23]
  wire [2:0] lsq_io_ldu_s3_loadIn_0_bits_uop_cf_ftqPtr_value; // @[MemBlock.scala 231:23]
  wire [2:0] lsq_io_ldu_s3_loadIn_0_bits_uop_cf_ftqOffset; // @[MemBlock.scala 231:23]
  wire [3:0] lsq_io_ldu_s3_loadIn_0_bits_uop_ctrl_fuType; // @[MemBlock.scala 231:23]
  wire [6:0] lsq_io_ldu_s3_loadIn_0_bits_uop_ctrl_fuOpType; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s3_loadIn_0_bits_uop_ctrl_rfWen; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s3_loadIn_0_bits_uop_ctrl_fpWen; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s3_loadIn_0_bits_uop_ctrl_replayInst; // @[MemBlock.scala 231:23]
  wire [5:0] lsq_io_ldu_s3_loadIn_0_bits_uop_pdest; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s3_loadIn_0_bits_uop_robIdx_flag; // @[MemBlock.scala 231:23]
  wire [4:0] lsq_io_ldu_s3_loadIn_0_bits_uop_robIdx_value; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s3_loadIn_0_bits_uop_lqIdx_flag; // @[MemBlock.scala 231:23]
  wire [3:0] lsq_io_ldu_s3_loadIn_0_bits_uop_lqIdx_value; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s3_loadIn_0_bits_uop_sqIdx_flag; // @[MemBlock.scala 231:23]
  wire [3:0] lsq_io_ldu_s3_loadIn_0_bits_uop_sqIdx_value; // @[MemBlock.scala 231:23]
  wire [38:0] lsq_io_ldu_s3_loadIn_0_bits_vaddr; // @[MemBlock.scala 231:23]
  wire [35:0] lsq_io_ldu_s3_loadIn_0_bits_paddr; // @[MemBlock.scala 231:23]
  wire [15:0] lsq_io_ldu_s3_loadIn_0_bits_mask; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s3_loadIn_0_bits_miss; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s3_loadIn_0_bits_tlbMiss; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s3_loadIn_0_bits_mmio; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s3_loadIn_0_bits_rarAllocated; // @[MemBlock.scala 231:23]
  wire [3:0] lsq_io_ldu_s3_loadIn_0_bits_rarIndex; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s3_loadIn_0_bits_rawAllocated; // @[MemBlock.scala 231:23]
  wire [2:0] lsq_io_ldu_s3_loadIn_0_bits_rawIndex; // @[MemBlock.scala 231:23]
  wire [1:0] lsq_io_ldu_s3_loadIn_0_bits_replayInfo_missMSHRId; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s3_loadIn_0_bits_replayInfo_canForwardFullData; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s3_loadIn_0_bits_replayInfo_dataInvalidSqIdx_flag; // @[MemBlock.scala 231:23]
  wire [3:0] lsq_io_ldu_s3_loadIn_0_bits_replayInfo_dataInvalidSqIdx_value; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s3_loadIn_0_bits_replayInfo_addrInvalidSqIdx_flag; // @[MemBlock.scala 231:23]
  wire [3:0] lsq_io_ldu_s3_loadIn_0_bits_replayInfo_addrInvalidSqIdx_value; // @[MemBlock.scala 231:23]
  wire [7:0] lsq_io_ldu_s3_loadIn_0_bits_replayInfo_replayCarry_real_way_en; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s3_loadIn_0_bits_replayInfo_replayCarry_valid; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s3_loadIn_0_bits_replayInfo_dataInLastBeat; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s3_loadIn_0_bits_replayInfo_cause_0; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s3_loadIn_0_bits_replayInfo_cause_1; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s3_loadIn_0_bits_replayInfo_cause_2; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s3_loadIn_0_bits_replayInfo_cause_3; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s3_loadIn_0_bits_replayInfo_cause_4; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s3_loadIn_0_bits_replayInfo_cause_5; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s3_loadIn_0_bits_replayInfo_cause_6; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s3_loadIn_0_bits_replayInfo_cause_7; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s3_loadIn_0_bits_lqDataWenDup_1; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s3_loadIn_0_bits_lqDataWenDup_2; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s3_loadIn_0_bits_lqDataWenDup_3; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s3_loadIn_0_bits_lqDataWenDup_5; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s3_loadIn_1_valid; // @[MemBlock.scala 231:23]
  wire [9:0] lsq_io_ldu_s3_loadIn_1_bits_uop_cf_foldpc; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s3_loadIn_1_bits_uop_cf_exceptionVec_4; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s3_loadIn_1_bits_uop_cf_exceptionVec_5; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s3_loadIn_1_bits_uop_cf_exceptionVec_13; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s3_loadIn_1_bits_uop_cf_trigger_backendEn_1; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s3_loadIn_1_bits_uop_cf_trigger_backendHit_0; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s3_loadIn_1_bits_uop_cf_trigger_backendHit_1; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s3_loadIn_1_bits_uop_cf_trigger_backendHit_4; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s3_loadIn_1_bits_uop_cf_waitForRobIdx_flag; // @[MemBlock.scala 231:23]
  wire [4:0] lsq_io_ldu_s3_loadIn_1_bits_uop_cf_waitForRobIdx_value; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s3_loadIn_1_bits_uop_cf_loadWaitBit; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s3_loadIn_1_bits_uop_cf_loadWaitStrict; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s3_loadIn_1_bits_uop_cf_ftqPtr_flag; // @[MemBlock.scala 231:23]
  wire [2:0] lsq_io_ldu_s3_loadIn_1_bits_uop_cf_ftqPtr_value; // @[MemBlock.scala 231:23]
  wire [2:0] lsq_io_ldu_s3_loadIn_1_bits_uop_cf_ftqOffset; // @[MemBlock.scala 231:23]
  wire [3:0] lsq_io_ldu_s3_loadIn_1_bits_uop_ctrl_fuType; // @[MemBlock.scala 231:23]
  wire [6:0] lsq_io_ldu_s3_loadIn_1_bits_uop_ctrl_fuOpType; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s3_loadIn_1_bits_uop_ctrl_rfWen; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s3_loadIn_1_bits_uop_ctrl_fpWen; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s3_loadIn_1_bits_uop_ctrl_replayInst; // @[MemBlock.scala 231:23]
  wire [5:0] lsq_io_ldu_s3_loadIn_1_bits_uop_pdest; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s3_loadIn_1_bits_uop_robIdx_flag; // @[MemBlock.scala 231:23]
  wire [4:0] lsq_io_ldu_s3_loadIn_1_bits_uop_robIdx_value; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s3_loadIn_1_bits_uop_lqIdx_flag; // @[MemBlock.scala 231:23]
  wire [3:0] lsq_io_ldu_s3_loadIn_1_bits_uop_lqIdx_value; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s3_loadIn_1_bits_uop_sqIdx_flag; // @[MemBlock.scala 231:23]
  wire [3:0] lsq_io_ldu_s3_loadIn_1_bits_uop_sqIdx_value; // @[MemBlock.scala 231:23]
  wire [38:0] lsq_io_ldu_s3_loadIn_1_bits_vaddr; // @[MemBlock.scala 231:23]
  wire [35:0] lsq_io_ldu_s3_loadIn_1_bits_paddr; // @[MemBlock.scala 231:23]
  wire [15:0] lsq_io_ldu_s3_loadIn_1_bits_mask; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s3_loadIn_1_bits_miss; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s3_loadIn_1_bits_tlbMiss; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s3_loadIn_1_bits_mmio; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s3_loadIn_1_bits_rarAllocated; // @[MemBlock.scala 231:23]
  wire [3:0] lsq_io_ldu_s3_loadIn_1_bits_rarIndex; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s3_loadIn_1_bits_rawAllocated; // @[MemBlock.scala 231:23]
  wire [2:0] lsq_io_ldu_s3_loadIn_1_bits_rawIndex; // @[MemBlock.scala 231:23]
  wire [1:0] lsq_io_ldu_s3_loadIn_1_bits_replayInfo_missMSHRId; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s3_loadIn_1_bits_replayInfo_canForwardFullData; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s3_loadIn_1_bits_replayInfo_dataInvalidSqIdx_flag; // @[MemBlock.scala 231:23]
  wire [3:0] lsq_io_ldu_s3_loadIn_1_bits_replayInfo_dataInvalidSqIdx_value; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s3_loadIn_1_bits_replayInfo_addrInvalidSqIdx_flag; // @[MemBlock.scala 231:23]
  wire [3:0] lsq_io_ldu_s3_loadIn_1_bits_replayInfo_addrInvalidSqIdx_value; // @[MemBlock.scala 231:23]
  wire [7:0] lsq_io_ldu_s3_loadIn_1_bits_replayInfo_replayCarry_real_way_en; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s3_loadIn_1_bits_replayInfo_replayCarry_valid; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s3_loadIn_1_bits_replayInfo_dataInLastBeat; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s3_loadIn_1_bits_replayInfo_cause_0; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s3_loadIn_1_bits_replayInfo_cause_1; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s3_loadIn_1_bits_replayInfo_cause_2; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s3_loadIn_1_bits_replayInfo_cause_3; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s3_loadIn_1_bits_replayInfo_cause_4; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s3_loadIn_1_bits_replayInfo_cause_5; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s3_loadIn_1_bits_replayInfo_cause_6; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s3_loadIn_1_bits_replayInfo_cause_7; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s3_loadIn_1_bits_lqDataWenDup_1; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s3_loadIn_1_bits_lqDataWenDup_2; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s3_loadIn_1_bits_lqDataWenDup_3; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldu_s3_loadIn_1_bits_lqDataWenDup_5; // @[MemBlock.scala 231:23]
  wire  lsq_io_sta_s0_storeMaskIn_0_valid; // @[MemBlock.scala 231:23]
  wire [3:0] lsq_io_sta_s0_storeMaskIn_0_bits_sqIdx_value; // @[MemBlock.scala 231:23]
  wire [15:0] lsq_io_sta_s0_storeMaskIn_0_bits_mask; // @[MemBlock.scala 231:23]
  wire  lsq_io_sta_s0_storeMaskIn_1_valid; // @[MemBlock.scala 231:23]
  wire [3:0] lsq_io_sta_s0_storeMaskIn_1_bits_sqIdx_value; // @[MemBlock.scala 231:23]
  wire [15:0] lsq_io_sta_s0_storeMaskIn_1_bits_mask; // @[MemBlock.scala 231:23]
  wire  lsq_io_sta_s1_storeAddrIn_0_valid; // @[MemBlock.scala 231:23]
  wire [2:0] lsq_io_sta_s1_storeAddrIn_0_bits_uop_cf_ftqPtr_value; // @[MemBlock.scala 231:23]
  wire [2:0] lsq_io_sta_s1_storeAddrIn_0_bits_uop_cf_ftqOffset; // @[MemBlock.scala 231:23]
  wire [6:0] lsq_io_sta_s1_storeAddrIn_0_bits_uop_ctrl_fuOpType; // @[MemBlock.scala 231:23]
  wire  lsq_io_sta_s1_storeAddrIn_0_bits_uop_robIdx_flag; // @[MemBlock.scala 231:23]
  wire [4:0] lsq_io_sta_s1_storeAddrIn_0_bits_uop_robIdx_value; // @[MemBlock.scala 231:23]
  wire  lsq_io_sta_s1_storeAddrIn_0_bits_uop_sqIdx_flag; // @[MemBlock.scala 231:23]
  wire [3:0] lsq_io_sta_s1_storeAddrIn_0_bits_uop_sqIdx_value; // @[MemBlock.scala 231:23]
  wire [38:0] lsq_io_sta_s1_storeAddrIn_0_bits_vaddr; // @[MemBlock.scala 231:23]
  wire [35:0] lsq_io_sta_s1_storeAddrIn_0_bits_paddr; // @[MemBlock.scala 231:23]
  wire [15:0] lsq_io_sta_s1_storeAddrIn_0_bits_mask; // @[MemBlock.scala 231:23]
  wire  lsq_io_sta_s1_storeAddrIn_0_bits_wlineflag; // @[MemBlock.scala 231:23]
  wire  lsq_io_sta_s1_storeAddrIn_0_bits_miss; // @[MemBlock.scala 231:23]
  wire  lsq_io_sta_s1_storeAddrIn_1_valid; // @[MemBlock.scala 231:23]
  wire [2:0] lsq_io_sta_s1_storeAddrIn_1_bits_uop_cf_ftqPtr_value; // @[MemBlock.scala 231:23]
  wire [2:0] lsq_io_sta_s1_storeAddrIn_1_bits_uop_cf_ftqOffset; // @[MemBlock.scala 231:23]
  wire [6:0] lsq_io_sta_s1_storeAddrIn_1_bits_uop_ctrl_fuOpType; // @[MemBlock.scala 231:23]
  wire  lsq_io_sta_s1_storeAddrIn_1_bits_uop_robIdx_flag; // @[MemBlock.scala 231:23]
  wire [4:0] lsq_io_sta_s1_storeAddrIn_1_bits_uop_robIdx_value; // @[MemBlock.scala 231:23]
  wire  lsq_io_sta_s1_storeAddrIn_1_bits_uop_sqIdx_flag; // @[MemBlock.scala 231:23]
  wire [3:0] lsq_io_sta_s1_storeAddrIn_1_bits_uop_sqIdx_value; // @[MemBlock.scala 231:23]
  wire [38:0] lsq_io_sta_s1_storeAddrIn_1_bits_vaddr; // @[MemBlock.scala 231:23]
  wire [35:0] lsq_io_sta_s1_storeAddrIn_1_bits_paddr; // @[MemBlock.scala 231:23]
  wire [15:0] lsq_io_sta_s1_storeAddrIn_1_bits_mask; // @[MemBlock.scala 231:23]
  wire  lsq_io_sta_s1_storeAddrIn_1_bits_wlineflag; // @[MemBlock.scala 231:23]
  wire  lsq_io_sta_s1_storeAddrIn_1_bits_miss; // @[MemBlock.scala 231:23]
  wire  lsq_io_sta_s2_storeAddrInRe_0_mmio; // @[MemBlock.scala 231:23]
  wire  lsq_io_sta_s2_storeAddrInRe_0_atomic; // @[MemBlock.scala 231:23]
  wire  lsq_io_sta_s2_storeAddrInRe_1_mmio; // @[MemBlock.scala 231:23]
  wire  lsq_io_sta_s2_storeAddrInRe_1_atomic; // @[MemBlock.scala 231:23]
  wire  lsq_io_std_s0_storeDataIn_0_valid; // @[MemBlock.scala 231:23]
  wire [6:0] lsq_io_std_s0_storeDataIn_0_bits_uop_ctrl_fuOpType; // @[MemBlock.scala 231:23]
  wire  lsq_io_std_s0_storeDataIn_0_bits_uop_sqIdx_flag; // @[MemBlock.scala 231:23]
  wire [3:0] lsq_io_std_s0_storeDataIn_0_bits_uop_sqIdx_value; // @[MemBlock.scala 231:23]
  wire [63:0] lsq_io_std_s0_storeDataIn_0_bits_data; // @[MemBlock.scala 231:23]
  wire  lsq_io_std_s0_storeDataIn_1_valid; // @[MemBlock.scala 231:23]
  wire [6:0] lsq_io_std_s0_storeDataIn_1_bits_uop_ctrl_fuOpType; // @[MemBlock.scala 231:23]
  wire  lsq_io_std_s0_storeDataIn_1_bits_uop_sqIdx_flag; // @[MemBlock.scala 231:23]
  wire [3:0] lsq_io_std_s0_storeDataIn_1_bits_uop_sqIdx_value; // @[MemBlock.scala 231:23]
  wire [63:0] lsq_io_std_s0_storeDataIn_1_bits_data; // @[MemBlock.scala 231:23]
  wire  lsq_io_loadOut_0_ready; // @[MemBlock.scala 231:23]
  wire  lsq_io_loadOut_0_valid; // @[MemBlock.scala 231:23]
  wire  lsq_io_loadOut_0_bits_uop_cf_exceptionVec_4; // @[MemBlock.scala 231:23]
  wire  lsq_io_loadOut_0_bits_uop_cf_exceptionVec_5; // @[MemBlock.scala 231:23]
  wire  lsq_io_loadOut_0_bits_uop_cf_exceptionVec_13; // @[MemBlock.scala 231:23]
  wire  lsq_io_loadOut_0_bits_uop_cf_trigger_backendEn_1; // @[MemBlock.scala 231:23]
  wire  lsq_io_loadOut_0_bits_uop_cf_trigger_backendHit_0; // @[MemBlock.scala 231:23]
  wire  lsq_io_loadOut_0_bits_uop_cf_trigger_backendHit_1; // @[MemBlock.scala 231:23]
  wire  lsq_io_loadOut_0_bits_uop_cf_trigger_backendHit_4; // @[MemBlock.scala 231:23]
  wire  lsq_io_loadOut_0_bits_uop_ctrl_rfWen; // @[MemBlock.scala 231:23]
  wire  lsq_io_loadOut_0_bits_uop_ctrl_fpWen; // @[MemBlock.scala 231:23]
  wire  lsq_io_loadOut_0_bits_uop_ctrl_flushPipe; // @[MemBlock.scala 231:23]
  wire  lsq_io_loadOut_0_bits_uop_ctrl_replayInst; // @[MemBlock.scala 231:23]
  wire [5:0] lsq_io_loadOut_0_bits_uop_pdest; // @[MemBlock.scala 231:23]
  wire  lsq_io_loadOut_0_bits_uop_robIdx_flag; // @[MemBlock.scala 231:23]
  wire [4:0] lsq_io_loadOut_0_bits_uop_robIdx_value; // @[MemBlock.scala 231:23]
  wire [63:0] lsq_io_ldRawDataOut_0_lqData; // @[MemBlock.scala 231:23]
  wire [6:0] lsq_io_ldRawDataOut_0_uop_ctrl_fuOpType; // @[MemBlock.scala 231:23]
  wire  lsq_io_ldRawDataOut_0_uop_ctrl_fpWen; // @[MemBlock.scala 231:23]
  wire [2:0] lsq_io_ldRawDataOut_0_addrOffset; // @[MemBlock.scala 231:23]
  wire  lsq_io_replay_0_ready; // @[MemBlock.scala 231:23]
  wire  lsq_io_replay_0_valid; // @[MemBlock.scala 231:23]
  wire [9:0] lsq_io_replay_0_bits_uop_cf_foldpc; // @[MemBlock.scala 231:23]
  wire  lsq_io_replay_0_bits_uop_cf_trigger_backendEn_1; // @[MemBlock.scala 231:23]
  wire  lsq_io_replay_0_bits_uop_cf_trigger_backendHit_0; // @[MemBlock.scala 231:23]
  wire  lsq_io_replay_0_bits_uop_cf_trigger_backendHit_1; // @[MemBlock.scala 231:23]
  wire  lsq_io_replay_0_bits_uop_cf_trigger_backendHit_4; // @[MemBlock.scala 231:23]
  wire  lsq_io_replay_0_bits_uop_cf_waitForRobIdx_flag; // @[MemBlock.scala 231:23]
  wire [4:0] lsq_io_replay_0_bits_uop_cf_waitForRobIdx_value; // @[MemBlock.scala 231:23]
  wire  lsq_io_replay_0_bits_uop_cf_loadWaitBit; // @[MemBlock.scala 231:23]
  wire  lsq_io_replay_0_bits_uop_cf_loadWaitStrict; // @[MemBlock.scala 231:23]
  wire  lsq_io_replay_0_bits_uop_cf_ftqPtr_flag; // @[MemBlock.scala 231:23]
  wire [2:0] lsq_io_replay_0_bits_uop_cf_ftqPtr_value; // @[MemBlock.scala 231:23]
  wire [2:0] lsq_io_replay_0_bits_uop_cf_ftqOffset; // @[MemBlock.scala 231:23]
  wire [3:0] lsq_io_replay_0_bits_uop_ctrl_fuType; // @[MemBlock.scala 231:23]
  wire [6:0] lsq_io_replay_0_bits_uop_ctrl_fuOpType; // @[MemBlock.scala 231:23]
  wire  lsq_io_replay_0_bits_uop_ctrl_rfWen; // @[MemBlock.scala 231:23]
  wire  lsq_io_replay_0_bits_uop_ctrl_fpWen; // @[MemBlock.scala 231:23]
  wire [5:0] lsq_io_replay_0_bits_uop_pdest; // @[MemBlock.scala 231:23]
  wire  lsq_io_replay_0_bits_uop_robIdx_flag; // @[MemBlock.scala 231:23]
  wire [4:0] lsq_io_replay_0_bits_uop_robIdx_value; // @[MemBlock.scala 231:23]
  wire  lsq_io_replay_0_bits_uop_lqIdx_flag; // @[MemBlock.scala 231:23]
  wire [3:0] lsq_io_replay_0_bits_uop_lqIdx_value; // @[MemBlock.scala 231:23]
  wire  lsq_io_replay_0_bits_uop_sqIdx_flag; // @[MemBlock.scala 231:23]
  wire [3:0] lsq_io_replay_0_bits_uop_sqIdx_value; // @[MemBlock.scala 231:23]
  wire [38:0] lsq_io_replay_0_bits_vaddr; // @[MemBlock.scala 231:23]
  wire  lsq_io_replay_0_bits_isFirstIssue; // @[MemBlock.scala 231:23]
  wire [7:0] lsq_io_replay_0_bits_replayCarry_real_way_en; // @[MemBlock.scala 231:23]
  wire  lsq_io_replay_0_bits_replayCarry_valid; // @[MemBlock.scala 231:23]
  wire [1:0] lsq_io_replay_0_bits_mshrid; // @[MemBlock.scala 231:23]
  wire  lsq_io_replay_0_bits_forward_tlDchannel; // @[MemBlock.scala 231:23]
  wire  lsq_io_replay_0_bits_rarAllocated; // @[MemBlock.scala 231:23]
  wire [3:0] lsq_io_replay_0_bits_rarIndex; // @[MemBlock.scala 231:23]
  wire  lsq_io_replay_0_bits_rawAllocated; // @[MemBlock.scala 231:23]
  wire [2:0] lsq_io_replay_0_bits_rawIndex; // @[MemBlock.scala 231:23]
  wire  lsq_io_replay_1_ready; // @[MemBlock.scala 231:23]
  wire  lsq_io_replay_1_valid; // @[MemBlock.scala 231:23]
  wire [9:0] lsq_io_replay_1_bits_uop_cf_foldpc; // @[MemBlock.scala 231:23]
  wire  lsq_io_replay_1_bits_uop_cf_trigger_backendEn_1; // @[MemBlock.scala 231:23]
  wire  lsq_io_replay_1_bits_uop_cf_trigger_backendHit_0; // @[MemBlock.scala 231:23]
  wire  lsq_io_replay_1_bits_uop_cf_trigger_backendHit_1; // @[MemBlock.scala 231:23]
  wire  lsq_io_replay_1_bits_uop_cf_trigger_backendHit_4; // @[MemBlock.scala 231:23]
  wire  lsq_io_replay_1_bits_uop_cf_waitForRobIdx_flag; // @[MemBlock.scala 231:23]
  wire [4:0] lsq_io_replay_1_bits_uop_cf_waitForRobIdx_value; // @[MemBlock.scala 231:23]
  wire  lsq_io_replay_1_bits_uop_cf_loadWaitBit; // @[MemBlock.scala 231:23]
  wire  lsq_io_replay_1_bits_uop_cf_loadWaitStrict; // @[MemBlock.scala 231:23]
  wire  lsq_io_replay_1_bits_uop_cf_ftqPtr_flag; // @[MemBlock.scala 231:23]
  wire [2:0] lsq_io_replay_1_bits_uop_cf_ftqPtr_value; // @[MemBlock.scala 231:23]
  wire [2:0] lsq_io_replay_1_bits_uop_cf_ftqOffset; // @[MemBlock.scala 231:23]
  wire [3:0] lsq_io_replay_1_bits_uop_ctrl_fuType; // @[MemBlock.scala 231:23]
  wire [6:0] lsq_io_replay_1_bits_uop_ctrl_fuOpType; // @[MemBlock.scala 231:23]
  wire  lsq_io_replay_1_bits_uop_ctrl_rfWen; // @[MemBlock.scala 231:23]
  wire  lsq_io_replay_1_bits_uop_ctrl_fpWen; // @[MemBlock.scala 231:23]
  wire [5:0] lsq_io_replay_1_bits_uop_pdest; // @[MemBlock.scala 231:23]
  wire  lsq_io_replay_1_bits_uop_robIdx_flag; // @[MemBlock.scala 231:23]
  wire [4:0] lsq_io_replay_1_bits_uop_robIdx_value; // @[MemBlock.scala 231:23]
  wire  lsq_io_replay_1_bits_uop_lqIdx_flag; // @[MemBlock.scala 231:23]
  wire [3:0] lsq_io_replay_1_bits_uop_lqIdx_value; // @[MemBlock.scala 231:23]
  wire  lsq_io_replay_1_bits_uop_sqIdx_flag; // @[MemBlock.scala 231:23]
  wire [3:0] lsq_io_replay_1_bits_uop_sqIdx_value; // @[MemBlock.scala 231:23]
  wire [38:0] lsq_io_replay_1_bits_vaddr; // @[MemBlock.scala 231:23]
  wire  lsq_io_replay_1_bits_isFirstIssue; // @[MemBlock.scala 231:23]
  wire [7:0] lsq_io_replay_1_bits_replayCarry_real_way_en; // @[MemBlock.scala 231:23]
  wire  lsq_io_replay_1_bits_replayCarry_valid; // @[MemBlock.scala 231:23]
  wire [1:0] lsq_io_replay_1_bits_mshrid; // @[MemBlock.scala 231:23]
  wire  lsq_io_replay_1_bits_forward_tlDchannel; // @[MemBlock.scala 231:23]
  wire  lsq_io_replay_1_bits_rarAllocated; // @[MemBlock.scala 231:23]
  wire [3:0] lsq_io_replay_1_bits_rarIndex; // @[MemBlock.scala 231:23]
  wire  lsq_io_replay_1_bits_rawAllocated; // @[MemBlock.scala 231:23]
  wire [2:0] lsq_io_replay_1_bits_rawIndex; // @[MemBlock.scala 231:23]
  wire  lsq_io_sbuffer_0_ready; // @[MemBlock.scala 231:23]
  wire  lsq_io_sbuffer_0_valid; // @[MemBlock.scala 231:23]
  wire [35:0] lsq_io_sbuffer_0_bits_addr; // @[MemBlock.scala 231:23]
  wire [127:0] lsq_io_sbuffer_0_bits_data; // @[MemBlock.scala 231:23]
  wire [15:0] lsq_io_sbuffer_0_bits_mask; // @[MemBlock.scala 231:23]
  wire [38:0] lsq_io_sbuffer_0_bits_vaddr; // @[MemBlock.scala 231:23]
  wire  lsq_io_sbuffer_0_bits_wline; // @[MemBlock.scala 231:23]
  wire  lsq_io_sbuffer_1_ready; // @[MemBlock.scala 231:23]
  wire  lsq_io_sbuffer_1_valid; // @[MemBlock.scala 231:23]
  wire [35:0] lsq_io_sbuffer_1_bits_addr; // @[MemBlock.scala 231:23]
  wire [127:0] lsq_io_sbuffer_1_bits_data; // @[MemBlock.scala 231:23]
  wire [15:0] lsq_io_sbuffer_1_bits_mask; // @[MemBlock.scala 231:23]
  wire [38:0] lsq_io_sbuffer_1_bits_vaddr; // @[MemBlock.scala 231:23]
  wire  lsq_io_sbuffer_1_bits_wline; // @[MemBlock.scala 231:23]
  wire [38:0] lsq_io_forward_0_vaddr; // @[MemBlock.scala 231:23]
  wire [35:0] lsq_io_forward_0_paddr; // @[MemBlock.scala 231:23]
  wire  lsq_io_forward_0_uop_cf_waitForRobIdx_flag; // @[MemBlock.scala 231:23]
  wire [4:0] lsq_io_forward_0_uop_cf_waitForRobIdx_value; // @[MemBlock.scala 231:23]
  wire  lsq_io_forward_0_uop_sqIdx_flag; // @[MemBlock.scala 231:23]
  wire [3:0] lsq_io_forward_0_uop_sqIdx_value; // @[MemBlock.scala 231:23]
  wire  lsq_io_forward_0_valid; // @[MemBlock.scala 231:23]
  wire  lsq_io_forward_0_forwardMask_0; // @[MemBlock.scala 231:23]
  wire  lsq_io_forward_0_forwardMask_1; // @[MemBlock.scala 231:23]
  wire  lsq_io_forward_0_forwardMask_2; // @[MemBlock.scala 231:23]
  wire  lsq_io_forward_0_forwardMask_3; // @[MemBlock.scala 231:23]
  wire  lsq_io_forward_0_forwardMask_4; // @[MemBlock.scala 231:23]
  wire  lsq_io_forward_0_forwardMask_5; // @[MemBlock.scala 231:23]
  wire  lsq_io_forward_0_forwardMask_6; // @[MemBlock.scala 231:23]
  wire  lsq_io_forward_0_forwardMask_7; // @[MemBlock.scala 231:23]
  wire  lsq_io_forward_0_forwardMask_8; // @[MemBlock.scala 231:23]
  wire  lsq_io_forward_0_forwardMask_9; // @[MemBlock.scala 231:23]
  wire  lsq_io_forward_0_forwardMask_10; // @[MemBlock.scala 231:23]
  wire  lsq_io_forward_0_forwardMask_11; // @[MemBlock.scala 231:23]
  wire  lsq_io_forward_0_forwardMask_12; // @[MemBlock.scala 231:23]
  wire  lsq_io_forward_0_forwardMask_13; // @[MemBlock.scala 231:23]
  wire  lsq_io_forward_0_forwardMask_14; // @[MemBlock.scala 231:23]
  wire  lsq_io_forward_0_forwardMask_15; // @[MemBlock.scala 231:23]
  wire [7:0] lsq_io_forward_0_forwardData_0; // @[MemBlock.scala 231:23]
  wire [7:0] lsq_io_forward_0_forwardData_1; // @[MemBlock.scala 231:23]
  wire [7:0] lsq_io_forward_0_forwardData_2; // @[MemBlock.scala 231:23]
  wire [7:0] lsq_io_forward_0_forwardData_3; // @[MemBlock.scala 231:23]
  wire [7:0] lsq_io_forward_0_forwardData_4; // @[MemBlock.scala 231:23]
  wire [7:0] lsq_io_forward_0_forwardData_5; // @[MemBlock.scala 231:23]
  wire [7:0] lsq_io_forward_0_forwardData_6; // @[MemBlock.scala 231:23]
  wire [7:0] lsq_io_forward_0_forwardData_7; // @[MemBlock.scala 231:23]
  wire [7:0] lsq_io_forward_0_forwardData_8; // @[MemBlock.scala 231:23]
  wire [7:0] lsq_io_forward_0_forwardData_9; // @[MemBlock.scala 231:23]
  wire [7:0] lsq_io_forward_0_forwardData_10; // @[MemBlock.scala 231:23]
  wire [7:0] lsq_io_forward_0_forwardData_11; // @[MemBlock.scala 231:23]
  wire [7:0] lsq_io_forward_0_forwardData_12; // @[MemBlock.scala 231:23]
  wire [7:0] lsq_io_forward_0_forwardData_13; // @[MemBlock.scala 231:23]
  wire [7:0] lsq_io_forward_0_forwardData_14; // @[MemBlock.scala 231:23]
  wire [7:0] lsq_io_forward_0_forwardData_15; // @[MemBlock.scala 231:23]
  wire  lsq_io_forward_0_sqIdx_flag; // @[MemBlock.scala 231:23]
  wire  lsq_io_forward_0_dataInvalid; // @[MemBlock.scala 231:23]
  wire  lsq_io_forward_0_matchInvalid; // @[MemBlock.scala 231:23]
  wire  lsq_io_forward_0_schedWait; // @[MemBlock.scala 231:23]
  wire [11:0] lsq_io_forward_0_sqIdxMask; // @[MemBlock.scala 231:23]
  wire  lsq_io_forward_0_dataInvalidSqIdx_flag; // @[MemBlock.scala 231:23]
  wire [3:0] lsq_io_forward_0_dataInvalidSqIdx_value; // @[MemBlock.scala 231:23]
  wire  lsq_io_forward_0_addrInvalidSqIdx_flag; // @[MemBlock.scala 231:23]
  wire [3:0] lsq_io_forward_0_addrInvalidSqIdx_value; // @[MemBlock.scala 231:23]
  wire [38:0] lsq_io_forward_1_vaddr; // @[MemBlock.scala 231:23]
  wire [35:0] lsq_io_forward_1_paddr; // @[MemBlock.scala 231:23]
  wire  lsq_io_forward_1_uop_cf_waitForRobIdx_flag; // @[MemBlock.scala 231:23]
  wire [4:0] lsq_io_forward_1_uop_cf_waitForRobIdx_value; // @[MemBlock.scala 231:23]
  wire  lsq_io_forward_1_uop_sqIdx_flag; // @[MemBlock.scala 231:23]
  wire [3:0] lsq_io_forward_1_uop_sqIdx_value; // @[MemBlock.scala 231:23]
  wire  lsq_io_forward_1_valid; // @[MemBlock.scala 231:23]
  wire  lsq_io_forward_1_forwardMask_0; // @[MemBlock.scala 231:23]
  wire  lsq_io_forward_1_forwardMask_1; // @[MemBlock.scala 231:23]
  wire  lsq_io_forward_1_forwardMask_2; // @[MemBlock.scala 231:23]
  wire  lsq_io_forward_1_forwardMask_3; // @[MemBlock.scala 231:23]
  wire  lsq_io_forward_1_forwardMask_4; // @[MemBlock.scala 231:23]
  wire  lsq_io_forward_1_forwardMask_5; // @[MemBlock.scala 231:23]
  wire  lsq_io_forward_1_forwardMask_6; // @[MemBlock.scala 231:23]
  wire  lsq_io_forward_1_forwardMask_7; // @[MemBlock.scala 231:23]
  wire  lsq_io_forward_1_forwardMask_8; // @[MemBlock.scala 231:23]
  wire  lsq_io_forward_1_forwardMask_9; // @[MemBlock.scala 231:23]
  wire  lsq_io_forward_1_forwardMask_10; // @[MemBlock.scala 231:23]
  wire  lsq_io_forward_1_forwardMask_11; // @[MemBlock.scala 231:23]
  wire  lsq_io_forward_1_forwardMask_12; // @[MemBlock.scala 231:23]
  wire  lsq_io_forward_1_forwardMask_13; // @[MemBlock.scala 231:23]
  wire  lsq_io_forward_1_forwardMask_14; // @[MemBlock.scala 231:23]
  wire  lsq_io_forward_1_forwardMask_15; // @[MemBlock.scala 231:23]
  wire [7:0] lsq_io_forward_1_forwardData_0; // @[MemBlock.scala 231:23]
  wire [7:0] lsq_io_forward_1_forwardData_1; // @[MemBlock.scala 231:23]
  wire [7:0] lsq_io_forward_1_forwardData_2; // @[MemBlock.scala 231:23]
  wire [7:0] lsq_io_forward_1_forwardData_3; // @[MemBlock.scala 231:23]
  wire [7:0] lsq_io_forward_1_forwardData_4; // @[MemBlock.scala 231:23]
  wire [7:0] lsq_io_forward_1_forwardData_5; // @[MemBlock.scala 231:23]
  wire [7:0] lsq_io_forward_1_forwardData_6; // @[MemBlock.scala 231:23]
  wire [7:0] lsq_io_forward_1_forwardData_7; // @[MemBlock.scala 231:23]
  wire [7:0] lsq_io_forward_1_forwardData_8; // @[MemBlock.scala 231:23]
  wire [7:0] lsq_io_forward_1_forwardData_9; // @[MemBlock.scala 231:23]
  wire [7:0] lsq_io_forward_1_forwardData_10; // @[MemBlock.scala 231:23]
  wire [7:0] lsq_io_forward_1_forwardData_11; // @[MemBlock.scala 231:23]
  wire [7:0] lsq_io_forward_1_forwardData_12; // @[MemBlock.scala 231:23]
  wire [7:0] lsq_io_forward_1_forwardData_13; // @[MemBlock.scala 231:23]
  wire [7:0] lsq_io_forward_1_forwardData_14; // @[MemBlock.scala 231:23]
  wire [7:0] lsq_io_forward_1_forwardData_15; // @[MemBlock.scala 231:23]
  wire  lsq_io_forward_1_sqIdx_flag; // @[MemBlock.scala 231:23]
  wire  lsq_io_forward_1_dataInvalid; // @[MemBlock.scala 231:23]
  wire  lsq_io_forward_1_matchInvalid; // @[MemBlock.scala 231:23]
  wire  lsq_io_forward_1_schedWait; // @[MemBlock.scala 231:23]
  wire [11:0] lsq_io_forward_1_sqIdxMask; // @[MemBlock.scala 231:23]
  wire  lsq_io_forward_1_dataInvalidSqIdx_flag; // @[MemBlock.scala 231:23]
  wire [3:0] lsq_io_forward_1_dataInvalidSqIdx_value; // @[MemBlock.scala 231:23]
  wire  lsq_io_forward_1_addrInvalidSqIdx_flag; // @[MemBlock.scala 231:23]
  wire [3:0] lsq_io_forward_1_addrInvalidSqIdx_value; // @[MemBlock.scala 231:23]
  wire [1:0] lsq_io_rob_scommit; // @[MemBlock.scala 231:23]
  wire  lsq_io_rob_pendingld; // @[MemBlock.scala 231:23]
  wire  lsq_io_rob_pendingst; // @[MemBlock.scala 231:23]
  wire  lsq_io_rob_commit; // @[MemBlock.scala 231:23]
  wire  lsq_io_rob_isMMIO_0; // @[MemBlock.scala 231:23]
  wire  lsq_io_rob_isMMIO_1; // @[MemBlock.scala 231:23]
  wire [4:0] lsq_io_rob_uop_0_robIdx_value; // @[MemBlock.scala 231:23]
  wire [4:0] lsq_io_rob_uop_1_robIdx_value; // @[MemBlock.scala 231:23]
  wire  lsq_io_rollback_valid; // @[MemBlock.scala 231:23]
  wire  lsq_io_rollback_bits_robIdx_flag; // @[MemBlock.scala 231:23]
  wire [4:0] lsq_io_rollback_bits_robIdx_value; // @[MemBlock.scala 231:23]
  wire  lsq_io_rollback_bits_ftqIdx_flag; // @[MemBlock.scala 231:23]
  wire [2:0] lsq_io_rollback_bits_ftqIdx_value; // @[MemBlock.scala 231:23]
  wire [2:0] lsq_io_rollback_bits_ftqOffset; // @[MemBlock.scala 231:23]
  wire [2:0] lsq_io_rollback_bits_stFtqIdx_value; // @[MemBlock.scala 231:23]
  wire [2:0] lsq_io_rollback_bits_stFtqOffset; // @[MemBlock.scala 231:23]
  wire  lsq_io_correctTableUpdate_valid; // @[MemBlock.scala 231:23]
  wire [9:0] lsq_io_correctTableUpdate_bits_addr; // @[MemBlock.scala 231:23]
  wire  lsq_io_release_valid; // @[MemBlock.scala 231:23]
  wire [35:0] lsq_io_release_bits_paddr; // @[MemBlock.scala 231:23]
  wire  lsq_io_refill_valid; // @[MemBlock.scala 231:23]
  wire [1:0] lsq_io_refill_bits_id; // @[MemBlock.scala 231:23]
  wire  lsq_io_uncacheOutstanding; // @[MemBlock.scala 231:23]
  wire  lsq_io_uncache_req_ready; // @[MemBlock.scala 231:23]
  wire  lsq_io_uncache_req_valid; // @[MemBlock.scala 231:23]
  wire [4:0] lsq_io_uncache_req_bits_cmd; // @[MemBlock.scala 231:23]
  wire [35:0] lsq_io_uncache_req_bits_addr; // @[MemBlock.scala 231:23]
  wire [63:0] lsq_io_uncache_req_bits_data; // @[MemBlock.scala 231:23]
  wire [7:0] lsq_io_uncache_req_bits_mask; // @[MemBlock.scala 231:23]
  wire  lsq_io_uncache_req_bits_atomic; // @[MemBlock.scala 231:23]
  wire  lsq_io_uncache_resp_ready; // @[MemBlock.scala 231:23]
  wire  lsq_io_uncache_resp_valid; // @[MemBlock.scala 231:23]
  wire [63:0] lsq_io_uncache_resp_bits_data; // @[MemBlock.scala 231:23]
  wire  lsq_io_mmioStout_ready; // @[MemBlock.scala 231:23]
  wire  lsq_io_mmioStout_valid; // @[MemBlock.scala 231:23]
  wire  lsq_io_mmioStout_bits_uop_cf_trigger_backendEn_0; // @[MemBlock.scala 231:23]
  wire  lsq_io_mmioStout_bits_uop_robIdx_flag; // @[MemBlock.scala 231:23]
  wire [4:0] lsq_io_mmioStout_bits_uop_robIdx_value; // @[MemBlock.scala 231:23]
  wire  lsq_io_sqEmpty; // @[MemBlock.scala 231:23]
  wire  lsq_io_lqReplayFull; // @[MemBlock.scala 231:23]
  wire [3:0] lsq_io_sqCancelCnt; // @[MemBlock.scala 231:23]
  wire [4:0] lsq_io_lqCancelCnt; // @[MemBlock.scala 231:23]
  wire [1:0] lsq_io_lqDeq; // @[MemBlock.scala 231:23]
  wire [1:0] lsq_io_sqDeq; // @[MemBlock.scala 231:23]
  wire  lsq_io_exceptionAddr_isStore; // @[MemBlock.scala 231:23]
  wire [38:0] lsq_io_exceptionAddr_vaddr; // @[MemBlock.scala 231:23]
  wire  lsq_io_trigger_0_hitLoadAddrTriggerHitVec_0; // @[MemBlock.scala 231:23]
  wire  lsq_io_trigger_0_hitLoadAddrTriggerHitVec_1; // @[MemBlock.scala 231:23]
  wire  lsq_io_trigger_0_hitLoadAddrTriggerHitVec_2; // @[MemBlock.scala 231:23]
  wire  lsq_io_trigger_0_lqLoadAddrTriggerHitVec_0; // @[MemBlock.scala 231:23]
  wire  lsq_io_trigger_0_lqLoadAddrTriggerHitVec_1; // @[MemBlock.scala 231:23]
  wire  lsq_io_trigger_0_lqLoadAddrTriggerHitVec_2; // @[MemBlock.scala 231:23]
  wire  lsq_io_trigger_1_hitLoadAddrTriggerHitVec_0; // @[MemBlock.scala 231:23]
  wire  lsq_io_trigger_1_hitLoadAddrTriggerHitVec_1; // @[MemBlock.scala 231:23]
  wire  lsq_io_trigger_1_hitLoadAddrTriggerHitVec_2; // @[MemBlock.scala 231:23]
  wire [5:0] lsq_io_perf_0_value; // @[MemBlock.scala 231:23]
  wire [5:0] lsq_io_perf_1_value; // @[MemBlock.scala 231:23]
  wire [5:0] lsq_io_perf_2_value; // @[MemBlock.scala 231:23]
  wire [5:0] lsq_io_perf_3_value; // @[MemBlock.scala 231:23]
  wire [5:0] lsq_io_perf_4_value; // @[MemBlock.scala 231:23]
  wire [5:0] lsq_io_perf_5_value; // @[MemBlock.scala 231:23]
  wire [5:0] lsq_io_perf_6_value; // @[MemBlock.scala 231:23]
  wire [5:0] lsq_io_perf_7_value; // @[MemBlock.scala 231:23]
  wire [5:0] lsq_io_perf_8_value; // @[MemBlock.scala 231:23]
  wire [5:0] lsq_io_perf_9_value; // @[MemBlock.scala 231:23]
  wire [5:0] lsq_io_perf_10_value; // @[MemBlock.scala 231:23]
  wire [5:0] lsq_io_perf_11_value; // @[MemBlock.scala 231:23]
  wire [5:0] lsq_io_perf_12_value; // @[MemBlock.scala 231:23]
  wire [5:0] lsq_io_perf_13_value; // @[MemBlock.scala 231:23]
  wire [5:0] lsq_io_perf_14_value; // @[MemBlock.scala 231:23]
  wire [5:0] lsq_io_perf_15_value; // @[MemBlock.scala 231:23]
  wire [5:0] lsq_io_perf_16_value; // @[MemBlock.scala 231:23]
  wire [5:0] lsq_io_perf_17_value; // @[MemBlock.scala 231:23]
  wire [5:0] lsq_io_perf_18_value; // @[MemBlock.scala 231:23]
  wire [5:0] lsq_io_perf_19_value; // @[MemBlock.scala 231:23]
  wire [5:0] lsq_io_perf_20_value; // @[MemBlock.scala 231:23]
  wire [5:0] lsq_io_perf_21_value; // @[MemBlock.scala 231:23]
  wire [5:0] lsq_io_perf_22_value; // @[MemBlock.scala 231:23]
  wire [5:0] lsq_io_perf_23_value; // @[MemBlock.scala 231:23]
  wire [5:0] lsq_io_perf_24_value; // @[MemBlock.scala 231:23]
  wire [5:0] lsq_io_perf_25_value; // @[MemBlock.scala 231:23]
  wire [5:0] lsq_io_perf_26_value; // @[MemBlock.scala 231:23]
  wire [5:0] lsq_io_perf_27_value; // @[MemBlock.scala 231:23]
  wire [5:0] lsq_io_perf_28_value; // @[MemBlock.scala 231:23]
  wire [5:0] lsq_io_perf_29_value; // @[MemBlock.scala 231:23]
  wire  sbuffer_clock; // @[MemBlock.scala 232:23]
  wire  sbuffer_reset; // @[MemBlock.scala 232:23]
  wire  sbuffer_io_in_0_ready; // @[MemBlock.scala 232:23]
  wire  sbuffer_io_in_0_valid; // @[MemBlock.scala 232:23]
  wire [35:0] sbuffer_io_in_0_bits_addr; // @[MemBlock.scala 232:23]
  wire [127:0] sbuffer_io_in_0_bits_data; // @[MemBlock.scala 232:23]
  wire [15:0] sbuffer_io_in_0_bits_mask; // @[MemBlock.scala 232:23]
  wire [38:0] sbuffer_io_in_0_bits_vaddr; // @[MemBlock.scala 232:23]
  wire  sbuffer_io_in_0_bits_wline; // @[MemBlock.scala 232:23]
  wire  sbuffer_io_in_1_ready; // @[MemBlock.scala 232:23]
  wire  sbuffer_io_in_1_valid; // @[MemBlock.scala 232:23]
  wire [35:0] sbuffer_io_in_1_bits_addr; // @[MemBlock.scala 232:23]
  wire [127:0] sbuffer_io_in_1_bits_data; // @[MemBlock.scala 232:23]
  wire [15:0] sbuffer_io_in_1_bits_mask; // @[MemBlock.scala 232:23]
  wire [38:0] sbuffer_io_in_1_bits_vaddr; // @[MemBlock.scala 232:23]
  wire  sbuffer_io_in_1_bits_wline; // @[MemBlock.scala 232:23]
  wire  sbuffer_io_dcache_req_ready; // @[MemBlock.scala 232:23]
  wire  sbuffer_io_dcache_req_valid; // @[MemBlock.scala 232:23]
  wire [38:0] sbuffer_io_dcache_req_bits_vaddr; // @[MemBlock.scala 232:23]
  wire [35:0] sbuffer_io_dcache_req_bits_addr; // @[MemBlock.scala 232:23]
  wire [511:0] sbuffer_io_dcache_req_bits_data; // @[MemBlock.scala 232:23]
  wire [63:0] sbuffer_io_dcache_req_bits_mask; // @[MemBlock.scala 232:23]
  wire [3:0] sbuffer_io_dcache_req_bits_id; // @[MemBlock.scala 232:23]
  wire  sbuffer_io_dcache_main_pipe_hit_resp_valid; // @[MemBlock.scala 232:23]
  wire [3:0] sbuffer_io_dcache_main_pipe_hit_resp_bits_id; // @[MemBlock.scala 232:23]
  wire  sbuffer_io_dcache_refill_hit_resp_valid; // @[MemBlock.scala 232:23]
  wire [3:0] sbuffer_io_dcache_refill_hit_resp_bits_id; // @[MemBlock.scala 232:23]
  wire  sbuffer_io_dcache_replay_resp_valid; // @[MemBlock.scala 232:23]
  wire [3:0] sbuffer_io_dcache_replay_resp_bits_id; // @[MemBlock.scala 232:23]
  wire [38:0] sbuffer_io_forward_0_vaddr; // @[MemBlock.scala 232:23]
  wire [35:0] sbuffer_io_forward_0_paddr; // @[MemBlock.scala 232:23]
  wire  sbuffer_io_forward_0_valid; // @[MemBlock.scala 232:23]
  wire  sbuffer_io_forward_0_forwardMask_0; // @[MemBlock.scala 232:23]
  wire  sbuffer_io_forward_0_forwardMask_1; // @[MemBlock.scala 232:23]
  wire  sbuffer_io_forward_0_forwardMask_2; // @[MemBlock.scala 232:23]
  wire  sbuffer_io_forward_0_forwardMask_3; // @[MemBlock.scala 232:23]
  wire  sbuffer_io_forward_0_forwardMask_4; // @[MemBlock.scala 232:23]
  wire  sbuffer_io_forward_0_forwardMask_5; // @[MemBlock.scala 232:23]
  wire  sbuffer_io_forward_0_forwardMask_6; // @[MemBlock.scala 232:23]
  wire  sbuffer_io_forward_0_forwardMask_7; // @[MemBlock.scala 232:23]
  wire  sbuffer_io_forward_0_forwardMask_8; // @[MemBlock.scala 232:23]
  wire  sbuffer_io_forward_0_forwardMask_9; // @[MemBlock.scala 232:23]
  wire  sbuffer_io_forward_0_forwardMask_10; // @[MemBlock.scala 232:23]
  wire  sbuffer_io_forward_0_forwardMask_11; // @[MemBlock.scala 232:23]
  wire  sbuffer_io_forward_0_forwardMask_12; // @[MemBlock.scala 232:23]
  wire  sbuffer_io_forward_0_forwardMask_13; // @[MemBlock.scala 232:23]
  wire  sbuffer_io_forward_0_forwardMask_14; // @[MemBlock.scala 232:23]
  wire  sbuffer_io_forward_0_forwardMask_15; // @[MemBlock.scala 232:23]
  wire [7:0] sbuffer_io_forward_0_forwardData_0; // @[MemBlock.scala 232:23]
  wire [7:0] sbuffer_io_forward_0_forwardData_1; // @[MemBlock.scala 232:23]
  wire [7:0] sbuffer_io_forward_0_forwardData_2; // @[MemBlock.scala 232:23]
  wire [7:0] sbuffer_io_forward_0_forwardData_3; // @[MemBlock.scala 232:23]
  wire [7:0] sbuffer_io_forward_0_forwardData_4; // @[MemBlock.scala 232:23]
  wire [7:0] sbuffer_io_forward_0_forwardData_5; // @[MemBlock.scala 232:23]
  wire [7:0] sbuffer_io_forward_0_forwardData_6; // @[MemBlock.scala 232:23]
  wire [7:0] sbuffer_io_forward_0_forwardData_7; // @[MemBlock.scala 232:23]
  wire [7:0] sbuffer_io_forward_0_forwardData_8; // @[MemBlock.scala 232:23]
  wire [7:0] sbuffer_io_forward_0_forwardData_9; // @[MemBlock.scala 232:23]
  wire [7:0] sbuffer_io_forward_0_forwardData_10; // @[MemBlock.scala 232:23]
  wire [7:0] sbuffer_io_forward_0_forwardData_11; // @[MemBlock.scala 232:23]
  wire [7:0] sbuffer_io_forward_0_forwardData_12; // @[MemBlock.scala 232:23]
  wire [7:0] sbuffer_io_forward_0_forwardData_13; // @[MemBlock.scala 232:23]
  wire [7:0] sbuffer_io_forward_0_forwardData_14; // @[MemBlock.scala 232:23]
  wire [7:0] sbuffer_io_forward_0_forwardData_15; // @[MemBlock.scala 232:23]
  wire  sbuffer_io_forward_0_matchInvalid; // @[MemBlock.scala 232:23]
  wire [38:0] sbuffer_io_forward_1_vaddr; // @[MemBlock.scala 232:23]
  wire [35:0] sbuffer_io_forward_1_paddr; // @[MemBlock.scala 232:23]
  wire  sbuffer_io_forward_1_valid; // @[MemBlock.scala 232:23]
  wire  sbuffer_io_forward_1_forwardMask_0; // @[MemBlock.scala 232:23]
  wire  sbuffer_io_forward_1_forwardMask_1; // @[MemBlock.scala 232:23]
  wire  sbuffer_io_forward_1_forwardMask_2; // @[MemBlock.scala 232:23]
  wire  sbuffer_io_forward_1_forwardMask_3; // @[MemBlock.scala 232:23]
  wire  sbuffer_io_forward_1_forwardMask_4; // @[MemBlock.scala 232:23]
  wire  sbuffer_io_forward_1_forwardMask_5; // @[MemBlock.scala 232:23]
  wire  sbuffer_io_forward_1_forwardMask_6; // @[MemBlock.scala 232:23]
  wire  sbuffer_io_forward_1_forwardMask_7; // @[MemBlock.scala 232:23]
  wire  sbuffer_io_forward_1_forwardMask_8; // @[MemBlock.scala 232:23]
  wire  sbuffer_io_forward_1_forwardMask_9; // @[MemBlock.scala 232:23]
  wire  sbuffer_io_forward_1_forwardMask_10; // @[MemBlock.scala 232:23]
  wire  sbuffer_io_forward_1_forwardMask_11; // @[MemBlock.scala 232:23]
  wire  sbuffer_io_forward_1_forwardMask_12; // @[MemBlock.scala 232:23]
  wire  sbuffer_io_forward_1_forwardMask_13; // @[MemBlock.scala 232:23]
  wire  sbuffer_io_forward_1_forwardMask_14; // @[MemBlock.scala 232:23]
  wire  sbuffer_io_forward_1_forwardMask_15; // @[MemBlock.scala 232:23]
  wire [7:0] sbuffer_io_forward_1_forwardData_0; // @[MemBlock.scala 232:23]
  wire [7:0] sbuffer_io_forward_1_forwardData_1; // @[MemBlock.scala 232:23]
  wire [7:0] sbuffer_io_forward_1_forwardData_2; // @[MemBlock.scala 232:23]
  wire [7:0] sbuffer_io_forward_1_forwardData_3; // @[MemBlock.scala 232:23]
  wire [7:0] sbuffer_io_forward_1_forwardData_4; // @[MemBlock.scala 232:23]
  wire [7:0] sbuffer_io_forward_1_forwardData_5; // @[MemBlock.scala 232:23]
  wire [7:0] sbuffer_io_forward_1_forwardData_6; // @[MemBlock.scala 232:23]
  wire [7:0] sbuffer_io_forward_1_forwardData_7; // @[MemBlock.scala 232:23]
  wire [7:0] sbuffer_io_forward_1_forwardData_8; // @[MemBlock.scala 232:23]
  wire [7:0] sbuffer_io_forward_1_forwardData_9; // @[MemBlock.scala 232:23]
  wire [7:0] sbuffer_io_forward_1_forwardData_10; // @[MemBlock.scala 232:23]
  wire [7:0] sbuffer_io_forward_1_forwardData_11; // @[MemBlock.scala 232:23]
  wire [7:0] sbuffer_io_forward_1_forwardData_12; // @[MemBlock.scala 232:23]
  wire [7:0] sbuffer_io_forward_1_forwardData_13; // @[MemBlock.scala 232:23]
  wire [7:0] sbuffer_io_forward_1_forwardData_14; // @[MemBlock.scala 232:23]
  wire [7:0] sbuffer_io_forward_1_forwardData_15; // @[MemBlock.scala 232:23]
  wire  sbuffer_io_forward_1_matchInvalid; // @[MemBlock.scala 232:23]
  wire  sbuffer_io_sqempty; // @[MemBlock.scala 232:23]
  wire  sbuffer_io_flush_valid; // @[MemBlock.scala 232:23]
  wire  sbuffer_io_flush_empty; // @[MemBlock.scala 232:23]
  wire [3:0] sbuffer_io_csrCtrl_sbuffer_threshold; // @[MemBlock.scala 232:23]
  wire [5:0] sbuffer_io_perf_0_value; // @[MemBlock.scala 232:23]
  wire [5:0] sbuffer_io_perf_1_value; // @[MemBlock.scala 232:23]
  wire [5:0] sbuffer_io_perf_2_value; // @[MemBlock.scala 232:23]
  wire [5:0] sbuffer_io_perf_3_value; // @[MemBlock.scala 232:23]
  wire [5:0] sbuffer_io_perf_4_value; // @[MemBlock.scala 232:23]
  wire [5:0] sbuffer_io_perf_5_value; // @[MemBlock.scala 232:23]
  wire [5:0] sbuffer_io_perf_6_value; // @[MemBlock.scala 232:23]
  wire [5:0] sbuffer_io_perf_7_value; // @[MemBlock.scala 232:23]
  wire [5:0] sbuffer_io_perf_8_value; // @[MemBlock.scala 232:23]
  wire [5:0] sbuffer_io_perf_9_value; // @[MemBlock.scala 232:23]
  wire [5:0] sbuffer_io_perf_10_value; // @[MemBlock.scala 232:23]
  wire [5:0] sbuffer_io_perf_11_value; // @[MemBlock.scala 232:23]
  wire [5:0] sbuffer_io_perf_12_value; // @[MemBlock.scala 232:23]
  wire [5:0] sbuffer_io_perf_13_value; // @[MemBlock.scala 232:23]
  wire [5:0] sbuffer_io_perf_14_value; // @[MemBlock.scala 232:23]
  wire [5:0] sbuffer_io_perf_15_value; // @[MemBlock.scala 232:23]
  wire [5:0] sbuffer_io_perf_16_value; // @[MemBlock.scala 232:23]
  wire  dtlb_ld_tlb_ld_clock; // @[MemBlock.scala 246:24]
  wire  dtlb_ld_tlb_ld_reset; // @[MemBlock.scala 246:24]
  wire  dtlb_ld_tlb_ld_io_sfence_valid; // @[MemBlock.scala 246:24]
  wire  dtlb_ld_tlb_ld_io_sfence_bits_rs1; // @[MemBlock.scala 246:24]
  wire  dtlb_ld_tlb_ld_io_sfence_bits_rs2; // @[MemBlock.scala 246:24]
  wire [38:0] dtlb_ld_tlb_ld_io_sfence_bits_addr; // @[MemBlock.scala 246:24]
  wire [15:0] dtlb_ld_tlb_ld_io_sfence_bits_asid; // @[MemBlock.scala 246:24]
  wire [3:0] dtlb_ld_tlb_ld_io_csr_satp_mode; // @[MemBlock.scala 246:24]
  wire [15:0] dtlb_ld_tlb_ld_io_csr_satp_asid; // @[MemBlock.scala 246:24]
  wire  dtlb_ld_tlb_ld_io_csr_satp_changed; // @[MemBlock.scala 246:24]
  wire  dtlb_ld_tlb_ld_io_csr_priv_mxr; // @[MemBlock.scala 246:24]
  wire  dtlb_ld_tlb_ld_io_csr_priv_sum; // @[MemBlock.scala 246:24]
  wire [1:0] dtlb_ld_tlb_ld_io_csr_priv_dmode; // @[MemBlock.scala 246:24]
  wire  dtlb_ld_tlb_ld_io_requestor_0_req_ready; // @[MemBlock.scala 246:24]
  wire  dtlb_ld_tlb_ld_io_requestor_0_req_valid; // @[MemBlock.scala 246:24]
  wire [38:0] dtlb_ld_tlb_ld_io_requestor_0_req_bits_vaddr; // @[MemBlock.scala 246:24]
  wire [2:0] dtlb_ld_tlb_ld_io_requestor_0_req_bits_cmd; // @[MemBlock.scala 246:24]
  wire  dtlb_ld_tlb_ld_io_requestor_0_req_bits_no_translate; // @[MemBlock.scala 246:24]
  wire  dtlb_ld_tlb_ld_io_requestor_0_req_kill; // @[MemBlock.scala 246:24]
  wire  dtlb_ld_tlb_ld_io_requestor_0_resp_valid; // @[MemBlock.scala 246:24]
  wire [35:0] dtlb_ld_tlb_ld_io_requestor_0_resp_bits_paddr_0; // @[MemBlock.scala 246:24]
  wire [35:0] dtlb_ld_tlb_ld_io_requestor_0_resp_bits_paddr_1; // @[MemBlock.scala 246:24]
  wire  dtlb_ld_tlb_ld_io_requestor_0_resp_bits_miss; // @[MemBlock.scala 246:24]
  wire  dtlb_ld_tlb_ld_io_requestor_0_resp_bits_excp_0_pf_ld; // @[MemBlock.scala 246:24]
  wire  dtlb_ld_tlb_ld_io_requestor_0_resp_bits_excp_0_pf_st; // @[MemBlock.scala 246:24]
  wire  dtlb_ld_tlb_ld_io_requestor_0_resp_bits_excp_0_af_ld; // @[MemBlock.scala 246:24]
  wire  dtlb_ld_tlb_ld_io_requestor_0_resp_bits_excp_0_af_st; // @[MemBlock.scala 246:24]
  wire  dtlb_ld_tlb_ld_io_requestor_0_resp_bits_static_pm_valid; // @[MemBlock.scala 246:24]
  wire  dtlb_ld_tlb_ld_io_requestor_0_resp_bits_static_pm_bits; // @[MemBlock.scala 246:24]
  wire  dtlb_ld_tlb_ld_io_requestor_1_req_ready; // @[MemBlock.scala 246:24]
  wire  dtlb_ld_tlb_ld_io_requestor_1_req_valid; // @[MemBlock.scala 246:24]
  wire [38:0] dtlb_ld_tlb_ld_io_requestor_1_req_bits_vaddr; // @[MemBlock.scala 246:24]
  wire [2:0] dtlb_ld_tlb_ld_io_requestor_1_req_bits_cmd; // @[MemBlock.scala 246:24]
  wire  dtlb_ld_tlb_ld_io_requestor_1_req_bits_no_translate; // @[MemBlock.scala 246:24]
  wire  dtlb_ld_tlb_ld_io_requestor_1_req_kill; // @[MemBlock.scala 246:24]
  wire  dtlb_ld_tlb_ld_io_requestor_1_resp_valid; // @[MemBlock.scala 246:24]
  wire [35:0] dtlb_ld_tlb_ld_io_requestor_1_resp_bits_paddr_0; // @[MemBlock.scala 246:24]
  wire [35:0] dtlb_ld_tlb_ld_io_requestor_1_resp_bits_paddr_1; // @[MemBlock.scala 246:24]
  wire  dtlb_ld_tlb_ld_io_requestor_1_resp_bits_miss; // @[MemBlock.scala 246:24]
  wire  dtlb_ld_tlb_ld_io_requestor_1_resp_bits_excp_0_pf_ld; // @[MemBlock.scala 246:24]
  wire  dtlb_ld_tlb_ld_io_requestor_1_resp_bits_excp_0_af_ld; // @[MemBlock.scala 246:24]
  wire  dtlb_ld_tlb_ld_io_requestor_1_resp_bits_static_pm_valid; // @[MemBlock.scala 246:24]
  wire  dtlb_ld_tlb_ld_io_requestor_1_resp_bits_static_pm_bits; // @[MemBlock.scala 246:24]
  wire  dtlb_ld_tlb_ld_io_ptw_req_0_valid; // @[MemBlock.scala 246:24]
  wire [26:0] dtlb_ld_tlb_ld_io_ptw_req_0_bits_vpn; // @[MemBlock.scala 246:24]
  wire  dtlb_ld_tlb_ld_io_ptw_req_1_valid; // @[MemBlock.scala 246:24]
  wire [26:0] dtlb_ld_tlb_ld_io_ptw_req_1_bits_vpn; // @[MemBlock.scala 246:24]
  wire  dtlb_ld_tlb_ld_io_ptw_resp_ready; // @[MemBlock.scala 246:24]
  wire  dtlb_ld_tlb_ld_io_ptw_resp_valid; // @[MemBlock.scala 246:24]
  wire [26:0] dtlb_ld_tlb_ld_io_ptw_resp_bits_entry_tag; // @[MemBlock.scala 246:24]
  wire [15:0] dtlb_ld_tlb_ld_io_ptw_resp_bits_entry_asid; // @[MemBlock.scala 246:24]
  wire [23:0] dtlb_ld_tlb_ld_io_ptw_resp_bits_entry_ppn; // @[MemBlock.scala 246:24]
  wire  dtlb_ld_tlb_ld_io_ptw_resp_bits_entry_perm_d; // @[MemBlock.scala 246:24]
  wire  dtlb_ld_tlb_ld_io_ptw_resp_bits_entry_perm_a; // @[MemBlock.scala 246:24]
  wire  dtlb_ld_tlb_ld_io_ptw_resp_bits_entry_perm_g; // @[MemBlock.scala 246:24]
  wire  dtlb_ld_tlb_ld_io_ptw_resp_bits_entry_perm_u; // @[MemBlock.scala 246:24]
  wire  dtlb_ld_tlb_ld_io_ptw_resp_bits_entry_perm_x; // @[MemBlock.scala 246:24]
  wire  dtlb_ld_tlb_ld_io_ptw_resp_bits_entry_perm_w; // @[MemBlock.scala 246:24]
  wire  dtlb_ld_tlb_ld_io_ptw_resp_bits_entry_perm_r; // @[MemBlock.scala 246:24]
  wire [1:0] dtlb_ld_tlb_ld_io_ptw_resp_bits_entry_level; // @[MemBlock.scala 246:24]
  wire  dtlb_ld_tlb_ld_io_ptw_resp_bits_pf; // @[MemBlock.scala 246:24]
  wire  dtlb_ld_tlb_ld_io_ptw_resp_bits_af; // @[MemBlock.scala 246:24]
  wire  dtlb_ld_tlb_ld_io_ptw_replenish_c; // @[MemBlock.scala 246:24]
  wire  dtlb_ld_tlb_ld_io_ptw_replenish_atomic; // @[MemBlock.scala 246:24]
  wire  dtlb_ld_tlb_ld_io_ptw_replenish_x; // @[MemBlock.scala 246:24]
  wire  dtlb_ld_tlb_ld_io_ptw_replenish_w; // @[MemBlock.scala 246:24]
  wire  dtlb_ld_tlb_ld_io_ptw_replenish_r; // @[MemBlock.scala 246:24]
  wire  dtlb_ld_tlb_ld_io_pmp_0_valid; // @[MemBlock.scala 246:24]
  wire [35:0] dtlb_ld_tlb_ld_io_pmp_0_bits_addr; // @[MemBlock.scala 246:24]
  wire [2:0] dtlb_ld_tlb_ld_io_pmp_0_bits_cmd; // @[MemBlock.scala 246:24]
  wire  dtlb_ld_tlb_ld_io_pmp_1_valid; // @[MemBlock.scala 246:24]
  wire [35:0] dtlb_ld_tlb_ld_io_pmp_1_bits_addr; // @[MemBlock.scala 246:24]
  wire [2:0] dtlb_ld_tlb_ld_io_pmp_1_bits_cmd; // @[MemBlock.scala 246:24]
  wire  dtlb_st_tlb_st_clock; // @[MemBlock.scala 250:24]
  wire  dtlb_st_tlb_st_reset; // @[MemBlock.scala 250:24]
  wire  dtlb_st_tlb_st_io_sfence_valid; // @[MemBlock.scala 250:24]
  wire  dtlb_st_tlb_st_io_sfence_bits_rs1; // @[MemBlock.scala 250:24]
  wire  dtlb_st_tlb_st_io_sfence_bits_rs2; // @[MemBlock.scala 250:24]
  wire [38:0] dtlb_st_tlb_st_io_sfence_bits_addr; // @[MemBlock.scala 250:24]
  wire [15:0] dtlb_st_tlb_st_io_sfence_bits_asid; // @[MemBlock.scala 250:24]
  wire [3:0] dtlb_st_tlb_st_io_csr_satp_mode; // @[MemBlock.scala 250:24]
  wire [15:0] dtlb_st_tlb_st_io_csr_satp_asid; // @[MemBlock.scala 250:24]
  wire  dtlb_st_tlb_st_io_csr_satp_changed; // @[MemBlock.scala 250:24]
  wire  dtlb_st_tlb_st_io_csr_priv_sum; // @[MemBlock.scala 250:24]
  wire [1:0] dtlb_st_tlb_st_io_csr_priv_dmode; // @[MemBlock.scala 250:24]
  wire  dtlb_st_tlb_st_io_requestor_0_req_ready; // @[MemBlock.scala 250:24]
  wire  dtlb_st_tlb_st_io_requestor_0_req_valid; // @[MemBlock.scala 250:24]
  wire [38:0] dtlb_st_tlb_st_io_requestor_0_req_bits_vaddr; // @[MemBlock.scala 250:24]
  wire  dtlb_st_tlb_st_io_requestor_0_resp_valid; // @[MemBlock.scala 250:24]
  wire [35:0] dtlb_st_tlb_st_io_requestor_0_resp_bits_paddr_0; // @[MemBlock.scala 250:24]
  wire  dtlb_st_tlb_st_io_requestor_0_resp_bits_miss; // @[MemBlock.scala 250:24]
  wire  dtlb_st_tlb_st_io_requestor_0_resp_bits_excp_0_pf_st; // @[MemBlock.scala 250:24]
  wire  dtlb_st_tlb_st_io_requestor_0_resp_bits_excp_0_af_st; // @[MemBlock.scala 250:24]
  wire  dtlb_st_tlb_st_io_requestor_0_resp_bits_static_pm_valid; // @[MemBlock.scala 250:24]
  wire  dtlb_st_tlb_st_io_requestor_0_resp_bits_static_pm_bits; // @[MemBlock.scala 250:24]
  wire  dtlb_st_tlb_st_io_requestor_1_req_ready; // @[MemBlock.scala 250:24]
  wire  dtlb_st_tlb_st_io_requestor_1_req_valid; // @[MemBlock.scala 250:24]
  wire [38:0] dtlb_st_tlb_st_io_requestor_1_req_bits_vaddr; // @[MemBlock.scala 250:24]
  wire  dtlb_st_tlb_st_io_requestor_1_resp_valid; // @[MemBlock.scala 250:24]
  wire [35:0] dtlb_st_tlb_st_io_requestor_1_resp_bits_paddr_0; // @[MemBlock.scala 250:24]
  wire  dtlb_st_tlb_st_io_requestor_1_resp_bits_miss; // @[MemBlock.scala 250:24]
  wire  dtlb_st_tlb_st_io_requestor_1_resp_bits_excp_0_pf_st; // @[MemBlock.scala 250:24]
  wire  dtlb_st_tlb_st_io_requestor_1_resp_bits_excp_0_af_st; // @[MemBlock.scala 250:24]
  wire  dtlb_st_tlb_st_io_requestor_1_resp_bits_static_pm_valid; // @[MemBlock.scala 250:24]
  wire  dtlb_st_tlb_st_io_requestor_1_resp_bits_static_pm_bits; // @[MemBlock.scala 250:24]
  wire  dtlb_st_tlb_st_io_ptw_req_0_valid; // @[MemBlock.scala 250:24]
  wire [26:0] dtlb_st_tlb_st_io_ptw_req_0_bits_vpn; // @[MemBlock.scala 250:24]
  wire  dtlb_st_tlb_st_io_ptw_req_1_valid; // @[MemBlock.scala 250:24]
  wire [26:0] dtlb_st_tlb_st_io_ptw_req_1_bits_vpn; // @[MemBlock.scala 250:24]
  wire  dtlb_st_tlb_st_io_ptw_resp_ready; // @[MemBlock.scala 250:24]
  wire  dtlb_st_tlb_st_io_ptw_resp_valid; // @[MemBlock.scala 250:24]
  wire [26:0] dtlb_st_tlb_st_io_ptw_resp_bits_entry_tag; // @[MemBlock.scala 250:24]
  wire [15:0] dtlb_st_tlb_st_io_ptw_resp_bits_entry_asid; // @[MemBlock.scala 250:24]
  wire [23:0] dtlb_st_tlb_st_io_ptw_resp_bits_entry_ppn; // @[MemBlock.scala 250:24]
  wire  dtlb_st_tlb_st_io_ptw_resp_bits_entry_perm_d; // @[MemBlock.scala 250:24]
  wire  dtlb_st_tlb_st_io_ptw_resp_bits_entry_perm_a; // @[MemBlock.scala 250:24]
  wire  dtlb_st_tlb_st_io_ptw_resp_bits_entry_perm_g; // @[MemBlock.scala 250:24]
  wire  dtlb_st_tlb_st_io_ptw_resp_bits_entry_perm_u; // @[MemBlock.scala 250:24]
  wire  dtlb_st_tlb_st_io_ptw_resp_bits_entry_perm_x; // @[MemBlock.scala 250:24]
  wire  dtlb_st_tlb_st_io_ptw_resp_bits_entry_perm_w; // @[MemBlock.scala 250:24]
  wire  dtlb_st_tlb_st_io_ptw_resp_bits_entry_perm_r; // @[MemBlock.scala 250:24]
  wire [1:0] dtlb_st_tlb_st_io_ptw_resp_bits_entry_level; // @[MemBlock.scala 250:24]
  wire  dtlb_st_tlb_st_io_ptw_resp_bits_pf; // @[MemBlock.scala 250:24]
  wire  dtlb_st_tlb_st_io_ptw_resp_bits_af; // @[MemBlock.scala 250:24]
  wire  dtlb_st_tlb_st_io_ptw_replenish_c; // @[MemBlock.scala 250:24]
  wire  dtlb_st_tlb_st_io_ptw_replenish_atomic; // @[MemBlock.scala 250:24]
  wire  dtlb_st_tlb_st_io_ptw_replenish_x; // @[MemBlock.scala 250:24]
  wire  dtlb_st_tlb_st_io_ptw_replenish_w; // @[MemBlock.scala 250:24]
  wire  dtlb_st_tlb_st_io_ptw_replenish_r; // @[MemBlock.scala 250:24]
  wire  dtlb_st_tlb_st_io_pmp_0_valid; // @[MemBlock.scala 250:24]
  wire [35:0] dtlb_st_tlb_st_io_pmp_0_bits_addr; // @[MemBlock.scala 250:24]
  wire  dtlb_st_tlb_st_io_pmp_1_valid; // @[MemBlock.scala 250:24]
  wire [35:0] dtlb_st_tlb_st_io_pmp_1_bits_addr; // @[MemBlock.scala 250:24]
  wire  dtlb_prefetch_tlb_prefetch_clock; // @[MemBlock.scala 254:30]
  wire  dtlb_prefetch_tlb_prefetch_io_sfence_valid; // @[MemBlock.scala 254:30]
  wire  dtlb_prefetch_tlb_prefetch_io_sfence_bits_rs1; // @[MemBlock.scala 254:30]
  wire  dtlb_prefetch_tlb_prefetch_io_sfence_bits_rs2; // @[MemBlock.scala 254:30]
  wire [38:0] dtlb_prefetch_tlb_prefetch_io_sfence_bits_addr; // @[MemBlock.scala 254:30]
  wire [15:0] dtlb_prefetch_tlb_prefetch_io_sfence_bits_asid; // @[MemBlock.scala 254:30]
  wire [3:0] dtlb_prefetch_tlb_prefetch_io_csr_satp_mode; // @[MemBlock.scala 254:30]
  wire [15:0] dtlb_prefetch_tlb_prefetch_io_csr_satp_asid; // @[MemBlock.scala 254:30]
  wire  dtlb_prefetch_tlb_prefetch_io_csr_satp_changed; // @[MemBlock.scala 254:30]
  wire [1:0] dtlb_prefetch_tlb_prefetch_io_csr_priv_dmode; // @[MemBlock.scala 254:30]
  wire  dtlb_prefetch_tlb_prefetch_io_requestor_0_resp_valid; // @[MemBlock.scala 254:30]
  wire  dtlb_prefetch_tlb_prefetch_io_ptw_resp_ready; // @[MemBlock.scala 254:30]
  wire  dtlb_prefetch_tlb_prefetch_io_ptw_resp_valid; // @[MemBlock.scala 254:30]
  wire [26:0] dtlb_prefetch_tlb_prefetch_io_ptw_resp_bits_entry_tag; // @[MemBlock.scala 254:30]
  wire [15:0] dtlb_prefetch_tlb_prefetch_io_ptw_resp_bits_entry_asid; // @[MemBlock.scala 254:30]
  wire [23:0] dtlb_prefetch_tlb_prefetch_io_ptw_resp_bits_entry_ppn; // @[MemBlock.scala 254:30]
  wire [1:0] dtlb_prefetch_tlb_prefetch_io_ptw_resp_bits_entry_level; // @[MemBlock.scala 254:30]
  wire  dtlb_prefetch_tlb_prefetch_io_pmp_0_valid; // @[MemBlock.scala 254:30]
  wire [35:0] dtlb_prefetch_tlb_prefetch_io_pmp_0_bits_addr; // @[MemBlock.scala 254:30]
  wire  pmp_clock; // @[MemBlock.scala 311:19]
  wire  pmp_reset; // @[MemBlock.scala 311:19]
  wire  pmp_io_distribute_csr_wvalid; // @[MemBlock.scala 311:19]
  wire [11:0] pmp_io_distribute_csr_waddr; // @[MemBlock.scala 311:19]
  wire [63:0] pmp_io_distribute_csr_wdata; // @[MemBlock.scala 311:19]
  wire  pmp_io_pmp_0_cfg_l; // @[MemBlock.scala 311:19]
  wire [1:0] pmp_io_pmp_0_cfg_a; // @[MemBlock.scala 311:19]
  wire  pmp_io_pmp_0_cfg_x; // @[MemBlock.scala 311:19]
  wire  pmp_io_pmp_0_cfg_w; // @[MemBlock.scala 311:19]
  wire  pmp_io_pmp_0_cfg_r; // @[MemBlock.scala 311:19]
  wire [33:0] pmp_io_pmp_0_addr; // @[MemBlock.scala 311:19]
  wire [35:0] pmp_io_pmp_0_mask; // @[MemBlock.scala 311:19]
  wire  pmp_io_pmp_1_cfg_l; // @[MemBlock.scala 311:19]
  wire [1:0] pmp_io_pmp_1_cfg_a; // @[MemBlock.scala 311:19]
  wire  pmp_io_pmp_1_cfg_x; // @[MemBlock.scala 311:19]
  wire  pmp_io_pmp_1_cfg_w; // @[MemBlock.scala 311:19]
  wire  pmp_io_pmp_1_cfg_r; // @[MemBlock.scala 311:19]
  wire [33:0] pmp_io_pmp_1_addr; // @[MemBlock.scala 311:19]
  wire [35:0] pmp_io_pmp_1_mask; // @[MemBlock.scala 311:19]
  wire  pmp_io_pmp_2_cfg_l; // @[MemBlock.scala 311:19]
  wire [1:0] pmp_io_pmp_2_cfg_a; // @[MemBlock.scala 311:19]
  wire  pmp_io_pmp_2_cfg_x; // @[MemBlock.scala 311:19]
  wire  pmp_io_pmp_2_cfg_w; // @[MemBlock.scala 311:19]
  wire  pmp_io_pmp_2_cfg_r; // @[MemBlock.scala 311:19]
  wire [33:0] pmp_io_pmp_2_addr; // @[MemBlock.scala 311:19]
  wire [35:0] pmp_io_pmp_2_mask; // @[MemBlock.scala 311:19]
  wire  pmp_io_pmp_3_cfg_l; // @[MemBlock.scala 311:19]
  wire [1:0] pmp_io_pmp_3_cfg_a; // @[MemBlock.scala 311:19]
  wire  pmp_io_pmp_3_cfg_x; // @[MemBlock.scala 311:19]
  wire  pmp_io_pmp_3_cfg_w; // @[MemBlock.scala 311:19]
  wire  pmp_io_pmp_3_cfg_r; // @[MemBlock.scala 311:19]
  wire [33:0] pmp_io_pmp_3_addr; // @[MemBlock.scala 311:19]
  wire [35:0] pmp_io_pmp_3_mask; // @[MemBlock.scala 311:19]
  wire  pmp_io_pmp_4_cfg_l; // @[MemBlock.scala 311:19]
  wire [1:0] pmp_io_pmp_4_cfg_a; // @[MemBlock.scala 311:19]
  wire  pmp_io_pmp_4_cfg_x; // @[MemBlock.scala 311:19]
  wire  pmp_io_pmp_4_cfg_w; // @[MemBlock.scala 311:19]
  wire  pmp_io_pmp_4_cfg_r; // @[MemBlock.scala 311:19]
  wire [33:0] pmp_io_pmp_4_addr; // @[MemBlock.scala 311:19]
  wire [35:0] pmp_io_pmp_4_mask; // @[MemBlock.scala 311:19]
  wire  pmp_io_pmp_5_cfg_l; // @[MemBlock.scala 311:19]
  wire [1:0] pmp_io_pmp_5_cfg_a; // @[MemBlock.scala 311:19]
  wire  pmp_io_pmp_5_cfg_x; // @[MemBlock.scala 311:19]
  wire  pmp_io_pmp_5_cfg_w; // @[MemBlock.scala 311:19]
  wire  pmp_io_pmp_5_cfg_r; // @[MemBlock.scala 311:19]
  wire [33:0] pmp_io_pmp_5_addr; // @[MemBlock.scala 311:19]
  wire [35:0] pmp_io_pmp_5_mask; // @[MemBlock.scala 311:19]
  wire  pmp_io_pmp_6_cfg_l; // @[MemBlock.scala 311:19]
  wire [1:0] pmp_io_pmp_6_cfg_a; // @[MemBlock.scala 311:19]
  wire  pmp_io_pmp_6_cfg_x; // @[MemBlock.scala 311:19]
  wire  pmp_io_pmp_6_cfg_w; // @[MemBlock.scala 311:19]
  wire  pmp_io_pmp_6_cfg_r; // @[MemBlock.scala 311:19]
  wire [33:0] pmp_io_pmp_6_addr; // @[MemBlock.scala 311:19]
  wire [35:0] pmp_io_pmp_6_mask; // @[MemBlock.scala 311:19]
  wire  pmp_io_pmp_7_cfg_l; // @[MemBlock.scala 311:19]
  wire [1:0] pmp_io_pmp_7_cfg_a; // @[MemBlock.scala 311:19]
  wire  pmp_io_pmp_7_cfg_x; // @[MemBlock.scala 311:19]
  wire  pmp_io_pmp_7_cfg_w; // @[MemBlock.scala 311:19]
  wire  pmp_io_pmp_7_cfg_r; // @[MemBlock.scala 311:19]
  wire [33:0] pmp_io_pmp_7_addr; // @[MemBlock.scala 311:19]
  wire [35:0] pmp_io_pmp_7_mask; // @[MemBlock.scala 311:19]
  wire  pmp_io_pmp_8_cfg_l; // @[MemBlock.scala 311:19]
  wire [1:0] pmp_io_pmp_8_cfg_a; // @[MemBlock.scala 311:19]
  wire  pmp_io_pmp_8_cfg_x; // @[MemBlock.scala 311:19]
  wire  pmp_io_pmp_8_cfg_w; // @[MemBlock.scala 311:19]
  wire  pmp_io_pmp_8_cfg_r; // @[MemBlock.scala 311:19]
  wire [33:0] pmp_io_pmp_8_addr; // @[MemBlock.scala 311:19]
  wire [35:0] pmp_io_pmp_8_mask; // @[MemBlock.scala 311:19]
  wire  pmp_io_pmp_9_cfg_l; // @[MemBlock.scala 311:19]
  wire [1:0] pmp_io_pmp_9_cfg_a; // @[MemBlock.scala 311:19]
  wire  pmp_io_pmp_9_cfg_x; // @[MemBlock.scala 311:19]
  wire  pmp_io_pmp_9_cfg_w; // @[MemBlock.scala 311:19]
  wire  pmp_io_pmp_9_cfg_r; // @[MemBlock.scala 311:19]
  wire [33:0] pmp_io_pmp_9_addr; // @[MemBlock.scala 311:19]
  wire [35:0] pmp_io_pmp_9_mask; // @[MemBlock.scala 311:19]
  wire  pmp_io_pmp_10_cfg_l; // @[MemBlock.scala 311:19]
  wire [1:0] pmp_io_pmp_10_cfg_a; // @[MemBlock.scala 311:19]
  wire  pmp_io_pmp_10_cfg_x; // @[MemBlock.scala 311:19]
  wire  pmp_io_pmp_10_cfg_w; // @[MemBlock.scala 311:19]
  wire  pmp_io_pmp_10_cfg_r; // @[MemBlock.scala 311:19]
  wire [33:0] pmp_io_pmp_10_addr; // @[MemBlock.scala 311:19]
  wire [35:0] pmp_io_pmp_10_mask; // @[MemBlock.scala 311:19]
  wire  pmp_io_pmp_11_cfg_l; // @[MemBlock.scala 311:19]
  wire [1:0] pmp_io_pmp_11_cfg_a; // @[MemBlock.scala 311:19]
  wire  pmp_io_pmp_11_cfg_x; // @[MemBlock.scala 311:19]
  wire  pmp_io_pmp_11_cfg_w; // @[MemBlock.scala 311:19]
  wire  pmp_io_pmp_11_cfg_r; // @[MemBlock.scala 311:19]
  wire [33:0] pmp_io_pmp_11_addr; // @[MemBlock.scala 311:19]
  wire [35:0] pmp_io_pmp_11_mask; // @[MemBlock.scala 311:19]
  wire  pmp_io_pmp_12_cfg_l; // @[MemBlock.scala 311:19]
  wire [1:0] pmp_io_pmp_12_cfg_a; // @[MemBlock.scala 311:19]
  wire  pmp_io_pmp_12_cfg_x; // @[MemBlock.scala 311:19]
  wire  pmp_io_pmp_12_cfg_w; // @[MemBlock.scala 311:19]
  wire  pmp_io_pmp_12_cfg_r; // @[MemBlock.scala 311:19]
  wire [33:0] pmp_io_pmp_12_addr; // @[MemBlock.scala 311:19]
  wire [35:0] pmp_io_pmp_12_mask; // @[MemBlock.scala 311:19]
  wire  pmp_io_pmp_13_cfg_l; // @[MemBlock.scala 311:19]
  wire [1:0] pmp_io_pmp_13_cfg_a; // @[MemBlock.scala 311:19]
  wire  pmp_io_pmp_13_cfg_x; // @[MemBlock.scala 311:19]
  wire  pmp_io_pmp_13_cfg_w; // @[MemBlock.scala 311:19]
  wire  pmp_io_pmp_13_cfg_r; // @[MemBlock.scala 311:19]
  wire [33:0] pmp_io_pmp_13_addr; // @[MemBlock.scala 311:19]
  wire [35:0] pmp_io_pmp_13_mask; // @[MemBlock.scala 311:19]
  wire  pmp_io_pmp_14_cfg_l; // @[MemBlock.scala 311:19]
  wire [1:0] pmp_io_pmp_14_cfg_a; // @[MemBlock.scala 311:19]
  wire  pmp_io_pmp_14_cfg_x; // @[MemBlock.scala 311:19]
  wire  pmp_io_pmp_14_cfg_w; // @[MemBlock.scala 311:19]
  wire  pmp_io_pmp_14_cfg_r; // @[MemBlock.scala 311:19]
  wire [33:0] pmp_io_pmp_14_addr; // @[MemBlock.scala 311:19]
  wire [35:0] pmp_io_pmp_14_mask; // @[MemBlock.scala 311:19]
  wire  pmp_io_pmp_15_cfg_l; // @[MemBlock.scala 311:19]
  wire [1:0] pmp_io_pmp_15_cfg_a; // @[MemBlock.scala 311:19]
  wire  pmp_io_pmp_15_cfg_x; // @[MemBlock.scala 311:19]
  wire  pmp_io_pmp_15_cfg_w; // @[MemBlock.scala 311:19]
  wire  pmp_io_pmp_15_cfg_r; // @[MemBlock.scala 311:19]
  wire [33:0] pmp_io_pmp_15_addr; // @[MemBlock.scala 311:19]
  wire [35:0] pmp_io_pmp_15_mask; // @[MemBlock.scala 311:19]
  wire  pmp_io_pma_0_cfg_c; // @[MemBlock.scala 311:19]
  wire  pmp_io_pma_0_cfg_atomic; // @[MemBlock.scala 311:19]
  wire [1:0] pmp_io_pma_0_cfg_a; // @[MemBlock.scala 311:19]
  wire  pmp_io_pma_0_cfg_x; // @[MemBlock.scala 311:19]
  wire  pmp_io_pma_0_cfg_w; // @[MemBlock.scala 311:19]
  wire  pmp_io_pma_0_cfg_r; // @[MemBlock.scala 311:19]
  wire [33:0] pmp_io_pma_0_addr; // @[MemBlock.scala 311:19]
  wire [35:0] pmp_io_pma_0_mask; // @[MemBlock.scala 311:19]
  wire  pmp_io_pma_1_cfg_c; // @[MemBlock.scala 311:19]
  wire  pmp_io_pma_1_cfg_atomic; // @[MemBlock.scala 311:19]
  wire [1:0] pmp_io_pma_1_cfg_a; // @[MemBlock.scala 311:19]
  wire  pmp_io_pma_1_cfg_x; // @[MemBlock.scala 311:19]
  wire  pmp_io_pma_1_cfg_w; // @[MemBlock.scala 311:19]
  wire  pmp_io_pma_1_cfg_r; // @[MemBlock.scala 311:19]
  wire [33:0] pmp_io_pma_1_addr; // @[MemBlock.scala 311:19]
  wire [35:0] pmp_io_pma_1_mask; // @[MemBlock.scala 311:19]
  wire  pmp_io_pma_2_cfg_c; // @[MemBlock.scala 311:19]
  wire  pmp_io_pma_2_cfg_atomic; // @[MemBlock.scala 311:19]
  wire [1:0] pmp_io_pma_2_cfg_a; // @[MemBlock.scala 311:19]
  wire  pmp_io_pma_2_cfg_x; // @[MemBlock.scala 311:19]
  wire  pmp_io_pma_2_cfg_w; // @[MemBlock.scala 311:19]
  wire  pmp_io_pma_2_cfg_r; // @[MemBlock.scala 311:19]
  wire [33:0] pmp_io_pma_2_addr; // @[MemBlock.scala 311:19]
  wire [35:0] pmp_io_pma_2_mask; // @[MemBlock.scala 311:19]
  wire  pmp_io_pma_3_cfg_c; // @[MemBlock.scala 311:19]
  wire  pmp_io_pma_3_cfg_atomic; // @[MemBlock.scala 311:19]
  wire [1:0] pmp_io_pma_3_cfg_a; // @[MemBlock.scala 311:19]
  wire  pmp_io_pma_3_cfg_x; // @[MemBlock.scala 311:19]
  wire  pmp_io_pma_3_cfg_w; // @[MemBlock.scala 311:19]
  wire  pmp_io_pma_3_cfg_r; // @[MemBlock.scala 311:19]
  wire [33:0] pmp_io_pma_3_addr; // @[MemBlock.scala 311:19]
  wire [35:0] pmp_io_pma_3_mask; // @[MemBlock.scala 311:19]
  wire  pmp_io_pma_4_cfg_c; // @[MemBlock.scala 311:19]
  wire  pmp_io_pma_4_cfg_atomic; // @[MemBlock.scala 311:19]
  wire [1:0] pmp_io_pma_4_cfg_a; // @[MemBlock.scala 311:19]
  wire  pmp_io_pma_4_cfg_x; // @[MemBlock.scala 311:19]
  wire  pmp_io_pma_4_cfg_w; // @[MemBlock.scala 311:19]
  wire  pmp_io_pma_4_cfg_r; // @[MemBlock.scala 311:19]
  wire [33:0] pmp_io_pma_4_addr; // @[MemBlock.scala 311:19]
  wire [35:0] pmp_io_pma_4_mask; // @[MemBlock.scala 311:19]
  wire  pmp_io_pma_5_cfg_c; // @[MemBlock.scala 311:19]
  wire  pmp_io_pma_5_cfg_atomic; // @[MemBlock.scala 311:19]
  wire [1:0] pmp_io_pma_5_cfg_a; // @[MemBlock.scala 311:19]
  wire  pmp_io_pma_5_cfg_x; // @[MemBlock.scala 311:19]
  wire  pmp_io_pma_5_cfg_w; // @[MemBlock.scala 311:19]
  wire  pmp_io_pma_5_cfg_r; // @[MemBlock.scala 311:19]
  wire [33:0] pmp_io_pma_5_addr; // @[MemBlock.scala 311:19]
  wire [35:0] pmp_io_pma_5_mask; // @[MemBlock.scala 311:19]
  wire  pmp_io_pma_6_cfg_c; // @[MemBlock.scala 311:19]
  wire  pmp_io_pma_6_cfg_atomic; // @[MemBlock.scala 311:19]
  wire [1:0] pmp_io_pma_6_cfg_a; // @[MemBlock.scala 311:19]
  wire  pmp_io_pma_6_cfg_x; // @[MemBlock.scala 311:19]
  wire  pmp_io_pma_6_cfg_w; // @[MemBlock.scala 311:19]
  wire  pmp_io_pma_6_cfg_r; // @[MemBlock.scala 311:19]
  wire [33:0] pmp_io_pma_6_addr; // @[MemBlock.scala 311:19]
  wire [35:0] pmp_io_pma_6_mask; // @[MemBlock.scala 311:19]
  wire  pmp_io_pma_7_cfg_c; // @[MemBlock.scala 311:19]
  wire  pmp_io_pma_7_cfg_atomic; // @[MemBlock.scala 311:19]
  wire [1:0] pmp_io_pma_7_cfg_a; // @[MemBlock.scala 311:19]
  wire  pmp_io_pma_7_cfg_x; // @[MemBlock.scala 311:19]
  wire  pmp_io_pma_7_cfg_w; // @[MemBlock.scala 311:19]
  wire  pmp_io_pma_7_cfg_r; // @[MemBlock.scala 311:19]
  wire [33:0] pmp_io_pma_7_addr; // @[MemBlock.scala 311:19]
  wire [35:0] pmp_io_pma_7_mask; // @[MemBlock.scala 311:19]
  wire  pmp_io_pma_8_cfg_c; // @[MemBlock.scala 311:19]
  wire  pmp_io_pma_8_cfg_atomic; // @[MemBlock.scala 311:19]
  wire [1:0] pmp_io_pma_8_cfg_a; // @[MemBlock.scala 311:19]
  wire  pmp_io_pma_8_cfg_x; // @[MemBlock.scala 311:19]
  wire  pmp_io_pma_8_cfg_w; // @[MemBlock.scala 311:19]
  wire  pmp_io_pma_8_cfg_r; // @[MemBlock.scala 311:19]
  wire [33:0] pmp_io_pma_8_addr; // @[MemBlock.scala 311:19]
  wire [35:0] pmp_io_pma_8_mask; // @[MemBlock.scala 311:19]
  wire  pmp_io_pma_9_cfg_c; // @[MemBlock.scala 311:19]
  wire  pmp_io_pma_9_cfg_atomic; // @[MemBlock.scala 311:19]
  wire [1:0] pmp_io_pma_9_cfg_a; // @[MemBlock.scala 311:19]
  wire  pmp_io_pma_9_cfg_x; // @[MemBlock.scala 311:19]
  wire  pmp_io_pma_9_cfg_w; // @[MemBlock.scala 311:19]
  wire  pmp_io_pma_9_cfg_r; // @[MemBlock.scala 311:19]
  wire [33:0] pmp_io_pma_9_addr; // @[MemBlock.scala 311:19]
  wire [35:0] pmp_io_pma_9_mask; // @[MemBlock.scala 311:19]
  wire  pmp_io_pma_10_cfg_c; // @[MemBlock.scala 311:19]
  wire  pmp_io_pma_10_cfg_atomic; // @[MemBlock.scala 311:19]
  wire [1:0] pmp_io_pma_10_cfg_a; // @[MemBlock.scala 311:19]
  wire  pmp_io_pma_10_cfg_x; // @[MemBlock.scala 311:19]
  wire  pmp_io_pma_10_cfg_w; // @[MemBlock.scala 311:19]
  wire  pmp_io_pma_10_cfg_r; // @[MemBlock.scala 311:19]
  wire [33:0] pmp_io_pma_10_addr; // @[MemBlock.scala 311:19]
  wire [35:0] pmp_io_pma_10_mask; // @[MemBlock.scala 311:19]
  wire  pmp_io_pma_11_cfg_c; // @[MemBlock.scala 311:19]
  wire  pmp_io_pma_11_cfg_atomic; // @[MemBlock.scala 311:19]
  wire [1:0] pmp_io_pma_11_cfg_a; // @[MemBlock.scala 311:19]
  wire  pmp_io_pma_11_cfg_x; // @[MemBlock.scala 311:19]
  wire  pmp_io_pma_11_cfg_w; // @[MemBlock.scala 311:19]
  wire  pmp_io_pma_11_cfg_r; // @[MemBlock.scala 311:19]
  wire [33:0] pmp_io_pma_11_addr; // @[MemBlock.scala 311:19]
  wire [35:0] pmp_io_pma_11_mask; // @[MemBlock.scala 311:19]
  wire  pmp_io_pma_12_cfg_c; // @[MemBlock.scala 311:19]
  wire  pmp_io_pma_12_cfg_atomic; // @[MemBlock.scala 311:19]
  wire [1:0] pmp_io_pma_12_cfg_a; // @[MemBlock.scala 311:19]
  wire  pmp_io_pma_12_cfg_x; // @[MemBlock.scala 311:19]
  wire  pmp_io_pma_12_cfg_w; // @[MemBlock.scala 311:19]
  wire  pmp_io_pma_12_cfg_r; // @[MemBlock.scala 311:19]
  wire [33:0] pmp_io_pma_12_addr; // @[MemBlock.scala 311:19]
  wire [35:0] pmp_io_pma_12_mask; // @[MemBlock.scala 311:19]
  wire  pmp_io_pma_13_cfg_c; // @[MemBlock.scala 311:19]
  wire  pmp_io_pma_13_cfg_atomic; // @[MemBlock.scala 311:19]
  wire [1:0] pmp_io_pma_13_cfg_a; // @[MemBlock.scala 311:19]
  wire  pmp_io_pma_13_cfg_x; // @[MemBlock.scala 311:19]
  wire  pmp_io_pma_13_cfg_w; // @[MemBlock.scala 311:19]
  wire  pmp_io_pma_13_cfg_r; // @[MemBlock.scala 311:19]
  wire [33:0] pmp_io_pma_13_addr; // @[MemBlock.scala 311:19]
  wire [35:0] pmp_io_pma_13_mask; // @[MemBlock.scala 311:19]
  wire  pmp_io_pma_14_cfg_c; // @[MemBlock.scala 311:19]
  wire  pmp_io_pma_14_cfg_atomic; // @[MemBlock.scala 311:19]
  wire [1:0] pmp_io_pma_14_cfg_a; // @[MemBlock.scala 311:19]
  wire  pmp_io_pma_14_cfg_x; // @[MemBlock.scala 311:19]
  wire  pmp_io_pma_14_cfg_w; // @[MemBlock.scala 311:19]
  wire  pmp_io_pma_14_cfg_r; // @[MemBlock.scala 311:19]
  wire [33:0] pmp_io_pma_14_addr; // @[MemBlock.scala 311:19]
  wire [35:0] pmp_io_pma_14_mask; // @[MemBlock.scala 311:19]
  wire  pmp_io_pma_15_cfg_c; // @[MemBlock.scala 311:19]
  wire  pmp_io_pma_15_cfg_atomic; // @[MemBlock.scala 311:19]
  wire [1:0] pmp_io_pma_15_cfg_a; // @[MemBlock.scala 311:19]
  wire  pmp_io_pma_15_cfg_x; // @[MemBlock.scala 311:19]
  wire  pmp_io_pma_15_cfg_w; // @[MemBlock.scala 311:19]
  wire  pmp_io_pma_15_cfg_r; // @[MemBlock.scala 311:19]
  wire [33:0] pmp_io_pma_15_addr; // @[MemBlock.scala 311:19]
  wire [35:0] pmp_io_pma_15_mask; // @[MemBlock.scala 311:19]
  wire  PMPChecker_clock; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_io_check_env_mode; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pmp_0_cfg_l; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_io_check_env_pmp_0_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pmp_0_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pmp_0_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_io_check_env_pmp_0_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_io_check_env_pmp_0_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pmp_1_cfg_l; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_io_check_env_pmp_1_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pmp_1_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pmp_1_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_io_check_env_pmp_1_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_io_check_env_pmp_1_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pmp_2_cfg_l; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_io_check_env_pmp_2_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pmp_2_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pmp_2_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_io_check_env_pmp_2_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_io_check_env_pmp_2_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pmp_3_cfg_l; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_io_check_env_pmp_3_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pmp_3_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pmp_3_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_io_check_env_pmp_3_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_io_check_env_pmp_3_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pmp_4_cfg_l; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_io_check_env_pmp_4_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pmp_4_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pmp_4_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_io_check_env_pmp_4_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_io_check_env_pmp_4_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pmp_5_cfg_l; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_io_check_env_pmp_5_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pmp_5_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pmp_5_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_io_check_env_pmp_5_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_io_check_env_pmp_5_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pmp_6_cfg_l; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_io_check_env_pmp_6_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pmp_6_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pmp_6_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_io_check_env_pmp_6_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_io_check_env_pmp_6_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pmp_7_cfg_l; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_io_check_env_pmp_7_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pmp_7_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pmp_7_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_io_check_env_pmp_7_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_io_check_env_pmp_7_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pmp_8_cfg_l; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_io_check_env_pmp_8_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pmp_8_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pmp_8_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_io_check_env_pmp_8_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_io_check_env_pmp_8_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pmp_9_cfg_l; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_io_check_env_pmp_9_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pmp_9_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pmp_9_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_io_check_env_pmp_9_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_io_check_env_pmp_9_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pmp_10_cfg_l; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_io_check_env_pmp_10_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pmp_10_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pmp_10_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_io_check_env_pmp_10_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_io_check_env_pmp_10_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pmp_11_cfg_l; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_io_check_env_pmp_11_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pmp_11_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pmp_11_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_io_check_env_pmp_11_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_io_check_env_pmp_11_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pmp_12_cfg_l; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_io_check_env_pmp_12_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pmp_12_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pmp_12_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_io_check_env_pmp_12_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_io_check_env_pmp_12_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pmp_13_cfg_l; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_io_check_env_pmp_13_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pmp_13_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pmp_13_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_io_check_env_pmp_13_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_io_check_env_pmp_13_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pmp_14_cfg_l; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_io_check_env_pmp_14_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pmp_14_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pmp_14_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_io_check_env_pmp_14_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_io_check_env_pmp_14_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pmp_15_cfg_l; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_io_check_env_pmp_15_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pmp_15_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pmp_15_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_io_check_env_pmp_15_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_io_check_env_pmp_15_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pma_0_cfg_c; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pma_0_cfg_atomic; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_io_check_env_pma_0_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pma_0_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pma_0_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_io_check_env_pma_0_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_io_check_env_pma_0_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pma_1_cfg_c; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pma_1_cfg_atomic; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_io_check_env_pma_1_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pma_1_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pma_1_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_io_check_env_pma_1_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_io_check_env_pma_1_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pma_2_cfg_c; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pma_2_cfg_atomic; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_io_check_env_pma_2_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pma_2_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pma_2_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_io_check_env_pma_2_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_io_check_env_pma_2_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pma_3_cfg_c; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pma_3_cfg_atomic; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_io_check_env_pma_3_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pma_3_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pma_3_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_io_check_env_pma_3_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_io_check_env_pma_3_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pma_4_cfg_c; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pma_4_cfg_atomic; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_io_check_env_pma_4_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pma_4_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pma_4_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_io_check_env_pma_4_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_io_check_env_pma_4_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pma_5_cfg_c; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pma_5_cfg_atomic; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_io_check_env_pma_5_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pma_5_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pma_5_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_io_check_env_pma_5_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_io_check_env_pma_5_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pma_6_cfg_c; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pma_6_cfg_atomic; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_io_check_env_pma_6_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pma_6_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pma_6_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_io_check_env_pma_6_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_io_check_env_pma_6_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pma_7_cfg_c; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pma_7_cfg_atomic; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_io_check_env_pma_7_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pma_7_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pma_7_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_io_check_env_pma_7_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_io_check_env_pma_7_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pma_8_cfg_c; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pma_8_cfg_atomic; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_io_check_env_pma_8_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pma_8_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pma_8_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_io_check_env_pma_8_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_io_check_env_pma_8_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pma_9_cfg_c; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pma_9_cfg_atomic; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_io_check_env_pma_9_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pma_9_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pma_9_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_io_check_env_pma_9_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_io_check_env_pma_9_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pma_10_cfg_c; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pma_10_cfg_atomic; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_io_check_env_pma_10_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pma_10_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pma_10_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_io_check_env_pma_10_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_io_check_env_pma_10_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pma_11_cfg_c; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pma_11_cfg_atomic; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_io_check_env_pma_11_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pma_11_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pma_11_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_io_check_env_pma_11_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_io_check_env_pma_11_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pma_12_cfg_c; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pma_12_cfg_atomic; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_io_check_env_pma_12_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pma_12_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pma_12_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_io_check_env_pma_12_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_io_check_env_pma_12_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pma_13_cfg_c; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pma_13_cfg_atomic; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_io_check_env_pma_13_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pma_13_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pma_13_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_io_check_env_pma_13_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_io_check_env_pma_13_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pma_14_cfg_c; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pma_14_cfg_atomic; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_io_check_env_pma_14_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pma_14_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pma_14_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_io_check_env_pma_14_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_io_check_env_pma_14_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pma_15_cfg_c; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pma_15_cfg_atomic; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_io_check_env_pma_15_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pma_15_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_check_env_pma_15_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_io_check_env_pma_15_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_io_check_env_pma_15_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_req_valid; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_io_req_bits_addr; // @[MemBlock.scala 314:91]
  wire [2:0] PMPChecker_io_req_bits_cmd; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_resp_ld; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_resp_st; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_resp_mmio; // @[MemBlock.scala 314:91]
  wire  PMPChecker_io_resp_atomic; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_clock; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_1_io_check_env_mode; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pmp_0_cfg_l; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_1_io_check_env_pmp_0_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pmp_0_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pmp_0_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_1_io_check_env_pmp_0_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_1_io_check_env_pmp_0_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pmp_1_cfg_l; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_1_io_check_env_pmp_1_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pmp_1_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pmp_1_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_1_io_check_env_pmp_1_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_1_io_check_env_pmp_1_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pmp_2_cfg_l; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_1_io_check_env_pmp_2_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pmp_2_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pmp_2_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_1_io_check_env_pmp_2_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_1_io_check_env_pmp_2_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pmp_3_cfg_l; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_1_io_check_env_pmp_3_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pmp_3_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pmp_3_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_1_io_check_env_pmp_3_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_1_io_check_env_pmp_3_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pmp_4_cfg_l; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_1_io_check_env_pmp_4_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pmp_4_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pmp_4_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_1_io_check_env_pmp_4_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_1_io_check_env_pmp_4_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pmp_5_cfg_l; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_1_io_check_env_pmp_5_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pmp_5_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pmp_5_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_1_io_check_env_pmp_5_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_1_io_check_env_pmp_5_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pmp_6_cfg_l; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_1_io_check_env_pmp_6_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pmp_6_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pmp_6_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_1_io_check_env_pmp_6_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_1_io_check_env_pmp_6_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pmp_7_cfg_l; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_1_io_check_env_pmp_7_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pmp_7_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pmp_7_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_1_io_check_env_pmp_7_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_1_io_check_env_pmp_7_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pmp_8_cfg_l; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_1_io_check_env_pmp_8_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pmp_8_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pmp_8_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_1_io_check_env_pmp_8_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_1_io_check_env_pmp_8_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pmp_9_cfg_l; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_1_io_check_env_pmp_9_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pmp_9_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pmp_9_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_1_io_check_env_pmp_9_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_1_io_check_env_pmp_9_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pmp_10_cfg_l; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_1_io_check_env_pmp_10_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pmp_10_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pmp_10_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_1_io_check_env_pmp_10_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_1_io_check_env_pmp_10_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pmp_11_cfg_l; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_1_io_check_env_pmp_11_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pmp_11_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pmp_11_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_1_io_check_env_pmp_11_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_1_io_check_env_pmp_11_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pmp_12_cfg_l; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_1_io_check_env_pmp_12_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pmp_12_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pmp_12_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_1_io_check_env_pmp_12_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_1_io_check_env_pmp_12_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pmp_13_cfg_l; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_1_io_check_env_pmp_13_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pmp_13_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pmp_13_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_1_io_check_env_pmp_13_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_1_io_check_env_pmp_13_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pmp_14_cfg_l; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_1_io_check_env_pmp_14_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pmp_14_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pmp_14_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_1_io_check_env_pmp_14_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_1_io_check_env_pmp_14_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pmp_15_cfg_l; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_1_io_check_env_pmp_15_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pmp_15_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pmp_15_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_1_io_check_env_pmp_15_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_1_io_check_env_pmp_15_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pma_0_cfg_c; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pma_0_cfg_atomic; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_1_io_check_env_pma_0_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pma_0_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pma_0_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_1_io_check_env_pma_0_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_1_io_check_env_pma_0_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pma_1_cfg_c; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pma_1_cfg_atomic; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_1_io_check_env_pma_1_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pma_1_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pma_1_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_1_io_check_env_pma_1_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_1_io_check_env_pma_1_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pma_2_cfg_c; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pma_2_cfg_atomic; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_1_io_check_env_pma_2_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pma_2_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pma_2_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_1_io_check_env_pma_2_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_1_io_check_env_pma_2_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pma_3_cfg_c; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pma_3_cfg_atomic; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_1_io_check_env_pma_3_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pma_3_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pma_3_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_1_io_check_env_pma_3_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_1_io_check_env_pma_3_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pma_4_cfg_c; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pma_4_cfg_atomic; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_1_io_check_env_pma_4_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pma_4_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pma_4_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_1_io_check_env_pma_4_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_1_io_check_env_pma_4_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pma_5_cfg_c; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pma_5_cfg_atomic; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_1_io_check_env_pma_5_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pma_5_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pma_5_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_1_io_check_env_pma_5_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_1_io_check_env_pma_5_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pma_6_cfg_c; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pma_6_cfg_atomic; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_1_io_check_env_pma_6_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pma_6_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pma_6_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_1_io_check_env_pma_6_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_1_io_check_env_pma_6_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pma_7_cfg_c; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pma_7_cfg_atomic; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_1_io_check_env_pma_7_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pma_7_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pma_7_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_1_io_check_env_pma_7_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_1_io_check_env_pma_7_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pma_8_cfg_c; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pma_8_cfg_atomic; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_1_io_check_env_pma_8_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pma_8_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pma_8_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_1_io_check_env_pma_8_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_1_io_check_env_pma_8_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pma_9_cfg_c; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pma_9_cfg_atomic; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_1_io_check_env_pma_9_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pma_9_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pma_9_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_1_io_check_env_pma_9_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_1_io_check_env_pma_9_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pma_10_cfg_c; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pma_10_cfg_atomic; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_1_io_check_env_pma_10_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pma_10_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pma_10_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_1_io_check_env_pma_10_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_1_io_check_env_pma_10_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pma_11_cfg_c; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pma_11_cfg_atomic; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_1_io_check_env_pma_11_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pma_11_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pma_11_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_1_io_check_env_pma_11_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_1_io_check_env_pma_11_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pma_12_cfg_c; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pma_12_cfg_atomic; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_1_io_check_env_pma_12_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pma_12_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pma_12_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_1_io_check_env_pma_12_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_1_io_check_env_pma_12_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pma_13_cfg_c; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pma_13_cfg_atomic; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_1_io_check_env_pma_13_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pma_13_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pma_13_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_1_io_check_env_pma_13_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_1_io_check_env_pma_13_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pma_14_cfg_c; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pma_14_cfg_atomic; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_1_io_check_env_pma_14_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pma_14_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pma_14_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_1_io_check_env_pma_14_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_1_io_check_env_pma_14_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pma_15_cfg_c; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pma_15_cfg_atomic; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_1_io_check_env_pma_15_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pma_15_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_check_env_pma_15_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_1_io_check_env_pma_15_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_1_io_check_env_pma_15_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_req_valid; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_1_io_req_bits_addr; // @[MemBlock.scala 314:91]
  wire [2:0] PMPChecker_1_io_req_bits_cmd; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_resp_ld; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_resp_st; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_resp_mmio; // @[MemBlock.scala 314:91]
  wire  PMPChecker_1_io_resp_atomic; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_clock; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_2_io_check_env_mode; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pmp_0_cfg_l; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_2_io_check_env_pmp_0_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pmp_0_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pmp_0_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_2_io_check_env_pmp_0_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_2_io_check_env_pmp_0_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pmp_1_cfg_l; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_2_io_check_env_pmp_1_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pmp_1_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pmp_1_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_2_io_check_env_pmp_1_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_2_io_check_env_pmp_1_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pmp_2_cfg_l; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_2_io_check_env_pmp_2_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pmp_2_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pmp_2_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_2_io_check_env_pmp_2_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_2_io_check_env_pmp_2_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pmp_3_cfg_l; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_2_io_check_env_pmp_3_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pmp_3_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pmp_3_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_2_io_check_env_pmp_3_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_2_io_check_env_pmp_3_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pmp_4_cfg_l; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_2_io_check_env_pmp_4_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pmp_4_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pmp_4_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_2_io_check_env_pmp_4_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_2_io_check_env_pmp_4_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pmp_5_cfg_l; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_2_io_check_env_pmp_5_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pmp_5_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pmp_5_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_2_io_check_env_pmp_5_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_2_io_check_env_pmp_5_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pmp_6_cfg_l; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_2_io_check_env_pmp_6_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pmp_6_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pmp_6_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_2_io_check_env_pmp_6_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_2_io_check_env_pmp_6_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pmp_7_cfg_l; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_2_io_check_env_pmp_7_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pmp_7_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pmp_7_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_2_io_check_env_pmp_7_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_2_io_check_env_pmp_7_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pmp_8_cfg_l; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_2_io_check_env_pmp_8_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pmp_8_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pmp_8_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_2_io_check_env_pmp_8_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_2_io_check_env_pmp_8_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pmp_9_cfg_l; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_2_io_check_env_pmp_9_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pmp_9_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pmp_9_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_2_io_check_env_pmp_9_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_2_io_check_env_pmp_9_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pmp_10_cfg_l; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_2_io_check_env_pmp_10_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pmp_10_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pmp_10_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_2_io_check_env_pmp_10_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_2_io_check_env_pmp_10_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pmp_11_cfg_l; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_2_io_check_env_pmp_11_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pmp_11_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pmp_11_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_2_io_check_env_pmp_11_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_2_io_check_env_pmp_11_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pmp_12_cfg_l; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_2_io_check_env_pmp_12_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pmp_12_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pmp_12_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_2_io_check_env_pmp_12_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_2_io_check_env_pmp_12_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pmp_13_cfg_l; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_2_io_check_env_pmp_13_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pmp_13_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pmp_13_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_2_io_check_env_pmp_13_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_2_io_check_env_pmp_13_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pmp_14_cfg_l; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_2_io_check_env_pmp_14_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pmp_14_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pmp_14_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_2_io_check_env_pmp_14_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_2_io_check_env_pmp_14_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pmp_15_cfg_l; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_2_io_check_env_pmp_15_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pmp_15_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pmp_15_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_2_io_check_env_pmp_15_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_2_io_check_env_pmp_15_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pma_0_cfg_c; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pma_0_cfg_atomic; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_2_io_check_env_pma_0_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pma_0_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pma_0_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_2_io_check_env_pma_0_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_2_io_check_env_pma_0_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pma_1_cfg_c; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pma_1_cfg_atomic; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_2_io_check_env_pma_1_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pma_1_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pma_1_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_2_io_check_env_pma_1_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_2_io_check_env_pma_1_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pma_2_cfg_c; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pma_2_cfg_atomic; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_2_io_check_env_pma_2_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pma_2_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pma_2_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_2_io_check_env_pma_2_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_2_io_check_env_pma_2_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pma_3_cfg_c; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pma_3_cfg_atomic; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_2_io_check_env_pma_3_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pma_3_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pma_3_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_2_io_check_env_pma_3_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_2_io_check_env_pma_3_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pma_4_cfg_c; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pma_4_cfg_atomic; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_2_io_check_env_pma_4_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pma_4_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pma_4_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_2_io_check_env_pma_4_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_2_io_check_env_pma_4_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pma_5_cfg_c; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pma_5_cfg_atomic; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_2_io_check_env_pma_5_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pma_5_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pma_5_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_2_io_check_env_pma_5_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_2_io_check_env_pma_5_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pma_6_cfg_c; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pma_6_cfg_atomic; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_2_io_check_env_pma_6_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pma_6_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pma_6_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_2_io_check_env_pma_6_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_2_io_check_env_pma_6_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pma_7_cfg_c; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pma_7_cfg_atomic; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_2_io_check_env_pma_7_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pma_7_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pma_7_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_2_io_check_env_pma_7_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_2_io_check_env_pma_7_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pma_8_cfg_c; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pma_8_cfg_atomic; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_2_io_check_env_pma_8_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pma_8_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pma_8_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_2_io_check_env_pma_8_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_2_io_check_env_pma_8_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pma_9_cfg_c; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pma_9_cfg_atomic; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_2_io_check_env_pma_9_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pma_9_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pma_9_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_2_io_check_env_pma_9_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_2_io_check_env_pma_9_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pma_10_cfg_c; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pma_10_cfg_atomic; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_2_io_check_env_pma_10_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pma_10_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pma_10_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_2_io_check_env_pma_10_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_2_io_check_env_pma_10_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pma_11_cfg_c; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pma_11_cfg_atomic; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_2_io_check_env_pma_11_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pma_11_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pma_11_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_2_io_check_env_pma_11_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_2_io_check_env_pma_11_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pma_12_cfg_c; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pma_12_cfg_atomic; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_2_io_check_env_pma_12_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pma_12_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pma_12_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_2_io_check_env_pma_12_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_2_io_check_env_pma_12_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pma_13_cfg_c; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pma_13_cfg_atomic; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_2_io_check_env_pma_13_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pma_13_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pma_13_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_2_io_check_env_pma_13_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_2_io_check_env_pma_13_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pma_14_cfg_c; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pma_14_cfg_atomic; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_2_io_check_env_pma_14_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pma_14_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pma_14_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_2_io_check_env_pma_14_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_2_io_check_env_pma_14_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pma_15_cfg_c; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pma_15_cfg_atomic; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_2_io_check_env_pma_15_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pma_15_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_check_env_pma_15_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_2_io_check_env_pma_15_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_2_io_check_env_pma_15_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_req_valid; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_2_io_req_bits_addr; // @[MemBlock.scala 314:91]
  wire [2:0] PMPChecker_2_io_req_bits_cmd; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_resp_ld; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_resp_st; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_resp_mmio; // @[MemBlock.scala 314:91]
  wire  PMPChecker_2_io_resp_atomic; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_clock; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_3_io_check_env_mode; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pmp_0_cfg_l; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_3_io_check_env_pmp_0_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pmp_0_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pmp_0_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_3_io_check_env_pmp_0_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_3_io_check_env_pmp_0_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pmp_1_cfg_l; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_3_io_check_env_pmp_1_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pmp_1_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pmp_1_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_3_io_check_env_pmp_1_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_3_io_check_env_pmp_1_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pmp_2_cfg_l; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_3_io_check_env_pmp_2_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pmp_2_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pmp_2_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_3_io_check_env_pmp_2_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_3_io_check_env_pmp_2_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pmp_3_cfg_l; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_3_io_check_env_pmp_3_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pmp_3_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pmp_3_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_3_io_check_env_pmp_3_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_3_io_check_env_pmp_3_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pmp_4_cfg_l; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_3_io_check_env_pmp_4_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pmp_4_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pmp_4_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_3_io_check_env_pmp_4_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_3_io_check_env_pmp_4_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pmp_5_cfg_l; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_3_io_check_env_pmp_5_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pmp_5_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pmp_5_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_3_io_check_env_pmp_5_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_3_io_check_env_pmp_5_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pmp_6_cfg_l; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_3_io_check_env_pmp_6_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pmp_6_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pmp_6_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_3_io_check_env_pmp_6_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_3_io_check_env_pmp_6_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pmp_7_cfg_l; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_3_io_check_env_pmp_7_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pmp_7_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pmp_7_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_3_io_check_env_pmp_7_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_3_io_check_env_pmp_7_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pmp_8_cfg_l; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_3_io_check_env_pmp_8_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pmp_8_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pmp_8_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_3_io_check_env_pmp_8_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_3_io_check_env_pmp_8_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pmp_9_cfg_l; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_3_io_check_env_pmp_9_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pmp_9_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pmp_9_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_3_io_check_env_pmp_9_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_3_io_check_env_pmp_9_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pmp_10_cfg_l; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_3_io_check_env_pmp_10_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pmp_10_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pmp_10_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_3_io_check_env_pmp_10_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_3_io_check_env_pmp_10_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pmp_11_cfg_l; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_3_io_check_env_pmp_11_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pmp_11_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pmp_11_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_3_io_check_env_pmp_11_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_3_io_check_env_pmp_11_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pmp_12_cfg_l; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_3_io_check_env_pmp_12_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pmp_12_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pmp_12_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_3_io_check_env_pmp_12_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_3_io_check_env_pmp_12_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pmp_13_cfg_l; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_3_io_check_env_pmp_13_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pmp_13_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pmp_13_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_3_io_check_env_pmp_13_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_3_io_check_env_pmp_13_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pmp_14_cfg_l; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_3_io_check_env_pmp_14_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pmp_14_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pmp_14_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_3_io_check_env_pmp_14_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_3_io_check_env_pmp_14_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pmp_15_cfg_l; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_3_io_check_env_pmp_15_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pmp_15_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pmp_15_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_3_io_check_env_pmp_15_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_3_io_check_env_pmp_15_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pma_0_cfg_c; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pma_0_cfg_atomic; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_3_io_check_env_pma_0_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pma_0_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pma_0_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_3_io_check_env_pma_0_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_3_io_check_env_pma_0_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pma_1_cfg_c; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pma_1_cfg_atomic; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_3_io_check_env_pma_1_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pma_1_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pma_1_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_3_io_check_env_pma_1_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_3_io_check_env_pma_1_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pma_2_cfg_c; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pma_2_cfg_atomic; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_3_io_check_env_pma_2_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pma_2_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pma_2_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_3_io_check_env_pma_2_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_3_io_check_env_pma_2_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pma_3_cfg_c; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pma_3_cfg_atomic; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_3_io_check_env_pma_3_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pma_3_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pma_3_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_3_io_check_env_pma_3_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_3_io_check_env_pma_3_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pma_4_cfg_c; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pma_4_cfg_atomic; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_3_io_check_env_pma_4_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pma_4_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pma_4_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_3_io_check_env_pma_4_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_3_io_check_env_pma_4_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pma_5_cfg_c; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pma_5_cfg_atomic; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_3_io_check_env_pma_5_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pma_5_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pma_5_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_3_io_check_env_pma_5_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_3_io_check_env_pma_5_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pma_6_cfg_c; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pma_6_cfg_atomic; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_3_io_check_env_pma_6_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pma_6_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pma_6_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_3_io_check_env_pma_6_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_3_io_check_env_pma_6_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pma_7_cfg_c; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pma_7_cfg_atomic; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_3_io_check_env_pma_7_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pma_7_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pma_7_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_3_io_check_env_pma_7_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_3_io_check_env_pma_7_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pma_8_cfg_c; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pma_8_cfg_atomic; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_3_io_check_env_pma_8_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pma_8_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pma_8_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_3_io_check_env_pma_8_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_3_io_check_env_pma_8_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pma_9_cfg_c; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pma_9_cfg_atomic; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_3_io_check_env_pma_9_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pma_9_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pma_9_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_3_io_check_env_pma_9_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_3_io_check_env_pma_9_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pma_10_cfg_c; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pma_10_cfg_atomic; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_3_io_check_env_pma_10_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pma_10_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pma_10_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_3_io_check_env_pma_10_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_3_io_check_env_pma_10_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pma_11_cfg_c; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pma_11_cfg_atomic; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_3_io_check_env_pma_11_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pma_11_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pma_11_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_3_io_check_env_pma_11_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_3_io_check_env_pma_11_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pma_12_cfg_c; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pma_12_cfg_atomic; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_3_io_check_env_pma_12_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pma_12_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pma_12_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_3_io_check_env_pma_12_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_3_io_check_env_pma_12_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pma_13_cfg_c; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pma_13_cfg_atomic; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_3_io_check_env_pma_13_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pma_13_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pma_13_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_3_io_check_env_pma_13_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_3_io_check_env_pma_13_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pma_14_cfg_c; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pma_14_cfg_atomic; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_3_io_check_env_pma_14_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pma_14_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pma_14_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_3_io_check_env_pma_14_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_3_io_check_env_pma_14_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pma_15_cfg_c; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pma_15_cfg_atomic; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_3_io_check_env_pma_15_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pma_15_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_check_env_pma_15_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_3_io_check_env_pma_15_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_3_io_check_env_pma_15_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_req_valid; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_3_io_req_bits_addr; // @[MemBlock.scala 314:91]
  wire [2:0] PMPChecker_3_io_req_bits_cmd; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_resp_ld; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_resp_st; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_resp_mmio; // @[MemBlock.scala 314:91]
  wire  PMPChecker_3_io_resp_atomic; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_clock; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_4_io_check_env_mode; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pmp_0_cfg_l; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_4_io_check_env_pmp_0_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pmp_0_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pmp_0_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_4_io_check_env_pmp_0_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_4_io_check_env_pmp_0_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pmp_1_cfg_l; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_4_io_check_env_pmp_1_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pmp_1_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pmp_1_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_4_io_check_env_pmp_1_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_4_io_check_env_pmp_1_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pmp_2_cfg_l; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_4_io_check_env_pmp_2_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pmp_2_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pmp_2_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_4_io_check_env_pmp_2_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_4_io_check_env_pmp_2_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pmp_3_cfg_l; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_4_io_check_env_pmp_3_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pmp_3_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pmp_3_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_4_io_check_env_pmp_3_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_4_io_check_env_pmp_3_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pmp_4_cfg_l; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_4_io_check_env_pmp_4_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pmp_4_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pmp_4_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_4_io_check_env_pmp_4_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_4_io_check_env_pmp_4_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pmp_5_cfg_l; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_4_io_check_env_pmp_5_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pmp_5_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pmp_5_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_4_io_check_env_pmp_5_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_4_io_check_env_pmp_5_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pmp_6_cfg_l; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_4_io_check_env_pmp_6_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pmp_6_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pmp_6_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_4_io_check_env_pmp_6_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_4_io_check_env_pmp_6_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pmp_7_cfg_l; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_4_io_check_env_pmp_7_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pmp_7_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pmp_7_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_4_io_check_env_pmp_7_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_4_io_check_env_pmp_7_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pmp_8_cfg_l; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_4_io_check_env_pmp_8_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pmp_8_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pmp_8_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_4_io_check_env_pmp_8_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_4_io_check_env_pmp_8_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pmp_9_cfg_l; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_4_io_check_env_pmp_9_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pmp_9_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pmp_9_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_4_io_check_env_pmp_9_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_4_io_check_env_pmp_9_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pmp_10_cfg_l; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_4_io_check_env_pmp_10_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pmp_10_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pmp_10_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_4_io_check_env_pmp_10_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_4_io_check_env_pmp_10_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pmp_11_cfg_l; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_4_io_check_env_pmp_11_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pmp_11_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pmp_11_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_4_io_check_env_pmp_11_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_4_io_check_env_pmp_11_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pmp_12_cfg_l; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_4_io_check_env_pmp_12_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pmp_12_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pmp_12_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_4_io_check_env_pmp_12_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_4_io_check_env_pmp_12_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pmp_13_cfg_l; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_4_io_check_env_pmp_13_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pmp_13_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pmp_13_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_4_io_check_env_pmp_13_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_4_io_check_env_pmp_13_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pmp_14_cfg_l; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_4_io_check_env_pmp_14_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pmp_14_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pmp_14_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_4_io_check_env_pmp_14_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_4_io_check_env_pmp_14_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pmp_15_cfg_l; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_4_io_check_env_pmp_15_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pmp_15_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pmp_15_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_4_io_check_env_pmp_15_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_4_io_check_env_pmp_15_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pma_0_cfg_c; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pma_0_cfg_atomic; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_4_io_check_env_pma_0_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pma_0_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pma_0_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_4_io_check_env_pma_0_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_4_io_check_env_pma_0_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pma_1_cfg_c; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pma_1_cfg_atomic; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_4_io_check_env_pma_1_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pma_1_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pma_1_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_4_io_check_env_pma_1_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_4_io_check_env_pma_1_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pma_2_cfg_c; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pma_2_cfg_atomic; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_4_io_check_env_pma_2_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pma_2_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pma_2_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_4_io_check_env_pma_2_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_4_io_check_env_pma_2_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pma_3_cfg_c; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pma_3_cfg_atomic; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_4_io_check_env_pma_3_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pma_3_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pma_3_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_4_io_check_env_pma_3_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_4_io_check_env_pma_3_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pma_4_cfg_c; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pma_4_cfg_atomic; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_4_io_check_env_pma_4_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pma_4_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pma_4_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_4_io_check_env_pma_4_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_4_io_check_env_pma_4_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pma_5_cfg_c; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pma_5_cfg_atomic; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_4_io_check_env_pma_5_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pma_5_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pma_5_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_4_io_check_env_pma_5_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_4_io_check_env_pma_5_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pma_6_cfg_c; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pma_6_cfg_atomic; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_4_io_check_env_pma_6_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pma_6_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pma_6_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_4_io_check_env_pma_6_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_4_io_check_env_pma_6_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pma_7_cfg_c; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pma_7_cfg_atomic; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_4_io_check_env_pma_7_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pma_7_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pma_7_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_4_io_check_env_pma_7_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_4_io_check_env_pma_7_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pma_8_cfg_c; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pma_8_cfg_atomic; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_4_io_check_env_pma_8_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pma_8_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pma_8_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_4_io_check_env_pma_8_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_4_io_check_env_pma_8_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pma_9_cfg_c; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pma_9_cfg_atomic; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_4_io_check_env_pma_9_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pma_9_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pma_9_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_4_io_check_env_pma_9_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_4_io_check_env_pma_9_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pma_10_cfg_c; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pma_10_cfg_atomic; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_4_io_check_env_pma_10_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pma_10_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pma_10_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_4_io_check_env_pma_10_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_4_io_check_env_pma_10_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pma_11_cfg_c; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pma_11_cfg_atomic; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_4_io_check_env_pma_11_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pma_11_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pma_11_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_4_io_check_env_pma_11_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_4_io_check_env_pma_11_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pma_12_cfg_c; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pma_12_cfg_atomic; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_4_io_check_env_pma_12_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pma_12_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pma_12_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_4_io_check_env_pma_12_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_4_io_check_env_pma_12_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pma_13_cfg_c; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pma_13_cfg_atomic; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_4_io_check_env_pma_13_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pma_13_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pma_13_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_4_io_check_env_pma_13_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_4_io_check_env_pma_13_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pma_14_cfg_c; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pma_14_cfg_atomic; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_4_io_check_env_pma_14_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pma_14_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pma_14_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_4_io_check_env_pma_14_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_4_io_check_env_pma_14_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pma_15_cfg_c; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pma_15_cfg_atomic; // @[MemBlock.scala 314:91]
  wire [1:0] PMPChecker_4_io_check_env_pma_15_cfg_a; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pma_15_cfg_w; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_check_env_pma_15_cfg_r; // @[MemBlock.scala 314:91]
  wire [33:0] PMPChecker_4_io_check_env_pma_15_addr; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_4_io_check_env_pma_15_mask; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_req_valid; // @[MemBlock.scala 314:91]
  wire [35:0] PMPChecker_4_io_req_bits_addr; // @[MemBlock.scala 314:91]
  wire [2:0] PMPChecker_4_io_req_bits_cmd; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_resp_ld; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_resp_st; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_resp_mmio; // @[MemBlock.scala 314:91]
  wire  PMPChecker_4_io_resp_atomic; // @[MemBlock.scala 314:91]
  wire  pmp_check_ptw_clock; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_reset; // @[MemBlock.scala 319:29]
  wire [1:0] pmp_check_ptw_io_check_env_mode; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pmp_0_cfg_l; // @[MemBlock.scala 319:29]
  wire [1:0] pmp_check_ptw_io_check_env_pmp_0_cfg_a; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pmp_0_cfg_x; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pmp_0_cfg_w; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pmp_0_cfg_r; // @[MemBlock.scala 319:29]
  wire [33:0] pmp_check_ptw_io_check_env_pmp_0_addr; // @[MemBlock.scala 319:29]
  wire [35:0] pmp_check_ptw_io_check_env_pmp_0_mask; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pmp_1_cfg_l; // @[MemBlock.scala 319:29]
  wire [1:0] pmp_check_ptw_io_check_env_pmp_1_cfg_a; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pmp_1_cfg_x; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pmp_1_cfg_w; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pmp_1_cfg_r; // @[MemBlock.scala 319:29]
  wire [33:0] pmp_check_ptw_io_check_env_pmp_1_addr; // @[MemBlock.scala 319:29]
  wire [35:0] pmp_check_ptw_io_check_env_pmp_1_mask; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pmp_2_cfg_l; // @[MemBlock.scala 319:29]
  wire [1:0] pmp_check_ptw_io_check_env_pmp_2_cfg_a; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pmp_2_cfg_x; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pmp_2_cfg_w; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pmp_2_cfg_r; // @[MemBlock.scala 319:29]
  wire [33:0] pmp_check_ptw_io_check_env_pmp_2_addr; // @[MemBlock.scala 319:29]
  wire [35:0] pmp_check_ptw_io_check_env_pmp_2_mask; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pmp_3_cfg_l; // @[MemBlock.scala 319:29]
  wire [1:0] pmp_check_ptw_io_check_env_pmp_3_cfg_a; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pmp_3_cfg_x; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pmp_3_cfg_w; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pmp_3_cfg_r; // @[MemBlock.scala 319:29]
  wire [33:0] pmp_check_ptw_io_check_env_pmp_3_addr; // @[MemBlock.scala 319:29]
  wire [35:0] pmp_check_ptw_io_check_env_pmp_3_mask; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pmp_4_cfg_l; // @[MemBlock.scala 319:29]
  wire [1:0] pmp_check_ptw_io_check_env_pmp_4_cfg_a; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pmp_4_cfg_x; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pmp_4_cfg_w; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pmp_4_cfg_r; // @[MemBlock.scala 319:29]
  wire [33:0] pmp_check_ptw_io_check_env_pmp_4_addr; // @[MemBlock.scala 319:29]
  wire [35:0] pmp_check_ptw_io_check_env_pmp_4_mask; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pmp_5_cfg_l; // @[MemBlock.scala 319:29]
  wire [1:0] pmp_check_ptw_io_check_env_pmp_5_cfg_a; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pmp_5_cfg_x; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pmp_5_cfg_w; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pmp_5_cfg_r; // @[MemBlock.scala 319:29]
  wire [33:0] pmp_check_ptw_io_check_env_pmp_5_addr; // @[MemBlock.scala 319:29]
  wire [35:0] pmp_check_ptw_io_check_env_pmp_5_mask; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pmp_6_cfg_l; // @[MemBlock.scala 319:29]
  wire [1:0] pmp_check_ptw_io_check_env_pmp_6_cfg_a; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pmp_6_cfg_x; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pmp_6_cfg_w; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pmp_6_cfg_r; // @[MemBlock.scala 319:29]
  wire [33:0] pmp_check_ptw_io_check_env_pmp_6_addr; // @[MemBlock.scala 319:29]
  wire [35:0] pmp_check_ptw_io_check_env_pmp_6_mask; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pmp_7_cfg_l; // @[MemBlock.scala 319:29]
  wire [1:0] pmp_check_ptw_io_check_env_pmp_7_cfg_a; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pmp_7_cfg_x; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pmp_7_cfg_w; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pmp_7_cfg_r; // @[MemBlock.scala 319:29]
  wire [33:0] pmp_check_ptw_io_check_env_pmp_7_addr; // @[MemBlock.scala 319:29]
  wire [35:0] pmp_check_ptw_io_check_env_pmp_7_mask; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pmp_8_cfg_l; // @[MemBlock.scala 319:29]
  wire [1:0] pmp_check_ptw_io_check_env_pmp_8_cfg_a; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pmp_8_cfg_x; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pmp_8_cfg_w; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pmp_8_cfg_r; // @[MemBlock.scala 319:29]
  wire [33:0] pmp_check_ptw_io_check_env_pmp_8_addr; // @[MemBlock.scala 319:29]
  wire [35:0] pmp_check_ptw_io_check_env_pmp_8_mask; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pmp_9_cfg_l; // @[MemBlock.scala 319:29]
  wire [1:0] pmp_check_ptw_io_check_env_pmp_9_cfg_a; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pmp_9_cfg_x; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pmp_9_cfg_w; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pmp_9_cfg_r; // @[MemBlock.scala 319:29]
  wire [33:0] pmp_check_ptw_io_check_env_pmp_9_addr; // @[MemBlock.scala 319:29]
  wire [35:0] pmp_check_ptw_io_check_env_pmp_9_mask; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pmp_10_cfg_l; // @[MemBlock.scala 319:29]
  wire [1:0] pmp_check_ptw_io_check_env_pmp_10_cfg_a; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pmp_10_cfg_x; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pmp_10_cfg_w; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pmp_10_cfg_r; // @[MemBlock.scala 319:29]
  wire [33:0] pmp_check_ptw_io_check_env_pmp_10_addr; // @[MemBlock.scala 319:29]
  wire [35:0] pmp_check_ptw_io_check_env_pmp_10_mask; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pmp_11_cfg_l; // @[MemBlock.scala 319:29]
  wire [1:0] pmp_check_ptw_io_check_env_pmp_11_cfg_a; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pmp_11_cfg_x; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pmp_11_cfg_w; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pmp_11_cfg_r; // @[MemBlock.scala 319:29]
  wire [33:0] pmp_check_ptw_io_check_env_pmp_11_addr; // @[MemBlock.scala 319:29]
  wire [35:0] pmp_check_ptw_io_check_env_pmp_11_mask; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pmp_12_cfg_l; // @[MemBlock.scala 319:29]
  wire [1:0] pmp_check_ptw_io_check_env_pmp_12_cfg_a; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pmp_12_cfg_x; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pmp_12_cfg_w; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pmp_12_cfg_r; // @[MemBlock.scala 319:29]
  wire [33:0] pmp_check_ptw_io_check_env_pmp_12_addr; // @[MemBlock.scala 319:29]
  wire [35:0] pmp_check_ptw_io_check_env_pmp_12_mask; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pmp_13_cfg_l; // @[MemBlock.scala 319:29]
  wire [1:0] pmp_check_ptw_io_check_env_pmp_13_cfg_a; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pmp_13_cfg_x; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pmp_13_cfg_w; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pmp_13_cfg_r; // @[MemBlock.scala 319:29]
  wire [33:0] pmp_check_ptw_io_check_env_pmp_13_addr; // @[MemBlock.scala 319:29]
  wire [35:0] pmp_check_ptw_io_check_env_pmp_13_mask; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pmp_14_cfg_l; // @[MemBlock.scala 319:29]
  wire [1:0] pmp_check_ptw_io_check_env_pmp_14_cfg_a; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pmp_14_cfg_x; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pmp_14_cfg_w; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pmp_14_cfg_r; // @[MemBlock.scala 319:29]
  wire [33:0] pmp_check_ptw_io_check_env_pmp_14_addr; // @[MemBlock.scala 319:29]
  wire [35:0] pmp_check_ptw_io_check_env_pmp_14_mask; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pmp_15_cfg_l; // @[MemBlock.scala 319:29]
  wire [1:0] pmp_check_ptw_io_check_env_pmp_15_cfg_a; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pmp_15_cfg_x; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pmp_15_cfg_w; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pmp_15_cfg_r; // @[MemBlock.scala 319:29]
  wire [33:0] pmp_check_ptw_io_check_env_pmp_15_addr; // @[MemBlock.scala 319:29]
  wire [35:0] pmp_check_ptw_io_check_env_pmp_15_mask; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pma_0_cfg_c; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pma_0_cfg_atomic; // @[MemBlock.scala 319:29]
  wire [1:0] pmp_check_ptw_io_check_env_pma_0_cfg_a; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pma_0_cfg_x; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pma_0_cfg_w; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pma_0_cfg_r; // @[MemBlock.scala 319:29]
  wire [33:0] pmp_check_ptw_io_check_env_pma_0_addr; // @[MemBlock.scala 319:29]
  wire [35:0] pmp_check_ptw_io_check_env_pma_0_mask; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pma_1_cfg_c; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pma_1_cfg_atomic; // @[MemBlock.scala 319:29]
  wire [1:0] pmp_check_ptw_io_check_env_pma_1_cfg_a; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pma_1_cfg_x; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pma_1_cfg_w; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pma_1_cfg_r; // @[MemBlock.scala 319:29]
  wire [33:0] pmp_check_ptw_io_check_env_pma_1_addr; // @[MemBlock.scala 319:29]
  wire [35:0] pmp_check_ptw_io_check_env_pma_1_mask; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pma_2_cfg_c; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pma_2_cfg_atomic; // @[MemBlock.scala 319:29]
  wire [1:0] pmp_check_ptw_io_check_env_pma_2_cfg_a; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pma_2_cfg_x; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pma_2_cfg_w; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pma_2_cfg_r; // @[MemBlock.scala 319:29]
  wire [33:0] pmp_check_ptw_io_check_env_pma_2_addr; // @[MemBlock.scala 319:29]
  wire [35:0] pmp_check_ptw_io_check_env_pma_2_mask; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pma_3_cfg_c; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pma_3_cfg_atomic; // @[MemBlock.scala 319:29]
  wire [1:0] pmp_check_ptw_io_check_env_pma_3_cfg_a; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pma_3_cfg_x; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pma_3_cfg_w; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pma_3_cfg_r; // @[MemBlock.scala 319:29]
  wire [33:0] pmp_check_ptw_io_check_env_pma_3_addr; // @[MemBlock.scala 319:29]
  wire [35:0] pmp_check_ptw_io_check_env_pma_3_mask; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pma_4_cfg_c; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pma_4_cfg_atomic; // @[MemBlock.scala 319:29]
  wire [1:0] pmp_check_ptw_io_check_env_pma_4_cfg_a; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pma_4_cfg_x; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pma_4_cfg_w; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pma_4_cfg_r; // @[MemBlock.scala 319:29]
  wire [33:0] pmp_check_ptw_io_check_env_pma_4_addr; // @[MemBlock.scala 319:29]
  wire [35:0] pmp_check_ptw_io_check_env_pma_4_mask; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pma_5_cfg_c; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pma_5_cfg_atomic; // @[MemBlock.scala 319:29]
  wire [1:0] pmp_check_ptw_io_check_env_pma_5_cfg_a; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pma_5_cfg_x; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pma_5_cfg_w; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pma_5_cfg_r; // @[MemBlock.scala 319:29]
  wire [33:0] pmp_check_ptw_io_check_env_pma_5_addr; // @[MemBlock.scala 319:29]
  wire [35:0] pmp_check_ptw_io_check_env_pma_5_mask; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pma_6_cfg_c; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pma_6_cfg_atomic; // @[MemBlock.scala 319:29]
  wire [1:0] pmp_check_ptw_io_check_env_pma_6_cfg_a; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pma_6_cfg_x; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pma_6_cfg_w; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pma_6_cfg_r; // @[MemBlock.scala 319:29]
  wire [33:0] pmp_check_ptw_io_check_env_pma_6_addr; // @[MemBlock.scala 319:29]
  wire [35:0] pmp_check_ptw_io_check_env_pma_6_mask; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pma_7_cfg_c; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pma_7_cfg_atomic; // @[MemBlock.scala 319:29]
  wire [1:0] pmp_check_ptw_io_check_env_pma_7_cfg_a; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pma_7_cfg_x; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pma_7_cfg_w; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pma_7_cfg_r; // @[MemBlock.scala 319:29]
  wire [33:0] pmp_check_ptw_io_check_env_pma_7_addr; // @[MemBlock.scala 319:29]
  wire [35:0] pmp_check_ptw_io_check_env_pma_7_mask; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pma_8_cfg_c; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pma_8_cfg_atomic; // @[MemBlock.scala 319:29]
  wire [1:0] pmp_check_ptw_io_check_env_pma_8_cfg_a; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pma_8_cfg_x; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pma_8_cfg_w; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pma_8_cfg_r; // @[MemBlock.scala 319:29]
  wire [33:0] pmp_check_ptw_io_check_env_pma_8_addr; // @[MemBlock.scala 319:29]
  wire [35:0] pmp_check_ptw_io_check_env_pma_8_mask; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pma_9_cfg_c; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pma_9_cfg_atomic; // @[MemBlock.scala 319:29]
  wire [1:0] pmp_check_ptw_io_check_env_pma_9_cfg_a; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pma_9_cfg_x; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pma_9_cfg_w; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pma_9_cfg_r; // @[MemBlock.scala 319:29]
  wire [33:0] pmp_check_ptw_io_check_env_pma_9_addr; // @[MemBlock.scala 319:29]
  wire [35:0] pmp_check_ptw_io_check_env_pma_9_mask; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pma_10_cfg_c; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pma_10_cfg_atomic; // @[MemBlock.scala 319:29]
  wire [1:0] pmp_check_ptw_io_check_env_pma_10_cfg_a; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pma_10_cfg_x; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pma_10_cfg_w; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pma_10_cfg_r; // @[MemBlock.scala 319:29]
  wire [33:0] pmp_check_ptw_io_check_env_pma_10_addr; // @[MemBlock.scala 319:29]
  wire [35:0] pmp_check_ptw_io_check_env_pma_10_mask; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pma_11_cfg_c; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pma_11_cfg_atomic; // @[MemBlock.scala 319:29]
  wire [1:0] pmp_check_ptw_io_check_env_pma_11_cfg_a; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pma_11_cfg_x; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pma_11_cfg_w; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pma_11_cfg_r; // @[MemBlock.scala 319:29]
  wire [33:0] pmp_check_ptw_io_check_env_pma_11_addr; // @[MemBlock.scala 319:29]
  wire [35:0] pmp_check_ptw_io_check_env_pma_11_mask; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pma_12_cfg_c; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pma_12_cfg_atomic; // @[MemBlock.scala 319:29]
  wire [1:0] pmp_check_ptw_io_check_env_pma_12_cfg_a; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pma_12_cfg_x; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pma_12_cfg_w; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pma_12_cfg_r; // @[MemBlock.scala 319:29]
  wire [33:0] pmp_check_ptw_io_check_env_pma_12_addr; // @[MemBlock.scala 319:29]
  wire [35:0] pmp_check_ptw_io_check_env_pma_12_mask; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pma_13_cfg_c; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pma_13_cfg_atomic; // @[MemBlock.scala 319:29]
  wire [1:0] pmp_check_ptw_io_check_env_pma_13_cfg_a; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pma_13_cfg_x; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pma_13_cfg_w; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pma_13_cfg_r; // @[MemBlock.scala 319:29]
  wire [33:0] pmp_check_ptw_io_check_env_pma_13_addr; // @[MemBlock.scala 319:29]
  wire [35:0] pmp_check_ptw_io_check_env_pma_13_mask; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pma_14_cfg_c; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pma_14_cfg_atomic; // @[MemBlock.scala 319:29]
  wire [1:0] pmp_check_ptw_io_check_env_pma_14_cfg_a; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pma_14_cfg_x; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pma_14_cfg_w; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pma_14_cfg_r; // @[MemBlock.scala 319:29]
  wire [33:0] pmp_check_ptw_io_check_env_pma_14_addr; // @[MemBlock.scala 319:29]
  wire [35:0] pmp_check_ptw_io_check_env_pma_14_mask; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pma_15_cfg_c; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pma_15_cfg_atomic; // @[MemBlock.scala 319:29]
  wire [1:0] pmp_check_ptw_io_check_env_pma_15_cfg_a; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pma_15_cfg_x; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pma_15_cfg_w; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_check_env_pma_15_cfg_r; // @[MemBlock.scala 319:29]
  wire [33:0] pmp_check_ptw_io_check_env_pma_15_addr; // @[MemBlock.scala 319:29]
  wire [35:0] pmp_check_ptw_io_check_env_pma_15_mask; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_req_valid; // @[MemBlock.scala 319:29]
  wire [35:0] pmp_check_ptw_io_req_bits_addr; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_resp_c; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_resp_atomic; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_resp_x; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_resp_w; // @[MemBlock.scala 319:29]
  wire  pmp_check_ptw_io_resp_r; // @[MemBlock.scala 319:29]
  wire  pipelineReg_clock; // @[MemCommon.scala 396:29]
  wire  pipelineReg_reset; // @[MemCommon.scala 396:29]
  wire  pipelineReg_io_in_ready; // @[MemCommon.scala 396:29]
  wire  pipelineReg_io_in_valid; // @[MemCommon.scala 396:29]
  wire [4:0] pipelineReg_io_in_bits_cmd; // @[MemCommon.scala 396:29]
  wire [35:0] pipelineReg_io_in_bits_addr; // @[MemCommon.scala 396:29]
  wire [63:0] pipelineReg_io_in_bits_data; // @[MemCommon.scala 396:29]
  wire [7:0] pipelineReg_io_in_bits_mask; // @[MemCommon.scala 396:29]
  wire  pipelineReg_io_in_bits_atomic; // @[MemCommon.scala 396:29]
  wire  pipelineReg_io_out_ready; // @[MemCommon.scala 396:29]
  wire  pipelineReg_io_out_valid; // @[MemCommon.scala 396:29]
  wire [4:0] pipelineReg_io_out_bits_cmd; // @[MemCommon.scala 396:29]
  wire [35:0] pipelineReg_io_out_bits_addr; // @[MemCommon.scala 396:29]
  wire [63:0] pipelineReg_io_out_bits_data; // @[MemCommon.scala 396:29]
  wire [7:0] pipelineReg_io_out_bits_mask; // @[MemCommon.scala 396:29]
  wire  pipelineReg_io_out_bits_atomic; // @[MemCommon.scala 396:29]
  wire  pipelineReg_1_clock; // @[MemCommon.scala 396:29]
  wire  pipelineReg_1_reset; // @[MemCommon.scala 396:29]
  wire  pipelineReg_1_io_in_ready; // @[MemCommon.scala 396:29]
  wire  pipelineReg_1_io_in_valid; // @[MemCommon.scala 396:29]
  wire [63:0] pipelineReg_1_io_in_bits_data; // @[MemCommon.scala 396:29]
  wire  pipelineReg_1_io_out_valid; // @[MemCommon.scala 396:29]
  wire [63:0] pipelineReg_1_io_out_bits_data; // @[MemCommon.scala 396:29]
  wire  delay_clock; // @[Hold.scala 97:23]
  wire  delay_io_in; // @[Hold.scala 97:23]
  wire  delay_io_out; // @[Hold.scala 97:23]
  wire  pfevent_clock; // @[MemBlock.scala 687:23]
  wire  pfevent_reset; // @[MemBlock.scala 687:23]
  wire  pfevent_io_distribute_csr_wvalid; // @[MemBlock.scala 687:23]
  wire [11:0] pfevent_io_distribute_csr_waddr; // @[MemBlock.scala 687:23]
  wire [63:0] pfevent_io_distribute_csr_wdata; // @[MemBlock.scala 687:23]
  wire [63:0] pfevent_io_hpmevent_0; // @[MemBlock.scala 687:23]
  wire [63:0] pfevent_io_hpmevent_1; // @[MemBlock.scala 687:23]
  wire [63:0] pfevent_io_hpmevent_2; // @[MemBlock.scala 687:23]
  wire [63:0] pfevent_io_hpmevent_3; // @[MemBlock.scala 687:23]
  wire [63:0] pfevent_io_hpmevent_4; // @[MemBlock.scala 687:23]
  wire [63:0] pfevent_io_hpmevent_5; // @[MemBlock.scala 687:23]
  wire [63:0] pfevent_io_hpmevent_6; // @[MemBlock.scala 687:23]
  wire [63:0] pfevent_io_hpmevent_7; // @[MemBlock.scala 687:23]
  wire [63:0] pfevent_io_hpmevent_8; // @[MemBlock.scala 687:23]
  wire [63:0] pfevent_io_hpmevent_9; // @[MemBlock.scala 687:23]
  wire [63:0] pfevent_io_hpmevent_10; // @[MemBlock.scala 687:23]
  wire [63:0] pfevent_io_hpmevent_11; // @[MemBlock.scala 687:23]
  wire [63:0] pfevent_io_hpmevent_12; // @[MemBlock.scala 687:23]
  wire [63:0] pfevent_io_hpmevent_13; // @[MemBlock.scala 687:23]
  wire [63:0] pfevent_io_hpmevent_14; // @[MemBlock.scala 687:23]
  wire [63:0] pfevent_io_hpmevent_15; // @[MemBlock.scala 687:23]
  wire [63:0] pfevent_io_hpmevent_16; // @[MemBlock.scala 687:23]
  wire [63:0] pfevent_io_hpmevent_17; // @[MemBlock.scala 687:23]
  wire [63:0] pfevent_io_hpmevent_18; // @[MemBlock.scala 687:23]
  wire [63:0] pfevent_io_hpmevent_19; // @[MemBlock.scala 687:23]
  wire [63:0] pfevent_io_hpmevent_20; // @[MemBlock.scala 687:23]
  wire [63:0] pfevent_io_hpmevent_21; // @[MemBlock.scala 687:23]
  wire [63:0] pfevent_io_hpmevent_22; // @[MemBlock.scala 687:23]
  wire [63:0] pfevent_io_hpmevent_23; // @[MemBlock.scala 687:23]
  wire  hpm_clock; // @[PerfCounterUtils.scala 255:21]
  wire [63:0] hpm_io_hpm_event_0; // @[PerfCounterUtils.scala 255:21]
  wire [63:0] hpm_io_hpm_event_1; // @[PerfCounterUtils.scala 255:21]
  wire [63:0] hpm_io_hpm_event_2; // @[PerfCounterUtils.scala 255:21]
  wire [63:0] hpm_io_hpm_event_3; // @[PerfCounterUtils.scala 255:21]
  wire [63:0] hpm_io_hpm_event_4; // @[PerfCounterUtils.scala 255:21]
  wire [63:0] hpm_io_hpm_event_5; // @[PerfCounterUtils.scala 255:21]
  wire [63:0] hpm_io_hpm_event_6; // @[PerfCounterUtils.scala 255:21]
  wire [63:0] hpm_io_hpm_event_7; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_0_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_1_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_2_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_3_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_4_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_5_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_6_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_7_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_8_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_9_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_10_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_11_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_12_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_13_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_14_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_15_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_16_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_17_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_18_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_19_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_20_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_21_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_22_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_23_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_24_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_25_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_26_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_27_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_28_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_29_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_30_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_31_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_32_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_33_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_34_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_35_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_36_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_37_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_38_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_39_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_40_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_41_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_42_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_43_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_44_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_45_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_46_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_47_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_48_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_49_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_50_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_51_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_52_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_53_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_54_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_55_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_56_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_57_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_58_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_59_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_60_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_61_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_62_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_63_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_64_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_65_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_66_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_67_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_68_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_69_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_70_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_71_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_72_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_73_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_74_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_75_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_76_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_77_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_78_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_79_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_80_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_81_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_82_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_83_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_84_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_85_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_86_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_87_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_88_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_89_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_90_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_91_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_92_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_93_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_94_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_95_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_96_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_97_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_98_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_99_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_100_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_101_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_102_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_103_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_104_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_105_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_106_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_107_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_events_sets_108_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_perf_0_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_perf_1_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_perf_2_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_perf_3_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_perf_4_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_perf_5_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_perf_6_value; // @[PerfCounterUtils.scala 255:21]
  wire [5:0] hpm_io_perf_7_value; // @[PerfCounterUtils.scala 255:21]
  reg  redirect_next_valid_REG; // @[BitUtils.scala 28:28]
  reg  redirect_next_bits_rrobIdx_flag; // @[Reg.scala 16:16]
  reg [4:0] redirect_next_bits_rrobIdx_value; // @[Reg.scala 16:16]
  reg  redirect_next_bits_rlevel; // @[Reg.scala 16:16]
  reg  delayedDcacheRefill_valid; // @[MemBlock.scala 127:36]
  reg [1:0] delayedDcacheRefill_bits_id; // @[MemBlock.scala 127:36]
  reg  io_csrUpdate_REG_wvalid; // @[MemBlock.scala 132:26]
  reg [11:0] io_csrUpdate_REG_waddr; // @[MemBlock.scala 132:26]
  reg [63:0] io_csrUpdate_REG_wdata; // @[MemBlock.scala 132:26]
  reg [35:0] io_error_REG_paddr; // @[MemBlock.scala 133:30]
  reg  io_error_REG_report_to_beu; // @[MemBlock.scala 133:30]
  reg [35:0] io_error_REG_1_paddr; // @[MemBlock.scala 133:22]
  reg  io_error_REG_1_report_to_beu; // @[MemBlock.scala 133:22]
  wire  loadWritebackOverride_uop_cf_exceptionVec_4 = atomicsUnit_io_out_valid ?
    atomicsUnit_io_out_bits_uop_cf_exceptionVec_4 : LoadUnit_0_io_loadOut_bits_uop_cf_exceptionVec_4; // @[MemBlock.scala 182:35]
  wire  loadWritebackOverride_uop_cf_exceptionVec_5 = atomicsUnit_io_out_valid ?
    atomicsUnit_io_out_bits_uop_cf_exceptionVec_5 : LoadUnit_0_io_loadOut_bits_uop_cf_exceptionVec_5; // @[MemBlock.scala 182:35]
  wire  loadWritebackOverride_uop_cf_exceptionVec_13 = atomicsUnit_io_out_valid ?
    atomicsUnit_io_out_bits_uop_cf_exceptionVec_13 : LoadUnit_0_io_loadOut_bits_uop_cf_exceptionVec_13; // @[MemBlock.scala 182:35]
  wire  loadWritebackOverride_uop_cf_trigger_backendHit_0 = atomicsUnit_io_out_valid ?
    atomicsUnit_io_out_bits_uop_cf_trigger_backendHit_0 : LoadUnit_0_io_loadOut_bits_uop_cf_trigger_backendHit_0; // @[MemBlock.scala 182:35]
  wire  loadWritebackOverride_uop_cf_trigger_backendHit_1 = atomicsUnit_io_out_valid ?
    atomicsUnit_io_out_bits_uop_cf_trigger_backendHit_1 : LoadUnit_0_io_loadOut_bits_uop_cf_trigger_backendHit_1; // @[MemBlock.scala 182:35]
  wire  loadWritebackOverride_uop_cf_trigger_backendHit_4 = atomicsUnit_io_out_valid ?
    atomicsUnit_io_out_bits_uop_cf_trigger_backendHit_4 : LoadUnit_0_io_loadOut_bits_uop_cf_trigger_backendHit_4; // @[MemBlock.scala 182:35]
  reg  sfence_REG_valid; // @[MemBlock.scala 243:31]
  reg  sfence_REG_bits_rs1; // @[MemBlock.scala 243:31]
  reg  sfence_REG_bits_rs2; // @[MemBlock.scala 243:31]
  reg [38:0] sfence_REG_bits_addr; // @[MemBlock.scala 243:31]
  reg [15:0] sfence_REG_bits_asid; // @[MemBlock.scala 243:31]
  reg  sfence_valid; // @[MemBlock.scala 243:23]
  reg  sfence_bits_rs1; // @[MemBlock.scala 243:23]
  reg  sfence_bits_rs2; // @[MemBlock.scala 243:23]
  reg [38:0] sfence_bits_addr; // @[MemBlock.scala 243:23]
  reg [15:0] sfence_bits_asid; // @[MemBlock.scala 243:23]
  reg [3:0] tlbcsr_REG_satp_mode; // @[MemBlock.scala 244:31]
  reg [15:0] tlbcsr_REG_satp_asid; // @[MemBlock.scala 244:31]
  reg  tlbcsr_REG_satp_changed; // @[MemBlock.scala 244:31]
  reg  tlbcsr_REG_priv_mxr; // @[MemBlock.scala 244:31]
  reg  tlbcsr_REG_priv_sum; // @[MemBlock.scala 244:31]
  reg [1:0] tlbcsr_REG_priv_dmode; // @[MemBlock.scala 244:31]
  reg [3:0] tlbcsr_satp_mode; // @[MemBlock.scala 244:23]
  reg [15:0] tlbcsr_satp_asid; // @[MemBlock.scala 244:23]
  reg  tlbcsr_satp_changed; // @[MemBlock.scala 244:23]
  reg  tlbcsr_priv_mxr; // @[MemBlock.scala 244:23]
  reg  tlbcsr_priv_sum; // @[MemBlock.scala 244:23]
  reg [1:0] tlbcsr_priv_dmode; // @[MemBlock.scala 244:23]
  reg [26:0] ptw_resp_next_data_entry_tag; // @[Reg.scala 16:16]
  reg [15:0] ptw_resp_next_data_entry_asid; // @[Reg.scala 16:16]
  reg [23:0] ptw_resp_next_data_entry_ppn; // @[Reg.scala 16:16]
  reg  ptw_resp_next_data_entry_perm_d; // @[Reg.scala 16:16]
  reg  ptw_resp_next_data_entry_perm_a; // @[Reg.scala 16:16]
  reg  ptw_resp_next_data_entry_perm_g; // @[Reg.scala 16:16]
  reg  ptw_resp_next_data_entry_perm_u; // @[Reg.scala 16:16]
  reg  ptw_resp_next_data_entry_perm_x; // @[Reg.scala 16:16]
  reg  ptw_resp_next_data_entry_perm_w; // @[Reg.scala 16:16]
  reg  ptw_resp_next_data_entry_perm_r; // @[Reg.scala 16:16]
  reg [1:0] ptw_resp_next_data_entry_level; // @[Reg.scala 16:16]
  reg  ptw_resp_next_data_pf; // @[Reg.scala 16:16]
  reg  ptw_resp_next_data_af; // @[Reg.scala 16:16]
  reg  ptw_resp_next_vector_0; // @[Reg.scala 16:16]
  reg  ptw_resp_next_vector_1; // @[Reg.scala 16:16]
  reg  ptw_resp_next_vector_2; // @[Reg.scala 16:16]
  reg  ptw_resp_next_vector_3; // @[Reg.scala 16:16]
  reg  ptw_resp_next_vector_4; // @[Reg.scala 16:16]
  reg  ptw_resp_v; // @[MemBlock.scala 281:27]
  wire [1:0] _vector_hit_T = {ptw_resp_next_vector_0,ptw_resp_next_vector_1}; // @[Cat.scala 31:58]
  wire  vector_hit = |_vector_hit_T; // @[MemBlock.scala 289:95]
  wire [26:0] dtlb_ld_0_ptw_req_0_bits_vpn = dtlb_ld_tlb_ld_io_ptw_req_0_bits_vpn; // @[MemBlock.scala 245:{24,24}]
  wire  io_ptw_req_0_valid_hit0 = ptw_resp_next_data_entry_tag[26:18] == dtlb_ld_0_ptw_req_0_bits_vpn[26:18]; // @[MMUBundle.scala 581:48]
  wire  io_ptw_req_0_valid_hit1 = ptw_resp_next_data_entry_tag[17:9] == dtlb_ld_0_ptw_req_0_bits_vpn[17:9]; // @[MMUBundle.scala 582:48]
  wire  io_ptw_req_0_valid_hit2 = ptw_resp_next_data_entry_tag[8:0] == dtlb_ld_0_ptw_req_0_bits_vpn[8:0]; // @[MMUBundle.scala 583:50]
  wire  _io_ptw_req_0_valid_T_6 = ptw_resp_next_data_entry_level == 2'h1 ? io_ptw_req_0_valid_hit1 &
    io_ptw_req_0_valid_hit0 : io_ptw_req_0_valid_hit0; // @[MMUBundle.scala 585:78]
  wire  _io_ptw_req_0_valid_T_7 = ptw_resp_next_data_entry_level == 2'h2 ? io_ptw_req_0_valid_hit2 &
    io_ptw_req_0_valid_hit1 & io_ptw_req_0_valid_hit0 : _io_ptw_req_0_valid_T_6; // @[MMUBundle.scala 585:22]
  wire  dtlb_ld_0_ptw_req_0_valid = dtlb_ld_tlb_ld_io_ptw_req_0_valid; // @[MemBlock.scala 245:{24,24}]
  wire [26:0] dtlb_ld_0_ptw_req_1_bits_vpn = dtlb_ld_tlb_ld_io_ptw_req_1_bits_vpn; // @[MemBlock.scala 245:{24,24}]
  wire  io_ptw_req_1_valid_hit0 = ptw_resp_next_data_entry_tag[26:18] == dtlb_ld_0_ptw_req_1_bits_vpn[26:18]; // @[MMUBundle.scala 581:48]
  wire  io_ptw_req_1_valid_hit1 = ptw_resp_next_data_entry_tag[17:9] == dtlb_ld_0_ptw_req_1_bits_vpn[17:9]; // @[MMUBundle.scala 582:48]
  wire  io_ptw_req_1_valid_hit2 = ptw_resp_next_data_entry_tag[8:0] == dtlb_ld_0_ptw_req_1_bits_vpn[8:0]; // @[MMUBundle.scala 583:50]
  wire  _io_ptw_req_1_valid_T_6 = ptw_resp_next_data_entry_level == 2'h1 ? io_ptw_req_1_valid_hit1 &
    io_ptw_req_1_valid_hit0 : io_ptw_req_1_valid_hit0; // @[MMUBundle.scala 585:78]
  wire  _io_ptw_req_1_valid_T_7 = ptw_resp_next_data_entry_level == 2'h2 ? io_ptw_req_1_valid_hit2 &
    io_ptw_req_1_valid_hit1 & io_ptw_req_1_valid_hit0 : _io_ptw_req_1_valid_T_6; // @[MMUBundle.scala 585:22]
  wire  dtlb_ld_0_ptw_req_1_valid = dtlb_ld_tlb_ld_io_ptw_req_1_valid; // @[MemBlock.scala 245:{24,24}]
  wire [1:0] vector_hit_hi = {ptw_resp_next_vector_2,ptw_resp_next_vector_3}; // @[Cat.scala 31:58]
  wire [2:0] _vector_hit_T_2 = {ptw_resp_next_vector_2,ptw_resp_next_vector_3,ptw_resp_next_vector_4}; // @[Cat.scala 31:58]
  wire  vector_hit_2 = |_vector_hit_T_2; // @[MemBlock.scala 290:65]
  wire [26:0] dtlb_st_0_ptw_req_0_bits_vpn = dtlb_st_tlb_st_io_ptw_req_0_bits_vpn; // @[MemBlock.scala 249:{24,24}]
  wire  io_ptw_req_2_valid_hit0 = ptw_resp_next_data_entry_tag[26:18] == dtlb_st_0_ptw_req_0_bits_vpn[26:18]; // @[MMUBundle.scala 581:48]
  wire  io_ptw_req_2_valid_hit1 = ptw_resp_next_data_entry_tag[17:9] == dtlb_st_0_ptw_req_0_bits_vpn[17:9]; // @[MMUBundle.scala 582:48]
  wire  io_ptw_req_2_valid_hit2 = ptw_resp_next_data_entry_tag[8:0] == dtlb_st_0_ptw_req_0_bits_vpn[8:0]; // @[MMUBundle.scala 583:50]
  wire  _io_ptw_req_2_valid_T_6 = ptw_resp_next_data_entry_level == 2'h1 ? io_ptw_req_2_valid_hit1 &
    io_ptw_req_2_valid_hit0 : io_ptw_req_2_valid_hit0; // @[MMUBundle.scala 585:78]
  wire  _io_ptw_req_2_valid_T_7 = ptw_resp_next_data_entry_level == 2'h2 ? io_ptw_req_2_valid_hit2 &
    io_ptw_req_2_valid_hit1 & io_ptw_req_2_valid_hit0 : _io_ptw_req_2_valid_T_6; // @[MMUBundle.scala 585:22]
  wire  dtlb_st_0_ptw_req_0_valid = dtlb_st_tlb_st_io_ptw_req_0_valid; // @[MemBlock.scala 249:{24,24}]
  wire [26:0] dtlb_st_0_ptw_req_1_bits_vpn = dtlb_st_tlb_st_io_ptw_req_1_bits_vpn; // @[MemBlock.scala 249:{24,24}]
  wire  io_ptw_req_3_valid_hit0 = ptw_resp_next_data_entry_tag[26:18] == dtlb_st_0_ptw_req_1_bits_vpn[26:18]; // @[MMUBundle.scala 581:48]
  wire  io_ptw_req_3_valid_hit1 = ptw_resp_next_data_entry_tag[17:9] == dtlb_st_0_ptw_req_1_bits_vpn[17:9]; // @[MMUBundle.scala 582:48]
  wire  io_ptw_req_3_valid_hit2 = ptw_resp_next_data_entry_tag[8:0] == dtlb_st_0_ptw_req_1_bits_vpn[8:0]; // @[MMUBundle.scala 583:50]
  wire  _io_ptw_req_3_valid_T_6 = ptw_resp_next_data_entry_level == 2'h1 ? io_ptw_req_3_valid_hit1 &
    io_ptw_req_3_valid_hit0 : io_ptw_req_3_valid_hit0; // @[MMUBundle.scala 585:78]
  wire  _io_ptw_req_3_valid_T_7 = ptw_resp_next_data_entry_level == 2'h2 ? io_ptw_req_3_valid_hit2 &
    io_ptw_req_3_valid_hit1 & io_ptw_req_3_valid_hit0 : _io_ptw_req_3_valid_T_6; // @[MMUBundle.scala 585:22]
  wire  dtlb_st_0_ptw_req_1_valid = dtlb_st_tlb_st_io_ptw_req_1_valid; // @[MemBlock.scala 249:{24,24}]
  reg [1:0] tdata_0_matchType; // @[MemBlock.scala 324:22]
  reg  tdata_0_select; // @[MemBlock.scala 324:22]
  reg  tdata_0_chain; // @[MemBlock.scala 324:22]
  reg [63:0] tdata_0_tdata2; // @[MemBlock.scala 324:22]
  reg [1:0] tdata_1_matchType; // @[MemBlock.scala 324:22]
  reg  tdata_1_select; // @[MemBlock.scala 324:22]
  reg [63:0] tdata_1_tdata2; // @[MemBlock.scala 324:22]
  reg [1:0] tdata_2_matchType; // @[MemBlock.scala 324:22]
  reg  tdata_2_select; // @[MemBlock.scala 324:22]
  reg  tdata_2_chain; // @[MemBlock.scala 324:22]
  reg [63:0] tdata_2_tdata2; // @[MemBlock.scala 324:22]
  reg [1:0] tdata_3_matchType; // @[MemBlock.scala 324:22]
  reg  tdata_3_select; // @[MemBlock.scala 324:22]
  reg [63:0] tdata_3_tdata2; // @[MemBlock.scala 324:22]
  reg [1:0] tdata_4_matchType; // @[MemBlock.scala 324:22]
  reg  tdata_4_select; // @[MemBlock.scala 324:22]
  reg [63:0] tdata_4_tdata2; // @[MemBlock.scala 324:22]
  reg [1:0] tdata_5_matchType; // @[MemBlock.scala 324:22]
  reg  tdata_5_select; // @[MemBlock.scala 324:22]
  reg [63:0] tdata_5_tdata2; // @[MemBlock.scala 324:22]
  reg  tEnable_0; // @[MemBlock.scala 325:24]
  reg  tEnable_1; // @[MemBlock.scala 325:24]
  reg  tEnable_2; // @[MemBlock.scala 325:24]
  reg  tEnable_3; // @[MemBlock.scala 325:24]
  reg  tEnable_4; // @[MemBlock.scala 325:24]
  reg  tEnable_5; // @[MemBlock.scala 325:24]
  wire [1:0] _tdata_csrCtrl_delay_io_out_mem_trigger_t_bits_addr_matchType =
    csrCtrl_delay_io_out_mem_trigger_t_bits_tdata_matchType; // @[MemBlock.scala 329:{44,44}]
  wire [63:0] _tdata_csrCtrl_delay_io_out_mem_trigger_t_bits_addr_tdata2 =
    csrCtrl_delay_io_out_mem_trigger_t_bits_tdata_tdata2; // @[MemBlock.scala 329:{44,44}]
  wire  fastMatchVec_0 = io_loadFastMatch_0[0]; // @[MemBlock.scala 390:65]
  wire  fastMatchVec_1 = io_loadFastMatch_0[1]; // @[MemBlock.scala 390:65]
  wire  _LoadUnit_0_io_fastpathIn_valid_WIRE_1 = LoadUnit_1_io_fastpathOut_valid; // @[MemBlock.scala 391:{48,48}]
  wire  _LoadUnit_0_io_fastpathIn_valid_WIRE_0 = LoadUnit_0_io_fastpathOut_valid; // @[MemBlock.scala 391:{48,48}]
  wire [1:0] _LoadUnit_0_io_fastpathIn_valid_T = {_LoadUnit_0_io_fastpathIn_valid_WIRE_1,
    _LoadUnit_0_io_fastpathIn_valid_WIRE_0}; // @[MemBlock.scala 391:63]
  wire  hit__0 = LoadUnit_0_io_trigger_0_addrHit & ~tdata_2_select; // @[MemBlock.scala 420:52]
  wire  hit__1 = LoadUnit_0_io_trigger_1_addrHit & ~tdata_3_select; // @[MemBlock.scala 420:52]
  wire  hit__2 = LoadUnit_0_io_trigger_2_addrHit & ~tdata_5_select; // @[MemBlock.scala 420:52]
  wire  _io_writeback_0_bits_uop_cf_trigger_backendHit_2_T = hit__0 & hit__1; // @[MemBlock.scala 426:67]
  wire  _GEN_188 = tdata_2_chain ? hit__0 & hit__1 : hit__0; // @[MemBlock.scala 425:26 426:57 421:74]
  wire  _GEN_189 = tdata_2_chain ? _io_writeback_0_bits_uop_cf_trigger_backendHit_2_T : hit__1; // @[MemBlock.scala 425:26 427:57 421:74]
  wire  _GEN_190 = ~io_writeback_0_bits_uop_cf_trigger_backendEn_1 ? 1'h0 : hit__2; // @[MemBlock.scala 429:61 430:57 421:74]
  wire  fastMatchVec_0_1 = io_loadFastMatch_1[1]; // @[MemBlock.scala 390:65]
  wire  fastMatchVec_1_1 = io_loadFastMatch_1[0]; // @[MemBlock.scala 390:65]
  wire [1:0] _LoadUnit_1_io_fastpathIn_valid_T = {_LoadUnit_0_io_fastpathIn_valid_WIRE_0,
    _LoadUnit_0_io_fastpathIn_valid_WIRE_1}; // @[MemBlock.scala 391:63]
  wire  hit_1_0 = LoadUnit_1_io_trigger_0_addrHit & ~tdata_2_select; // @[MemBlock.scala 420:52]
  wire  hit_1_1 = LoadUnit_1_io_trigger_1_addrHit & ~tdata_3_select; // @[MemBlock.scala 420:52]
  wire  hit_1_2 = LoadUnit_1_io_trigger_2_addrHit & ~tdata_5_select; // @[MemBlock.scala 420:52]
  wire  _io_writeback_1_bits_uop_cf_trigger_backendHit_2_T = hit_1_0 & hit_1_1; // @[MemBlock.scala 426:67]
  wire  _GEN_191 = tdata_2_chain ? hit_1_0 & hit_1_1 : hit_1_0; // @[MemBlock.scala 425:26 426:57 421:74]
  wire  _GEN_192 = tdata_2_chain ? _io_writeback_1_bits_uop_cf_trigger_backendHit_2_T : hit_1_1; // @[MemBlock.scala 425:26 427:57 421:74]
  wire  _GEN_193 = ~io_writeback_1_bits_uop_cf_trigger_backendEn_1 ? 1'h0 : hit_1_2; // @[MemBlock.scala 429:61 430:57 421:74]
  wire [63:0] _GEN_673 = {{25'd0}, io_writeback_2_bits_debug_vaddr}; // @[Trigger.scala 27:24]
  wire  hit_0_equal = _GEN_673 == tdata_0_tdata2; // @[Trigger.scala 27:24]
  wire  hit_0_greater = _GEN_673 >= tdata_0_tdata2; // @[Trigger.scala 28:26]
  wire  hit_0_less = _GEN_673 <= tdata_0_tdata2; // @[Trigger.scala 29:23]
  wire  _hit_0_res_T_3 = 2'h2 == tdata_0_matchType ? hit_0_greater : 2'h0 == tdata_0_matchType & hit_0_equal; // @[Mux.scala 81:58]
  wire  hit_0_res = 2'h3 == tdata_0_matchType ? hit_0_less : _hit_0_res_T_3; // @[Mux.scala 81:58]
  wire  _hit_0_T_5 = hit_0_res & tEnable_0; // @[Trigger.scala 34:9]
  wire  hit_2_0 = ~tdata_0_select & _hit_0_T_5; // @[MemBlock.scala 492:54]
  wire  hit_1_equal = _GEN_673 == tdata_1_tdata2; // @[Trigger.scala 27:24]
  wire  hit_1_greater = _GEN_673 >= tdata_1_tdata2; // @[Trigger.scala 28:26]
  wire  hit_1_less = _GEN_673 <= tdata_1_tdata2; // @[Trigger.scala 29:23]
  wire  _hit_1_res_T_3 = 2'h2 == tdata_1_matchType ? hit_1_greater : 2'h0 == tdata_1_matchType & hit_1_equal; // @[Mux.scala 81:58]
  wire  hit_1_res = 2'h3 == tdata_1_matchType ? hit_1_less : _hit_1_res_T_3; // @[Mux.scala 81:58]
  wire  _hit_1_T_5 = hit_1_res & tEnable_1; // @[Trigger.scala 34:9]
  wire  hit_2_1 = ~tdata_1_select & _hit_1_T_5; // @[MemBlock.scala 492:54]
  wire  hit_2_equal = _GEN_673 == tdata_4_tdata2; // @[Trigger.scala 27:24]
  wire  hit_2_greater = _GEN_673 >= tdata_4_tdata2; // @[Trigger.scala 28:26]
  wire  hit_2_less = _GEN_673 <= tdata_4_tdata2; // @[Trigger.scala 29:23]
  wire  _hit_2_res_T_3 = 2'h2 == tdata_4_matchType ? hit_2_greater : 2'h0 == tdata_4_matchType & hit_2_equal; // @[Mux.scala 81:58]
  wire  hit_2_res = 2'h3 == tdata_4_matchType ? hit_2_less : _hit_2_res_T_3; // @[Mux.scala 81:58]
  wire  _hit_2_T_5 = hit_2_res & tEnable_4; // @[Trigger.scala 34:9]
  wire  hit_2_2 = ~tdata_4_select & _hit_2_T_5; // @[MemBlock.scala 492:54]
  wire  _io_writeback_0_bits_uop_cf_trigger_backendHit_0_T = hit_2_0 & hit_2_1; // @[MemBlock.scala 502:68]
  wire  _GEN_194 = tdata_0_chain ? hit_2_0 & hit_2_1 : loadWritebackOverride_uop_cf_trigger_backendHit_0; // @[MemBlock.scala 193:16 501:27 502:58]
  wire  _GEN_195 = tdata_0_chain ? _io_writeback_0_bits_uop_cf_trigger_backendHit_0_T :
    loadWritebackOverride_uop_cf_trigger_backendHit_1; // @[MemBlock.scala 193:16 501:27 503:58]
  wire  _GEN_196 = ~io_writeback_2_bits_uop_cf_trigger_backendEn_0 ? 1'h0 : hit_2_2; // @[MemBlock.scala 506:55 507:51 498:68]
  wire  _GEN_197 = io_writeback_2_valid & hit_2_0; // @[MemBlock.scala 193:16 489:26 498:68]
  wire  _GEN_198 = io_writeback_2_valid & hit_2_1; // @[MemBlock.scala 193:16 489:26 498:68]
  wire  _GEN_199 = io_writeback_2_valid & _GEN_196; // @[MemBlock.scala 193:16 489:26]
  wire  _GEN_200 = io_writeback_2_valid ? _GEN_194 : loadWritebackOverride_uop_cf_trigger_backendHit_0; // @[MemBlock.scala 193:16 489:26]
  wire  _GEN_201 = io_writeback_2_valid ? _GEN_195 : loadWritebackOverride_uop_cf_trigger_backendHit_1; // @[MemBlock.scala 193:16 489:26]
  wire [63:0] _GEN_682 = {{25'd0}, io_writeback_3_bits_debug_vaddr}; // @[Trigger.scala 27:24]
  wire  hit_0_equal_1 = _GEN_682 == tdata_0_tdata2; // @[Trigger.scala 27:24]
  wire  hit_0_greater_1 = _GEN_682 >= tdata_0_tdata2; // @[Trigger.scala 28:26]
  wire  hit_0_less_1 = _GEN_682 <= tdata_0_tdata2; // @[Trigger.scala 29:23]
  wire  _hit_0_res_T_8 = 2'h2 == tdata_0_matchType ? hit_0_greater_1 : 2'h0 == tdata_0_matchType & hit_0_equal_1; // @[Mux.scala 81:58]
  wire  hit_0_res_1 = 2'h3 == tdata_0_matchType ? hit_0_less_1 : _hit_0_res_T_8; // @[Mux.scala 81:58]
  wire  _hit_0_T_8 = hit_0_res_1 & tEnable_0; // @[Trigger.scala 34:9]
  wire  hit_3_0 = ~tdata_0_select & _hit_0_T_8; // @[MemBlock.scala 492:54]
  wire  hit_1_equal_1 = _GEN_682 == tdata_1_tdata2; // @[Trigger.scala 27:24]
  wire  hit_1_greater_1 = _GEN_682 >= tdata_1_tdata2; // @[Trigger.scala 28:26]
  wire  hit_1_less_1 = _GEN_682 <= tdata_1_tdata2; // @[Trigger.scala 29:23]
  wire  _hit_1_res_T_8 = 2'h2 == tdata_1_matchType ? hit_1_greater_1 : 2'h0 == tdata_1_matchType & hit_1_equal_1; // @[Mux.scala 81:58]
  wire  hit_1_res_1 = 2'h3 == tdata_1_matchType ? hit_1_less_1 : _hit_1_res_T_8; // @[Mux.scala 81:58]
  wire  _hit_1_T_8 = hit_1_res_1 & tEnable_1; // @[Trigger.scala 34:9]
  wire  hit_3_1 = ~tdata_1_select & _hit_1_T_8; // @[MemBlock.scala 492:54]
  wire  hit_2_equal_1 = _GEN_682 == tdata_4_tdata2; // @[Trigger.scala 27:24]
  wire  hit_2_greater_1 = _GEN_682 >= tdata_4_tdata2; // @[Trigger.scala 28:26]
  wire  hit_2_less_1 = _GEN_682 <= tdata_4_tdata2; // @[Trigger.scala 29:23]
  wire  _hit_2_res_T_8 = 2'h2 == tdata_4_matchType ? hit_2_greater_1 : 2'h0 == tdata_4_matchType & hit_2_equal_1; // @[Mux.scala 81:58]
  wire  hit_2_res_1 = 2'h3 == tdata_4_matchType ? hit_2_less_1 : _hit_2_res_T_8; // @[Mux.scala 81:58]
  wire  _hit_2_T_8 = hit_2_res_1 & tEnable_4; // @[Trigger.scala 34:9]
  wire  hit_3_2 = ~tdata_4_select & _hit_2_T_8; // @[MemBlock.scala 492:54]
  wire  _io_writeback_1_bits_uop_cf_trigger_backendHit_0_T = hit_3_0 & hit_3_1; // @[MemBlock.scala 502:68]
  wire  _GEN_202 = tdata_0_chain ? hit_3_0 & hit_3_1 : LoadUnit_1_io_loadOut_bits_uop_cf_trigger_backendHit_0; // @[MemBlock.scala 193:16 501:27 502:58]
  wire  _GEN_203 = tdata_0_chain ? _io_writeback_1_bits_uop_cf_trigger_backendHit_0_T :
    LoadUnit_1_io_loadOut_bits_uop_cf_trigger_backendHit_1; // @[MemBlock.scala 193:16 501:27 503:58]
  wire  _GEN_204 = ~io_writeback_3_bits_uop_cf_trigger_backendEn_0 ? 1'h0 : hit_3_2; // @[MemBlock.scala 506:55 507:51 498:68]
  wire  _GEN_208 = io_writeback_3_valid ? _GEN_202 : LoadUnit_1_io_loadOut_bits_uop_cf_trigger_backendHit_0; // @[MemBlock.scala 193:16 489:26]
  wire  _GEN_209 = io_writeback_3_valid ? _GEN_203 : LoadUnit_1_io_loadOut_bits_uop_cf_trigger_backendHit_1; // @[MemBlock.scala 193:16 489:26]
  wire  _GEN_210 = lsq_io_mmioStout_valid & ~StoreUnit_0_io_stout_valid | StoreUnit_0_io_stout_valid; // @[MemBlock.scala 193:16 514:66 515:20]
  wire  _GEN_220 = lsq_io_mmioStout_valid & ~StoreUnit_0_io_stout_valid ? 1'h0 :
    StoreUnit_0_io_stout_bits_uop_cf_exceptionVec_6; // @[MemBlock.scala 193:16 514:66 516:20]
  wire  _GEN_221 = lsq_io_mmioStout_valid & ~StoreUnit_0_io_stout_valid ? 1'h0 :
    StoreUnit_0_io_stout_bits_uop_cf_exceptionVec_7; // @[MemBlock.scala 193:16 514:66 516:20]
  wire  _GEN_229 = lsq_io_mmioStout_valid & ~StoreUnit_0_io_stout_valid ? 1'h0 :
    StoreUnit_0_io_stout_bits_uop_cf_exceptionVec_15; // @[MemBlock.scala 193:16 514:66 516:20]
  wire  _GEN_234 = lsq_io_mmioStout_valid & ~StoreUnit_0_io_stout_valid ?
    lsq_io_mmioStout_bits_uop_cf_trigger_backendEn_0 : StoreUnit_0_io_stout_bits_uop_cf_trigger_backendEn_0; // @[MemBlock.scala 193:16 514:66 516:20]
  wire  _GEN_236 = lsq_io_mmioStout_valid & ~StoreUnit_0_io_stout_valid ? 1'h0 : _GEN_197; // @[MemBlock.scala 514:66 516:20]
  wire  _GEN_237 = lsq_io_mmioStout_valid & ~StoreUnit_0_io_stout_valid ? 1'h0 : _GEN_198; // @[MemBlock.scala 514:66 516:20]
  wire  _GEN_240 = lsq_io_mmioStout_valid & ~StoreUnit_0_io_stout_valid ? 1'h0 : _GEN_199; // @[MemBlock.scala 514:66 516:20]
  wire  _GEN_302 = lsq_io_mmioStout_valid & ~StoreUnit_0_io_stout_valid ? lsq_io_mmioStout_bits_uop_robIdx_flag :
    StoreUnit_0_io_stout_bits_uop_robIdx_flag; // @[MemBlock.scala 193:16 514:66 516:20]
  wire [4:0] _WIRE__0_bits_uop_robIdx_value = StoreUnit_0_io_stout_bits_uop_robIdx_value; // @[MemBlock.scala 193:{41,41}]
  wire [4:0] _GEN_303 = lsq_io_mmioStout_valid & ~StoreUnit_0_io_stout_valid ? lsq_io_mmioStout_bits_uop_robIdx_value :
    _WIRE__0_bits_uop_robIdx_value; // @[MemBlock.scala 193:16 514:66 516:20]
  wire  _GEN_397 = lsq_io_mmioStout_valid & ~StoreUnit_0_io_stout_valid | StoreUnit_0_io_stout_bits_debug_isMMIO; // @[MemBlock.scala 193:16 514:66 516:20]
  wire [38:0] _WIRE__0_bits_debug_vaddr = StoreUnit_0_io_stout_bits_debug_vaddr; // @[MemBlock.scala 193:{41,41}]
  wire [38:0] _GEN_400 = lsq_io_mmioStout_valid & ~StoreUnit_0_io_stout_valid ? 39'h0 : _WIRE__0_bits_debug_vaddr; // @[MemBlock.scala 193:16 514:66 516:20]
  reg  io_fenceToSbuffer_sbIsEmpty_REG; // @[MemBlock.scala 567:41]
  reg  sbuffer_io_flush_valid_REG; // @[MemBlock.scala 572:36]
  reg [1:0] state; // @[MemBlock.scala 590:22]
  wire  st_atomics_0 = io_issue_2_valid & io_issue_2_bits_uop_ctrl_fuType[1]; // @[MemBlock.scala 595:34]
  wire  st_atomics_1 = io_issue_3_valid & io_issue_3_bits_uop_ctrl_fuType[1]; // @[MemBlock.scala 595:34]
  wire  st_data_atomics_0 = stdExeUnits_0_io_out_valid & stdExeUnits_0_io_out_bits_uop_ctrl_fuType[1]; // @[MemBlock.scala 599:21]
  wire  st_data_atomics_1 = stdExeUnits_1_io_out_valid & stdExeUnits_1_io_out_bits_uop_ctrl_fuType[1]; // @[MemBlock.scala 599:21]
  wire  _T_43 = state == 2'h1; // @[MemBlock.scala 611:53]
  wire  _T_44 = state == 2'h2; // @[MemBlock.scala 611:53]
  wire [63:0] _atomicsUnit_io_in_bits_T = st_atomics_0 ? io_issue_2_bits_src_0 : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _atomicsUnit_io_in_bits_T_1 = st_atomics_1 ? io_issue_3_bits_src_0 : 64'h0; // @[Mux.scala 27:73]
  wire [4:0] _atomicsUnit_io_in_bits_T_54 = st_atomics_0 ? io_issue_2_bits_uop_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [4:0] _atomicsUnit_io_in_bits_T_55 = st_atomics_1 ? io_issue_3_bits_uop_robIdx_value : 5'h0; // @[Mux.scala 27:73]
  wire [5:0] _atomicsUnit_io_in_bits_T_63 = st_atomics_0 ? io_issue_2_bits_uop_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [5:0] _atomicsUnit_io_in_bits_T_64 = st_atomics_1 ? io_issue_3_bits_uop_pdest : 6'h0; // @[Mux.scala 27:73]
  wire [6:0] _atomicsUnit_io_in_bits_T_162 = st_atomics_0 ? io_issue_2_bits_uop_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [6:0] _atomicsUnit_io_in_bits_T_163 = st_atomics_1 ? io_issue_3_bits_uop_ctrl_fuOpType : 7'h0; // @[Mux.scala 27:73]
  wire [63:0] _atomicsUnit_io_storeDataIn_bits_T_243 = st_data_atomics_0 ? stdExeUnits_0_io_out_bits_data : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _atomicsUnit_io_storeDataIn_bits_T_244 = st_data_atomics_1 ? stdExeUnits_1_io_out_bits_data : 64'h0; // @[Mux.scala 27:73]
  wire [3:0] _atomicsUnit_io_rsIdx_T = st_atomics_0 ? io_rsfeedback_0_rsIdx : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _atomicsUnit_io_rsIdx_T_1 = st_atomics_1 ? io_rsfeedback_1_rsIdx : 4'h0; // @[Mux.scala 27:73]
  wire  dtlb_ld_0_requestor_0_resp_valid = dtlb_ld_tlb_ld_io_requestor_0_resp_valid; // @[MemBlock.scala 245:{24,24}]
  reg  atomicsException; // @[MemBlock.scala 661:33]
  wire  _GEN_670 = atomicsUnit_io_exceptionAddr_valid | atomicsException; // @[MemBlock.scala 664:51 665:22 661:33]
  reg [38:0] atomicsExceptionAddress; // @[Reg.scala 16:16]
  reg [38:0] io_lsqio_exceptionAddr_vaddr_REG; // @[MemBlock.scala 668:42]
  wire [1:0] ldDeqCount = io_issue_0_valid + io_issue_1_valid; // @[Bitwise.scala 48:55]
  wire [1:0] _stDeqCount_T = io_issue_2_valid + io_issue_3_valid; // @[Bitwise.scala 48:55]
  wire [1:0] _stDeqCount_T_2 = io_issue_4_valid + io_issue_5_valid; // @[Bitwise.scala 48:55]
  wire [2:0] stDeqCount = _stDeqCount_T + _stDeqCount_T_2; // @[Bitwise.scala 48:55]
  reg [5:0] io_perf_0_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg [5:0] io_perf_0_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  reg [5:0] io_perf_1_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg [5:0] io_perf_1_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  reg [5:0] io_perf_2_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg [5:0] io_perf_2_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  reg [5:0] io_perf_3_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg [5:0] io_perf_3_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  reg [5:0] io_perf_4_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg [5:0] io_perf_4_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  reg [5:0] io_perf_5_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg [5:0] io_perf_5_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  reg [5:0] io_perf_6_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg [5:0] io_perf_6_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  reg [5:0] io_perf_7_value_REG; // @[PerfCounterUtils.scala 188:35]
  reg [5:0] io_perf_7_value_REG_1; // @[PerfCounterUtils.scala 188:27]
  DCacheWrapper dcache ( // @[MemBlock.scala 47:26]
    .clock(dcache_clock),
    .reset(dcache_reset),
    .auto_client_out_a_ready(dcache_auto_client_out_a_ready),
    .auto_client_out_a_valid(dcache_auto_client_out_a_valid),
    .auto_client_out_a_bits_opcode(dcache_auto_client_out_a_bits_opcode),
    .auto_client_out_a_bits_param(dcache_auto_client_out_a_bits_param),
    .auto_client_out_a_bits_size(dcache_auto_client_out_a_bits_size),
    .auto_client_out_a_bits_source(dcache_auto_client_out_a_bits_source),
    .auto_client_out_a_bits_address(dcache_auto_client_out_a_bits_address),
    .auto_client_out_a_bits_mask(dcache_auto_client_out_a_bits_mask),
    .auto_client_out_bready(dcache_auto_client_out_bready),
    .auto_client_out_bvalid(dcache_auto_client_out_bvalid),
    .auto_client_out_bparam(dcache_auto_client_out_bparam),
    .auto_client_out_baddress(dcache_auto_client_out_baddress),
    .auto_client_out_bdata(dcache_auto_client_out_bdata),
    .auto_client_out_c_ready(dcache_auto_client_out_c_ready),
    .auto_client_out_c_valid(dcache_auto_client_out_c_valid),
    .auto_client_out_c_bits_opcode(dcache_auto_client_out_c_bits_opcode),
    .auto_client_out_c_bits_param(dcache_auto_client_out_c_bits_param),
    .auto_client_out_c_bits_size(dcache_auto_client_out_c_bits_size),
    .auto_client_out_c_bits_source(dcache_auto_client_out_c_bits_source),
    .auto_client_out_c_bits_address(dcache_auto_client_out_c_bits_address),
    .auto_client_out_c_bits_echo_blockisdirty(dcache_auto_client_out_c_bits_echo_blockisdirty),
    .auto_client_out_c_bits_data(dcache_auto_client_out_c_bits_data),
    .auto_client_out_d_ready(dcache_auto_client_out_d_ready),
    .auto_client_out_d_valid(dcache_auto_client_out_d_valid),
    .auto_client_out_d_bits_opcode(dcache_auto_client_out_d_bits_opcode),
    .auto_client_out_d_bits_param(dcache_auto_client_out_d_bits_param),
    .auto_client_out_d_bits_size(dcache_auto_client_out_d_bits_size),
    .auto_client_out_d_bits_source(dcache_auto_client_out_d_bits_source),
    .auto_client_out_d_bits_sink(dcache_auto_client_out_d_bits_sink),
    .auto_client_out_d_bits_denied(dcache_auto_client_out_d_bits_denied),
    .auto_client_out_d_bits_echo_blockisdirty(dcache_auto_client_out_d_bits_echo_blockisdirty),
    .auto_client_out_d_bits_data(dcache_auto_client_out_d_bits_data),
    .auto_client_out_d_bits_corrupt(dcache_auto_client_out_d_bits_corrupt),
    .auto_client_out_e_ready(dcache_auto_client_out_e_ready),
    .auto_client_out_e_valid(dcache_auto_client_out_e_valid),
    .auto_client_out_e_bits_sink(dcache_auto_client_out_e_bits_sink),
    .io_lsu_load_0_req_ready(dcache_io_lsu_load_0_req_ready),
    .io_lsu_load_0_req_valid(dcache_io_lsu_load_0_req_valid),
    .io_lsu_load_0_req_bits_cmd(dcache_io_lsu_load_0_req_bits_cmd),
    .io_lsu_load_0_req_bits_addr(dcache_io_lsu_load_0_req_bits_addr),
    .io_lsu_load_0_req_bits_instrtype(dcache_io_lsu_load_0_req_bits_instrtype),
    .io_lsu_load_0_req_bits_replayCarry_real_way_en(dcache_io_lsu_load_0_req_bits_replayCarry_real_way_en),
    .io_lsu_load_0_req_bits_replayCarry_valid(dcache_io_lsu_load_0_req_bits_replayCarry_valid),
    .io_lsu_load_0_resp_bits_data_delayed(dcache_io_lsu_load_0_resp_bits_data_delayed),
    .io_lsu_load_0_resp_bits_miss(dcache_io_lsu_load_0_resp_bits_miss),
    .io_lsu_load_0_resp_bits_replay(dcache_io_lsu_load_0_resp_bits_replay),
    .io_lsu_load_0_resp_bits_replayCarry_real_way_en(dcache_io_lsu_load_0_resp_bits_replayCarry_real_way_en),
    .io_lsu_load_0_resp_bits_replayCarry_valid(dcache_io_lsu_load_0_resp_bits_replayCarry_valid),
    .io_lsu_load_0_resp_bits_tag_error(dcache_io_lsu_load_0_resp_bits_tag_error),
    .io_lsu_load_0_resp_bits_mshr_id(dcache_io_lsu_load_0_resp_bits_mshr_id),
    .io_lsu_load_0_resp_bits_error_delayed(dcache_io_lsu_load_0_resp_bits_error_delayed),
    .io_lsu_load_0_s1_kill(dcache_io_lsu_load_0_s1_kill),
    .io_lsu_load_0_s2_kill(dcache_io_lsu_load_0_s2_kill),
    .io_lsu_load_0_s1_paddr_dup_lsu(dcache_io_lsu_load_0_s1_paddr_dup_lsu),
    .io_lsu_load_0_s1_paddr_dup_dcache(dcache_io_lsu_load_0_s1_paddr_dup_dcache),
    .io_lsu_load_0_s1_bank_conflict(dcache_io_lsu_load_0_s1_bank_conflict),
    .io_lsu_load_1_req_ready(dcache_io_lsu_load_1_req_ready),
    .io_lsu_load_1_req_valid(dcache_io_lsu_load_1_req_valid),
    .io_lsu_load_1_req_bits_cmd(dcache_io_lsu_load_1_req_bits_cmd),
    .io_lsu_load_1_req_bits_addr(dcache_io_lsu_load_1_req_bits_addr),
    .io_lsu_load_1_req_bits_instrtype(dcache_io_lsu_load_1_req_bits_instrtype),
    .io_lsu_load_1_req_bits_replayCarry_real_way_en(dcache_io_lsu_load_1_req_bits_replayCarry_real_way_en),
    .io_lsu_load_1_req_bits_replayCarry_valid(dcache_io_lsu_load_1_req_bits_replayCarry_valid),
    .io_lsu_load_1_resp_bits_data_delayed(dcache_io_lsu_load_1_resp_bits_data_delayed),
    .io_lsu_load_1_resp_bits_miss(dcache_io_lsu_load_1_resp_bits_miss),
    .io_lsu_load_1_resp_bits_replay(dcache_io_lsu_load_1_resp_bits_replay),
    .io_lsu_load_1_resp_bits_replayCarry_real_way_en(dcache_io_lsu_load_1_resp_bits_replayCarry_real_way_en),
    .io_lsu_load_1_resp_bits_replayCarry_valid(dcache_io_lsu_load_1_resp_bits_replayCarry_valid),
    .io_lsu_load_1_resp_bits_tag_error(dcache_io_lsu_load_1_resp_bits_tag_error),
    .io_lsu_load_1_resp_bits_mshr_id(dcache_io_lsu_load_1_resp_bits_mshr_id),
    .io_lsu_load_1_resp_bits_error_delayed(dcache_io_lsu_load_1_resp_bits_error_delayed),
    .io_lsu_load_1_s1_kill(dcache_io_lsu_load_1_s1_kill),
    .io_lsu_load_1_s2_kill(dcache_io_lsu_load_1_s2_kill),
    .io_lsu_load_1_s1_paddr_dup_lsu(dcache_io_lsu_load_1_s1_paddr_dup_lsu),
    .io_lsu_load_1_s1_paddr_dup_dcache(dcache_io_lsu_load_1_s1_paddr_dup_dcache),
    .io_lsu_load_1_s1_bank_conflict(dcache_io_lsu_load_1_s1_bank_conflict),
    .io_lsu_lsq_valid(dcache_io_lsu_lsq_valid),
    .io_lsu_lsq_bits_id(dcache_io_lsu_lsq_bits_id),
    .io_lsu_store_req_ready(dcache_io_lsu_store_req_ready),
    .io_lsu_store_req_valid(dcache_io_lsu_store_req_valid),
    .io_lsu_store_req_bits_vaddr(dcache_io_lsu_store_req_bits_vaddr),
    .io_lsu_store_req_bits_addr(dcache_io_lsu_store_req_bits_addr),
    .io_lsu_store_req_bits_data(dcache_io_lsu_store_req_bits_data),
    .io_lsu_store_req_bits_mask(dcache_io_lsu_store_req_bits_mask),
    .io_lsu_store_req_bits_id(dcache_io_lsu_store_req_bits_id),
    .io_lsu_store_main_pipe_hit_resp_valid(dcache_io_lsu_store_main_pipe_hit_resp_valid),
    .io_lsu_store_main_pipe_hit_resp_bits_id(dcache_io_lsu_store_main_pipe_hit_resp_bits_id),
    .io_lsu_store_refill_hit_resp_valid(dcache_io_lsu_store_refill_hit_resp_valid),
    .io_lsu_store_refill_hit_resp_bits_id(dcache_io_lsu_store_refill_hit_resp_bits_id),
    .io_lsu_store_replay_resp_valid(dcache_io_lsu_store_replay_resp_valid),
    .io_lsu_store_replay_resp_bits_id(dcache_io_lsu_store_replay_resp_bits_id),
    .io_lsu_atomics_req_ready(dcache_io_lsu_atomics_req_ready),
    .io_lsu_atomics_req_valid(dcache_io_lsu_atomics_req_valid),
    .io_lsu_atomics_req_bits_cmd(dcache_io_lsu_atomics_req_bits_cmd),
    .io_lsu_atomics_req_bits_vaddr(dcache_io_lsu_atomics_req_bits_vaddr),
    .io_lsu_atomics_req_bits_addr(dcache_io_lsu_atomics_req_bits_addr),
    .io_lsu_atomics_req_bits_word_idx(dcache_io_lsu_atomics_req_bits_word_idx),
    .io_lsu_atomics_req_bits_amo_data(dcache_io_lsu_atomics_req_bits_amo_data),
    .io_lsu_atomics_req_bits_amo_mask(dcache_io_lsu_atomics_req_bits_amo_mask),
    .io_lsu_atomics_resp_valid(dcache_io_lsu_atomics_resp_valid),
    .io_lsu_atomics_resp_bits_data(dcache_io_lsu_atomics_resp_bits_data),
    .io_lsu_atomics_resp_bits_miss(dcache_io_lsu_atomics_resp_bits_miss),
    .io_lsu_atomics_resp_bits_replay(dcache_io_lsu_atomics_resp_bits_replay),
    .io_lsu_atomics_resp_bits_error(dcache_io_lsu_atomics_resp_bits_error),
    .io_lsu_atomics_resp_bits_id(dcache_io_lsu_atomics_resp_bits_id),
    .io_lsu_atomics_block_lr(dcache_io_lsu_atomics_block_lr),
    .io_lsu_release_valid(dcache_io_lsu_release_valid),
    .io_lsu_release_bits_paddr(dcache_io_lsu_release_bits_paddr),
    .io_lsu_forward_D_0_valid(dcache_io_lsu_forward_D_0_valid),
    .io_lsu_forward_D_0_data(dcache_io_lsu_forward_D_0_data),
    .io_lsu_forward_D_0_mshrid(dcache_io_lsu_forward_D_0_mshrid),
    .io_lsu_forward_D_0_last(dcache_io_lsu_forward_D_0_last),
    .io_lsu_forward_D_1_valid(dcache_io_lsu_forward_D_1_valid),
    .io_lsu_forward_D_1_data(dcache_io_lsu_forward_D_1_data),
    .io_lsu_forward_D_1_mshrid(dcache_io_lsu_forward_D_1_mshrid),
    .io_lsu_forward_D_1_last(dcache_io_lsu_forward_D_1_last),
    .io_lsu_forward_mshr_0_valid(dcache_io_lsu_forward_mshr_0_valid),
    .io_lsu_forward_mshr_0_mshrid(dcache_io_lsu_forward_mshr_0_mshrid),
    .io_lsu_forward_mshr_0_paddr(dcache_io_lsu_forward_mshr_0_paddr),
    .io_lsu_forward_mshr_0_forward_mshr(dcache_io_lsu_forward_mshr_0_forward_mshr),
    .io_lsu_forward_mshr_0_forwardData_0(dcache_io_lsu_forward_mshr_0_forwardData_0),
    .io_lsu_forward_mshr_0_forwardData_1(dcache_io_lsu_forward_mshr_0_forwardData_1),
    .io_lsu_forward_mshr_0_forwardData_2(dcache_io_lsu_forward_mshr_0_forwardData_2),
    .io_lsu_forward_mshr_0_forwardData_3(dcache_io_lsu_forward_mshr_0_forwardData_3),
    .io_lsu_forward_mshr_0_forwardData_4(dcache_io_lsu_forward_mshr_0_forwardData_4),
    .io_lsu_forward_mshr_0_forwardData_5(dcache_io_lsu_forward_mshr_0_forwardData_5),
    .io_lsu_forward_mshr_0_forwardData_6(dcache_io_lsu_forward_mshr_0_forwardData_6),
    .io_lsu_forward_mshr_0_forwardData_7(dcache_io_lsu_forward_mshr_0_forwardData_7),
    .io_lsu_forward_mshr_0_forwardData_8(dcache_io_lsu_forward_mshr_0_forwardData_8),
    .io_lsu_forward_mshr_0_forwardData_9(dcache_io_lsu_forward_mshr_0_forwardData_9),
    .io_lsu_forward_mshr_0_forwardData_10(dcache_io_lsu_forward_mshr_0_forwardData_10),
    .io_lsu_forward_mshr_0_forwardData_11(dcache_io_lsu_forward_mshr_0_forwardData_11),
    .io_lsu_forward_mshr_0_forwardData_12(dcache_io_lsu_forward_mshr_0_forwardData_12),
    .io_lsu_forward_mshr_0_forwardData_13(dcache_io_lsu_forward_mshr_0_forwardData_13),
    .io_lsu_forward_mshr_0_forwardData_14(dcache_io_lsu_forward_mshr_0_forwardData_14),
    .io_lsu_forward_mshr_0_forwardData_15(dcache_io_lsu_forward_mshr_0_forwardData_15),
    .io_lsu_forward_mshr_0_forward_result_valid(dcache_io_lsu_forward_mshr_0_forward_result_valid),
    .io_lsu_forward_mshr_1_valid(dcache_io_lsu_forward_mshr_1_valid),
    .io_lsu_forward_mshr_1_mshrid(dcache_io_lsu_forward_mshr_1_mshrid),
    .io_lsu_forward_mshr_1_paddr(dcache_io_lsu_forward_mshr_1_paddr),
    .io_lsu_forward_mshr_1_forward_mshr(dcache_io_lsu_forward_mshr_1_forward_mshr),
    .io_lsu_forward_mshr_1_forwardData_0(dcache_io_lsu_forward_mshr_1_forwardData_0),
    .io_lsu_forward_mshr_1_forwardData_1(dcache_io_lsu_forward_mshr_1_forwardData_1),
    .io_lsu_forward_mshr_1_forwardData_2(dcache_io_lsu_forward_mshr_1_forwardData_2),
    .io_lsu_forward_mshr_1_forwardData_3(dcache_io_lsu_forward_mshr_1_forwardData_3),
    .io_lsu_forward_mshr_1_forwardData_4(dcache_io_lsu_forward_mshr_1_forwardData_4),
    .io_lsu_forward_mshr_1_forwardData_5(dcache_io_lsu_forward_mshr_1_forwardData_5),
    .io_lsu_forward_mshr_1_forwardData_6(dcache_io_lsu_forward_mshr_1_forwardData_6),
    .io_lsu_forward_mshr_1_forwardData_7(dcache_io_lsu_forward_mshr_1_forwardData_7),
    .io_lsu_forward_mshr_1_forwardData_8(dcache_io_lsu_forward_mshr_1_forwardData_8),
    .io_lsu_forward_mshr_1_forwardData_9(dcache_io_lsu_forward_mshr_1_forwardData_9),
    .io_lsu_forward_mshr_1_forwardData_10(dcache_io_lsu_forward_mshr_1_forwardData_10),
    .io_lsu_forward_mshr_1_forwardData_11(dcache_io_lsu_forward_mshr_1_forwardData_11),
    .io_lsu_forward_mshr_1_forwardData_12(dcache_io_lsu_forward_mshr_1_forwardData_12),
    .io_lsu_forward_mshr_1_forwardData_13(dcache_io_lsu_forward_mshr_1_forwardData_13),
    .io_lsu_forward_mshr_1_forwardData_14(dcache_io_lsu_forward_mshr_1_forwardData_14),
    .io_lsu_forward_mshr_1_forwardData_15(dcache_io_lsu_forward_mshr_1_forwardData_15),
    .io_lsu_forward_mshr_1_forward_result_valid(dcache_io_lsu_forward_mshr_1_forward_result_valid),
    .io_csr_distribute_csr_wvalid(dcache_io_csr_distribute_csr_wvalid),
    .io_csr_distribute_csr_waddr(dcache_io_csr_distribute_csr_waddr),
    .io_csr_distribute_csr_wdata(dcache_io_csr_distribute_csr_wdata),
    .io_csr_update_wvalid(dcache_io_csr_update_wvalid),
    .io_csr_update_waddr(dcache_io_csr_update_waddr),
    .io_csr_update_wdata(dcache_io_csr_update_wdata),
    .io_error_paddr(dcache_io_error_paddr),
    .io_error_report_to_beu(dcache_io_error_report_to_beu),
    .io_perf_0_value(dcache_io_perf_0_value),
    .io_perf_1_value(dcache_io_perf_1_value),
    .io_perf_2_value(dcache_io_perf_2_value),
    .io_perf_3_value(dcache_io_perf_3_value),
    .io_perf_4_value(dcache_io_perf_4_value),
    .io_perf_5_value(dcache_io_perf_5_value),
    .io_perf_6_value(dcache_io_perf_6_value),
    .io_perf_7_value(dcache_io_perf_7_value),
    .io_perf_8_value(dcache_io_perf_8_value),
    .io_perf_9_value(dcache_io_perf_9_value),
    .io_perf_10_value(dcache_io_perf_10_value),
    .io_perf_11_value(dcache_io_perf_11_value),
    .io_perf_12_value(dcache_io_perf_12_value),
    .io_perf_13_value(dcache_io_perf_13_value),
    .io_perf_14_value(dcache_io_perf_14_value),
    .io_perf_15_value(dcache_io_perf_15_value),
    .io_perf_16_value(dcache_io_perf_16_value),
    .io_perf_17_value(dcache_io_perf_17_value),
    .io_perf_18_value(dcache_io_perf_18_value),
    .io_perf_19_value(dcache_io_perf_19_value),
    .io_perf_20_value(dcache_io_perf_20_value),
    .io_perf_21_value(dcache_io_perf_21_value),
    .io_perf_22_value(dcache_io_perf_22_value),
    .io_perf_23_value(dcache_io_perf_23_value),
    .io_perf_24_value(dcache_io_perf_24_value),
    .io_perf_25_value(dcache_io_perf_25_value),
    .io_perf_26_value(dcache_io_perf_26_value)
  );
  Uncache uncache ( // @[MemBlock.scala 48:27]
    .clock(uncache_clock),
    .reset(uncache_reset),
    .auto_client_out_a_ready(uncache_auto_client_out_a_ready),
    .auto_client_out_a_valid(uncache_auto_client_out_a_valid),
    .auto_client_out_a_bits_opcode(uncache_auto_client_out_a_bits_opcode),
    .auto_client_out_a_bits_size(uncache_auto_client_out_a_bits_size),
    .auto_client_out_a_bits_source(uncache_auto_client_out_a_bits_source),
    .auto_client_out_a_bits_address(uncache_auto_client_out_a_bits_address),
    .auto_client_out_a_bits_mask(uncache_auto_client_out_a_bits_mask),
    .auto_client_out_a_bits_data(uncache_auto_client_out_a_bits_data),
    .auto_client_out_d_ready(uncache_auto_client_out_d_ready),
    .auto_client_out_d_valid(uncache_auto_client_out_d_valid),
    .auto_client_out_d_bits_opcode(uncache_auto_client_out_d_bits_opcode),
    .auto_client_out_d_bits_data(uncache_auto_client_out_d_bits_data),
    .io_hartId(uncache_io_hartId),
    .io_enableOutstanding(uncache_io_enableOutstanding),
    .io_flush_empty(uncache_io_flush_empty),
    .io_lsq_req_ready(uncache_io_lsq_req_ready),
    .io_lsq_req_valid(uncache_io_lsq_req_valid),
    .io_lsq_req_bits_cmd(uncache_io_lsq_req_bits_cmd),
    .io_lsq_req_bits_addr(uncache_io_lsq_req_bits_addr),
    .io_lsq_req_bits_data(uncache_io_lsq_req_bits_data),
    .io_lsq_req_bits_mask(uncache_io_lsq_req_bits_mask),
    .io_lsq_req_bits_atomic(uncache_io_lsq_req_bits_atomic),
    .io_lsq_resp_valid(uncache_io_lsq_resp_valid),
    .io_lsq_resp_bits_data(uncache_io_lsq_resp_bits_data)
  );
  DelayN_18 csrCtrl_delay ( // @[Hold.scala 97:23]
    .clock(csrCtrl_delay_clock),
    .io_in_icache_parity_enable(csrCtrl_delay_io_in_icache_parity_enable),
    .io_in_lvpred_disable(csrCtrl_delay_io_in_lvpred_disable),
    .io_in_no_spec_load(csrCtrl_delay_io_in_no_spec_load),
    .io_in_storeset_wait_store(csrCtrl_delay_io_in_storeset_wait_store),
    .io_in_lvpred_timeout(csrCtrl_delay_io_in_lvpred_timeout),
    .io_in_bp_ctrl_ubtb_enable(csrCtrl_delay_io_in_bp_ctrl_ubtb_enable),
    .io_in_bp_ctrl_btb_enable(csrCtrl_delay_io_in_bp_ctrl_btb_enable),
    .io_in_bp_ctrl_tage_enable(csrCtrl_delay_io_in_bp_ctrl_tage_enable),
    .io_in_bp_ctrl_sc_enable(csrCtrl_delay_io_in_bp_ctrl_sc_enable),
    .io_in_bp_ctrl_ras_enable(csrCtrl_delay_io_in_bp_ctrl_ras_enable),
    .io_in_sbuffer_threshold(csrCtrl_delay_io_in_sbuffer_threshold),
    .io_in_ldld_vio_check_enable(csrCtrl_delay_io_in_ldld_vio_check_enable),
    .io_in_cache_error_enable(csrCtrl_delay_io_in_cache_error_enable),
    .io_in_uncache_write_outstanding_enable(csrCtrl_delay_io_in_uncache_write_outstanding_enable),
    .io_in_fusion_enable(csrCtrl_delay_io_in_fusion_enable),
    .io_in_wfi_enable(csrCtrl_delay_io_in_wfi_enable),
    .io_in_svinval_enable(csrCtrl_delay_io_in_svinval_enable),
    .io_in_distribute_csr_wvalid(csrCtrl_delay_io_in_distribute_csr_wvalid),
    .io_in_distribute_csr_waddr(csrCtrl_delay_io_in_distribute_csr_waddr),
    .io_in_distribute_csr_wdata(csrCtrl_delay_io_in_distribute_csr_wdata),
    .io_in_singlestep(csrCtrl_delay_io_in_singlestep),
    .io_in_frontend_trigger_t_valid(csrCtrl_delay_io_in_frontend_trigger_t_valid),
    .io_in_frontend_trigger_t_bits_addr(csrCtrl_delay_io_in_frontend_trigger_t_bits_addr),
    .io_in_frontend_trigger_t_bits_tdata_matchType(csrCtrl_delay_io_in_frontend_trigger_t_bits_tdata_matchType),
    .io_in_frontend_trigger_t_bits_tdata_select(csrCtrl_delay_io_in_frontend_trigger_t_bits_tdata_select),
    .io_in_frontend_trigger_t_bits_tdata_timing(csrCtrl_delay_io_in_frontend_trigger_t_bits_tdata_timing),
    .io_in_frontend_trigger_t_bits_tdata_chain(csrCtrl_delay_io_in_frontend_trigger_t_bits_tdata_chain),
    .io_in_frontend_trigger_t_bits_tdata_tdata2(csrCtrl_delay_io_in_frontend_trigger_t_bits_tdata_tdata2),
    .io_in_mem_trigger_t_valid(csrCtrl_delay_io_in_mem_trigger_t_valid),
    .io_in_mem_trigger_t_bits_addr(csrCtrl_delay_io_in_mem_trigger_t_bits_addr),
    .io_in_mem_trigger_t_bits_tdata_matchType(csrCtrl_delay_io_in_mem_trigger_t_bits_tdata_matchType),
    .io_in_mem_trigger_t_bits_tdata_select(csrCtrl_delay_io_in_mem_trigger_t_bits_tdata_select),
    .io_in_mem_trigger_t_bits_tdata_chain(csrCtrl_delay_io_in_mem_trigger_t_bits_tdata_chain),
    .io_in_mem_trigger_t_bits_tdata_tdata2(csrCtrl_delay_io_in_mem_trigger_t_bits_tdata_tdata2),
    .io_in_trigger_enable_0(csrCtrl_delay_io_in_trigger_enable_0),
    .io_in_trigger_enable_1(csrCtrl_delay_io_in_trigger_enable_1),
    .io_in_trigger_enable_2(csrCtrl_delay_io_in_trigger_enable_2),
    .io_in_trigger_enable_3(csrCtrl_delay_io_in_trigger_enable_3),
    .io_in_trigger_enable_4(csrCtrl_delay_io_in_trigger_enable_4),
    .io_in_trigger_enable_5(csrCtrl_delay_io_in_trigger_enable_5),
    .io_in_trigger_enable_6(csrCtrl_delay_io_in_trigger_enable_6),
    .io_in_trigger_enable_7(csrCtrl_delay_io_in_trigger_enable_7),
    .io_in_trigger_enable_8(csrCtrl_delay_io_in_trigger_enable_8),
    .io_in_trigger_enable_9(csrCtrl_delay_io_in_trigger_enable_9),
    .io_out_icache_parity_enable(csrCtrl_delay_io_out_icache_parity_enable),
    .io_out_lvpred_disable(csrCtrl_delay_io_out_lvpred_disable),
    .io_out_no_spec_load(csrCtrl_delay_io_out_no_spec_load),
    .io_out_storeset_wait_store(csrCtrl_delay_io_out_storeset_wait_store),
    .io_out_lvpred_timeout(csrCtrl_delay_io_out_lvpred_timeout),
    .io_out_bp_ctrl_ubtb_enable(csrCtrl_delay_io_out_bp_ctrl_ubtb_enable),
    .io_out_bp_ctrl_btb_enable(csrCtrl_delay_io_out_bp_ctrl_btb_enable),
    .io_out_bp_ctrl_tage_enable(csrCtrl_delay_io_out_bp_ctrl_tage_enable),
    .io_out_bp_ctrl_sc_enable(csrCtrl_delay_io_out_bp_ctrl_sc_enable),
    .io_out_bp_ctrl_ras_enable(csrCtrl_delay_io_out_bp_ctrl_ras_enable),
    .io_out_sbuffer_threshold(csrCtrl_delay_io_out_sbuffer_threshold),
    .io_out_ldld_vio_check_enable(csrCtrl_delay_io_out_ldld_vio_check_enable),
    .io_out_cache_error_enable(csrCtrl_delay_io_out_cache_error_enable),
    .io_out_uncache_write_outstanding_enable(csrCtrl_delay_io_out_uncache_write_outstanding_enable),
    .io_out_fusion_enable(csrCtrl_delay_io_out_fusion_enable),
    .io_out_wfi_enable(csrCtrl_delay_io_out_wfi_enable),
    .io_out_svinval_enable(csrCtrl_delay_io_out_svinval_enable),
    .io_out_distribute_csr_wvalid(csrCtrl_delay_io_out_distribute_csr_wvalid),
    .io_out_distribute_csr_waddr(csrCtrl_delay_io_out_distribute_csr_waddr),
    .io_out_distribute_csr_wdata(csrCtrl_delay_io_out_distribute_csr_wdata),
    .io_out_singlestep(csrCtrl_delay_io_out_singlestep),
    .io_out_frontend_trigger_t_valid(csrCtrl_delay_io_out_frontend_trigger_t_valid),
    .io_out_frontend_trigger_t_bits_addr(csrCtrl_delay_io_out_frontend_trigger_t_bits_addr),
    .io_out_frontend_trigger_t_bits_tdata_matchType(csrCtrl_delay_io_out_frontend_trigger_t_bits_tdata_matchType),
    .io_out_frontend_trigger_t_bits_tdata_select(csrCtrl_delay_io_out_frontend_trigger_t_bits_tdata_select),
    .io_out_frontend_trigger_t_bits_tdata_timing(csrCtrl_delay_io_out_frontend_trigger_t_bits_tdata_timing),
    .io_out_frontend_trigger_t_bits_tdata_chain(csrCtrl_delay_io_out_frontend_trigger_t_bits_tdata_chain),
    .io_out_frontend_trigger_t_bits_tdata_tdata2(csrCtrl_delay_io_out_frontend_trigger_t_bits_tdata_tdata2),
    .io_out_mem_trigger_t_valid(csrCtrl_delay_io_out_mem_trigger_t_valid),
    .io_out_mem_trigger_t_bits_addr(csrCtrl_delay_io_out_mem_trigger_t_bits_addr),
    .io_out_mem_trigger_t_bits_tdata_matchType(csrCtrl_delay_io_out_mem_trigger_t_bits_tdata_matchType),
    .io_out_mem_trigger_t_bits_tdata_select(csrCtrl_delay_io_out_mem_trigger_t_bits_tdata_select),
    .io_out_mem_trigger_t_bits_tdata_chain(csrCtrl_delay_io_out_mem_trigger_t_bits_tdata_chain),
    .io_out_mem_trigger_t_bits_tdata_tdata2(csrCtrl_delay_io_out_mem_trigger_t_bits_tdata_tdata2),
    .io_out_trigger_enable_0(csrCtrl_delay_io_out_trigger_enable_0),
    .io_out_trigger_enable_1(csrCtrl_delay_io_out_trigger_enable_1),
    .io_out_trigger_enable_2(csrCtrl_delay_io_out_trigger_enable_2),
    .io_out_trigger_enable_3(csrCtrl_delay_io_out_trigger_enable_3),
    .io_out_trigger_enable_4(csrCtrl_delay_io_out_trigger_enable_4),
    .io_out_trigger_enable_5(csrCtrl_delay_io_out_trigger_enable_5),
    .io_out_trigger_enable_6(csrCtrl_delay_io_out_trigger_enable_6),
    .io_out_trigger_enable_7(csrCtrl_delay_io_out_trigger_enable_7),
    .io_out_trigger_enable_8(csrCtrl_delay_io_out_trigger_enable_8),
    .io_out_trigger_enable_9(csrCtrl_delay_io_out_trigger_enable_9)
  );
  LoadUnit LoadUnit_0 ( // @[MemBlock.scala 139:56]
    .clock(LoadUnit_0_clock),
    .reset(LoadUnit_0_reset),
    .io_loadIn_ready(LoadUnit_0_io_loadIn_ready),
    .io_loadIn_valid(LoadUnit_0_io_loadIn_valid),
    .io_loadIn_bits_uop_cf_foldpc(LoadUnit_0_io_loadIn_bits_uop_cf_foldpc),
    .io_loadIn_bits_uop_cf_trigger_backendEn_1(LoadUnit_0_io_loadIn_bits_uop_cf_trigger_backendEn_1),
    .io_loadIn_bits_uop_cf_waitForRobIdx_flag(LoadUnit_0_io_loadIn_bits_uop_cf_waitForRobIdx_flag),
    .io_loadIn_bits_uop_cf_waitForRobIdx_value(LoadUnit_0_io_loadIn_bits_uop_cf_waitForRobIdx_value),
    .io_loadIn_bits_uop_cf_loadWaitBit(LoadUnit_0_io_loadIn_bits_uop_cf_loadWaitBit),
    .io_loadIn_bits_uop_cf_loadWaitStrict(LoadUnit_0_io_loadIn_bits_uop_cf_loadWaitStrict),
    .io_loadIn_bits_uop_cf_ftqPtr_flag(LoadUnit_0_io_loadIn_bits_uop_cf_ftqPtr_flag),
    .io_loadIn_bits_uop_cf_ftqPtr_value(LoadUnit_0_io_loadIn_bits_uop_cf_ftqPtr_value),
    .io_loadIn_bits_uop_cf_ftqOffset(LoadUnit_0_io_loadIn_bits_uop_cf_ftqOffset),
    .io_loadIn_bits_uop_ctrl_fuType(LoadUnit_0_io_loadIn_bits_uop_ctrl_fuType),
    .io_loadIn_bits_uop_ctrl_fuOpType(LoadUnit_0_io_loadIn_bits_uop_ctrl_fuOpType),
    .io_loadIn_bits_uop_ctrl_rfWen(LoadUnit_0_io_loadIn_bits_uop_ctrl_rfWen),
    .io_loadIn_bits_uop_ctrl_fpWen(LoadUnit_0_io_loadIn_bits_uop_ctrl_fpWen),
    .io_loadIn_bits_uop_ctrl_imm(LoadUnit_0_io_loadIn_bits_uop_ctrl_imm),
    .io_loadIn_bits_uop_pdest(LoadUnit_0_io_loadIn_bits_uop_pdest),
    .io_loadIn_bits_uop_robIdx_flag(LoadUnit_0_io_loadIn_bits_uop_robIdx_flag),
    .io_loadIn_bits_uop_robIdx_value(LoadUnit_0_io_loadIn_bits_uop_robIdx_value),
    .io_loadIn_bits_uop_lqIdx_flag(LoadUnit_0_io_loadIn_bits_uop_lqIdx_flag),
    .io_loadIn_bits_uop_lqIdx_value(LoadUnit_0_io_loadIn_bits_uop_lqIdx_value),
    .io_loadIn_bits_uop_sqIdx_flag(LoadUnit_0_io_loadIn_bits_uop_sqIdx_flag),
    .io_loadIn_bits_uop_sqIdx_value(LoadUnit_0_io_loadIn_bits_uop_sqIdx_value),
    .io_loadIn_bits_src_0(LoadUnit_0_io_loadIn_bits_src_0),
    .io_VecloadIn_ready(LoadUnit_0_io_VecloadIn_ready),
    .io_VecloadIn_valid(LoadUnit_0_io_VecloadIn_valid),
    .io_VecloadIn_bits_vaddr(LoadUnit_0_io_VecloadIn_bits_vaddr),
    .io_loadOut_valid(LoadUnit_0_io_loadOut_valid),
    .io_loadOut_bits_uop_cf_exceptionVec_4(LoadUnit_0_io_loadOut_bits_uop_cf_exceptionVec_4),
    .io_loadOut_bits_uop_cf_exceptionVec_5(LoadUnit_0_io_loadOut_bits_uop_cf_exceptionVec_5),
    .io_loadOut_bits_uop_cf_exceptionVec_13(LoadUnit_0_io_loadOut_bits_uop_cf_exceptionVec_13),
    .io_loadOut_bits_uop_cf_trigger_backendEn_1(LoadUnit_0_io_loadOut_bits_uop_cf_trigger_backendEn_1),
    .io_loadOut_bits_uop_cf_trigger_backendHit_0(LoadUnit_0_io_loadOut_bits_uop_cf_trigger_backendHit_0),
    .io_loadOut_bits_uop_cf_trigger_backendHit_1(LoadUnit_0_io_loadOut_bits_uop_cf_trigger_backendHit_1),
    .io_loadOut_bits_uop_cf_trigger_backendHit_4(LoadUnit_0_io_loadOut_bits_uop_cf_trigger_backendHit_4),
    .io_loadOut_bits_uop_ctrl_rfWen(LoadUnit_0_io_loadOut_bits_uop_ctrl_rfWen),
    .io_loadOut_bits_uop_ctrl_fpWen(LoadUnit_0_io_loadOut_bits_uop_ctrl_fpWen),
    .io_loadOut_bits_uop_ctrl_flushPipe(LoadUnit_0_io_loadOut_bits_uop_ctrl_flushPipe),
    .io_loadOut_bits_uop_ctrl_replayInst(LoadUnit_0_io_loadOut_bits_uop_ctrl_replayInst),
    .io_loadOut_bits_uop_pdest(LoadUnit_0_io_loadOut_bits_uop_pdest),
    .io_loadOut_bits_uop_robIdx_flag(LoadUnit_0_io_loadOut_bits_uop_robIdx_flag),
    .io_loadOut_bits_uop_robIdx_value(LoadUnit_0_io_loadOut_bits_uop_robIdx_value),
    .io_loadOut_bits_data(LoadUnit_0_io_loadOut_bits_data),
    .io_loadOut_bits_debug_isMMIO(LoadUnit_0_io_loadOut_bits_debug_isMMIO),
    .io_redirect_valid(LoadUnit_0_io_redirect_valid),
    .io_redirect_bits_robIdx_flag(LoadUnit_0_io_redirect_bits_robIdx_flag),
    .io_redirect_bits_robIdx_value(LoadUnit_0_io_redirect_bits_robIdx_value),
    .io_redirect_bits_level(LoadUnit_0_io_redirect_bits_level),
    .io_dcache_req_ready(LoadUnit_0_io_dcache_req_ready),
    .io_dcache_req_valid(LoadUnit_0_io_dcache_req_valid),
    .io_dcache_req_bits_cmd(LoadUnit_0_io_dcache_req_bits_cmd),
    .io_dcache_req_bits_addr(LoadUnit_0_io_dcache_req_bits_addr),
    .io_dcache_req_bits_instrtype(LoadUnit_0_io_dcache_req_bits_instrtype),
    .io_dcache_req_bits_replayCarry_real_way_en(LoadUnit_0_io_dcache_req_bits_replayCarry_real_way_en),
    .io_dcache_req_bits_replayCarry_valid(LoadUnit_0_io_dcache_req_bits_replayCarry_valid),
    .io_dcache_resp_bits_data_delayed(LoadUnit_0_io_dcache_resp_bits_data_delayed),
    .io_dcache_resp_bits_miss(LoadUnit_0_io_dcache_resp_bits_miss),
    .io_dcache_resp_bits_replay(LoadUnit_0_io_dcache_resp_bits_replay),
    .io_dcache_resp_bits_replayCarry_real_way_en(LoadUnit_0_io_dcache_resp_bits_replayCarry_real_way_en),
    .io_dcache_resp_bits_replayCarry_valid(LoadUnit_0_io_dcache_resp_bits_replayCarry_valid),
    .io_dcache_resp_bits_tag_error(LoadUnit_0_io_dcache_resp_bits_tag_error),
    .io_dcache_resp_bits_mshr_id(LoadUnit_0_io_dcache_resp_bits_mshr_id),
    .io_dcache_resp_bits_error_delayed(LoadUnit_0_io_dcache_resp_bits_error_delayed),
    .io_dcache_s1_kill(LoadUnit_0_io_dcache_s1_kill),
    .io_dcache_s2_kill(LoadUnit_0_io_dcache_s2_kill),
    .io_dcache_s1_paddr_dup_lsu(LoadUnit_0_io_dcache_s1_paddr_dup_lsu),
    .io_dcache_s1_paddr_dup_dcache(LoadUnit_0_io_dcache_s1_paddr_dup_dcache),
    .io_dcache_s1_bank_conflict(LoadUnit_0_io_dcache_s1_bank_conflict),
    .io_sbuffer_vaddr(LoadUnit_0_io_sbuffer_vaddr),
    .io_sbuffer_paddr(LoadUnit_0_io_sbuffer_paddr),
    .io_sbuffer_valid(LoadUnit_0_io_sbuffer_valid),
    .io_sbuffer_forwardMask_0(LoadUnit_0_io_sbuffer_forwardMask_0),
    .io_sbuffer_forwardMask_1(LoadUnit_0_io_sbuffer_forwardMask_1),
    .io_sbuffer_forwardMask_2(LoadUnit_0_io_sbuffer_forwardMask_2),
    .io_sbuffer_forwardMask_3(LoadUnit_0_io_sbuffer_forwardMask_3),
    .io_sbuffer_forwardMask_4(LoadUnit_0_io_sbuffer_forwardMask_4),
    .io_sbuffer_forwardMask_5(LoadUnit_0_io_sbuffer_forwardMask_5),
    .io_sbuffer_forwardMask_6(LoadUnit_0_io_sbuffer_forwardMask_6),
    .io_sbuffer_forwardMask_7(LoadUnit_0_io_sbuffer_forwardMask_7),
    .io_sbuffer_forwardMask_8(LoadUnit_0_io_sbuffer_forwardMask_8),
    .io_sbuffer_forwardMask_9(LoadUnit_0_io_sbuffer_forwardMask_9),
    .io_sbuffer_forwardMask_10(LoadUnit_0_io_sbuffer_forwardMask_10),
    .io_sbuffer_forwardMask_11(LoadUnit_0_io_sbuffer_forwardMask_11),
    .io_sbuffer_forwardMask_12(LoadUnit_0_io_sbuffer_forwardMask_12),
    .io_sbuffer_forwardMask_13(LoadUnit_0_io_sbuffer_forwardMask_13),
    .io_sbuffer_forwardMask_14(LoadUnit_0_io_sbuffer_forwardMask_14),
    .io_sbuffer_forwardMask_15(LoadUnit_0_io_sbuffer_forwardMask_15),
    .io_sbuffer_forwardData_0(LoadUnit_0_io_sbuffer_forwardData_0),
    .io_sbuffer_forwardData_1(LoadUnit_0_io_sbuffer_forwardData_1),
    .io_sbuffer_forwardData_2(LoadUnit_0_io_sbuffer_forwardData_2),
    .io_sbuffer_forwardData_3(LoadUnit_0_io_sbuffer_forwardData_3),
    .io_sbuffer_forwardData_4(LoadUnit_0_io_sbuffer_forwardData_4),
    .io_sbuffer_forwardData_5(LoadUnit_0_io_sbuffer_forwardData_5),
    .io_sbuffer_forwardData_6(LoadUnit_0_io_sbuffer_forwardData_6),
    .io_sbuffer_forwardData_7(LoadUnit_0_io_sbuffer_forwardData_7),
    .io_sbuffer_forwardData_8(LoadUnit_0_io_sbuffer_forwardData_8),
    .io_sbuffer_forwardData_9(LoadUnit_0_io_sbuffer_forwardData_9),
    .io_sbuffer_forwardData_10(LoadUnit_0_io_sbuffer_forwardData_10),
    .io_sbuffer_forwardData_11(LoadUnit_0_io_sbuffer_forwardData_11),
    .io_sbuffer_forwardData_12(LoadUnit_0_io_sbuffer_forwardData_12),
    .io_sbuffer_forwardData_13(LoadUnit_0_io_sbuffer_forwardData_13),
    .io_sbuffer_forwardData_14(LoadUnit_0_io_sbuffer_forwardData_14),
    .io_sbuffer_forwardData_15(LoadUnit_0_io_sbuffer_forwardData_15),
    .io_sbuffer_matchInvalid(LoadUnit_0_io_sbuffer_matchInvalid),
    .io_lsq_loadIn_valid(LoadUnit_0_io_lsq_loadIn_valid),
    .io_lsq_loadIn_bits_uop_cf_foldpc(LoadUnit_0_io_lsq_loadIn_bits_uop_cf_foldpc),
    .io_lsq_loadIn_bits_uop_cf_exceptionVec_4(LoadUnit_0_io_lsq_loadIn_bits_uop_cf_exceptionVec_4),
    .io_lsq_loadIn_bits_uop_cf_exceptionVec_5(LoadUnit_0_io_lsq_loadIn_bits_uop_cf_exceptionVec_5),
    .io_lsq_loadIn_bits_uop_cf_exceptionVec_13(LoadUnit_0_io_lsq_loadIn_bits_uop_cf_exceptionVec_13),
    .io_lsq_loadIn_bits_uop_cf_trigger_backendEn_1(LoadUnit_0_io_lsq_loadIn_bits_uop_cf_trigger_backendEn_1),
    .io_lsq_loadIn_bits_uop_cf_trigger_backendHit_0(LoadUnit_0_io_lsq_loadIn_bits_uop_cf_trigger_backendHit_0),
    .io_lsq_loadIn_bits_uop_cf_trigger_backendHit_1(LoadUnit_0_io_lsq_loadIn_bits_uop_cf_trigger_backendHit_1),
    .io_lsq_loadIn_bits_uop_cf_trigger_backendHit_4(LoadUnit_0_io_lsq_loadIn_bits_uop_cf_trigger_backendHit_4),
    .io_lsq_loadIn_bits_uop_cf_waitForRobIdx_flag(LoadUnit_0_io_lsq_loadIn_bits_uop_cf_waitForRobIdx_flag),
    .io_lsq_loadIn_bits_uop_cf_waitForRobIdx_value(LoadUnit_0_io_lsq_loadIn_bits_uop_cf_waitForRobIdx_value),
    .io_lsq_loadIn_bits_uop_cf_loadWaitBit(LoadUnit_0_io_lsq_loadIn_bits_uop_cf_loadWaitBit),
    .io_lsq_loadIn_bits_uop_cf_loadWaitStrict(LoadUnit_0_io_lsq_loadIn_bits_uop_cf_loadWaitStrict),
    .io_lsq_loadIn_bits_uop_cf_ftqPtr_flag(LoadUnit_0_io_lsq_loadIn_bits_uop_cf_ftqPtr_flag),
    .io_lsq_loadIn_bits_uop_cf_ftqPtr_value(LoadUnit_0_io_lsq_loadIn_bits_uop_cf_ftqPtr_value),
    .io_lsq_loadIn_bits_uop_cf_ftqOffset(LoadUnit_0_io_lsq_loadIn_bits_uop_cf_ftqOffset),
    .io_lsq_loadIn_bits_uop_ctrl_fuType(LoadUnit_0_io_lsq_loadIn_bits_uop_ctrl_fuType),
    .io_lsq_loadIn_bits_uop_ctrl_fuOpType(LoadUnit_0_io_lsq_loadIn_bits_uop_ctrl_fuOpType),
    .io_lsq_loadIn_bits_uop_ctrl_rfWen(LoadUnit_0_io_lsq_loadIn_bits_uop_ctrl_rfWen),
    .io_lsq_loadIn_bits_uop_ctrl_fpWen(LoadUnit_0_io_lsq_loadIn_bits_uop_ctrl_fpWen),
    .io_lsq_loadIn_bits_uop_ctrl_replayInst(LoadUnit_0_io_lsq_loadIn_bits_uop_ctrl_replayInst),
    .io_lsq_loadIn_bits_uop_pdest(LoadUnit_0_io_lsq_loadIn_bits_uop_pdest),
    .io_lsq_loadIn_bits_uop_robIdx_flag(LoadUnit_0_io_lsq_loadIn_bits_uop_robIdx_flag),
    .io_lsq_loadIn_bits_uop_robIdx_value(LoadUnit_0_io_lsq_loadIn_bits_uop_robIdx_value),
    .io_lsq_loadIn_bits_uop_lqIdx_flag(LoadUnit_0_io_lsq_loadIn_bits_uop_lqIdx_flag),
    .io_lsq_loadIn_bits_uop_lqIdx_value(LoadUnit_0_io_lsq_loadIn_bits_uop_lqIdx_value),
    .io_lsq_loadIn_bits_uop_sqIdx_flag(LoadUnit_0_io_lsq_loadIn_bits_uop_sqIdx_flag),
    .io_lsq_loadIn_bits_uop_sqIdx_value(LoadUnit_0_io_lsq_loadIn_bits_uop_sqIdx_value),
    .io_lsq_loadIn_bits_vaddr(LoadUnit_0_io_lsq_loadIn_bits_vaddr),
    .io_lsq_loadIn_bits_paddr(LoadUnit_0_io_lsq_loadIn_bits_paddr),
    .io_lsq_loadIn_bits_mask(LoadUnit_0_io_lsq_loadIn_bits_mask),
    .io_lsq_loadIn_bits_miss(LoadUnit_0_io_lsq_loadIn_bits_miss),
    .io_lsq_loadIn_bits_tlbMiss(LoadUnit_0_io_lsq_loadIn_bits_tlbMiss),
    .io_lsq_loadIn_bits_mmio(LoadUnit_0_io_lsq_loadIn_bits_mmio),
    .io_lsq_loadIn_bits_rarAllocated(LoadUnit_0_io_lsq_loadIn_bits_rarAllocated),
    .io_lsq_loadIn_bits_rarIndex(LoadUnit_0_io_lsq_loadIn_bits_rarIndex),
    .io_lsq_loadIn_bits_rawAllocated(LoadUnit_0_io_lsq_loadIn_bits_rawAllocated),
    .io_lsq_loadIn_bits_rawIndex(LoadUnit_0_io_lsq_loadIn_bits_rawIndex),
    .io_lsq_loadIn_bits_canAccept(LoadUnit_0_io_lsq_loadIn_bits_canAccept),
    .io_lsq_loadIn_bits_replayInfo_missMSHRId(LoadUnit_0_io_lsq_loadIn_bits_replayInfo_missMSHRId),
    .io_lsq_loadIn_bits_replayInfo_canForwardFullData(LoadUnit_0_io_lsq_loadIn_bits_replayInfo_canForwardFullData),
    .io_lsq_loadIn_bits_replayInfo_dataInvalidSqIdx_flag(LoadUnit_0_io_lsq_loadIn_bits_replayInfo_dataInvalidSqIdx_flag)
      ,
    .io_lsq_loadIn_bits_replayInfo_dataInvalidSqIdx_value(
      LoadUnit_0_io_lsq_loadIn_bits_replayInfo_dataInvalidSqIdx_value),
    .io_lsq_loadIn_bits_replayInfo_addrInvalidSqIdx_flag(LoadUnit_0_io_lsq_loadIn_bits_replayInfo_addrInvalidSqIdx_flag)
      ,
    .io_lsq_loadIn_bits_replayInfo_addrInvalidSqIdx_value(
      LoadUnit_0_io_lsq_loadIn_bits_replayInfo_addrInvalidSqIdx_value),
    .io_lsq_loadIn_bits_replayInfo_replayCarry_real_way_en(
      LoadUnit_0_io_lsq_loadIn_bits_replayInfo_replayCarry_real_way_en),
    .io_lsq_loadIn_bits_replayInfo_replayCarry_valid(LoadUnit_0_io_lsq_loadIn_bits_replayInfo_replayCarry_valid),
    .io_lsq_loadIn_bits_replayInfo_dataInLastBeat(LoadUnit_0_io_lsq_loadIn_bits_replayInfo_dataInLastBeat),
    .io_lsq_loadIn_bits_replayInfo_cause_0(LoadUnit_0_io_lsq_loadIn_bits_replayInfo_cause_0),
    .io_lsq_loadIn_bits_replayInfo_cause_1(LoadUnit_0_io_lsq_loadIn_bits_replayInfo_cause_1),
    .io_lsq_loadIn_bits_replayInfo_cause_2(LoadUnit_0_io_lsq_loadIn_bits_replayInfo_cause_2),
    .io_lsq_loadIn_bits_replayInfo_cause_3(LoadUnit_0_io_lsq_loadIn_bits_replayInfo_cause_3),
    .io_lsq_loadIn_bits_replayInfo_cause_4(LoadUnit_0_io_lsq_loadIn_bits_replayInfo_cause_4),
    .io_lsq_loadIn_bits_replayInfo_cause_5(LoadUnit_0_io_lsq_loadIn_bits_replayInfo_cause_5),
    .io_lsq_loadIn_bits_replayInfo_cause_6(LoadUnit_0_io_lsq_loadIn_bits_replayInfo_cause_6),
    .io_lsq_loadIn_bits_replayInfo_cause_7(LoadUnit_0_io_lsq_loadIn_bits_replayInfo_cause_7),
    .io_lsq_loadIn_bits_lqDataWenDup_1(LoadUnit_0_io_lsq_loadIn_bits_lqDataWenDup_1),
    .io_lsq_loadIn_bits_lqDataWenDup_2(LoadUnit_0_io_lsq_loadIn_bits_lqDataWenDup_2),
    .io_lsq_loadIn_bits_lqDataWenDup_3(LoadUnit_0_io_lsq_loadIn_bits_lqDataWenDup_3),
    .io_lsq_loadIn_bits_lqDataWenDup_5(LoadUnit_0_io_lsq_loadIn_bits_lqDataWenDup_5),
    .io_lsq_loadOut_ready(LoadUnit_0_io_lsq_loadOut_ready),
    .io_lsq_loadOut_valid(LoadUnit_0_io_lsq_loadOut_valid),
    .io_lsq_loadOut_bits_uop_cf_exceptionVec_4(LoadUnit_0_io_lsq_loadOut_bits_uop_cf_exceptionVec_4),
    .io_lsq_loadOut_bits_uop_cf_exceptionVec_5(LoadUnit_0_io_lsq_loadOut_bits_uop_cf_exceptionVec_5),
    .io_lsq_loadOut_bits_uop_cf_exceptionVec_13(LoadUnit_0_io_lsq_loadOut_bits_uop_cf_exceptionVec_13),
    .io_lsq_loadOut_bits_uop_cf_trigger_backendEn_1(LoadUnit_0_io_lsq_loadOut_bits_uop_cf_trigger_backendEn_1),
    .io_lsq_loadOut_bits_uop_cf_trigger_backendHit_0(LoadUnit_0_io_lsq_loadOut_bits_uop_cf_trigger_backendHit_0),
    .io_lsq_loadOut_bits_uop_cf_trigger_backendHit_1(LoadUnit_0_io_lsq_loadOut_bits_uop_cf_trigger_backendHit_1),
    .io_lsq_loadOut_bits_uop_cf_trigger_backendHit_4(LoadUnit_0_io_lsq_loadOut_bits_uop_cf_trigger_backendHit_4),
    .io_lsq_loadOut_bits_uop_ctrl_rfWen(LoadUnit_0_io_lsq_loadOut_bits_uop_ctrl_rfWen),
    .io_lsq_loadOut_bits_uop_ctrl_fpWen(LoadUnit_0_io_lsq_loadOut_bits_uop_ctrl_fpWen),
    .io_lsq_loadOut_bits_uop_ctrl_flushPipe(LoadUnit_0_io_lsq_loadOut_bits_uop_ctrl_flushPipe),
    .io_lsq_loadOut_bits_uop_ctrl_replayInst(LoadUnit_0_io_lsq_loadOut_bits_uop_ctrl_replayInst),
    .io_lsq_loadOut_bits_uop_pdest(LoadUnit_0_io_lsq_loadOut_bits_uop_pdest),
    .io_lsq_loadOut_bits_uop_robIdx_flag(LoadUnit_0_io_lsq_loadOut_bits_uop_robIdx_flag),
    .io_lsq_loadOut_bits_uop_robIdx_value(LoadUnit_0_io_lsq_loadOut_bits_uop_robIdx_value),
    .io_lsq_loadOut_bits_debug_isMMIO(LoadUnit_0_io_lsq_loadOut_bits_debug_isMMIO),
    .io_lsq_ldRawData_lqData(LoadUnit_0_io_lsq_ldRawData_lqData),
    .io_lsq_ldRawData_uop_ctrl_fuOpType(LoadUnit_0_io_lsq_ldRawData_uop_ctrl_fuOpType),
    .io_lsq_ldRawData_uop_ctrl_fpWen(LoadUnit_0_io_lsq_ldRawData_uop_ctrl_fpWen),
    .io_lsq_ldRawData_addrOffset(LoadUnit_0_io_lsq_ldRawData_addrOffset),
    .io_lsq_forward_vaddr(LoadUnit_0_io_lsq_forward_vaddr),
    .io_lsq_forward_paddr(LoadUnit_0_io_lsq_forward_paddr),
    .io_lsq_forward_uop_cf_waitForRobIdx_flag(LoadUnit_0_io_lsq_forward_uop_cf_waitForRobIdx_flag),
    .io_lsq_forward_uop_cf_waitForRobIdx_value(LoadUnit_0_io_lsq_forward_uop_cf_waitForRobIdx_value),
    .io_lsq_forward_uop_sqIdx_flag(LoadUnit_0_io_lsq_forward_uop_sqIdx_flag),
    .io_lsq_forward_uop_sqIdx_value(LoadUnit_0_io_lsq_forward_uop_sqIdx_value),
    .io_lsq_forward_valid(LoadUnit_0_io_lsq_forward_valid),
    .io_lsq_forward_forwardMask_0(LoadUnit_0_io_lsq_forward_forwardMask_0),
    .io_lsq_forward_forwardMask_1(LoadUnit_0_io_lsq_forward_forwardMask_1),
    .io_lsq_forward_forwardMask_2(LoadUnit_0_io_lsq_forward_forwardMask_2),
    .io_lsq_forward_forwardMask_3(LoadUnit_0_io_lsq_forward_forwardMask_3),
    .io_lsq_forward_forwardMask_4(LoadUnit_0_io_lsq_forward_forwardMask_4),
    .io_lsq_forward_forwardMask_5(LoadUnit_0_io_lsq_forward_forwardMask_5),
    .io_lsq_forward_forwardMask_6(LoadUnit_0_io_lsq_forward_forwardMask_6),
    .io_lsq_forward_forwardMask_7(LoadUnit_0_io_lsq_forward_forwardMask_7),
    .io_lsq_forward_forwardMask_8(LoadUnit_0_io_lsq_forward_forwardMask_8),
    .io_lsq_forward_forwardMask_9(LoadUnit_0_io_lsq_forward_forwardMask_9),
    .io_lsq_forward_forwardMask_10(LoadUnit_0_io_lsq_forward_forwardMask_10),
    .io_lsq_forward_forwardMask_11(LoadUnit_0_io_lsq_forward_forwardMask_11),
    .io_lsq_forward_forwardMask_12(LoadUnit_0_io_lsq_forward_forwardMask_12),
    .io_lsq_forward_forwardMask_13(LoadUnit_0_io_lsq_forward_forwardMask_13),
    .io_lsq_forward_forwardMask_14(LoadUnit_0_io_lsq_forward_forwardMask_14),
    .io_lsq_forward_forwardMask_15(LoadUnit_0_io_lsq_forward_forwardMask_15),
    .io_lsq_forward_forwardData_0(LoadUnit_0_io_lsq_forward_forwardData_0),
    .io_lsq_forward_forwardData_1(LoadUnit_0_io_lsq_forward_forwardData_1),
    .io_lsq_forward_forwardData_2(LoadUnit_0_io_lsq_forward_forwardData_2),
    .io_lsq_forward_forwardData_3(LoadUnit_0_io_lsq_forward_forwardData_3),
    .io_lsq_forward_forwardData_4(LoadUnit_0_io_lsq_forward_forwardData_4),
    .io_lsq_forward_forwardData_5(LoadUnit_0_io_lsq_forward_forwardData_5),
    .io_lsq_forward_forwardData_6(LoadUnit_0_io_lsq_forward_forwardData_6),
    .io_lsq_forward_forwardData_7(LoadUnit_0_io_lsq_forward_forwardData_7),
    .io_lsq_forward_forwardData_8(LoadUnit_0_io_lsq_forward_forwardData_8),
    .io_lsq_forward_forwardData_9(LoadUnit_0_io_lsq_forward_forwardData_9),
    .io_lsq_forward_forwardData_10(LoadUnit_0_io_lsq_forward_forwardData_10),
    .io_lsq_forward_forwardData_11(LoadUnit_0_io_lsq_forward_forwardData_11),
    .io_lsq_forward_forwardData_12(LoadUnit_0_io_lsq_forward_forwardData_12),
    .io_lsq_forward_forwardData_13(LoadUnit_0_io_lsq_forward_forwardData_13),
    .io_lsq_forward_forwardData_14(LoadUnit_0_io_lsq_forward_forwardData_14),
    .io_lsq_forward_forwardData_15(LoadUnit_0_io_lsq_forward_forwardData_15),
    .io_lsq_forward_sqIdx_flag(LoadUnit_0_io_lsq_forward_sqIdx_flag),
    .io_lsq_forward_dataInvalid(LoadUnit_0_io_lsq_forward_dataInvalid),
    .io_lsq_forward_matchInvalid(LoadUnit_0_io_lsq_forward_matchInvalid),
    .io_lsq_forward_schedWait(LoadUnit_0_io_lsq_forward_schedWait),
    .io_lsq_forward_sqIdxMask(LoadUnit_0_io_lsq_forward_sqIdxMask),
    .io_lsq_forward_dataInvalidSqIdx_flag(LoadUnit_0_io_lsq_forward_dataInvalidSqIdx_flag),
    .io_lsq_forward_dataInvalidSqIdx_value(LoadUnit_0_io_lsq_forward_dataInvalidSqIdx_value),
    .io_lsq_forward_addrInvalidSqIdx_flag(LoadUnit_0_io_lsq_forward_addrInvalidSqIdx_flag),
    .io_lsq_forward_addrInvalidSqIdx_value(LoadUnit_0_io_lsq_forward_addrInvalidSqIdx_value),
    .io_lsq_storeLoadViolationQuery_req_valid(LoadUnit_0_io_lsq_storeLoadViolationQuery_req_valid),
    .io_lsq_storeLoadViolationQuery_req_bits_uop_cf_foldpc(
      LoadUnit_0_io_lsq_storeLoadViolationQuery_req_bits_uop_cf_foldpc),
    .io_lsq_storeLoadViolationQuery_req_bits_uop_cf_ftqPtr_flag(
      LoadUnit_0_io_lsq_storeLoadViolationQuery_req_bits_uop_cf_ftqPtr_flag),
    .io_lsq_storeLoadViolationQuery_req_bits_uop_cf_ftqPtr_value(
      LoadUnit_0_io_lsq_storeLoadViolationQuery_req_bits_uop_cf_ftqPtr_value),
    .io_lsq_storeLoadViolationQuery_req_bits_uop_cf_ftqOffset(
      LoadUnit_0_io_lsq_storeLoadViolationQuery_req_bits_uop_cf_ftqOffset),
    .io_lsq_storeLoadViolationQuery_req_bits_uop_robIdx_flag(
      LoadUnit_0_io_lsq_storeLoadViolationQuery_req_bits_uop_robIdx_flag),
    .io_lsq_storeLoadViolationQuery_req_bits_uop_robIdx_value(
      LoadUnit_0_io_lsq_storeLoadViolationQuery_req_bits_uop_robIdx_value),
    .io_lsq_storeLoadViolationQuery_req_bits_uop_sqIdx_flag(
      LoadUnit_0_io_lsq_storeLoadViolationQuery_req_bits_uop_sqIdx_flag),
    .io_lsq_storeLoadViolationQuery_req_bits_uop_sqIdx_value(
      LoadUnit_0_io_lsq_storeLoadViolationQuery_req_bits_uop_sqIdx_value),
    .io_lsq_storeLoadViolationQuery_req_bits_index(LoadUnit_0_io_lsq_storeLoadViolationQuery_req_bits_index),
    .io_lsq_storeLoadViolationQuery_req_bits_allocated(LoadUnit_0_io_lsq_storeLoadViolationQuery_req_bits_allocated),
    .io_lsq_storeLoadViolationQuery_req_bits_datavalid(LoadUnit_0_io_lsq_storeLoadViolationQuery_req_bits_datavalid),
    .io_lsq_storeLoadViolationQuery_req_bits_mask(LoadUnit_0_io_lsq_storeLoadViolationQuery_req_bits_mask),
    .io_lsq_storeLoadViolationQuery_req_bits_paddr(LoadUnit_0_io_lsq_storeLoadViolationQuery_req_bits_paddr),
    .io_lsq_storeLoadViolationQuery_resp_bits_index(LoadUnit_0_io_lsq_storeLoadViolationQuery_resp_bits_index),
    .io_lsq_storeLoadViolationQuery_resp_bits_canAccept(LoadUnit_0_io_lsq_storeLoadViolationQuery_resp_bits_canAccept),
    .io_lsq_storeLoadViolationQuery_resp_bits_allocated(LoadUnit_0_io_lsq_storeLoadViolationQuery_resp_bits_allocated),
    .io_lsq_loadLoadViolationQuery_req_valid(LoadUnit_0_io_lsq_loadLoadViolationQuery_req_valid),
    .io_lsq_loadLoadViolationQuery_req_bits_uop_robIdx_flag(
      LoadUnit_0_io_lsq_loadLoadViolationQuery_req_bits_uop_robIdx_flag),
    .io_lsq_loadLoadViolationQuery_req_bits_uop_robIdx_value(
      LoadUnit_0_io_lsq_loadLoadViolationQuery_req_bits_uop_robIdx_value),
    .io_lsq_loadLoadViolationQuery_req_bits_uop_lqIdx_flag(
      LoadUnit_0_io_lsq_loadLoadViolationQuery_req_bits_uop_lqIdx_flag),
    .io_lsq_loadLoadViolationQuery_req_bits_uop_lqIdx_value(
      LoadUnit_0_io_lsq_loadLoadViolationQuery_req_bits_uop_lqIdx_value),
    .io_lsq_loadLoadViolationQuery_req_bits_index(LoadUnit_0_io_lsq_loadLoadViolationQuery_req_bits_index),
    .io_lsq_loadLoadViolationQuery_req_bits_allocated(LoadUnit_0_io_lsq_loadLoadViolationQuery_req_bits_allocated),
    .io_lsq_loadLoadViolationQuery_req_bits_datavalid(LoadUnit_0_io_lsq_loadLoadViolationQuery_req_bits_datavalid),
    .io_lsq_loadLoadViolationQuery_req_bits_miss(LoadUnit_0_io_lsq_loadLoadViolationQuery_req_bits_miss),
    .io_lsq_loadLoadViolationQuery_req_bits_paddr(LoadUnit_0_io_lsq_loadLoadViolationQuery_req_bits_paddr),
    .io_lsq_loadLoadViolationQuery_resp_valid(LoadUnit_0_io_lsq_loadLoadViolationQuery_resp_valid),
    .io_lsq_loadLoadViolationQuery_resp_bits_index(LoadUnit_0_io_lsq_loadLoadViolationQuery_resp_bits_index),
    .io_lsq_loadLoadViolationQuery_resp_bits_canAccept(LoadUnit_0_io_lsq_loadLoadViolationQuery_resp_bits_canAccept),
    .io_lsq_loadLoadViolationQuery_resp_bits_allocated(LoadUnit_0_io_lsq_loadLoadViolationQuery_resp_bits_allocated),
    .io_lsq_loadLoadViolationQuery_resp_bits_replayFromFetch(
      LoadUnit_0_io_lsq_loadLoadViolationQuery_resp_bits_replayFromFetch),
    .io_lsq_trigger_hitLoadAddrTriggerHitVec_0(LoadUnit_0_io_lsq_trigger_hitLoadAddrTriggerHitVec_0),
    .io_lsq_trigger_hitLoadAddrTriggerHitVec_1(LoadUnit_0_io_lsq_trigger_hitLoadAddrTriggerHitVec_1),
    .io_lsq_trigger_hitLoadAddrTriggerHitVec_2(LoadUnit_0_io_lsq_trigger_hitLoadAddrTriggerHitVec_2),
    .io_lsq_trigger_lqLoadAddrTriggerHitVec_0(LoadUnit_0_io_lsq_trigger_lqLoadAddrTriggerHitVec_0),
    .io_lsq_trigger_lqLoadAddrTriggerHitVec_1(LoadUnit_0_io_lsq_trigger_lqLoadAddrTriggerHitVec_1),
    .io_lsq_trigger_lqLoadAddrTriggerHitVec_2(LoadUnit_0_io_lsq_trigger_lqLoadAddrTriggerHitVec_2),
    .io_tlDchannel_valid(LoadUnit_0_io_tlDchannel_valid),
    .io_tlDchannel_data(LoadUnit_0_io_tlDchannel_data),
    .io_tlDchannel_mshrid(LoadUnit_0_io_tlDchannel_mshrid),
    .io_tlDchannel_last(LoadUnit_0_io_tlDchannel_last),
    .io_forward_mshr_valid(LoadUnit_0_io_forward_mshr_valid),
    .io_forward_mshr_mshrid(LoadUnit_0_io_forward_mshr_mshrid),
    .io_forward_mshr_paddr(LoadUnit_0_io_forward_mshr_paddr),
    .io_forward_mshr_forward_mshr(LoadUnit_0_io_forward_mshr_forward_mshr),
    .io_forward_mshr_forwardData_0(LoadUnit_0_io_forward_mshr_forwardData_0),
    .io_forward_mshr_forwardData_1(LoadUnit_0_io_forward_mshr_forwardData_1),
    .io_forward_mshr_forwardData_2(LoadUnit_0_io_forward_mshr_forwardData_2),
    .io_forward_mshr_forwardData_3(LoadUnit_0_io_forward_mshr_forwardData_3),
    .io_forward_mshr_forwardData_4(LoadUnit_0_io_forward_mshr_forwardData_4),
    .io_forward_mshr_forwardData_5(LoadUnit_0_io_forward_mshr_forwardData_5),
    .io_forward_mshr_forwardData_6(LoadUnit_0_io_forward_mshr_forwardData_6),
    .io_forward_mshr_forwardData_7(LoadUnit_0_io_forward_mshr_forwardData_7),
    .io_forward_mshr_forwardData_8(LoadUnit_0_io_forward_mshr_forwardData_8),
    .io_forward_mshr_forwardData_9(LoadUnit_0_io_forward_mshr_forwardData_9),
    .io_forward_mshr_forwardData_10(LoadUnit_0_io_forward_mshr_forwardData_10),
    .io_forward_mshr_forwardData_11(LoadUnit_0_io_forward_mshr_forwardData_11),
    .io_forward_mshr_forwardData_12(LoadUnit_0_io_forward_mshr_forwardData_12),
    .io_forward_mshr_forwardData_13(LoadUnit_0_io_forward_mshr_forwardData_13),
    .io_forward_mshr_forwardData_14(LoadUnit_0_io_forward_mshr_forwardData_14),
    .io_forward_mshr_forwardData_15(LoadUnit_0_io_forward_mshr_forwardData_15),
    .io_forward_mshr_forward_result_valid(LoadUnit_0_io_forward_mshr_forward_result_valid),
    .io_trigger_0_tdata2(LoadUnit_0_io_trigger_0_tdata2),
    .io_trigger_0_matchType(LoadUnit_0_io_trigger_0_matchType),
    .io_trigger_0_tEnable(LoadUnit_0_io_trigger_0_tEnable),
    .io_trigger_0_addrHit(LoadUnit_0_io_trigger_0_addrHit),
    .io_trigger_1_tdata2(LoadUnit_0_io_trigger_1_tdata2),
    .io_trigger_1_matchType(LoadUnit_0_io_trigger_1_matchType),
    .io_trigger_1_tEnable(LoadUnit_0_io_trigger_1_tEnable),
    .io_trigger_1_addrHit(LoadUnit_0_io_trigger_1_addrHit),
    .io_trigger_2_tdata2(LoadUnit_0_io_trigger_2_tdata2),
    .io_trigger_2_matchType(LoadUnit_0_io_trigger_2_matchType),
    .io_trigger_2_tEnable(LoadUnit_0_io_trigger_2_tEnable),
    .io_trigger_2_addrHit(LoadUnit_0_io_trigger_2_addrHit),
    .io_tlb_req_valid(LoadUnit_0_io_tlb_req_valid),
    .io_tlb_req_bits_vaddr(LoadUnit_0_io_tlb_req_bits_vaddr),
    .io_tlb_req_bits_cmd(LoadUnit_0_io_tlb_req_bits_cmd),
    .io_tlb_req_bits_no_translate(LoadUnit_0_io_tlb_req_bits_no_translate),
    .io_tlb_req_kill(LoadUnit_0_io_tlb_req_kill),
    .io_tlb_resp_bits_paddr_0(LoadUnit_0_io_tlb_resp_bits_paddr_0),
    .io_tlb_resp_bits_paddr_1(LoadUnit_0_io_tlb_resp_bits_paddr_1),
    .io_tlb_resp_bits_miss(LoadUnit_0_io_tlb_resp_bits_miss),
    .io_tlb_resp_bits_excp_0_pf_ld(LoadUnit_0_io_tlb_resp_bits_excp_0_pf_ld),
    .io_tlb_resp_bits_excp_0_af_ld(LoadUnit_0_io_tlb_resp_bits_excp_0_af_ld),
    .io_tlb_resp_bits_static_pm_valid(LoadUnit_0_io_tlb_resp_bits_static_pm_valid),
    .io_tlb_resp_bits_static_pm_bits(LoadUnit_0_io_tlb_resp_bits_static_pm_bits),
    .io_pmp_ld(LoadUnit_0_io_pmp_ld),
    .io_pmp_mmio(LoadUnit_0_io_pmp_mmio),
    .io_fastpathOut_data(LoadUnit_0_io_fastpathOut_data),
    .io_fastpathOut_valid(LoadUnit_0_io_fastpathOut_valid),
    .io_fastpathIn_data(LoadUnit_0_io_fastpathIn_data),
    .io_fastpathIn_valid(LoadUnit_0_io_fastpathIn_valid),
    .io_loadFastMatch(LoadUnit_0_io_loadFastMatch),
    .io_loadFastImm(LoadUnit_0_io_loadFastImm),
    .io_csrCtrl_ldld_vio_check_enable(LoadUnit_0_io_csrCtrl_ldld_vio_check_enable),
    .io_csrCtrl_cache_error_enable(LoadUnit_0_io_csrCtrl_cache_error_enable),
    .io_correctTableQuery_req_addr(LoadUnit_0_io_correctTableQuery_req_addr),
    .io_correctTableQuery_resp_strict(LoadUnit_0_io_correctTableQuery_resp_strict),
    .io_correctTableUpdate_valid(LoadUnit_0_io_correctTableUpdate_valid),
    .io_correctTableUpdate_bits_addr(LoadUnit_0_io_correctTableUpdate_bits_addr),
    .io_correctTableUpdate_bits_strict(LoadUnit_0_io_correctTableUpdate_bits_strict),
    .io_correctTableUpdate_bits_violation(LoadUnit_0_io_correctTableUpdate_bits_violation),
    .io_reExecuteQuery_0_valid(LoadUnit_0_io_reExecuteQuery_0_valid),
    .io_reExecuteQuery_0_bits_robIdx_flag(LoadUnit_0_io_reExecuteQuery_0_bits_robIdx_flag),
    .io_reExecuteQuery_0_bits_robIdx_value(LoadUnit_0_io_reExecuteQuery_0_bits_robIdx_value),
    .io_reExecuteQuery_0_bits_paddr(LoadUnit_0_io_reExecuteQuery_0_bits_paddr),
    .io_reExecuteQuery_0_bits_mask(LoadUnit_0_io_reExecuteQuery_0_bits_mask),
    .io_reExecuteQuery_1_valid(LoadUnit_0_io_reExecuteQuery_1_valid),
    .io_reExecuteQuery_1_bits_robIdx_flag(LoadUnit_0_io_reExecuteQuery_1_bits_robIdx_flag),
    .io_reExecuteQuery_1_bits_robIdx_value(LoadUnit_0_io_reExecuteQuery_1_bits_robIdx_value),
    .io_reExecuteQuery_1_bits_paddr(LoadUnit_0_io_reExecuteQuery_1_bits_paddr),
    .io_reExecuteQuery_1_bits_mask(LoadUnit_0_io_reExecuteQuery_1_bits_mask),
    .io_replay_ready(LoadUnit_0_io_replay_ready),
    .io_replay_valid(LoadUnit_0_io_replay_valid),
    .io_replay_bits_uop_cf_foldpc(LoadUnit_0_io_replay_bits_uop_cf_foldpc),
    .io_replay_bits_uop_cf_trigger_backendEn_1(LoadUnit_0_io_replay_bits_uop_cf_trigger_backendEn_1),
    .io_replay_bits_uop_cf_trigger_backendHit_0(LoadUnit_0_io_replay_bits_uop_cf_trigger_backendHit_0),
    .io_replay_bits_uop_cf_trigger_backendHit_1(LoadUnit_0_io_replay_bits_uop_cf_trigger_backendHit_1),
    .io_replay_bits_uop_cf_trigger_backendHit_4(LoadUnit_0_io_replay_bits_uop_cf_trigger_backendHit_4),
    .io_replay_bits_uop_cf_waitForRobIdx_flag(LoadUnit_0_io_replay_bits_uop_cf_waitForRobIdx_flag),
    .io_replay_bits_uop_cf_waitForRobIdx_value(LoadUnit_0_io_replay_bits_uop_cf_waitForRobIdx_value),
    .io_replay_bits_uop_cf_loadWaitBit(LoadUnit_0_io_replay_bits_uop_cf_loadWaitBit),
    .io_replay_bits_uop_cf_loadWaitStrict(LoadUnit_0_io_replay_bits_uop_cf_loadWaitStrict),
    .io_replay_bits_uop_cf_ftqPtr_flag(LoadUnit_0_io_replay_bits_uop_cf_ftqPtr_flag),
    .io_replay_bits_uop_cf_ftqPtr_value(LoadUnit_0_io_replay_bits_uop_cf_ftqPtr_value),
    .io_replay_bits_uop_cf_ftqOffset(LoadUnit_0_io_replay_bits_uop_cf_ftqOffset),
    .io_replay_bits_uop_ctrl_fuType(LoadUnit_0_io_replay_bits_uop_ctrl_fuType),
    .io_replay_bits_uop_ctrl_fuOpType(LoadUnit_0_io_replay_bits_uop_ctrl_fuOpType),
    .io_replay_bits_uop_ctrl_rfWen(LoadUnit_0_io_replay_bits_uop_ctrl_rfWen),
    .io_replay_bits_uop_ctrl_fpWen(LoadUnit_0_io_replay_bits_uop_ctrl_fpWen),
    .io_replay_bits_uop_pdest(LoadUnit_0_io_replay_bits_uop_pdest),
    .io_replay_bits_uop_robIdx_flag(LoadUnit_0_io_replay_bits_uop_robIdx_flag),
    .io_replay_bits_uop_robIdx_value(LoadUnit_0_io_replay_bits_uop_robIdx_value),
    .io_replay_bits_uop_lqIdx_flag(LoadUnit_0_io_replay_bits_uop_lqIdx_flag),
    .io_replay_bits_uop_lqIdx_value(LoadUnit_0_io_replay_bits_uop_lqIdx_value),
    .io_replay_bits_uop_sqIdx_flag(LoadUnit_0_io_replay_bits_uop_sqIdx_flag),
    .io_replay_bits_uop_sqIdx_value(LoadUnit_0_io_replay_bits_uop_sqIdx_value),
    .io_replay_bits_vaddr(LoadUnit_0_io_replay_bits_vaddr),
    .io_replay_bits_isFirstIssue(LoadUnit_0_io_replay_bits_isFirstIssue),
    .io_replay_bits_replayCarry_real_way_en(LoadUnit_0_io_replay_bits_replayCarry_real_way_en),
    .io_replay_bits_replayCarry_valid(LoadUnit_0_io_replay_bits_replayCarry_valid),
    .io_replay_bits_mshrid(LoadUnit_0_io_replay_bits_mshrid),
    .io_replay_bits_forward_tlDchannel(LoadUnit_0_io_replay_bits_forward_tlDchannel),
    .io_replay_bits_rarAllocated(LoadUnit_0_io_replay_bits_rarAllocated),
    .io_replay_bits_rarIndex(LoadUnit_0_io_replay_bits_rarIndex),
    .io_replay_bits_rawAllocated(LoadUnit_0_io_replay_bits_rawAllocated),
    .io_replay_bits_rawIndex(LoadUnit_0_io_replay_bits_rawIndex),
    .io_lqReplayFull(LoadUnit_0_io_lqReplayFull),
    .io_perf_0_value(LoadUnit_0_io_perf_0_value),
    .io_perf_1_value(LoadUnit_0_io_perf_1_value),
    .io_perf_2_value(LoadUnit_0_io_perf_2_value),
    .io_perf_3_value(LoadUnit_0_io_perf_3_value),
    .io_perf_4_value(LoadUnit_0_io_perf_4_value),
    .io_perf_5_value(LoadUnit_0_io_perf_5_value),
    .io_perf_6_value(LoadUnit_0_io_perf_6_value)
  );
  LoadUnit LoadUnit_1 ( // @[MemBlock.scala 139:56]
    .clock(LoadUnit_1_clock),
    .reset(LoadUnit_1_reset),
    .io_loadIn_ready(LoadUnit_1_io_loadIn_ready),
    .io_loadIn_valid(LoadUnit_1_io_loadIn_valid),
    .io_loadIn_bits_uop_cf_foldpc(LoadUnit_1_io_loadIn_bits_uop_cf_foldpc),
    .io_loadIn_bits_uop_cf_trigger_backendEn_1(LoadUnit_1_io_loadIn_bits_uop_cf_trigger_backendEn_1),
    .io_loadIn_bits_uop_cf_waitForRobIdx_flag(LoadUnit_1_io_loadIn_bits_uop_cf_waitForRobIdx_flag),
    .io_loadIn_bits_uop_cf_waitForRobIdx_value(LoadUnit_1_io_loadIn_bits_uop_cf_waitForRobIdx_value),
    .io_loadIn_bits_uop_cf_loadWaitBit(LoadUnit_1_io_loadIn_bits_uop_cf_loadWaitBit),
    .io_loadIn_bits_uop_cf_loadWaitStrict(LoadUnit_1_io_loadIn_bits_uop_cf_loadWaitStrict),
    .io_loadIn_bits_uop_cf_ftqPtr_flag(LoadUnit_1_io_loadIn_bits_uop_cf_ftqPtr_flag),
    .io_loadIn_bits_uop_cf_ftqPtr_value(LoadUnit_1_io_loadIn_bits_uop_cf_ftqPtr_value),
    .io_loadIn_bits_uop_cf_ftqOffset(LoadUnit_1_io_loadIn_bits_uop_cf_ftqOffset),
    .io_loadIn_bits_uop_ctrl_fuType(LoadUnit_1_io_loadIn_bits_uop_ctrl_fuType),
    .io_loadIn_bits_uop_ctrl_fuOpType(LoadUnit_1_io_loadIn_bits_uop_ctrl_fuOpType),
    .io_loadIn_bits_uop_ctrl_rfWen(LoadUnit_1_io_loadIn_bits_uop_ctrl_rfWen),
    .io_loadIn_bits_uop_ctrl_fpWen(LoadUnit_1_io_loadIn_bits_uop_ctrl_fpWen),
    .io_loadIn_bits_uop_ctrl_imm(LoadUnit_1_io_loadIn_bits_uop_ctrl_imm),
    .io_loadIn_bits_uop_pdest(LoadUnit_1_io_loadIn_bits_uop_pdest),
    .io_loadIn_bits_uop_robIdx_flag(LoadUnit_1_io_loadIn_bits_uop_robIdx_flag),
    .io_loadIn_bits_uop_robIdx_value(LoadUnit_1_io_loadIn_bits_uop_robIdx_value),
    .io_loadIn_bits_uop_lqIdx_flag(LoadUnit_1_io_loadIn_bits_uop_lqIdx_flag),
    .io_loadIn_bits_uop_lqIdx_value(LoadUnit_1_io_loadIn_bits_uop_lqIdx_value),
    .io_loadIn_bits_uop_sqIdx_flag(LoadUnit_1_io_loadIn_bits_uop_sqIdx_flag),
    .io_loadIn_bits_uop_sqIdx_value(LoadUnit_1_io_loadIn_bits_uop_sqIdx_value),
    .io_loadIn_bits_src_0(LoadUnit_1_io_loadIn_bits_src_0),
    .io_VecloadIn_ready(LoadUnit_1_io_VecloadIn_ready),
    .io_VecloadIn_valid(LoadUnit_1_io_VecloadIn_valid),
    .io_VecloadIn_bits_vaddr(LoadUnit_1_io_VecloadIn_bits_vaddr),
    .io_loadOut_valid(LoadUnit_1_io_loadOut_valid),
    .io_loadOut_bits_uop_cf_exceptionVec_4(LoadUnit_1_io_loadOut_bits_uop_cf_exceptionVec_4),
    .io_loadOut_bits_uop_cf_exceptionVec_5(LoadUnit_1_io_loadOut_bits_uop_cf_exceptionVec_5),
    .io_loadOut_bits_uop_cf_exceptionVec_13(LoadUnit_1_io_loadOut_bits_uop_cf_exceptionVec_13),
    .io_loadOut_bits_uop_cf_trigger_backendEn_1(LoadUnit_1_io_loadOut_bits_uop_cf_trigger_backendEn_1),
    .io_loadOut_bits_uop_cf_trigger_backendHit_0(LoadUnit_1_io_loadOut_bits_uop_cf_trigger_backendHit_0),
    .io_loadOut_bits_uop_cf_trigger_backendHit_1(LoadUnit_1_io_loadOut_bits_uop_cf_trigger_backendHit_1),
    .io_loadOut_bits_uop_cf_trigger_backendHit_4(LoadUnit_1_io_loadOut_bits_uop_cf_trigger_backendHit_4),
    .io_loadOut_bits_uop_ctrl_rfWen(LoadUnit_1_io_loadOut_bits_uop_ctrl_rfWen),
    .io_loadOut_bits_uop_ctrl_fpWen(LoadUnit_1_io_loadOut_bits_uop_ctrl_fpWen),
    .io_loadOut_bits_uop_ctrl_flushPipe(LoadUnit_1_io_loadOut_bits_uop_ctrl_flushPipe),
    .io_loadOut_bits_uop_ctrl_replayInst(LoadUnit_1_io_loadOut_bits_uop_ctrl_replayInst),
    .io_loadOut_bits_uop_pdest(LoadUnit_1_io_loadOut_bits_uop_pdest),
    .io_loadOut_bits_uop_robIdx_flag(LoadUnit_1_io_loadOut_bits_uop_robIdx_flag),
    .io_loadOut_bits_uop_robIdx_value(LoadUnit_1_io_loadOut_bits_uop_robIdx_value),
    .io_loadOut_bits_data(LoadUnit_1_io_loadOut_bits_data),
    .io_loadOut_bits_debug_isMMIO(LoadUnit_1_io_loadOut_bits_debug_isMMIO),
    .io_redirect_valid(LoadUnit_1_io_redirect_valid),
    .io_redirect_bits_robIdx_flag(LoadUnit_1_io_redirect_bits_robIdx_flag),
    .io_redirect_bits_robIdx_value(LoadUnit_1_io_redirect_bits_robIdx_value),
    .io_redirect_bits_level(LoadUnit_1_io_redirect_bits_level),
    .io_dcache_req_ready(LoadUnit_1_io_dcache_req_ready),
    .io_dcache_req_valid(LoadUnit_1_io_dcache_req_valid),
    .io_dcache_req_bits_cmd(LoadUnit_1_io_dcache_req_bits_cmd),
    .io_dcache_req_bits_addr(LoadUnit_1_io_dcache_req_bits_addr),
    .io_dcache_req_bits_instrtype(LoadUnit_1_io_dcache_req_bits_instrtype),
    .io_dcache_req_bits_replayCarry_real_way_en(LoadUnit_1_io_dcache_req_bits_replayCarry_real_way_en),
    .io_dcache_req_bits_replayCarry_valid(LoadUnit_1_io_dcache_req_bits_replayCarry_valid),
    .io_dcache_resp_bits_data_delayed(LoadUnit_1_io_dcache_resp_bits_data_delayed),
    .io_dcache_resp_bits_miss(LoadUnit_1_io_dcache_resp_bits_miss),
    .io_dcache_resp_bits_replay(LoadUnit_1_io_dcache_resp_bits_replay),
    .io_dcache_resp_bits_replayCarry_real_way_en(LoadUnit_1_io_dcache_resp_bits_replayCarry_real_way_en),
    .io_dcache_resp_bits_replayCarry_valid(LoadUnit_1_io_dcache_resp_bits_replayCarry_valid),
    .io_dcache_resp_bits_tag_error(LoadUnit_1_io_dcache_resp_bits_tag_error),
    .io_dcache_resp_bits_mshr_id(LoadUnit_1_io_dcache_resp_bits_mshr_id),
    .io_dcache_resp_bits_error_delayed(LoadUnit_1_io_dcache_resp_bits_error_delayed),
    .io_dcache_s1_kill(LoadUnit_1_io_dcache_s1_kill),
    .io_dcache_s2_kill(LoadUnit_1_io_dcache_s2_kill),
    .io_dcache_s1_paddr_dup_lsu(LoadUnit_1_io_dcache_s1_paddr_dup_lsu),
    .io_dcache_s1_paddr_dup_dcache(LoadUnit_1_io_dcache_s1_paddr_dup_dcache),
    .io_dcache_s1_bank_conflict(LoadUnit_1_io_dcache_s1_bank_conflict),
    .io_sbuffer_vaddr(LoadUnit_1_io_sbuffer_vaddr),
    .io_sbuffer_paddr(LoadUnit_1_io_sbuffer_paddr),
    .io_sbuffer_valid(LoadUnit_1_io_sbuffer_valid),
    .io_sbuffer_forwardMask_0(LoadUnit_1_io_sbuffer_forwardMask_0),
    .io_sbuffer_forwardMask_1(LoadUnit_1_io_sbuffer_forwardMask_1),
    .io_sbuffer_forwardMask_2(LoadUnit_1_io_sbuffer_forwardMask_2),
    .io_sbuffer_forwardMask_3(LoadUnit_1_io_sbuffer_forwardMask_3),
    .io_sbuffer_forwardMask_4(LoadUnit_1_io_sbuffer_forwardMask_4),
    .io_sbuffer_forwardMask_5(LoadUnit_1_io_sbuffer_forwardMask_5),
    .io_sbuffer_forwardMask_6(LoadUnit_1_io_sbuffer_forwardMask_6),
    .io_sbuffer_forwardMask_7(LoadUnit_1_io_sbuffer_forwardMask_7),
    .io_sbuffer_forwardMask_8(LoadUnit_1_io_sbuffer_forwardMask_8),
    .io_sbuffer_forwardMask_9(LoadUnit_1_io_sbuffer_forwardMask_9),
    .io_sbuffer_forwardMask_10(LoadUnit_1_io_sbuffer_forwardMask_10),
    .io_sbuffer_forwardMask_11(LoadUnit_1_io_sbuffer_forwardMask_11),
    .io_sbuffer_forwardMask_12(LoadUnit_1_io_sbuffer_forwardMask_12),
    .io_sbuffer_forwardMask_13(LoadUnit_1_io_sbuffer_forwardMask_13),
    .io_sbuffer_forwardMask_14(LoadUnit_1_io_sbuffer_forwardMask_14),
    .io_sbuffer_forwardMask_15(LoadUnit_1_io_sbuffer_forwardMask_15),
    .io_sbuffer_forwardData_0(LoadUnit_1_io_sbuffer_forwardData_0),
    .io_sbuffer_forwardData_1(LoadUnit_1_io_sbuffer_forwardData_1),
    .io_sbuffer_forwardData_2(LoadUnit_1_io_sbuffer_forwardData_2),
    .io_sbuffer_forwardData_3(LoadUnit_1_io_sbuffer_forwardData_3),
    .io_sbuffer_forwardData_4(LoadUnit_1_io_sbuffer_forwardData_4),
    .io_sbuffer_forwardData_5(LoadUnit_1_io_sbuffer_forwardData_5),
    .io_sbuffer_forwardData_6(LoadUnit_1_io_sbuffer_forwardData_6),
    .io_sbuffer_forwardData_7(LoadUnit_1_io_sbuffer_forwardData_7),
    .io_sbuffer_forwardData_8(LoadUnit_1_io_sbuffer_forwardData_8),
    .io_sbuffer_forwardData_9(LoadUnit_1_io_sbuffer_forwardData_9),
    .io_sbuffer_forwardData_10(LoadUnit_1_io_sbuffer_forwardData_10),
    .io_sbuffer_forwardData_11(LoadUnit_1_io_sbuffer_forwardData_11),
    .io_sbuffer_forwardData_12(LoadUnit_1_io_sbuffer_forwardData_12),
    .io_sbuffer_forwardData_13(LoadUnit_1_io_sbuffer_forwardData_13),
    .io_sbuffer_forwardData_14(LoadUnit_1_io_sbuffer_forwardData_14),
    .io_sbuffer_forwardData_15(LoadUnit_1_io_sbuffer_forwardData_15),
    .io_sbuffer_matchInvalid(LoadUnit_1_io_sbuffer_matchInvalid),
    .io_lsq_loadIn_valid(LoadUnit_1_io_lsq_loadIn_valid),
    .io_lsq_loadIn_bits_uop_cf_foldpc(LoadUnit_1_io_lsq_loadIn_bits_uop_cf_foldpc),
    .io_lsq_loadIn_bits_uop_cf_exceptionVec_4(LoadUnit_1_io_lsq_loadIn_bits_uop_cf_exceptionVec_4),
    .io_lsq_loadIn_bits_uop_cf_exceptionVec_5(LoadUnit_1_io_lsq_loadIn_bits_uop_cf_exceptionVec_5),
    .io_lsq_loadIn_bits_uop_cf_exceptionVec_13(LoadUnit_1_io_lsq_loadIn_bits_uop_cf_exceptionVec_13),
    .io_lsq_loadIn_bits_uop_cf_trigger_backendEn_1(LoadUnit_1_io_lsq_loadIn_bits_uop_cf_trigger_backendEn_1),
    .io_lsq_loadIn_bits_uop_cf_trigger_backendHit_0(LoadUnit_1_io_lsq_loadIn_bits_uop_cf_trigger_backendHit_0),
    .io_lsq_loadIn_bits_uop_cf_trigger_backendHit_1(LoadUnit_1_io_lsq_loadIn_bits_uop_cf_trigger_backendHit_1),
    .io_lsq_loadIn_bits_uop_cf_trigger_backendHit_4(LoadUnit_1_io_lsq_loadIn_bits_uop_cf_trigger_backendHit_4),
    .io_lsq_loadIn_bits_uop_cf_waitForRobIdx_flag(LoadUnit_1_io_lsq_loadIn_bits_uop_cf_waitForRobIdx_flag),
    .io_lsq_loadIn_bits_uop_cf_waitForRobIdx_value(LoadUnit_1_io_lsq_loadIn_bits_uop_cf_waitForRobIdx_value),
    .io_lsq_loadIn_bits_uop_cf_loadWaitBit(LoadUnit_1_io_lsq_loadIn_bits_uop_cf_loadWaitBit),
    .io_lsq_loadIn_bits_uop_cf_loadWaitStrict(LoadUnit_1_io_lsq_loadIn_bits_uop_cf_loadWaitStrict),
    .io_lsq_loadIn_bits_uop_cf_ftqPtr_flag(LoadUnit_1_io_lsq_loadIn_bits_uop_cf_ftqPtr_flag),
    .io_lsq_loadIn_bits_uop_cf_ftqPtr_value(LoadUnit_1_io_lsq_loadIn_bits_uop_cf_ftqPtr_value),
    .io_lsq_loadIn_bits_uop_cf_ftqOffset(LoadUnit_1_io_lsq_loadIn_bits_uop_cf_ftqOffset),
    .io_lsq_loadIn_bits_uop_ctrl_fuType(LoadUnit_1_io_lsq_loadIn_bits_uop_ctrl_fuType),
    .io_lsq_loadIn_bits_uop_ctrl_fuOpType(LoadUnit_1_io_lsq_loadIn_bits_uop_ctrl_fuOpType),
    .io_lsq_loadIn_bits_uop_ctrl_rfWen(LoadUnit_1_io_lsq_loadIn_bits_uop_ctrl_rfWen),
    .io_lsq_loadIn_bits_uop_ctrl_fpWen(LoadUnit_1_io_lsq_loadIn_bits_uop_ctrl_fpWen),
    .io_lsq_loadIn_bits_uop_ctrl_replayInst(LoadUnit_1_io_lsq_loadIn_bits_uop_ctrl_replayInst),
    .io_lsq_loadIn_bits_uop_pdest(LoadUnit_1_io_lsq_loadIn_bits_uop_pdest),
    .io_lsq_loadIn_bits_uop_robIdx_flag(LoadUnit_1_io_lsq_loadIn_bits_uop_robIdx_flag),
    .io_lsq_loadIn_bits_uop_robIdx_value(LoadUnit_1_io_lsq_loadIn_bits_uop_robIdx_value),
    .io_lsq_loadIn_bits_uop_lqIdx_flag(LoadUnit_1_io_lsq_loadIn_bits_uop_lqIdx_flag),
    .io_lsq_loadIn_bits_uop_lqIdx_value(LoadUnit_1_io_lsq_loadIn_bits_uop_lqIdx_value),
    .io_lsq_loadIn_bits_uop_sqIdx_flag(LoadUnit_1_io_lsq_loadIn_bits_uop_sqIdx_flag),
    .io_lsq_loadIn_bits_uop_sqIdx_value(LoadUnit_1_io_lsq_loadIn_bits_uop_sqIdx_value),
    .io_lsq_loadIn_bits_vaddr(LoadUnit_1_io_lsq_loadIn_bits_vaddr),
    .io_lsq_loadIn_bits_paddr(LoadUnit_1_io_lsq_loadIn_bits_paddr),
    .io_lsq_loadIn_bits_mask(LoadUnit_1_io_lsq_loadIn_bits_mask),
    .io_lsq_loadIn_bits_miss(LoadUnit_1_io_lsq_loadIn_bits_miss),
    .io_lsq_loadIn_bits_tlbMiss(LoadUnit_1_io_lsq_loadIn_bits_tlbMiss),
    .io_lsq_loadIn_bits_mmio(LoadUnit_1_io_lsq_loadIn_bits_mmio),
    .io_lsq_loadIn_bits_rarAllocated(LoadUnit_1_io_lsq_loadIn_bits_rarAllocated),
    .io_lsq_loadIn_bits_rarIndex(LoadUnit_1_io_lsq_loadIn_bits_rarIndex),
    .io_lsq_loadIn_bits_rawAllocated(LoadUnit_1_io_lsq_loadIn_bits_rawAllocated),
    .io_lsq_loadIn_bits_rawIndex(LoadUnit_1_io_lsq_loadIn_bits_rawIndex),
    .io_lsq_loadIn_bits_canAccept(LoadUnit_1_io_lsq_loadIn_bits_canAccept),
    .io_lsq_loadIn_bits_replayInfo_missMSHRId(LoadUnit_1_io_lsq_loadIn_bits_replayInfo_missMSHRId),
    .io_lsq_loadIn_bits_replayInfo_canForwardFullData(LoadUnit_1_io_lsq_loadIn_bits_replayInfo_canForwardFullData),
    .io_lsq_loadIn_bits_replayInfo_dataInvalidSqIdx_flag(LoadUnit_1_io_lsq_loadIn_bits_replayInfo_dataInvalidSqIdx_flag)
      ,
    .io_lsq_loadIn_bits_replayInfo_dataInvalidSqIdx_value(
      LoadUnit_1_io_lsq_loadIn_bits_replayInfo_dataInvalidSqIdx_value),
    .io_lsq_loadIn_bits_replayInfo_addrInvalidSqIdx_flag(LoadUnit_1_io_lsq_loadIn_bits_replayInfo_addrInvalidSqIdx_flag)
      ,
    .io_lsq_loadIn_bits_replayInfo_addrInvalidSqIdx_value(
      LoadUnit_1_io_lsq_loadIn_bits_replayInfo_addrInvalidSqIdx_value),
    .io_lsq_loadIn_bits_replayInfo_replayCarry_real_way_en(
      LoadUnit_1_io_lsq_loadIn_bits_replayInfo_replayCarry_real_way_en),
    .io_lsq_loadIn_bits_replayInfo_replayCarry_valid(LoadUnit_1_io_lsq_loadIn_bits_replayInfo_replayCarry_valid),
    .io_lsq_loadIn_bits_replayInfo_dataInLastBeat(LoadUnit_1_io_lsq_loadIn_bits_replayInfo_dataInLastBeat),
    .io_lsq_loadIn_bits_replayInfo_cause_0(LoadUnit_1_io_lsq_loadIn_bits_replayInfo_cause_0),
    .io_lsq_loadIn_bits_replayInfo_cause_1(LoadUnit_1_io_lsq_loadIn_bits_replayInfo_cause_1),
    .io_lsq_loadIn_bits_replayInfo_cause_2(LoadUnit_1_io_lsq_loadIn_bits_replayInfo_cause_2),
    .io_lsq_loadIn_bits_replayInfo_cause_3(LoadUnit_1_io_lsq_loadIn_bits_replayInfo_cause_3),
    .io_lsq_loadIn_bits_replayInfo_cause_4(LoadUnit_1_io_lsq_loadIn_bits_replayInfo_cause_4),
    .io_lsq_loadIn_bits_replayInfo_cause_5(LoadUnit_1_io_lsq_loadIn_bits_replayInfo_cause_5),
    .io_lsq_loadIn_bits_replayInfo_cause_6(LoadUnit_1_io_lsq_loadIn_bits_replayInfo_cause_6),
    .io_lsq_loadIn_bits_replayInfo_cause_7(LoadUnit_1_io_lsq_loadIn_bits_replayInfo_cause_7),
    .io_lsq_loadIn_bits_lqDataWenDup_1(LoadUnit_1_io_lsq_loadIn_bits_lqDataWenDup_1),
    .io_lsq_loadIn_bits_lqDataWenDup_2(LoadUnit_1_io_lsq_loadIn_bits_lqDataWenDup_2),
    .io_lsq_loadIn_bits_lqDataWenDup_3(LoadUnit_1_io_lsq_loadIn_bits_lqDataWenDup_3),
    .io_lsq_loadIn_bits_lqDataWenDup_5(LoadUnit_1_io_lsq_loadIn_bits_lqDataWenDup_5),
    .io_lsq_loadOut_ready(LoadUnit_1_io_lsq_loadOut_ready),
    .io_lsq_loadOut_valid(LoadUnit_1_io_lsq_loadOut_valid),
    .io_lsq_loadOut_bits_uop_cf_exceptionVec_4(LoadUnit_1_io_lsq_loadOut_bits_uop_cf_exceptionVec_4),
    .io_lsq_loadOut_bits_uop_cf_exceptionVec_5(LoadUnit_1_io_lsq_loadOut_bits_uop_cf_exceptionVec_5),
    .io_lsq_loadOut_bits_uop_cf_exceptionVec_13(LoadUnit_1_io_lsq_loadOut_bits_uop_cf_exceptionVec_13),
    .io_lsq_loadOut_bits_uop_cf_trigger_backendEn_1(LoadUnit_1_io_lsq_loadOut_bits_uop_cf_trigger_backendEn_1),
    .io_lsq_loadOut_bits_uop_cf_trigger_backendHit_0(LoadUnit_1_io_lsq_loadOut_bits_uop_cf_trigger_backendHit_0),
    .io_lsq_loadOut_bits_uop_cf_trigger_backendHit_1(LoadUnit_1_io_lsq_loadOut_bits_uop_cf_trigger_backendHit_1),
    .io_lsq_loadOut_bits_uop_cf_trigger_backendHit_4(LoadUnit_1_io_lsq_loadOut_bits_uop_cf_trigger_backendHit_4),
    .io_lsq_loadOut_bits_uop_ctrl_rfWen(LoadUnit_1_io_lsq_loadOut_bits_uop_ctrl_rfWen),
    .io_lsq_loadOut_bits_uop_ctrl_fpWen(LoadUnit_1_io_lsq_loadOut_bits_uop_ctrl_fpWen),
    .io_lsq_loadOut_bits_uop_ctrl_flushPipe(LoadUnit_1_io_lsq_loadOut_bits_uop_ctrl_flushPipe),
    .io_lsq_loadOut_bits_uop_ctrl_replayInst(LoadUnit_1_io_lsq_loadOut_bits_uop_ctrl_replayInst),
    .io_lsq_loadOut_bits_uop_pdest(LoadUnit_1_io_lsq_loadOut_bits_uop_pdest),
    .io_lsq_loadOut_bits_uop_robIdx_flag(LoadUnit_1_io_lsq_loadOut_bits_uop_robIdx_flag),
    .io_lsq_loadOut_bits_uop_robIdx_value(LoadUnit_1_io_lsq_loadOut_bits_uop_robIdx_value),
    .io_lsq_loadOut_bits_debug_isMMIO(LoadUnit_1_io_lsq_loadOut_bits_debug_isMMIO),
    .io_lsq_ldRawData_lqData(LoadUnit_1_io_lsq_ldRawData_lqData),
    .io_lsq_ldRawData_uop_ctrl_fuOpType(LoadUnit_1_io_lsq_ldRawData_uop_ctrl_fuOpType),
    .io_lsq_ldRawData_uop_ctrl_fpWen(LoadUnit_1_io_lsq_ldRawData_uop_ctrl_fpWen),
    .io_lsq_ldRawData_addrOffset(LoadUnit_1_io_lsq_ldRawData_addrOffset),
    .io_lsq_forward_vaddr(LoadUnit_1_io_lsq_forward_vaddr),
    .io_lsq_forward_paddr(LoadUnit_1_io_lsq_forward_paddr),
    .io_lsq_forward_uop_cf_waitForRobIdx_flag(LoadUnit_1_io_lsq_forward_uop_cf_waitForRobIdx_flag),
    .io_lsq_forward_uop_cf_waitForRobIdx_value(LoadUnit_1_io_lsq_forward_uop_cf_waitForRobIdx_value),
    .io_lsq_forward_uop_sqIdx_flag(LoadUnit_1_io_lsq_forward_uop_sqIdx_flag),
    .io_lsq_forward_uop_sqIdx_value(LoadUnit_1_io_lsq_forward_uop_sqIdx_value),
    .io_lsq_forward_valid(LoadUnit_1_io_lsq_forward_valid),
    .io_lsq_forward_forwardMask_0(LoadUnit_1_io_lsq_forward_forwardMask_0),
    .io_lsq_forward_forwardMask_1(LoadUnit_1_io_lsq_forward_forwardMask_1),
    .io_lsq_forward_forwardMask_2(LoadUnit_1_io_lsq_forward_forwardMask_2),
    .io_lsq_forward_forwardMask_3(LoadUnit_1_io_lsq_forward_forwardMask_3),
    .io_lsq_forward_forwardMask_4(LoadUnit_1_io_lsq_forward_forwardMask_4),
    .io_lsq_forward_forwardMask_5(LoadUnit_1_io_lsq_forward_forwardMask_5),
    .io_lsq_forward_forwardMask_6(LoadUnit_1_io_lsq_forward_forwardMask_6),
    .io_lsq_forward_forwardMask_7(LoadUnit_1_io_lsq_forward_forwardMask_7),
    .io_lsq_forward_forwardMask_8(LoadUnit_1_io_lsq_forward_forwardMask_8),
    .io_lsq_forward_forwardMask_9(LoadUnit_1_io_lsq_forward_forwardMask_9),
    .io_lsq_forward_forwardMask_10(LoadUnit_1_io_lsq_forward_forwardMask_10),
    .io_lsq_forward_forwardMask_11(LoadUnit_1_io_lsq_forward_forwardMask_11),
    .io_lsq_forward_forwardMask_12(LoadUnit_1_io_lsq_forward_forwardMask_12),
    .io_lsq_forward_forwardMask_13(LoadUnit_1_io_lsq_forward_forwardMask_13),
    .io_lsq_forward_forwardMask_14(LoadUnit_1_io_lsq_forward_forwardMask_14),
    .io_lsq_forward_forwardMask_15(LoadUnit_1_io_lsq_forward_forwardMask_15),
    .io_lsq_forward_forwardData_0(LoadUnit_1_io_lsq_forward_forwardData_0),
    .io_lsq_forward_forwardData_1(LoadUnit_1_io_lsq_forward_forwardData_1),
    .io_lsq_forward_forwardData_2(LoadUnit_1_io_lsq_forward_forwardData_2),
    .io_lsq_forward_forwardData_3(LoadUnit_1_io_lsq_forward_forwardData_3),
    .io_lsq_forward_forwardData_4(LoadUnit_1_io_lsq_forward_forwardData_4),
    .io_lsq_forward_forwardData_5(LoadUnit_1_io_lsq_forward_forwardData_5),
    .io_lsq_forward_forwardData_6(LoadUnit_1_io_lsq_forward_forwardData_6),
    .io_lsq_forward_forwardData_7(LoadUnit_1_io_lsq_forward_forwardData_7),
    .io_lsq_forward_forwardData_8(LoadUnit_1_io_lsq_forward_forwardData_8),
    .io_lsq_forward_forwardData_9(LoadUnit_1_io_lsq_forward_forwardData_9),
    .io_lsq_forward_forwardData_10(LoadUnit_1_io_lsq_forward_forwardData_10),
    .io_lsq_forward_forwardData_11(LoadUnit_1_io_lsq_forward_forwardData_11),
    .io_lsq_forward_forwardData_12(LoadUnit_1_io_lsq_forward_forwardData_12),
    .io_lsq_forward_forwardData_13(LoadUnit_1_io_lsq_forward_forwardData_13),
    .io_lsq_forward_forwardData_14(LoadUnit_1_io_lsq_forward_forwardData_14),
    .io_lsq_forward_forwardData_15(LoadUnit_1_io_lsq_forward_forwardData_15),
    .io_lsq_forward_sqIdx_flag(LoadUnit_1_io_lsq_forward_sqIdx_flag),
    .io_lsq_forward_dataInvalid(LoadUnit_1_io_lsq_forward_dataInvalid),
    .io_lsq_forward_matchInvalid(LoadUnit_1_io_lsq_forward_matchInvalid),
    .io_lsq_forward_schedWait(LoadUnit_1_io_lsq_forward_schedWait),
    .io_lsq_forward_sqIdxMask(LoadUnit_1_io_lsq_forward_sqIdxMask),
    .io_lsq_forward_dataInvalidSqIdx_flag(LoadUnit_1_io_lsq_forward_dataInvalidSqIdx_flag),
    .io_lsq_forward_dataInvalidSqIdx_value(LoadUnit_1_io_lsq_forward_dataInvalidSqIdx_value),
    .io_lsq_forward_addrInvalidSqIdx_flag(LoadUnit_1_io_lsq_forward_addrInvalidSqIdx_flag),
    .io_lsq_forward_addrInvalidSqIdx_value(LoadUnit_1_io_lsq_forward_addrInvalidSqIdx_value),
    .io_lsq_storeLoadViolationQuery_req_valid(LoadUnit_1_io_lsq_storeLoadViolationQuery_req_valid),
    .io_lsq_storeLoadViolationQuery_req_bits_uop_cf_foldpc(
      LoadUnit_1_io_lsq_storeLoadViolationQuery_req_bits_uop_cf_foldpc),
    .io_lsq_storeLoadViolationQuery_req_bits_uop_cf_ftqPtr_flag(
      LoadUnit_1_io_lsq_storeLoadViolationQuery_req_bits_uop_cf_ftqPtr_flag),
    .io_lsq_storeLoadViolationQuery_req_bits_uop_cf_ftqPtr_value(
      LoadUnit_1_io_lsq_storeLoadViolationQuery_req_bits_uop_cf_ftqPtr_value),
    .io_lsq_storeLoadViolationQuery_req_bits_uop_cf_ftqOffset(
      LoadUnit_1_io_lsq_storeLoadViolationQuery_req_bits_uop_cf_ftqOffset),
    .io_lsq_storeLoadViolationQuery_req_bits_uop_robIdx_flag(
      LoadUnit_1_io_lsq_storeLoadViolationQuery_req_bits_uop_robIdx_flag),
    .io_lsq_storeLoadViolationQuery_req_bits_uop_robIdx_value(
      LoadUnit_1_io_lsq_storeLoadViolationQuery_req_bits_uop_robIdx_value),
    .io_lsq_storeLoadViolationQuery_req_bits_uop_sqIdx_flag(
      LoadUnit_1_io_lsq_storeLoadViolationQuery_req_bits_uop_sqIdx_flag),
    .io_lsq_storeLoadViolationQuery_req_bits_uop_sqIdx_value(
      LoadUnit_1_io_lsq_storeLoadViolationQuery_req_bits_uop_sqIdx_value),
    .io_lsq_storeLoadViolationQuery_req_bits_index(LoadUnit_1_io_lsq_storeLoadViolationQuery_req_bits_index),
    .io_lsq_storeLoadViolationQuery_req_bits_allocated(LoadUnit_1_io_lsq_storeLoadViolationQuery_req_bits_allocated),
    .io_lsq_storeLoadViolationQuery_req_bits_datavalid(LoadUnit_1_io_lsq_storeLoadViolationQuery_req_bits_datavalid),
    .io_lsq_storeLoadViolationQuery_req_bits_mask(LoadUnit_1_io_lsq_storeLoadViolationQuery_req_bits_mask),
    .io_lsq_storeLoadViolationQuery_req_bits_paddr(LoadUnit_1_io_lsq_storeLoadViolationQuery_req_bits_paddr),
    .io_lsq_storeLoadViolationQuery_resp_bits_index(LoadUnit_1_io_lsq_storeLoadViolationQuery_resp_bits_index),
    .io_lsq_storeLoadViolationQuery_resp_bits_canAccept(LoadUnit_1_io_lsq_storeLoadViolationQuery_resp_bits_canAccept),
    .io_lsq_storeLoadViolationQuery_resp_bits_allocated(LoadUnit_1_io_lsq_storeLoadViolationQuery_resp_bits_allocated),
    .io_lsq_loadLoadViolationQuery_req_valid(LoadUnit_1_io_lsq_loadLoadViolationQuery_req_valid),
    .io_lsq_loadLoadViolationQuery_req_bits_uop_robIdx_flag(
      LoadUnit_1_io_lsq_loadLoadViolationQuery_req_bits_uop_robIdx_flag),
    .io_lsq_loadLoadViolationQuery_req_bits_uop_robIdx_value(
      LoadUnit_1_io_lsq_loadLoadViolationQuery_req_bits_uop_robIdx_value),
    .io_lsq_loadLoadViolationQuery_req_bits_uop_lqIdx_flag(
      LoadUnit_1_io_lsq_loadLoadViolationQuery_req_bits_uop_lqIdx_flag),
    .io_lsq_loadLoadViolationQuery_req_bits_uop_lqIdx_value(
      LoadUnit_1_io_lsq_loadLoadViolationQuery_req_bits_uop_lqIdx_value),
    .io_lsq_loadLoadViolationQuery_req_bits_index(LoadUnit_1_io_lsq_loadLoadViolationQuery_req_bits_index),
    .io_lsq_loadLoadViolationQuery_req_bits_allocated(LoadUnit_1_io_lsq_loadLoadViolationQuery_req_bits_allocated),
    .io_lsq_loadLoadViolationQuery_req_bits_datavalid(LoadUnit_1_io_lsq_loadLoadViolationQuery_req_bits_datavalid),
    .io_lsq_loadLoadViolationQuery_req_bits_miss(LoadUnit_1_io_lsq_loadLoadViolationQuery_req_bits_miss),
    .io_lsq_loadLoadViolationQuery_req_bits_paddr(LoadUnit_1_io_lsq_loadLoadViolationQuery_req_bits_paddr),
    .io_lsq_loadLoadViolationQuery_resp_valid(LoadUnit_1_io_lsq_loadLoadViolationQuery_resp_valid),
    .io_lsq_loadLoadViolationQuery_resp_bits_index(LoadUnit_1_io_lsq_loadLoadViolationQuery_resp_bits_index),
    .io_lsq_loadLoadViolationQuery_resp_bits_canAccept(LoadUnit_1_io_lsq_loadLoadViolationQuery_resp_bits_canAccept),
    .io_lsq_loadLoadViolationQuery_resp_bits_allocated(LoadUnit_1_io_lsq_loadLoadViolationQuery_resp_bits_allocated),
    .io_lsq_loadLoadViolationQuery_resp_bits_replayFromFetch(
      LoadUnit_1_io_lsq_loadLoadViolationQuery_resp_bits_replayFromFetch),
    .io_lsq_trigger_hitLoadAddrTriggerHitVec_0(LoadUnit_1_io_lsq_trigger_hitLoadAddrTriggerHitVec_0),
    .io_lsq_trigger_hitLoadAddrTriggerHitVec_1(LoadUnit_1_io_lsq_trigger_hitLoadAddrTriggerHitVec_1),
    .io_lsq_trigger_hitLoadAddrTriggerHitVec_2(LoadUnit_1_io_lsq_trigger_hitLoadAddrTriggerHitVec_2),
    .io_lsq_trigger_lqLoadAddrTriggerHitVec_0(LoadUnit_1_io_lsq_trigger_lqLoadAddrTriggerHitVec_0),
    .io_lsq_trigger_lqLoadAddrTriggerHitVec_1(LoadUnit_1_io_lsq_trigger_lqLoadAddrTriggerHitVec_1),
    .io_lsq_trigger_lqLoadAddrTriggerHitVec_2(LoadUnit_1_io_lsq_trigger_lqLoadAddrTriggerHitVec_2),
    .io_tlDchannel_valid(LoadUnit_1_io_tlDchannel_valid),
    .io_tlDchannel_data(LoadUnit_1_io_tlDchannel_data),
    .io_tlDchannel_mshrid(LoadUnit_1_io_tlDchannel_mshrid),
    .io_tlDchannel_last(LoadUnit_1_io_tlDchannel_last),
    .io_forward_mshr_valid(LoadUnit_1_io_forward_mshr_valid),
    .io_forward_mshr_mshrid(LoadUnit_1_io_forward_mshr_mshrid),
    .io_forward_mshr_paddr(LoadUnit_1_io_forward_mshr_paddr),
    .io_forward_mshr_forward_mshr(LoadUnit_1_io_forward_mshr_forward_mshr),
    .io_forward_mshr_forwardData_0(LoadUnit_1_io_forward_mshr_forwardData_0),
    .io_forward_mshr_forwardData_1(LoadUnit_1_io_forward_mshr_forwardData_1),
    .io_forward_mshr_forwardData_2(LoadUnit_1_io_forward_mshr_forwardData_2),
    .io_forward_mshr_forwardData_3(LoadUnit_1_io_forward_mshr_forwardData_3),
    .io_forward_mshr_forwardData_4(LoadUnit_1_io_forward_mshr_forwardData_4),
    .io_forward_mshr_forwardData_5(LoadUnit_1_io_forward_mshr_forwardData_5),
    .io_forward_mshr_forwardData_6(LoadUnit_1_io_forward_mshr_forwardData_6),
    .io_forward_mshr_forwardData_7(LoadUnit_1_io_forward_mshr_forwardData_7),
    .io_forward_mshr_forwardData_8(LoadUnit_1_io_forward_mshr_forwardData_8),
    .io_forward_mshr_forwardData_9(LoadUnit_1_io_forward_mshr_forwardData_9),
    .io_forward_mshr_forwardData_10(LoadUnit_1_io_forward_mshr_forwardData_10),
    .io_forward_mshr_forwardData_11(LoadUnit_1_io_forward_mshr_forwardData_11),
    .io_forward_mshr_forwardData_12(LoadUnit_1_io_forward_mshr_forwardData_12),
    .io_forward_mshr_forwardData_13(LoadUnit_1_io_forward_mshr_forwardData_13),
    .io_forward_mshr_forwardData_14(LoadUnit_1_io_forward_mshr_forwardData_14),
    .io_forward_mshr_forwardData_15(LoadUnit_1_io_forward_mshr_forwardData_15),
    .io_forward_mshr_forward_result_valid(LoadUnit_1_io_forward_mshr_forward_result_valid),
    .io_trigger_0_tdata2(LoadUnit_1_io_trigger_0_tdata2),
    .io_trigger_0_matchType(LoadUnit_1_io_trigger_0_matchType),
    .io_trigger_0_tEnable(LoadUnit_1_io_trigger_0_tEnable),
    .io_trigger_0_addrHit(LoadUnit_1_io_trigger_0_addrHit),
    .io_trigger_1_tdata2(LoadUnit_1_io_trigger_1_tdata2),
    .io_trigger_1_matchType(LoadUnit_1_io_trigger_1_matchType),
    .io_trigger_1_tEnable(LoadUnit_1_io_trigger_1_tEnable),
    .io_trigger_1_addrHit(LoadUnit_1_io_trigger_1_addrHit),
    .io_trigger_2_tdata2(LoadUnit_1_io_trigger_2_tdata2),
    .io_trigger_2_matchType(LoadUnit_1_io_trigger_2_matchType),
    .io_trigger_2_tEnable(LoadUnit_1_io_trigger_2_tEnable),
    .io_trigger_2_addrHit(LoadUnit_1_io_trigger_2_addrHit),
    .io_tlb_req_valid(LoadUnit_1_io_tlb_req_valid),
    .io_tlb_req_bits_vaddr(LoadUnit_1_io_tlb_req_bits_vaddr),
    .io_tlb_req_bits_cmd(LoadUnit_1_io_tlb_req_bits_cmd),
    .io_tlb_req_bits_no_translate(LoadUnit_1_io_tlb_req_bits_no_translate),
    .io_tlb_req_kill(LoadUnit_1_io_tlb_req_kill),
    .io_tlb_resp_bits_paddr_0(LoadUnit_1_io_tlb_resp_bits_paddr_0),
    .io_tlb_resp_bits_paddr_1(LoadUnit_1_io_tlb_resp_bits_paddr_1),
    .io_tlb_resp_bits_miss(LoadUnit_1_io_tlb_resp_bits_miss),
    .io_tlb_resp_bits_excp_0_pf_ld(LoadUnit_1_io_tlb_resp_bits_excp_0_pf_ld),
    .io_tlb_resp_bits_excp_0_af_ld(LoadUnit_1_io_tlb_resp_bits_excp_0_af_ld),
    .io_tlb_resp_bits_static_pm_valid(LoadUnit_1_io_tlb_resp_bits_static_pm_valid),
    .io_tlb_resp_bits_static_pm_bits(LoadUnit_1_io_tlb_resp_bits_static_pm_bits),
    .io_pmp_ld(LoadUnit_1_io_pmp_ld),
    .io_pmp_mmio(LoadUnit_1_io_pmp_mmio),
    .io_fastpathOut_data(LoadUnit_1_io_fastpathOut_data),
    .io_fastpathOut_valid(LoadUnit_1_io_fastpathOut_valid),
    .io_fastpathIn_data(LoadUnit_1_io_fastpathIn_data),
    .io_fastpathIn_valid(LoadUnit_1_io_fastpathIn_valid),
    .io_loadFastMatch(LoadUnit_1_io_loadFastMatch),
    .io_loadFastImm(LoadUnit_1_io_loadFastImm),
    .io_csrCtrl_ldld_vio_check_enable(LoadUnit_1_io_csrCtrl_ldld_vio_check_enable),
    .io_csrCtrl_cache_error_enable(LoadUnit_1_io_csrCtrl_cache_error_enable),
    .io_correctTableQuery_req_addr(LoadUnit_1_io_correctTableQuery_req_addr),
    .io_correctTableQuery_resp_strict(LoadUnit_1_io_correctTableQuery_resp_strict),
    .io_correctTableUpdate_valid(LoadUnit_1_io_correctTableUpdate_valid),
    .io_correctTableUpdate_bits_addr(LoadUnit_1_io_correctTableUpdate_bits_addr),
    .io_correctTableUpdate_bits_strict(LoadUnit_1_io_correctTableUpdate_bits_strict),
    .io_correctTableUpdate_bits_violation(LoadUnit_1_io_correctTableUpdate_bits_violation),
    .io_reExecuteQuery_0_valid(LoadUnit_1_io_reExecuteQuery_0_valid),
    .io_reExecuteQuery_0_bits_robIdx_flag(LoadUnit_1_io_reExecuteQuery_0_bits_robIdx_flag),
    .io_reExecuteQuery_0_bits_robIdx_value(LoadUnit_1_io_reExecuteQuery_0_bits_robIdx_value),
    .io_reExecuteQuery_0_bits_paddr(LoadUnit_1_io_reExecuteQuery_0_bits_paddr),
    .io_reExecuteQuery_0_bits_mask(LoadUnit_1_io_reExecuteQuery_0_bits_mask),
    .io_reExecuteQuery_1_valid(LoadUnit_1_io_reExecuteQuery_1_valid),
    .io_reExecuteQuery_1_bits_robIdx_flag(LoadUnit_1_io_reExecuteQuery_1_bits_robIdx_flag),
    .io_reExecuteQuery_1_bits_robIdx_value(LoadUnit_1_io_reExecuteQuery_1_bits_robIdx_value),
    .io_reExecuteQuery_1_bits_paddr(LoadUnit_1_io_reExecuteQuery_1_bits_paddr),
    .io_reExecuteQuery_1_bits_mask(LoadUnit_1_io_reExecuteQuery_1_bits_mask),
    .io_replay_ready(LoadUnit_1_io_replay_ready),
    .io_replay_valid(LoadUnit_1_io_replay_valid),
    .io_replay_bits_uop_cf_foldpc(LoadUnit_1_io_replay_bits_uop_cf_foldpc),
    .io_replay_bits_uop_cf_trigger_backendEn_1(LoadUnit_1_io_replay_bits_uop_cf_trigger_backendEn_1),
    .io_replay_bits_uop_cf_trigger_backendHit_0(LoadUnit_1_io_replay_bits_uop_cf_trigger_backendHit_0),
    .io_replay_bits_uop_cf_trigger_backendHit_1(LoadUnit_1_io_replay_bits_uop_cf_trigger_backendHit_1),
    .io_replay_bits_uop_cf_trigger_backendHit_4(LoadUnit_1_io_replay_bits_uop_cf_trigger_backendHit_4),
    .io_replay_bits_uop_cf_waitForRobIdx_flag(LoadUnit_1_io_replay_bits_uop_cf_waitForRobIdx_flag),
    .io_replay_bits_uop_cf_waitForRobIdx_value(LoadUnit_1_io_replay_bits_uop_cf_waitForRobIdx_value),
    .io_replay_bits_uop_cf_loadWaitBit(LoadUnit_1_io_replay_bits_uop_cf_loadWaitBit),
    .io_replay_bits_uop_cf_loadWaitStrict(LoadUnit_1_io_replay_bits_uop_cf_loadWaitStrict),
    .io_replay_bits_uop_cf_ftqPtr_flag(LoadUnit_1_io_replay_bits_uop_cf_ftqPtr_flag),
    .io_replay_bits_uop_cf_ftqPtr_value(LoadUnit_1_io_replay_bits_uop_cf_ftqPtr_value),
    .io_replay_bits_uop_cf_ftqOffset(LoadUnit_1_io_replay_bits_uop_cf_ftqOffset),
    .io_replay_bits_uop_ctrl_fuType(LoadUnit_1_io_replay_bits_uop_ctrl_fuType),
    .io_replay_bits_uop_ctrl_fuOpType(LoadUnit_1_io_replay_bits_uop_ctrl_fuOpType),
    .io_replay_bits_uop_ctrl_rfWen(LoadUnit_1_io_replay_bits_uop_ctrl_rfWen),
    .io_replay_bits_uop_ctrl_fpWen(LoadUnit_1_io_replay_bits_uop_ctrl_fpWen),
    .io_replay_bits_uop_pdest(LoadUnit_1_io_replay_bits_uop_pdest),
    .io_replay_bits_uop_robIdx_flag(LoadUnit_1_io_replay_bits_uop_robIdx_flag),
    .io_replay_bits_uop_robIdx_value(LoadUnit_1_io_replay_bits_uop_robIdx_value),
    .io_replay_bits_uop_lqIdx_flag(LoadUnit_1_io_replay_bits_uop_lqIdx_flag),
    .io_replay_bits_uop_lqIdx_value(LoadUnit_1_io_replay_bits_uop_lqIdx_value),
    .io_replay_bits_uop_sqIdx_flag(LoadUnit_1_io_replay_bits_uop_sqIdx_flag),
    .io_replay_bits_uop_sqIdx_value(LoadUnit_1_io_replay_bits_uop_sqIdx_value),
    .io_replay_bits_vaddr(LoadUnit_1_io_replay_bits_vaddr),
    .io_replay_bits_isFirstIssue(LoadUnit_1_io_replay_bits_isFirstIssue),
    .io_replay_bits_replayCarry_real_way_en(LoadUnit_1_io_replay_bits_replayCarry_real_way_en),
    .io_replay_bits_replayCarry_valid(LoadUnit_1_io_replay_bits_replayCarry_valid),
    .io_replay_bits_mshrid(LoadUnit_1_io_replay_bits_mshrid),
    .io_replay_bits_forward_tlDchannel(LoadUnit_1_io_replay_bits_forward_tlDchannel),
    .io_replay_bits_rarAllocated(LoadUnit_1_io_replay_bits_rarAllocated),
    .io_replay_bits_rarIndex(LoadUnit_1_io_replay_bits_rarIndex),
    .io_replay_bits_rawAllocated(LoadUnit_1_io_replay_bits_rawAllocated),
    .io_replay_bits_rawIndex(LoadUnit_1_io_replay_bits_rawIndex),
    .io_lqReplayFull(LoadUnit_1_io_lqReplayFull),
    .io_perf_0_value(LoadUnit_1_io_perf_0_value),
    .io_perf_1_value(LoadUnit_1_io_perf_1_value),
    .io_perf_2_value(LoadUnit_1_io_perf_2_value),
    .io_perf_3_value(LoadUnit_1_io_perf_3_value),
    .io_perf_4_value(LoadUnit_1_io_perf_4_value),
    .io_perf_5_value(LoadUnit_1_io_perf_5_value),
    .io_perf_6_value(LoadUnit_1_io_perf_6_value)
  );
  StoreUnit StoreUnit_0 ( // @[MemBlock.scala 140:57]
    .clock(StoreUnit_0_clock),
    .reset(StoreUnit_0_reset),
    .io_stin_valid(StoreUnit_0_io_stin_valid),
    .io_stin_bits_uop_cf_trigger_backendEn_0(StoreUnit_0_io_stin_bits_uop_cf_trigger_backendEn_0),
    .io_stin_bits_uop_cf_storeSetHit(StoreUnit_0_io_stin_bits_uop_cf_storeSetHit),
    .io_stin_bits_uop_cf_ssid(StoreUnit_0_io_stin_bits_uop_cf_ssid),
    .io_stin_bits_uop_cf_ftqPtr_value(StoreUnit_0_io_stin_bits_uop_cf_ftqPtr_value),
    .io_stin_bits_uop_cf_ftqOffset(StoreUnit_0_io_stin_bits_uop_cf_ftqOffset),
    .io_stin_bits_uop_ctrl_fuOpType(StoreUnit_0_io_stin_bits_uop_ctrl_fuOpType),
    .io_stin_bits_uop_ctrl_imm(StoreUnit_0_io_stin_bits_uop_ctrl_imm),
    .io_stin_bits_uop_robIdx_flag(StoreUnit_0_io_stin_bits_uop_robIdx_flag),
    .io_stin_bits_uop_robIdx_value(StoreUnit_0_io_stin_bits_uop_robIdx_value),
    .io_stin_bits_uop_sqIdx_flag(StoreUnit_0_io_stin_bits_uop_sqIdx_flag),
    .io_stin_bits_uop_sqIdx_value(StoreUnit_0_io_stin_bits_uop_sqIdx_value),
    .io_stin_bits_src_0(StoreUnit_0_io_stin_bits_src_0),
    .io_redirect_valid(StoreUnit_0_io_redirect_valid),
    .io_redirect_bits_robIdx_flag(StoreUnit_0_io_redirect_bits_robIdx_flag),
    .io_redirect_bits_robIdx_value(StoreUnit_0_io_redirect_bits_robIdx_value),
    .io_redirect_bits_level(StoreUnit_0_io_redirect_bits_level),
    .io_feedbackSlow_valid(StoreUnit_0_io_feedbackSlow_valid),
    .io_feedbackSlow_bits_rsIdx(StoreUnit_0_io_feedbackSlow_bits_rsIdx),
    .io_feedbackSlow_bits_hit(StoreUnit_0_io_feedbackSlow_bits_hit),
    .io_tlb_req_valid(StoreUnit_0_io_tlb_req_valid),
    .io_tlb_req_bits_vaddr(StoreUnit_0_io_tlb_req_bits_vaddr),
    .io_tlb_resp_bits_paddr_0(StoreUnit_0_io_tlb_resp_bits_paddr_0),
    .io_tlb_resp_bits_miss(StoreUnit_0_io_tlb_resp_bits_miss),
    .io_tlb_resp_bits_excp_0_pf_st(StoreUnit_0_io_tlb_resp_bits_excp_0_pf_st),
    .io_tlb_resp_bits_excp_0_af_st(StoreUnit_0_io_tlb_resp_bits_excp_0_af_st),
    .io_tlb_resp_bits_static_pm_valid(StoreUnit_0_io_tlb_resp_bits_static_pm_valid),
    .io_tlb_resp_bits_static_pm_bits(StoreUnit_0_io_tlb_resp_bits_static_pm_bits),
    .io_pmp_st(StoreUnit_0_io_pmp_st),
    .io_pmp_mmio(StoreUnit_0_io_pmp_mmio),
    .io_pmp_atomic(StoreUnit_0_io_pmp_atomic),
    .io_rsIdx(StoreUnit_0_io_rsIdx),
    .io_lsq_valid(StoreUnit_0_io_lsq_valid),
    .io_lsq_bits_uop_cf_ftqPtr_value(StoreUnit_0_io_lsq_bits_uop_cf_ftqPtr_value),
    .io_lsq_bits_uop_cf_ftqOffset(StoreUnit_0_io_lsq_bits_uop_cf_ftqOffset),
    .io_lsq_bits_uop_ctrl_fuOpType(StoreUnit_0_io_lsq_bits_uop_ctrl_fuOpType),
    .io_lsq_bits_uop_robIdx_flag(StoreUnit_0_io_lsq_bits_uop_robIdx_flag),
    .io_lsq_bits_uop_robIdx_value(StoreUnit_0_io_lsq_bits_uop_robIdx_value),
    .io_lsq_bits_uop_sqIdx_flag(StoreUnit_0_io_lsq_bits_uop_sqIdx_flag),
    .io_lsq_bits_uop_sqIdx_value(StoreUnit_0_io_lsq_bits_uop_sqIdx_value),
    .io_lsq_bits_vaddr(StoreUnit_0_io_lsq_bits_vaddr),
    .io_lsq_bits_paddr(StoreUnit_0_io_lsq_bits_paddr),
    .io_lsq_bits_mask(StoreUnit_0_io_lsq_bits_mask),
    .io_lsq_bits_wlineflag(StoreUnit_0_io_lsq_bits_wlineflag),
    .io_lsq_bits_miss(StoreUnit_0_io_lsq_bits_miss),
    .io_lsq_replenish_mmio(StoreUnit_0_io_lsq_replenish_mmio),
    .io_lsq_replenish_atomic(StoreUnit_0_io_lsq_replenish_atomic),
    .io_stout_valid(StoreUnit_0_io_stout_valid),
    .io_stout_bits_uop_cf_exceptionVec_6(StoreUnit_0_io_stout_bits_uop_cf_exceptionVec_6),
    .io_stout_bits_uop_cf_exceptionVec_7(StoreUnit_0_io_stout_bits_uop_cf_exceptionVec_7),
    .io_stout_bits_uop_cf_exceptionVec_15(StoreUnit_0_io_stout_bits_uop_cf_exceptionVec_15),
    .io_stout_bits_uop_cf_trigger_backendEn_0(StoreUnit_0_io_stout_bits_uop_cf_trigger_backendEn_0),
    .io_stout_bits_uop_robIdx_flag(StoreUnit_0_io_stout_bits_uop_robIdx_flag),
    .io_stout_bits_uop_robIdx_value(StoreUnit_0_io_stout_bits_uop_robIdx_value),
    .io_stout_bits_debug_isMMIO(StoreUnit_0_io_stout_bits_debug_isMMIO),
    .io_stout_bits_debug_vaddr(StoreUnit_0_io_stout_bits_debug_vaddr),
    .io_storeMaskOut_valid(StoreUnit_0_io_storeMaskOut_valid),
    .io_storeMaskOut_bits_sqIdx_value(StoreUnit_0_io_storeMaskOut_bits_sqIdx_value),
    .io_storeMaskOut_bits_mask(StoreUnit_0_io_storeMaskOut_bits_mask),
    .io_reExecuteQuery_valid(StoreUnit_0_io_reExecuteQuery_valid),
    .io_reExecuteQuery_bits_robIdx_flag(StoreUnit_0_io_reExecuteQuery_bits_robIdx_flag),
    .io_reExecuteQuery_bits_robIdx_value(StoreUnit_0_io_reExecuteQuery_bits_robIdx_value),
    .io_reExecuteQuery_bits_paddr(StoreUnit_0_io_reExecuteQuery_bits_paddr),
    .io_reExecuteQuery_bits_mask(StoreUnit_0_io_reExecuteQuery_bits_mask),
    .io_issue_valid(StoreUnit_0_io_issue_valid),
    .io_issue_bits_uop_cf_storeSetHit(StoreUnit_0_io_issue_bits_uop_cf_storeSetHit),
    .io_issue_bits_uop_cf_ssid(StoreUnit_0_io_issue_bits_uop_cf_ssid),
    .io_issue_bits_uop_robIdx_value(StoreUnit_0_io_issue_bits_uop_robIdx_value)
  );
  StoreUnit StoreUnit_1 ( // @[MemBlock.scala 140:57]
    .clock(StoreUnit_1_clock),
    .reset(StoreUnit_1_reset),
    .io_stin_valid(StoreUnit_1_io_stin_valid),
    .io_stin_bits_uop_cf_trigger_backendEn_0(StoreUnit_1_io_stin_bits_uop_cf_trigger_backendEn_0),
    .io_stin_bits_uop_cf_storeSetHit(StoreUnit_1_io_stin_bits_uop_cf_storeSetHit),
    .io_stin_bits_uop_cf_ssid(StoreUnit_1_io_stin_bits_uop_cf_ssid),
    .io_stin_bits_uop_cf_ftqPtr_value(StoreUnit_1_io_stin_bits_uop_cf_ftqPtr_value),
    .io_stin_bits_uop_cf_ftqOffset(StoreUnit_1_io_stin_bits_uop_cf_ftqOffset),
    .io_stin_bits_uop_ctrl_fuOpType(StoreUnit_1_io_stin_bits_uop_ctrl_fuOpType),
    .io_stin_bits_uop_ctrl_imm(StoreUnit_1_io_stin_bits_uop_ctrl_imm),
    .io_stin_bits_uop_robIdx_flag(StoreUnit_1_io_stin_bits_uop_robIdx_flag),
    .io_stin_bits_uop_robIdx_value(StoreUnit_1_io_stin_bits_uop_robIdx_value),
    .io_stin_bits_uop_sqIdx_flag(StoreUnit_1_io_stin_bits_uop_sqIdx_flag),
    .io_stin_bits_uop_sqIdx_value(StoreUnit_1_io_stin_bits_uop_sqIdx_value),
    .io_stin_bits_src_0(StoreUnit_1_io_stin_bits_src_0),
    .io_redirect_valid(StoreUnit_1_io_redirect_valid),
    .io_redirect_bits_robIdx_flag(StoreUnit_1_io_redirect_bits_robIdx_flag),
    .io_redirect_bits_robIdx_value(StoreUnit_1_io_redirect_bits_robIdx_value),
    .io_redirect_bits_level(StoreUnit_1_io_redirect_bits_level),
    .io_feedbackSlow_valid(StoreUnit_1_io_feedbackSlow_valid),
    .io_feedbackSlow_bits_rsIdx(StoreUnit_1_io_feedbackSlow_bits_rsIdx),
    .io_feedbackSlow_bits_hit(StoreUnit_1_io_feedbackSlow_bits_hit),
    .io_tlb_req_valid(StoreUnit_1_io_tlb_req_valid),
    .io_tlb_req_bits_vaddr(StoreUnit_1_io_tlb_req_bits_vaddr),
    .io_tlb_resp_bits_paddr_0(StoreUnit_1_io_tlb_resp_bits_paddr_0),
    .io_tlb_resp_bits_miss(StoreUnit_1_io_tlb_resp_bits_miss),
    .io_tlb_resp_bits_excp_0_pf_st(StoreUnit_1_io_tlb_resp_bits_excp_0_pf_st),
    .io_tlb_resp_bits_excp_0_af_st(StoreUnit_1_io_tlb_resp_bits_excp_0_af_st),
    .io_tlb_resp_bits_static_pm_valid(StoreUnit_1_io_tlb_resp_bits_static_pm_valid),
    .io_tlb_resp_bits_static_pm_bits(StoreUnit_1_io_tlb_resp_bits_static_pm_bits),
    .io_pmp_st(StoreUnit_1_io_pmp_st),
    .io_pmp_mmio(StoreUnit_1_io_pmp_mmio),
    .io_pmp_atomic(StoreUnit_1_io_pmp_atomic),
    .io_rsIdx(StoreUnit_1_io_rsIdx),
    .io_lsq_valid(StoreUnit_1_io_lsq_valid),
    .io_lsq_bits_uop_cf_ftqPtr_value(StoreUnit_1_io_lsq_bits_uop_cf_ftqPtr_value),
    .io_lsq_bits_uop_cf_ftqOffset(StoreUnit_1_io_lsq_bits_uop_cf_ftqOffset),
    .io_lsq_bits_uop_ctrl_fuOpType(StoreUnit_1_io_lsq_bits_uop_ctrl_fuOpType),
    .io_lsq_bits_uop_robIdx_flag(StoreUnit_1_io_lsq_bits_uop_robIdx_flag),
    .io_lsq_bits_uop_robIdx_value(StoreUnit_1_io_lsq_bits_uop_robIdx_value),
    .io_lsq_bits_uop_sqIdx_flag(StoreUnit_1_io_lsq_bits_uop_sqIdx_flag),
    .io_lsq_bits_uop_sqIdx_value(StoreUnit_1_io_lsq_bits_uop_sqIdx_value),
    .io_lsq_bits_vaddr(StoreUnit_1_io_lsq_bits_vaddr),
    .io_lsq_bits_paddr(StoreUnit_1_io_lsq_bits_paddr),
    .io_lsq_bits_mask(StoreUnit_1_io_lsq_bits_mask),
    .io_lsq_bits_wlineflag(StoreUnit_1_io_lsq_bits_wlineflag),
    .io_lsq_bits_miss(StoreUnit_1_io_lsq_bits_miss),
    .io_lsq_replenish_mmio(StoreUnit_1_io_lsq_replenish_mmio),
    .io_lsq_replenish_atomic(StoreUnit_1_io_lsq_replenish_atomic),
    .io_stout_valid(StoreUnit_1_io_stout_valid),
    .io_stout_bits_uop_cf_exceptionVec_6(StoreUnit_1_io_stout_bits_uop_cf_exceptionVec_6),
    .io_stout_bits_uop_cf_exceptionVec_7(StoreUnit_1_io_stout_bits_uop_cf_exceptionVec_7),
    .io_stout_bits_uop_cf_exceptionVec_15(StoreUnit_1_io_stout_bits_uop_cf_exceptionVec_15),
    .io_stout_bits_uop_cf_trigger_backendEn_0(StoreUnit_1_io_stout_bits_uop_cf_trigger_backendEn_0),
    .io_stout_bits_uop_robIdx_flag(StoreUnit_1_io_stout_bits_uop_robIdx_flag),
    .io_stout_bits_uop_robIdx_value(StoreUnit_1_io_stout_bits_uop_robIdx_value),
    .io_stout_bits_debug_isMMIO(StoreUnit_1_io_stout_bits_debug_isMMIO),
    .io_stout_bits_debug_vaddr(StoreUnit_1_io_stout_bits_debug_vaddr),
    .io_storeMaskOut_valid(StoreUnit_1_io_storeMaskOut_valid),
    .io_storeMaskOut_bits_sqIdx_value(StoreUnit_1_io_storeMaskOut_bits_sqIdx_value),
    .io_storeMaskOut_bits_mask(StoreUnit_1_io_storeMaskOut_bits_mask),
    .io_reExecuteQuery_valid(StoreUnit_1_io_reExecuteQuery_valid),
    .io_reExecuteQuery_bits_robIdx_flag(StoreUnit_1_io_reExecuteQuery_bits_robIdx_flag),
    .io_reExecuteQuery_bits_robIdx_value(StoreUnit_1_io_reExecuteQuery_bits_robIdx_value),
    .io_reExecuteQuery_bits_paddr(StoreUnit_1_io_reExecuteQuery_bits_paddr),
    .io_reExecuteQuery_bits_mask(StoreUnit_1_io_reExecuteQuery_bits_mask),
    .io_issue_valid(StoreUnit_1_io_issue_valid),
    .io_issue_bits_uop_cf_storeSetHit(StoreUnit_1_io_issue_bits_uop_cf_storeSetHit),
    .io_issue_bits_uop_cf_ssid(StoreUnit_1_io_issue_bits_uop_cf_ssid),
    .io_issue_bits_uop_robIdx_value(StoreUnit_1_io_issue_bits_uop_robIdx_value)
  );
  StdExeUnit stdExeUnits_0 ( // @[MemBlock.scala 141:58]
    .io_fromInt_ready(stdExeUnits_0_io_fromInt_ready),
    .io_fromInt_valid(stdExeUnits_0_io_fromInt_valid),
    .io_fromInt_bits_uop_ctrl_fuType(stdExeUnits_0_io_fromInt_bits_uop_ctrl_fuType),
    .io_fromInt_bits_uop_ctrl_fuOpType(stdExeUnits_0_io_fromInt_bits_uop_ctrl_fuOpType),
    .io_fromInt_bits_uop_robIdx_flag(stdExeUnits_0_io_fromInt_bits_uop_robIdx_flag),
    .io_fromInt_bits_uop_robIdx_value(stdExeUnits_0_io_fromInt_bits_uop_robIdx_value),
    .io_fromInt_bits_uop_sqIdx_flag(stdExeUnits_0_io_fromInt_bits_uop_sqIdx_flag),
    .io_fromInt_bits_uop_sqIdx_value(stdExeUnits_0_io_fromInt_bits_uop_sqIdx_value),
    .io_fromInt_bits_src_0(stdExeUnits_0_io_fromInt_bits_src_0),
    .io_out_valid(stdExeUnits_0_io_out_valid),
    .io_out_bits_uop_ctrl_fuType(stdExeUnits_0_io_out_bits_uop_ctrl_fuType),
    .io_out_bits_uop_ctrl_fuOpType(stdExeUnits_0_io_out_bits_uop_ctrl_fuOpType),
    .io_out_bits_uop_robIdx_flag(stdExeUnits_0_io_out_bits_uop_robIdx_flag),
    .io_out_bits_uop_robIdx_value(stdExeUnits_0_io_out_bits_uop_robIdx_value),
    .io_out_bits_uop_sqIdx_flag(stdExeUnits_0_io_out_bits_uop_sqIdx_flag),
    .io_out_bits_uop_sqIdx_value(stdExeUnits_0_io_out_bits_uop_sqIdx_value),
    .io_out_bits_data(stdExeUnits_0_io_out_bits_data)
  );
  StdExeUnit stdExeUnits_1 ( // @[MemBlock.scala 141:58]
    .io_fromInt_ready(stdExeUnits_1_io_fromInt_ready),
    .io_fromInt_valid(stdExeUnits_1_io_fromInt_valid),
    .io_fromInt_bits_uop_ctrl_fuType(stdExeUnits_1_io_fromInt_bits_uop_ctrl_fuType),
    .io_fromInt_bits_uop_ctrl_fuOpType(stdExeUnits_1_io_fromInt_bits_uop_ctrl_fuOpType),
    .io_fromInt_bits_uop_robIdx_flag(stdExeUnits_1_io_fromInt_bits_uop_robIdx_flag),
    .io_fromInt_bits_uop_robIdx_value(stdExeUnits_1_io_fromInt_bits_uop_robIdx_value),
    .io_fromInt_bits_uop_sqIdx_flag(stdExeUnits_1_io_fromInt_bits_uop_sqIdx_flag),
    .io_fromInt_bits_uop_sqIdx_value(stdExeUnits_1_io_fromInt_bits_uop_sqIdx_value),
    .io_fromInt_bits_src_0(stdExeUnits_1_io_fromInt_bits_src_0),
    .io_out_valid(stdExeUnits_1_io_out_valid),
    .io_out_bits_uop_ctrl_fuType(stdExeUnits_1_io_out_bits_uop_ctrl_fuType),
    .io_out_bits_uop_ctrl_fuOpType(stdExeUnits_1_io_out_bits_uop_ctrl_fuOpType),
    .io_out_bits_uop_robIdx_flag(stdExeUnits_1_io_out_bits_uop_robIdx_flag),
    .io_out_bits_uop_robIdx_value(stdExeUnits_1_io_out_bits_uop_robIdx_value),
    .io_out_bits_uop_sqIdx_flag(stdExeUnits_1_io_out_bits_uop_sqIdx_flag),
    .io_out_bits_uop_sqIdx_value(stdExeUnits_1_io_out_bits_uop_sqIdx_value),
    .io_out_bits_data(stdExeUnits_1_io_out_bits_data)
  );
  CorrectTable correctTable ( // @[MemBlock.scala 144:28]
    .clock(correctTable_clock),
    .io_issue_0_req_addr(correctTable_io_issue_0_req_addr),
    .io_issue_0_resp_strict(correctTable_io_issue_0_resp_strict),
    .io_issue_1_req_addr(correctTable_io_issue_1_req_addr),
    .io_issue_1_resp_strict(correctTable_io_issue_1_resp_strict),
    .io_update_0_valid(correctTable_io_update_0_valid),
    .io_update_0_bits_addr(correctTable_io_update_0_bits_addr),
    .io_update_0_bits_strict(correctTable_io_update_0_bits_strict),
    .io_update_0_bits_violation(correctTable_io_update_0_bits_violation),
    .io_update_1_valid(correctTable_io_update_1_valid),
    .io_update_1_bits_addr(correctTable_io_update_1_bits_addr),
    .io_update_1_bits_strict(correctTable_io_update_1_bits_strict),
    .io_update_1_bits_violation(correctTable_io_update_1_bits_violation),
    .io_update_2_valid(correctTable_io_update_2_valid),
    .io_update_2_bits_addr(correctTable_io_update_2_bits_addr)
  );
  AtomicsUnit atomicsUnit ( // @[MemBlock.scala 174:27]
    .clock(atomicsUnit_clock),
    .reset(atomicsUnit_reset),
    .io_hartId(atomicsUnit_io_hartId),
    .io_in_ready(atomicsUnit_io_in_ready),
    .io_in_valid(atomicsUnit_io_in_valid),
    .io_in_bits_uop_cf_trigger_backendEn_0(atomicsUnit_io_in_bits_uop_cf_trigger_backendEn_0),
    .io_in_bits_uop_cf_trigger_backendEn_1(atomicsUnit_io_in_bits_uop_cf_trigger_backendEn_1),
    .io_in_bits_uop_ctrl_fuOpType(atomicsUnit_io_in_bits_uop_ctrl_fuOpType),
    .io_in_bits_uop_ctrl_rfWen(atomicsUnit_io_in_bits_uop_ctrl_rfWen),
    .io_in_bits_uop_ctrl_fpWen(atomicsUnit_io_in_bits_uop_ctrl_fpWen),
    .io_in_bits_uop_pdest(atomicsUnit_io_in_bits_uop_pdest),
    .io_in_bits_uop_robIdx_flag(atomicsUnit_io_in_bits_uop_robIdx_flag),
    .io_in_bits_uop_robIdx_value(atomicsUnit_io_in_bits_uop_robIdx_value),
    .io_in_bits_src_0(atomicsUnit_io_in_bits_src_0),
    .io_storeDataIn_valid(atomicsUnit_io_storeDataIn_valid),
    .io_storeDataIn_bits_data(atomicsUnit_io_storeDataIn_bits_data),
    .io_out_valid(atomicsUnit_io_out_valid),
    .io_out_bits_uop_cf_exceptionVec_4(atomicsUnit_io_out_bits_uop_cf_exceptionVec_4),
    .io_out_bits_uop_cf_exceptionVec_5(atomicsUnit_io_out_bits_uop_cf_exceptionVec_5),
    .io_out_bits_uop_cf_exceptionVec_6(atomicsUnit_io_out_bits_uop_cf_exceptionVec_6),
    .io_out_bits_uop_cf_exceptionVec_7(atomicsUnit_io_out_bits_uop_cf_exceptionVec_7),
    .io_out_bits_uop_cf_exceptionVec_13(atomicsUnit_io_out_bits_uop_cf_exceptionVec_13),
    .io_out_bits_uop_cf_exceptionVec_15(atomicsUnit_io_out_bits_uop_cf_exceptionVec_15),
    .io_out_bits_uop_cf_trigger_backendEn_0(atomicsUnit_io_out_bits_uop_cf_trigger_backendEn_0),
    .io_out_bits_uop_cf_trigger_backendEn_1(atomicsUnit_io_out_bits_uop_cf_trigger_backendEn_1),
    .io_out_bits_uop_cf_trigger_backendHit_0(atomicsUnit_io_out_bits_uop_cf_trigger_backendHit_0),
    .io_out_bits_uop_cf_trigger_backendHit_1(atomicsUnit_io_out_bits_uop_cf_trigger_backendHit_1),
    .io_out_bits_uop_cf_trigger_backendHit_2(atomicsUnit_io_out_bits_uop_cf_trigger_backendHit_2),
    .io_out_bits_uop_cf_trigger_backendHit_3(atomicsUnit_io_out_bits_uop_cf_trigger_backendHit_3),
    .io_out_bits_uop_cf_trigger_backendHit_4(atomicsUnit_io_out_bits_uop_cf_trigger_backendHit_4),
    .io_out_bits_uop_cf_trigger_backendHit_5(atomicsUnit_io_out_bits_uop_cf_trigger_backendHit_5),
    .io_out_bits_uop_ctrl_fuOpType(atomicsUnit_io_out_bits_uop_ctrl_fuOpType),
    .io_out_bits_uop_ctrl_rfWen(atomicsUnit_io_out_bits_uop_ctrl_rfWen),
    .io_out_bits_uop_ctrl_fpWen(atomicsUnit_io_out_bits_uop_ctrl_fpWen),
    .io_out_bits_uop_pdest(atomicsUnit_io_out_bits_uop_pdest),
    .io_out_bits_uop_robIdx_flag(atomicsUnit_io_out_bits_uop_robIdx_flag),
    .io_out_bits_uop_robIdx_value(atomicsUnit_io_out_bits_uop_robIdx_value),
    .io_out_bits_data(atomicsUnit_io_out_bits_data),
    .io_out_bits_debug_isMMIO(atomicsUnit_io_out_bits_debug_isMMIO),
    .io_dcache_req_ready(atomicsUnit_io_dcache_req_ready),
    .io_dcache_req_valid(atomicsUnit_io_dcache_req_valid),
    .io_dcache_req_bits_cmd(atomicsUnit_io_dcache_req_bits_cmd),
    .io_dcache_req_bits_vaddr(atomicsUnit_io_dcache_req_bits_vaddr),
    .io_dcache_req_bits_addr(atomicsUnit_io_dcache_req_bits_addr),
    .io_dcache_req_bits_word_idx(atomicsUnit_io_dcache_req_bits_word_idx),
    .io_dcache_req_bits_amo_data(atomicsUnit_io_dcache_req_bits_amo_data),
    .io_dcache_req_bits_amo_mask(atomicsUnit_io_dcache_req_bits_amo_mask),
    .io_dcache_resp_valid(atomicsUnit_io_dcache_resp_valid),
    .io_dcache_resp_bits_data(atomicsUnit_io_dcache_resp_bits_data),
    .io_dcache_resp_bits_miss(atomicsUnit_io_dcache_resp_bits_miss),
    .io_dcache_resp_bits_replay(atomicsUnit_io_dcache_resp_bits_replay),
    .io_dcache_resp_bits_error(atomicsUnit_io_dcache_resp_bits_error),
    .io_dcache_resp_bits_id(atomicsUnit_io_dcache_resp_bits_id),
    .io_dcache_block_lr(atomicsUnit_io_dcache_block_lr),
    .io_dtlb_req_valid(atomicsUnit_io_dtlb_req_valid),
    .io_dtlb_req_bits_vaddr(atomicsUnit_io_dtlb_req_bits_vaddr),
    .io_dtlb_req_bits_cmd(atomicsUnit_io_dtlb_req_bits_cmd),
    .io_dtlb_resp_ready(atomicsUnit_io_dtlb_resp_ready),
    .io_dtlb_resp_valid(atomicsUnit_io_dtlb_resp_valid),
    .io_dtlb_resp_bits_paddr_0(atomicsUnit_io_dtlb_resp_bits_paddr_0),
    .io_dtlb_resp_bits_miss(atomicsUnit_io_dtlb_resp_bits_miss),
    .io_dtlb_resp_bits_excp_0_pf_ld(atomicsUnit_io_dtlb_resp_bits_excp_0_pf_ld),
    .io_dtlb_resp_bits_excp_0_pf_st(atomicsUnit_io_dtlb_resp_bits_excp_0_pf_st),
    .io_dtlb_resp_bits_excp_0_af_ld(atomicsUnit_io_dtlb_resp_bits_excp_0_af_ld),
    .io_dtlb_resp_bits_excp_0_af_st(atomicsUnit_io_dtlb_resp_bits_excp_0_af_st),
    .io_dtlb_resp_bits_static_pm_valid(atomicsUnit_io_dtlb_resp_bits_static_pm_valid),
    .io_dtlb_resp_bits_static_pm_bits(atomicsUnit_io_dtlb_resp_bits_static_pm_bits),
    .io_pmpResp_ld(atomicsUnit_io_pmpResp_ld),
    .io_pmpResp_st(atomicsUnit_io_pmpResp_st),
    .io_pmpResp_mmio(atomicsUnit_io_pmpResp_mmio),
    .io_rsIdx(atomicsUnit_io_rsIdx),
    .io_flush_sbuffer_valid(atomicsUnit_io_flush_sbuffer_valid),
    .io_flush_sbuffer_empty(atomicsUnit_io_flush_sbuffer_empty),
    .io_feedbackSlow_valid(atomicsUnit_io_feedbackSlow_valid),
    .io_feedbackSlow_bits_rsIdx(atomicsUnit_io_feedbackSlow_bits_rsIdx),
    .io_redirect_valid(atomicsUnit_io_redirect_valid),
    .io_exceptionAddr_valid(atomicsUnit_io_exceptionAddr_valid),
    .io_exceptionAddr_bits(atomicsUnit_io_exceptionAddr_bits),
    .io_csrCtrl_cache_error_enable(atomicsUnit_io_csrCtrl_cache_error_enable),
    .io_csrCtrl_mem_trigger_t_valid(atomicsUnit_io_csrCtrl_mem_trigger_t_valid),
    .io_csrCtrl_mem_trigger_t_bits_addr(atomicsUnit_io_csrCtrl_mem_trigger_t_bits_addr),
    .io_csrCtrl_mem_trigger_t_bits_tdata_matchType(atomicsUnit_io_csrCtrl_mem_trigger_t_bits_tdata_matchType),
    .io_csrCtrl_mem_trigger_t_bits_tdata_select(atomicsUnit_io_csrCtrl_mem_trigger_t_bits_tdata_select),
    .io_csrCtrl_mem_trigger_t_bits_tdata_chain(atomicsUnit_io_csrCtrl_mem_trigger_t_bits_tdata_chain),
    .io_csrCtrl_mem_trigger_t_bits_tdata_tdata2(atomicsUnit_io_csrCtrl_mem_trigger_t_bits_tdata_tdata2),
    .io_csrCtrl_trigger_enable_2(atomicsUnit_io_csrCtrl_trigger_enable_2),
    .io_csrCtrl_trigger_enable_3(atomicsUnit_io_csrCtrl_trigger_enable_3),
    .io_csrCtrl_trigger_enable_4(atomicsUnit_io_csrCtrl_trigger_enable_4),
    .io_csrCtrl_trigger_enable_5(atomicsUnit_io_csrCtrl_trigger_enable_5),
    .io_csrCtrl_trigger_enable_7(atomicsUnit_io_csrCtrl_trigger_enable_7),
    .io_csrCtrl_trigger_enable_9(atomicsUnit_io_csrCtrl_trigger_enable_9)
  );
  VlflowQueue vlflowqueue ( // @[MemBlock.scala 226:27]
    .clock(vlflowqueue_clock),
    .reset(vlflowqueue_reset),
    .io_loadRegIn_0_valid(vlflowqueue_io_loadRegIn_0_valid),
    .io_loadRegIn_0_bits_uop_robIdx_value(vlflowqueue_io_loadRegIn_0_bits_uop_robIdx_value),
    .io_loadRegIn_0_bits_baseaddr(vlflowqueue_io_loadRegIn_0_bits_baseaddr),
    .io_loadRegIn_1_valid(vlflowqueue_io_loadRegIn_1_valid),
    .io_loadRegIn_1_bits_uop_robIdx_value(vlflowqueue_io_loadRegIn_1_bits_uop_robIdx_value),
    .io_loadRegIn_1_bits_baseaddr(vlflowqueue_io_loadRegIn_1_bits_baseaddr),
    .io_loadPipeOut_0_ready(vlflowqueue_io_loadPipeOut_0_ready),
    .io_loadPipeOut_0_valid(vlflowqueue_io_loadPipeOut_0_valid),
    .io_loadPipeOut_0_bits_vaddr(vlflowqueue_io_loadPipeOut_0_bits_vaddr),
    .io_loadPipeOut_1_ready(vlflowqueue_io_loadPipeOut_1_ready),
    .io_loadPipeOut_1_valid(vlflowqueue_io_loadPipeOut_1_valid),
    .io_loadPipeOut_1_bits_vaddr(vlflowqueue_io_loadPipeOut_1_bits_vaddr)
  );
  VlExcSignal vlExcSignal ( // @[MemBlock.scala 228:27]
    .clock(vlExcSignal_clock),
    .reset(vlExcSignal_reset),
    .io_vecloadRegIn_0_valid(vlExcSignal_io_vecloadRegIn_0_valid),
    .io_vecloadRegIn_0_bits_uop_robIdx_value(vlExcSignal_io_vecloadRegIn_0_bits_uop_robIdx_value),
    .io_vecloadRegIn_0_bits_baseaddr(vlExcSignal_io_vecloadRegIn_0_bits_baseaddr),
    .io_vecloadRegIn_1_valid(vlExcSignal_io_vecloadRegIn_1_valid),
    .io_vecloadRegIn_1_bits_uop_robIdx_value(vlExcSignal_io_vecloadRegIn_1_bits_uop_robIdx_value),
    .io_vecloadRegIn_1_bits_baseaddr(vlExcSignal_io_vecloadRegIn_1_bits_baseaddr)
  );
  LsqWrapper lsq ( // @[MemBlock.scala 231:23]
    .clock(lsq_clock),
    .reset(lsq_reset),
    .io_brqRedirect_valid(lsq_io_brqRedirect_valid),
    .io_brqRedirect_bits_robIdx_flag(lsq_io_brqRedirect_bits_robIdx_flag),
    .io_brqRedirect_bits_robIdx_value(lsq_io_brqRedirect_bits_robIdx_value),
    .io_brqRedirect_bits_level(lsq_io_brqRedirect_bits_level),
    .io_enq_needAlloc_0(lsq_io_enq_needAlloc_0),
    .io_enq_needAlloc_1(lsq_io_enq_needAlloc_1),
    .io_enq_needAlloc_2(lsq_io_enq_needAlloc_2),
    .io_enq_needAlloc_3(lsq_io_enq_needAlloc_3),
    .io_enq_req_0_valid(lsq_io_enq_req_0_valid),
    .io_enq_req_0_bits_cf_trigger_backendEn_0(lsq_io_enq_req_0_bits_cf_trigger_backendEn_0),
    .io_enq_req_0_bits_cf_trigger_backendEn_1(lsq_io_enq_req_0_bits_cf_trigger_backendEn_1),
    .io_enq_req_0_bits_ctrl_fuOpType(lsq_io_enq_req_0_bits_ctrl_fuOpType),
    .io_enq_req_0_bits_ctrl_rfWen(lsq_io_enq_req_0_bits_ctrl_rfWen),
    .io_enq_req_0_bits_ctrl_fpWen(lsq_io_enq_req_0_bits_ctrl_fpWen),
    .io_enq_req_0_bits_ctrl_flushPipe(lsq_io_enq_req_0_bits_ctrl_flushPipe),
    .io_enq_req_0_bits_ctrl_replayInst(lsq_io_enq_req_0_bits_ctrl_replayInst),
    .io_enq_req_0_bits_pdest(lsq_io_enq_req_0_bits_pdest),
    .io_enq_req_0_bits_robIdx_flag(lsq_io_enq_req_0_bits_robIdx_flag),
    .io_enq_req_0_bits_robIdx_value(lsq_io_enq_req_0_bits_robIdx_value),
    .io_enq_req_0_bits_lqIdx_value(lsq_io_enq_req_0_bits_lqIdx_value),
    .io_enq_req_0_bits_sqIdx_value(lsq_io_enq_req_0_bits_sqIdx_value),
    .io_enq_req_1_valid(lsq_io_enq_req_1_valid),
    .io_enq_req_1_bits_cf_trigger_backendEn_0(lsq_io_enq_req_1_bits_cf_trigger_backendEn_0),
    .io_enq_req_1_bits_cf_trigger_backendEn_1(lsq_io_enq_req_1_bits_cf_trigger_backendEn_1),
    .io_enq_req_1_bits_ctrl_fuOpType(lsq_io_enq_req_1_bits_ctrl_fuOpType),
    .io_enq_req_1_bits_ctrl_rfWen(lsq_io_enq_req_1_bits_ctrl_rfWen),
    .io_enq_req_1_bits_ctrl_fpWen(lsq_io_enq_req_1_bits_ctrl_fpWen),
    .io_enq_req_1_bits_ctrl_flushPipe(lsq_io_enq_req_1_bits_ctrl_flushPipe),
    .io_enq_req_1_bits_ctrl_replayInst(lsq_io_enq_req_1_bits_ctrl_replayInst),
    .io_enq_req_1_bits_pdest(lsq_io_enq_req_1_bits_pdest),
    .io_enq_req_1_bits_robIdx_flag(lsq_io_enq_req_1_bits_robIdx_flag),
    .io_enq_req_1_bits_robIdx_value(lsq_io_enq_req_1_bits_robIdx_value),
    .io_enq_req_1_bits_lqIdx_value(lsq_io_enq_req_1_bits_lqIdx_value),
    .io_enq_req_1_bits_sqIdx_value(lsq_io_enq_req_1_bits_sqIdx_value),
    .io_enq_req_2_valid(lsq_io_enq_req_2_valid),
    .io_enq_req_2_bits_cf_trigger_backendEn_0(lsq_io_enq_req_2_bits_cf_trigger_backendEn_0),
    .io_enq_req_2_bits_cf_trigger_backendEn_1(lsq_io_enq_req_2_bits_cf_trigger_backendEn_1),
    .io_enq_req_2_bits_ctrl_fuOpType(lsq_io_enq_req_2_bits_ctrl_fuOpType),
    .io_enq_req_2_bits_ctrl_rfWen(lsq_io_enq_req_2_bits_ctrl_rfWen),
    .io_enq_req_2_bits_ctrl_fpWen(lsq_io_enq_req_2_bits_ctrl_fpWen),
    .io_enq_req_2_bits_ctrl_flushPipe(lsq_io_enq_req_2_bits_ctrl_flushPipe),
    .io_enq_req_2_bits_ctrl_replayInst(lsq_io_enq_req_2_bits_ctrl_replayInst),
    .io_enq_req_2_bits_pdest(lsq_io_enq_req_2_bits_pdest),
    .io_enq_req_2_bits_robIdx_flag(lsq_io_enq_req_2_bits_robIdx_flag),
    .io_enq_req_2_bits_robIdx_value(lsq_io_enq_req_2_bits_robIdx_value),
    .io_enq_req_2_bits_lqIdx_value(lsq_io_enq_req_2_bits_lqIdx_value),
    .io_enq_req_2_bits_sqIdx_value(lsq_io_enq_req_2_bits_sqIdx_value),
    .io_enq_req_3_valid(lsq_io_enq_req_3_valid),
    .io_enq_req_3_bits_cf_trigger_backendEn_0(lsq_io_enq_req_3_bits_cf_trigger_backendEn_0),
    .io_enq_req_3_bits_cf_trigger_backendEn_1(lsq_io_enq_req_3_bits_cf_trigger_backendEn_1),
    .io_enq_req_3_bits_ctrl_fuOpType(lsq_io_enq_req_3_bits_ctrl_fuOpType),
    .io_enq_req_3_bits_ctrl_rfWen(lsq_io_enq_req_3_bits_ctrl_rfWen),
    .io_enq_req_3_bits_ctrl_fpWen(lsq_io_enq_req_3_bits_ctrl_fpWen),
    .io_enq_req_3_bits_ctrl_flushPipe(lsq_io_enq_req_3_bits_ctrl_flushPipe),
    .io_enq_req_3_bits_ctrl_replayInst(lsq_io_enq_req_3_bits_ctrl_replayInst),
    .io_enq_req_3_bits_pdest(lsq_io_enq_req_3_bits_pdest),
    .io_enq_req_3_bits_robIdx_flag(lsq_io_enq_req_3_bits_robIdx_flag),
    .io_enq_req_3_bits_robIdx_value(lsq_io_enq_req_3_bits_robIdx_value),
    .io_enq_req_3_bits_lqIdx_value(lsq_io_enq_req_3_bits_lqIdx_value),
    .io_enq_req_3_bits_sqIdx_value(lsq_io_enq_req_3_bits_sqIdx_value),
    .io_ldu_s2_storeLoadViolationQuery_0_req_valid(lsq_io_ldu_s2_storeLoadViolationQuery_0_req_valid),
    .io_ldu_s2_storeLoadViolationQuery_0_req_bits_uop_cf_foldpc(
      lsq_io_ldu_s2_storeLoadViolationQuery_0_req_bits_uop_cf_foldpc),
    .io_ldu_s2_storeLoadViolationQuery_0_req_bits_uop_cf_ftqPtr_flag(
      lsq_io_ldu_s2_storeLoadViolationQuery_0_req_bits_uop_cf_ftqPtr_flag),
    .io_ldu_s2_storeLoadViolationQuery_0_req_bits_uop_cf_ftqPtr_value(
      lsq_io_ldu_s2_storeLoadViolationQuery_0_req_bits_uop_cf_ftqPtr_value),
    .io_ldu_s2_storeLoadViolationQuery_0_req_bits_uop_cf_ftqOffset(
      lsq_io_ldu_s2_storeLoadViolationQuery_0_req_bits_uop_cf_ftqOffset),
    .io_ldu_s2_storeLoadViolationQuery_0_req_bits_uop_robIdx_flag(
      lsq_io_ldu_s2_storeLoadViolationQuery_0_req_bits_uop_robIdx_flag),
    .io_ldu_s2_storeLoadViolationQuery_0_req_bits_uop_robIdx_value(
      lsq_io_ldu_s2_storeLoadViolationQuery_0_req_bits_uop_robIdx_value),
    .io_ldu_s2_storeLoadViolationQuery_0_req_bits_uop_sqIdx_flag(
      lsq_io_ldu_s2_storeLoadViolationQuery_0_req_bits_uop_sqIdx_flag),
    .io_ldu_s2_storeLoadViolationQuery_0_req_bits_uop_sqIdx_value(
      lsq_io_ldu_s2_storeLoadViolationQuery_0_req_bits_uop_sqIdx_value),
    .io_ldu_s2_storeLoadViolationQuery_0_req_bits_index(lsq_io_ldu_s2_storeLoadViolationQuery_0_req_bits_index),
    .io_ldu_s2_storeLoadViolationQuery_0_req_bits_allocated(lsq_io_ldu_s2_storeLoadViolationQuery_0_req_bits_allocated),
    .io_ldu_s2_storeLoadViolationQuery_0_req_bits_datavalid(lsq_io_ldu_s2_storeLoadViolationQuery_0_req_bits_datavalid),
    .io_ldu_s2_storeLoadViolationQuery_0_req_bits_mask(lsq_io_ldu_s2_storeLoadViolationQuery_0_req_bits_mask),
    .io_ldu_s2_storeLoadViolationQuery_0_req_bits_paddr(lsq_io_ldu_s2_storeLoadViolationQuery_0_req_bits_paddr),
    .io_ldu_s2_storeLoadViolationQuery_0_resp_bits_index(lsq_io_ldu_s2_storeLoadViolationQuery_0_resp_bits_index),
    .io_ldu_s2_storeLoadViolationQuery_0_resp_bits_canAccept(lsq_io_ldu_s2_storeLoadViolationQuery_0_resp_bits_canAccept
      ),
    .io_ldu_s2_storeLoadViolationQuery_0_resp_bits_allocated(lsq_io_ldu_s2_storeLoadViolationQuery_0_resp_bits_allocated
      ),
    .io_ldu_s2_storeLoadViolationQuery_1_req_valid(lsq_io_ldu_s2_storeLoadViolationQuery_1_req_valid),
    .io_ldu_s2_storeLoadViolationQuery_1_req_bits_uop_cf_foldpc(
      lsq_io_ldu_s2_storeLoadViolationQuery_1_req_bits_uop_cf_foldpc),
    .io_ldu_s2_storeLoadViolationQuery_1_req_bits_uop_cf_ftqPtr_flag(
      lsq_io_ldu_s2_storeLoadViolationQuery_1_req_bits_uop_cf_ftqPtr_flag),
    .io_ldu_s2_storeLoadViolationQuery_1_req_bits_uop_cf_ftqPtr_value(
      lsq_io_ldu_s2_storeLoadViolationQuery_1_req_bits_uop_cf_ftqPtr_value),
    .io_ldu_s2_storeLoadViolationQuery_1_req_bits_uop_cf_ftqOffset(
      lsq_io_ldu_s2_storeLoadViolationQuery_1_req_bits_uop_cf_ftqOffset),
    .io_ldu_s2_storeLoadViolationQuery_1_req_bits_uop_robIdx_flag(
      lsq_io_ldu_s2_storeLoadViolationQuery_1_req_bits_uop_robIdx_flag),
    .io_ldu_s2_storeLoadViolationQuery_1_req_bits_uop_robIdx_value(
      lsq_io_ldu_s2_storeLoadViolationQuery_1_req_bits_uop_robIdx_value),
    .io_ldu_s2_storeLoadViolationQuery_1_req_bits_uop_sqIdx_flag(
      lsq_io_ldu_s2_storeLoadViolationQuery_1_req_bits_uop_sqIdx_flag),
    .io_ldu_s2_storeLoadViolationQuery_1_req_bits_uop_sqIdx_value(
      lsq_io_ldu_s2_storeLoadViolationQuery_1_req_bits_uop_sqIdx_value),
    .io_ldu_s2_storeLoadViolationQuery_1_req_bits_index(lsq_io_ldu_s2_storeLoadViolationQuery_1_req_bits_index),
    .io_ldu_s2_storeLoadViolationQuery_1_req_bits_allocated(lsq_io_ldu_s2_storeLoadViolationQuery_1_req_bits_allocated),
    .io_ldu_s2_storeLoadViolationQuery_1_req_bits_datavalid(lsq_io_ldu_s2_storeLoadViolationQuery_1_req_bits_datavalid),
    .io_ldu_s2_storeLoadViolationQuery_1_req_bits_mask(lsq_io_ldu_s2_storeLoadViolationQuery_1_req_bits_mask),
    .io_ldu_s2_storeLoadViolationQuery_1_req_bits_paddr(lsq_io_ldu_s2_storeLoadViolationQuery_1_req_bits_paddr),
    .io_ldu_s2_storeLoadViolationQuery_1_resp_bits_index(lsq_io_ldu_s2_storeLoadViolationQuery_1_resp_bits_index),
    .io_ldu_s2_storeLoadViolationQuery_1_resp_bits_canAccept(lsq_io_ldu_s2_storeLoadViolationQuery_1_resp_bits_canAccept
      ),
    .io_ldu_s2_storeLoadViolationQuery_1_resp_bits_allocated(lsq_io_ldu_s2_storeLoadViolationQuery_1_resp_bits_allocated
      ),
    .io_ldu_s2_loadLoadViolationQuery_0_req_valid(lsq_io_ldu_s2_loadLoadViolationQuery_0_req_valid),
    .io_ldu_s2_loadLoadViolationQuery_0_req_bits_uop_robIdx_flag(
      lsq_io_ldu_s2_loadLoadViolationQuery_0_req_bits_uop_robIdx_flag),
    .io_ldu_s2_loadLoadViolationQuery_0_req_bits_uop_robIdx_value(
      lsq_io_ldu_s2_loadLoadViolationQuery_0_req_bits_uop_robIdx_value),
    .io_ldu_s2_loadLoadViolationQuery_0_req_bits_uop_lqIdx_flag(
      lsq_io_ldu_s2_loadLoadViolationQuery_0_req_bits_uop_lqIdx_flag),
    .io_ldu_s2_loadLoadViolationQuery_0_req_bits_uop_lqIdx_value(
      lsq_io_ldu_s2_loadLoadViolationQuery_0_req_bits_uop_lqIdx_value),
    .io_ldu_s2_loadLoadViolationQuery_0_req_bits_index(lsq_io_ldu_s2_loadLoadViolationQuery_0_req_bits_index),
    .io_ldu_s2_loadLoadViolationQuery_0_req_bits_allocated(lsq_io_ldu_s2_loadLoadViolationQuery_0_req_bits_allocated),
    .io_ldu_s2_loadLoadViolationQuery_0_req_bits_datavalid(lsq_io_ldu_s2_loadLoadViolationQuery_0_req_bits_datavalid),
    .io_ldu_s2_loadLoadViolationQuery_0_req_bits_miss(lsq_io_ldu_s2_loadLoadViolationQuery_0_req_bits_miss),
    .io_ldu_s2_loadLoadViolationQuery_0_req_bits_paddr(lsq_io_ldu_s2_loadLoadViolationQuery_0_req_bits_paddr),
    .io_ldu_s2_loadLoadViolationQuery_0_resp_valid(lsq_io_ldu_s2_loadLoadViolationQuery_0_resp_valid),
    .io_ldu_s2_loadLoadViolationQuery_0_resp_bits_index(lsq_io_ldu_s2_loadLoadViolationQuery_0_resp_bits_index),
    .io_ldu_s2_loadLoadViolationQuery_0_resp_bits_canAccept(lsq_io_ldu_s2_loadLoadViolationQuery_0_resp_bits_canAccept),
    .io_ldu_s2_loadLoadViolationQuery_0_resp_bits_allocated(lsq_io_ldu_s2_loadLoadViolationQuery_0_resp_bits_allocated),
    .io_ldu_s2_loadLoadViolationQuery_0_resp_bits_replayFromFetch(
      lsq_io_ldu_s2_loadLoadViolationQuery_0_resp_bits_replayFromFetch),
    .io_ldu_s2_loadLoadViolationQuery_1_req_valid(lsq_io_ldu_s2_loadLoadViolationQuery_1_req_valid),
    .io_ldu_s2_loadLoadViolationQuery_1_req_bits_uop_robIdx_flag(
      lsq_io_ldu_s2_loadLoadViolationQuery_1_req_bits_uop_robIdx_flag),
    .io_ldu_s2_loadLoadViolationQuery_1_req_bits_uop_robIdx_value(
      lsq_io_ldu_s2_loadLoadViolationQuery_1_req_bits_uop_robIdx_value),
    .io_ldu_s2_loadLoadViolationQuery_1_req_bits_uop_lqIdx_flag(
      lsq_io_ldu_s2_loadLoadViolationQuery_1_req_bits_uop_lqIdx_flag),
    .io_ldu_s2_loadLoadViolationQuery_1_req_bits_uop_lqIdx_value(
      lsq_io_ldu_s2_loadLoadViolationQuery_1_req_bits_uop_lqIdx_value),
    .io_ldu_s2_loadLoadViolationQuery_1_req_bits_index(lsq_io_ldu_s2_loadLoadViolationQuery_1_req_bits_index),
    .io_ldu_s2_loadLoadViolationQuery_1_req_bits_allocated(lsq_io_ldu_s2_loadLoadViolationQuery_1_req_bits_allocated),
    .io_ldu_s2_loadLoadViolationQuery_1_req_bits_datavalid(lsq_io_ldu_s2_loadLoadViolationQuery_1_req_bits_datavalid),
    .io_ldu_s2_loadLoadViolationQuery_1_req_bits_miss(lsq_io_ldu_s2_loadLoadViolationQuery_1_req_bits_miss),
    .io_ldu_s2_loadLoadViolationQuery_1_req_bits_paddr(lsq_io_ldu_s2_loadLoadViolationQuery_1_req_bits_paddr),
    .io_ldu_s2_loadLoadViolationQuery_1_resp_valid(lsq_io_ldu_s2_loadLoadViolationQuery_1_resp_valid),
    .io_ldu_s2_loadLoadViolationQuery_1_resp_bits_index(lsq_io_ldu_s2_loadLoadViolationQuery_1_resp_bits_index),
    .io_ldu_s2_loadLoadViolationQuery_1_resp_bits_canAccept(lsq_io_ldu_s2_loadLoadViolationQuery_1_resp_bits_canAccept),
    .io_ldu_s2_loadLoadViolationQuery_1_resp_bits_allocated(lsq_io_ldu_s2_loadLoadViolationQuery_1_resp_bits_allocated),
    .io_ldu_s2_loadLoadViolationQuery_1_resp_bits_replayFromFetch(
      lsq_io_ldu_s2_loadLoadViolationQuery_1_resp_bits_replayFromFetch),
    .io_ldu_s3_loadIn_0_valid(lsq_io_ldu_s3_loadIn_0_valid),
    .io_ldu_s3_loadIn_0_bits_uop_cf_foldpc(lsq_io_ldu_s3_loadIn_0_bits_uop_cf_foldpc),
    .io_ldu_s3_loadIn_0_bits_uop_cf_exceptionVec_4(lsq_io_ldu_s3_loadIn_0_bits_uop_cf_exceptionVec_4),
    .io_ldu_s3_loadIn_0_bits_uop_cf_exceptionVec_5(lsq_io_ldu_s3_loadIn_0_bits_uop_cf_exceptionVec_5),
    .io_ldu_s3_loadIn_0_bits_uop_cf_exceptionVec_13(lsq_io_ldu_s3_loadIn_0_bits_uop_cf_exceptionVec_13),
    .io_ldu_s3_loadIn_0_bits_uop_cf_trigger_backendEn_1(lsq_io_ldu_s3_loadIn_0_bits_uop_cf_trigger_backendEn_1),
    .io_ldu_s3_loadIn_0_bits_uop_cf_trigger_backendHit_0(lsq_io_ldu_s3_loadIn_0_bits_uop_cf_trigger_backendHit_0),
    .io_ldu_s3_loadIn_0_bits_uop_cf_trigger_backendHit_1(lsq_io_ldu_s3_loadIn_0_bits_uop_cf_trigger_backendHit_1),
    .io_ldu_s3_loadIn_0_bits_uop_cf_trigger_backendHit_4(lsq_io_ldu_s3_loadIn_0_bits_uop_cf_trigger_backendHit_4),
    .io_ldu_s3_loadIn_0_bits_uop_cf_waitForRobIdx_flag(lsq_io_ldu_s3_loadIn_0_bits_uop_cf_waitForRobIdx_flag),
    .io_ldu_s3_loadIn_0_bits_uop_cf_waitForRobIdx_value(lsq_io_ldu_s3_loadIn_0_bits_uop_cf_waitForRobIdx_value),
    .io_ldu_s3_loadIn_0_bits_uop_cf_loadWaitBit(lsq_io_ldu_s3_loadIn_0_bits_uop_cf_loadWaitBit),
    .io_ldu_s3_loadIn_0_bits_uop_cf_loadWaitStrict(lsq_io_ldu_s3_loadIn_0_bits_uop_cf_loadWaitStrict),
    .io_ldu_s3_loadIn_0_bits_uop_cf_ftqPtr_flag(lsq_io_ldu_s3_loadIn_0_bits_uop_cf_ftqPtr_flag),
    .io_ldu_s3_loadIn_0_bits_uop_cf_ftqPtr_value(lsq_io_ldu_s3_loadIn_0_bits_uop_cf_ftqPtr_value),
    .io_ldu_s3_loadIn_0_bits_uop_cf_ftqOffset(lsq_io_ldu_s3_loadIn_0_bits_uop_cf_ftqOffset),
    .io_ldu_s3_loadIn_0_bits_uop_ctrl_fuType(lsq_io_ldu_s3_loadIn_0_bits_uop_ctrl_fuType),
    .io_ldu_s3_loadIn_0_bits_uop_ctrl_fuOpType(lsq_io_ldu_s3_loadIn_0_bits_uop_ctrl_fuOpType),
    .io_ldu_s3_loadIn_0_bits_uop_ctrl_rfWen(lsq_io_ldu_s3_loadIn_0_bits_uop_ctrl_rfWen),
    .io_ldu_s3_loadIn_0_bits_uop_ctrl_fpWen(lsq_io_ldu_s3_loadIn_0_bits_uop_ctrl_fpWen),
    .io_ldu_s3_loadIn_0_bits_uop_ctrl_replayInst(lsq_io_ldu_s3_loadIn_0_bits_uop_ctrl_replayInst),
    .io_ldu_s3_loadIn_0_bits_uop_pdest(lsq_io_ldu_s3_loadIn_0_bits_uop_pdest),
    .io_ldu_s3_loadIn_0_bits_uop_robIdx_flag(lsq_io_ldu_s3_loadIn_0_bits_uop_robIdx_flag),
    .io_ldu_s3_loadIn_0_bits_uop_robIdx_value(lsq_io_ldu_s3_loadIn_0_bits_uop_robIdx_value),
    .io_ldu_s3_loadIn_0_bits_uop_lqIdx_flag(lsq_io_ldu_s3_loadIn_0_bits_uop_lqIdx_flag),
    .io_ldu_s3_loadIn_0_bits_uop_lqIdx_value(lsq_io_ldu_s3_loadIn_0_bits_uop_lqIdx_value),
    .io_ldu_s3_loadIn_0_bits_uop_sqIdx_flag(lsq_io_ldu_s3_loadIn_0_bits_uop_sqIdx_flag),
    .io_ldu_s3_loadIn_0_bits_uop_sqIdx_value(lsq_io_ldu_s3_loadIn_0_bits_uop_sqIdx_value),
    .io_ldu_s3_loadIn_0_bits_vaddr(lsq_io_ldu_s3_loadIn_0_bits_vaddr),
    .io_ldu_s3_loadIn_0_bits_paddr(lsq_io_ldu_s3_loadIn_0_bits_paddr),
    .io_ldu_s3_loadIn_0_bits_mask(lsq_io_ldu_s3_loadIn_0_bits_mask),
    .io_ldu_s3_loadIn_0_bits_miss(lsq_io_ldu_s3_loadIn_0_bits_miss),
    .io_ldu_s3_loadIn_0_bits_tlbMiss(lsq_io_ldu_s3_loadIn_0_bits_tlbMiss),
    .io_ldu_s3_loadIn_0_bits_mmio(lsq_io_ldu_s3_loadIn_0_bits_mmio),
    .io_ldu_s3_loadIn_0_bits_rarAllocated(lsq_io_ldu_s3_loadIn_0_bits_rarAllocated),
    .io_ldu_s3_loadIn_0_bits_rarIndex(lsq_io_ldu_s3_loadIn_0_bits_rarIndex),
    .io_ldu_s3_loadIn_0_bits_rawAllocated(lsq_io_ldu_s3_loadIn_0_bits_rawAllocated),
    .io_ldu_s3_loadIn_0_bits_rawIndex(lsq_io_ldu_s3_loadIn_0_bits_rawIndex),
    .io_ldu_s3_loadIn_0_bits_replayInfo_missMSHRId(lsq_io_ldu_s3_loadIn_0_bits_replayInfo_missMSHRId),
    .io_ldu_s3_loadIn_0_bits_replayInfo_canForwardFullData(lsq_io_ldu_s3_loadIn_0_bits_replayInfo_canForwardFullData),
    .io_ldu_s3_loadIn_0_bits_replayInfo_dataInvalidSqIdx_flag(
      lsq_io_ldu_s3_loadIn_0_bits_replayInfo_dataInvalidSqIdx_flag),
    .io_ldu_s3_loadIn_0_bits_replayInfo_dataInvalidSqIdx_value(
      lsq_io_ldu_s3_loadIn_0_bits_replayInfo_dataInvalidSqIdx_value),
    .io_ldu_s3_loadIn_0_bits_replayInfo_addrInvalidSqIdx_flag(
      lsq_io_ldu_s3_loadIn_0_bits_replayInfo_addrInvalidSqIdx_flag),
    .io_ldu_s3_loadIn_0_bits_replayInfo_addrInvalidSqIdx_value(
      lsq_io_ldu_s3_loadIn_0_bits_replayInfo_addrInvalidSqIdx_value),
    .io_ldu_s3_loadIn_0_bits_replayInfo_replayCarry_real_way_en(
      lsq_io_ldu_s3_loadIn_0_bits_replayInfo_replayCarry_real_way_en),
    .io_ldu_s3_loadIn_0_bits_replayInfo_replayCarry_valid(lsq_io_ldu_s3_loadIn_0_bits_replayInfo_replayCarry_valid),
    .io_ldu_s3_loadIn_0_bits_replayInfo_dataInLastBeat(lsq_io_ldu_s3_loadIn_0_bits_replayInfo_dataInLastBeat),
    .io_ldu_s3_loadIn_0_bits_replayInfo_cause_0(lsq_io_ldu_s3_loadIn_0_bits_replayInfo_cause_0),
    .io_ldu_s3_loadIn_0_bits_replayInfo_cause_1(lsq_io_ldu_s3_loadIn_0_bits_replayInfo_cause_1),
    .io_ldu_s3_loadIn_0_bits_replayInfo_cause_2(lsq_io_ldu_s3_loadIn_0_bits_replayInfo_cause_2),
    .io_ldu_s3_loadIn_0_bits_replayInfo_cause_3(lsq_io_ldu_s3_loadIn_0_bits_replayInfo_cause_3),
    .io_ldu_s3_loadIn_0_bits_replayInfo_cause_4(lsq_io_ldu_s3_loadIn_0_bits_replayInfo_cause_4),
    .io_ldu_s3_loadIn_0_bits_replayInfo_cause_5(lsq_io_ldu_s3_loadIn_0_bits_replayInfo_cause_5),
    .io_ldu_s3_loadIn_0_bits_replayInfo_cause_6(lsq_io_ldu_s3_loadIn_0_bits_replayInfo_cause_6),
    .io_ldu_s3_loadIn_0_bits_replayInfo_cause_7(lsq_io_ldu_s3_loadIn_0_bits_replayInfo_cause_7),
    .io_ldu_s3_loadIn_0_bits_lqDataWenDup_1(lsq_io_ldu_s3_loadIn_0_bits_lqDataWenDup_1),
    .io_ldu_s3_loadIn_0_bits_lqDataWenDup_2(lsq_io_ldu_s3_loadIn_0_bits_lqDataWenDup_2),
    .io_ldu_s3_loadIn_0_bits_lqDataWenDup_3(lsq_io_ldu_s3_loadIn_0_bits_lqDataWenDup_3),
    .io_ldu_s3_loadIn_0_bits_lqDataWenDup_5(lsq_io_ldu_s3_loadIn_0_bits_lqDataWenDup_5),
    .io_ldu_s3_loadIn_1_valid(lsq_io_ldu_s3_loadIn_1_valid),
    .io_ldu_s3_loadIn_1_bits_uop_cf_foldpc(lsq_io_ldu_s3_loadIn_1_bits_uop_cf_foldpc),
    .io_ldu_s3_loadIn_1_bits_uop_cf_exceptionVec_4(lsq_io_ldu_s3_loadIn_1_bits_uop_cf_exceptionVec_4),
    .io_ldu_s3_loadIn_1_bits_uop_cf_exceptionVec_5(lsq_io_ldu_s3_loadIn_1_bits_uop_cf_exceptionVec_5),
    .io_ldu_s3_loadIn_1_bits_uop_cf_exceptionVec_13(lsq_io_ldu_s3_loadIn_1_bits_uop_cf_exceptionVec_13),
    .io_ldu_s3_loadIn_1_bits_uop_cf_trigger_backendEn_1(lsq_io_ldu_s3_loadIn_1_bits_uop_cf_trigger_backendEn_1),
    .io_ldu_s3_loadIn_1_bits_uop_cf_trigger_backendHit_0(lsq_io_ldu_s3_loadIn_1_bits_uop_cf_trigger_backendHit_0),
    .io_ldu_s3_loadIn_1_bits_uop_cf_trigger_backendHit_1(lsq_io_ldu_s3_loadIn_1_bits_uop_cf_trigger_backendHit_1),
    .io_ldu_s3_loadIn_1_bits_uop_cf_trigger_backendHit_4(lsq_io_ldu_s3_loadIn_1_bits_uop_cf_trigger_backendHit_4),
    .io_ldu_s3_loadIn_1_bits_uop_cf_waitForRobIdx_flag(lsq_io_ldu_s3_loadIn_1_bits_uop_cf_waitForRobIdx_flag),
    .io_ldu_s3_loadIn_1_bits_uop_cf_waitForRobIdx_value(lsq_io_ldu_s3_loadIn_1_bits_uop_cf_waitForRobIdx_value),
    .io_ldu_s3_loadIn_1_bits_uop_cf_loadWaitBit(lsq_io_ldu_s3_loadIn_1_bits_uop_cf_loadWaitBit),
    .io_ldu_s3_loadIn_1_bits_uop_cf_loadWaitStrict(lsq_io_ldu_s3_loadIn_1_bits_uop_cf_loadWaitStrict),
    .io_ldu_s3_loadIn_1_bits_uop_cf_ftqPtr_flag(lsq_io_ldu_s3_loadIn_1_bits_uop_cf_ftqPtr_flag),
    .io_ldu_s3_loadIn_1_bits_uop_cf_ftqPtr_value(lsq_io_ldu_s3_loadIn_1_bits_uop_cf_ftqPtr_value),
    .io_ldu_s3_loadIn_1_bits_uop_cf_ftqOffset(lsq_io_ldu_s3_loadIn_1_bits_uop_cf_ftqOffset),
    .io_ldu_s3_loadIn_1_bits_uop_ctrl_fuType(lsq_io_ldu_s3_loadIn_1_bits_uop_ctrl_fuType),
    .io_ldu_s3_loadIn_1_bits_uop_ctrl_fuOpType(lsq_io_ldu_s3_loadIn_1_bits_uop_ctrl_fuOpType),
    .io_ldu_s3_loadIn_1_bits_uop_ctrl_rfWen(lsq_io_ldu_s3_loadIn_1_bits_uop_ctrl_rfWen),
    .io_ldu_s3_loadIn_1_bits_uop_ctrl_fpWen(lsq_io_ldu_s3_loadIn_1_bits_uop_ctrl_fpWen),
    .io_ldu_s3_loadIn_1_bits_uop_ctrl_replayInst(lsq_io_ldu_s3_loadIn_1_bits_uop_ctrl_replayInst),
    .io_ldu_s3_loadIn_1_bits_uop_pdest(lsq_io_ldu_s3_loadIn_1_bits_uop_pdest),
    .io_ldu_s3_loadIn_1_bits_uop_robIdx_flag(lsq_io_ldu_s3_loadIn_1_bits_uop_robIdx_flag),
    .io_ldu_s3_loadIn_1_bits_uop_robIdx_value(lsq_io_ldu_s3_loadIn_1_bits_uop_robIdx_value),
    .io_ldu_s3_loadIn_1_bits_uop_lqIdx_flag(lsq_io_ldu_s3_loadIn_1_bits_uop_lqIdx_flag),
    .io_ldu_s3_loadIn_1_bits_uop_lqIdx_value(lsq_io_ldu_s3_loadIn_1_bits_uop_lqIdx_value),
    .io_ldu_s3_loadIn_1_bits_uop_sqIdx_flag(lsq_io_ldu_s3_loadIn_1_bits_uop_sqIdx_flag),
    .io_ldu_s3_loadIn_1_bits_uop_sqIdx_value(lsq_io_ldu_s3_loadIn_1_bits_uop_sqIdx_value),
    .io_ldu_s3_loadIn_1_bits_vaddr(lsq_io_ldu_s3_loadIn_1_bits_vaddr),
    .io_ldu_s3_loadIn_1_bits_paddr(lsq_io_ldu_s3_loadIn_1_bits_paddr),
    .io_ldu_s3_loadIn_1_bits_mask(lsq_io_ldu_s3_loadIn_1_bits_mask),
    .io_ldu_s3_loadIn_1_bits_miss(lsq_io_ldu_s3_loadIn_1_bits_miss),
    .io_ldu_s3_loadIn_1_bits_tlbMiss(lsq_io_ldu_s3_loadIn_1_bits_tlbMiss),
    .io_ldu_s3_loadIn_1_bits_mmio(lsq_io_ldu_s3_loadIn_1_bits_mmio),
    .io_ldu_s3_loadIn_1_bits_rarAllocated(lsq_io_ldu_s3_loadIn_1_bits_rarAllocated),
    .io_ldu_s3_loadIn_1_bits_rarIndex(lsq_io_ldu_s3_loadIn_1_bits_rarIndex),
    .io_ldu_s3_loadIn_1_bits_rawAllocated(lsq_io_ldu_s3_loadIn_1_bits_rawAllocated),
    .io_ldu_s3_loadIn_1_bits_rawIndex(lsq_io_ldu_s3_loadIn_1_bits_rawIndex),
    .io_ldu_s3_loadIn_1_bits_replayInfo_missMSHRId(lsq_io_ldu_s3_loadIn_1_bits_replayInfo_missMSHRId),
    .io_ldu_s3_loadIn_1_bits_replayInfo_canForwardFullData(lsq_io_ldu_s3_loadIn_1_bits_replayInfo_canForwardFullData),
    .io_ldu_s3_loadIn_1_bits_replayInfo_dataInvalidSqIdx_flag(
      lsq_io_ldu_s3_loadIn_1_bits_replayInfo_dataInvalidSqIdx_flag),
    .io_ldu_s3_loadIn_1_bits_replayInfo_dataInvalidSqIdx_value(
      lsq_io_ldu_s3_loadIn_1_bits_replayInfo_dataInvalidSqIdx_value),
    .io_ldu_s3_loadIn_1_bits_replayInfo_addrInvalidSqIdx_flag(
      lsq_io_ldu_s3_loadIn_1_bits_replayInfo_addrInvalidSqIdx_flag),
    .io_ldu_s3_loadIn_1_bits_replayInfo_addrInvalidSqIdx_value(
      lsq_io_ldu_s3_loadIn_1_bits_replayInfo_addrInvalidSqIdx_value),
    .io_ldu_s3_loadIn_1_bits_replayInfo_replayCarry_real_way_en(
      lsq_io_ldu_s3_loadIn_1_bits_replayInfo_replayCarry_real_way_en),
    .io_ldu_s3_loadIn_1_bits_replayInfo_replayCarry_valid(lsq_io_ldu_s3_loadIn_1_bits_replayInfo_replayCarry_valid),
    .io_ldu_s3_loadIn_1_bits_replayInfo_dataInLastBeat(lsq_io_ldu_s3_loadIn_1_bits_replayInfo_dataInLastBeat),
    .io_ldu_s3_loadIn_1_bits_replayInfo_cause_0(lsq_io_ldu_s3_loadIn_1_bits_replayInfo_cause_0),
    .io_ldu_s3_loadIn_1_bits_replayInfo_cause_1(lsq_io_ldu_s3_loadIn_1_bits_replayInfo_cause_1),
    .io_ldu_s3_loadIn_1_bits_replayInfo_cause_2(lsq_io_ldu_s3_loadIn_1_bits_replayInfo_cause_2),
    .io_ldu_s3_loadIn_1_bits_replayInfo_cause_3(lsq_io_ldu_s3_loadIn_1_bits_replayInfo_cause_3),
    .io_ldu_s3_loadIn_1_bits_replayInfo_cause_4(lsq_io_ldu_s3_loadIn_1_bits_replayInfo_cause_4),
    .io_ldu_s3_loadIn_1_bits_replayInfo_cause_5(lsq_io_ldu_s3_loadIn_1_bits_replayInfo_cause_5),
    .io_ldu_s3_loadIn_1_bits_replayInfo_cause_6(lsq_io_ldu_s3_loadIn_1_bits_replayInfo_cause_6),
    .io_ldu_s3_loadIn_1_bits_replayInfo_cause_7(lsq_io_ldu_s3_loadIn_1_bits_replayInfo_cause_7),
    .io_ldu_s3_loadIn_1_bits_lqDataWenDup_1(lsq_io_ldu_s3_loadIn_1_bits_lqDataWenDup_1),
    .io_ldu_s3_loadIn_1_bits_lqDataWenDup_2(lsq_io_ldu_s3_loadIn_1_bits_lqDataWenDup_2),
    .io_ldu_s3_loadIn_1_bits_lqDataWenDup_3(lsq_io_ldu_s3_loadIn_1_bits_lqDataWenDup_3),
    .io_ldu_s3_loadIn_1_bits_lqDataWenDup_5(lsq_io_ldu_s3_loadIn_1_bits_lqDataWenDup_5),
    .io_sta_s0_storeMaskIn_0_valid(lsq_io_sta_s0_storeMaskIn_0_valid),
    .io_sta_s0_storeMaskIn_0_bits_sqIdx_value(lsq_io_sta_s0_storeMaskIn_0_bits_sqIdx_value),
    .io_sta_s0_storeMaskIn_0_bits_mask(lsq_io_sta_s0_storeMaskIn_0_bits_mask),
    .io_sta_s0_storeMaskIn_1_valid(lsq_io_sta_s0_storeMaskIn_1_valid),
    .io_sta_s0_storeMaskIn_1_bits_sqIdx_value(lsq_io_sta_s0_storeMaskIn_1_bits_sqIdx_value),
    .io_sta_s0_storeMaskIn_1_bits_mask(lsq_io_sta_s0_storeMaskIn_1_bits_mask),
    .io_sta_s1_storeAddrIn_0_valid(lsq_io_sta_s1_storeAddrIn_0_valid),
    .io_sta_s1_storeAddrIn_0_bits_uop_cf_ftqPtr_value(lsq_io_sta_s1_storeAddrIn_0_bits_uop_cf_ftqPtr_value),
    .io_sta_s1_storeAddrIn_0_bits_uop_cf_ftqOffset(lsq_io_sta_s1_storeAddrIn_0_bits_uop_cf_ftqOffset),
    .io_sta_s1_storeAddrIn_0_bits_uop_ctrl_fuOpType(lsq_io_sta_s1_storeAddrIn_0_bits_uop_ctrl_fuOpType),
    .io_sta_s1_storeAddrIn_0_bits_uop_robIdx_flag(lsq_io_sta_s1_storeAddrIn_0_bits_uop_robIdx_flag),
    .io_sta_s1_storeAddrIn_0_bits_uop_robIdx_value(lsq_io_sta_s1_storeAddrIn_0_bits_uop_robIdx_value),
    .io_sta_s1_storeAddrIn_0_bits_uop_sqIdx_flag(lsq_io_sta_s1_storeAddrIn_0_bits_uop_sqIdx_flag),
    .io_sta_s1_storeAddrIn_0_bits_uop_sqIdx_value(lsq_io_sta_s1_storeAddrIn_0_bits_uop_sqIdx_value),
    .io_sta_s1_storeAddrIn_0_bits_vaddr(lsq_io_sta_s1_storeAddrIn_0_bits_vaddr),
    .io_sta_s1_storeAddrIn_0_bits_paddr(lsq_io_sta_s1_storeAddrIn_0_bits_paddr),
    .io_sta_s1_storeAddrIn_0_bits_mask(lsq_io_sta_s1_storeAddrIn_0_bits_mask),
    .io_sta_s1_storeAddrIn_0_bits_wlineflag(lsq_io_sta_s1_storeAddrIn_0_bits_wlineflag),
    .io_sta_s1_storeAddrIn_0_bits_miss(lsq_io_sta_s1_storeAddrIn_0_bits_miss),
    .io_sta_s1_storeAddrIn_1_valid(lsq_io_sta_s1_storeAddrIn_1_valid),
    .io_sta_s1_storeAddrIn_1_bits_uop_cf_ftqPtr_value(lsq_io_sta_s1_storeAddrIn_1_bits_uop_cf_ftqPtr_value),
    .io_sta_s1_storeAddrIn_1_bits_uop_cf_ftqOffset(lsq_io_sta_s1_storeAddrIn_1_bits_uop_cf_ftqOffset),
    .io_sta_s1_storeAddrIn_1_bits_uop_ctrl_fuOpType(lsq_io_sta_s1_storeAddrIn_1_bits_uop_ctrl_fuOpType),
    .io_sta_s1_storeAddrIn_1_bits_uop_robIdx_flag(lsq_io_sta_s1_storeAddrIn_1_bits_uop_robIdx_flag),
    .io_sta_s1_storeAddrIn_1_bits_uop_robIdx_value(lsq_io_sta_s1_storeAddrIn_1_bits_uop_robIdx_value),
    .io_sta_s1_storeAddrIn_1_bits_uop_sqIdx_flag(lsq_io_sta_s1_storeAddrIn_1_bits_uop_sqIdx_flag),
    .io_sta_s1_storeAddrIn_1_bits_uop_sqIdx_value(lsq_io_sta_s1_storeAddrIn_1_bits_uop_sqIdx_value),
    .io_sta_s1_storeAddrIn_1_bits_vaddr(lsq_io_sta_s1_storeAddrIn_1_bits_vaddr),
    .io_sta_s1_storeAddrIn_1_bits_paddr(lsq_io_sta_s1_storeAddrIn_1_bits_paddr),
    .io_sta_s1_storeAddrIn_1_bits_mask(lsq_io_sta_s1_storeAddrIn_1_bits_mask),
    .io_sta_s1_storeAddrIn_1_bits_wlineflag(lsq_io_sta_s1_storeAddrIn_1_bits_wlineflag),
    .io_sta_s1_storeAddrIn_1_bits_miss(lsq_io_sta_s1_storeAddrIn_1_bits_miss),
    .io_sta_s2_storeAddrInRe_0_mmio(lsq_io_sta_s2_storeAddrInRe_0_mmio),
    .io_sta_s2_storeAddrInRe_0_atomic(lsq_io_sta_s2_storeAddrInRe_0_atomic),
    .io_sta_s2_storeAddrInRe_1_mmio(lsq_io_sta_s2_storeAddrInRe_1_mmio),
    .io_sta_s2_storeAddrInRe_1_atomic(lsq_io_sta_s2_storeAddrInRe_1_atomic),
    .io_std_s0_storeDataIn_0_valid(lsq_io_std_s0_storeDataIn_0_valid),
    .io_std_s0_storeDataIn_0_bits_uop_ctrl_fuOpType(lsq_io_std_s0_storeDataIn_0_bits_uop_ctrl_fuOpType),
    .io_std_s0_storeDataIn_0_bits_uop_sqIdx_flag(lsq_io_std_s0_storeDataIn_0_bits_uop_sqIdx_flag),
    .io_std_s0_storeDataIn_0_bits_uop_sqIdx_value(lsq_io_std_s0_storeDataIn_0_bits_uop_sqIdx_value),
    .io_std_s0_storeDataIn_0_bits_data(lsq_io_std_s0_storeDataIn_0_bits_data),
    .io_std_s0_storeDataIn_1_valid(lsq_io_std_s0_storeDataIn_1_valid),
    .io_std_s0_storeDataIn_1_bits_uop_ctrl_fuOpType(lsq_io_std_s0_storeDataIn_1_bits_uop_ctrl_fuOpType),
    .io_std_s0_storeDataIn_1_bits_uop_sqIdx_flag(lsq_io_std_s0_storeDataIn_1_bits_uop_sqIdx_flag),
    .io_std_s0_storeDataIn_1_bits_uop_sqIdx_value(lsq_io_std_s0_storeDataIn_1_bits_uop_sqIdx_value),
    .io_std_s0_storeDataIn_1_bits_data(lsq_io_std_s0_storeDataIn_1_bits_data),
    .io_loadOut_0_ready(lsq_io_loadOut_0_ready),
    .io_loadOut_0_valid(lsq_io_loadOut_0_valid),
    .io_loadOut_0_bits_uop_cf_exceptionVec_4(lsq_io_loadOut_0_bits_uop_cf_exceptionVec_4),
    .io_loadOut_0_bits_uop_cf_exceptionVec_5(lsq_io_loadOut_0_bits_uop_cf_exceptionVec_5),
    .io_loadOut_0_bits_uop_cf_exceptionVec_13(lsq_io_loadOut_0_bits_uop_cf_exceptionVec_13),
    .io_loadOut_0_bits_uop_cf_trigger_backendEn_1(lsq_io_loadOut_0_bits_uop_cf_trigger_backendEn_1),
    .io_loadOut_0_bits_uop_cf_trigger_backendHit_0(lsq_io_loadOut_0_bits_uop_cf_trigger_backendHit_0),
    .io_loadOut_0_bits_uop_cf_trigger_backendHit_1(lsq_io_loadOut_0_bits_uop_cf_trigger_backendHit_1),
    .io_loadOut_0_bits_uop_cf_trigger_backendHit_4(lsq_io_loadOut_0_bits_uop_cf_trigger_backendHit_4),
    .io_loadOut_0_bits_uop_ctrl_rfWen(lsq_io_loadOut_0_bits_uop_ctrl_rfWen),
    .io_loadOut_0_bits_uop_ctrl_fpWen(lsq_io_loadOut_0_bits_uop_ctrl_fpWen),
    .io_loadOut_0_bits_uop_ctrl_flushPipe(lsq_io_loadOut_0_bits_uop_ctrl_flushPipe),
    .io_loadOut_0_bits_uop_ctrl_replayInst(lsq_io_loadOut_0_bits_uop_ctrl_replayInst),
    .io_loadOut_0_bits_uop_pdest(lsq_io_loadOut_0_bits_uop_pdest),
    .io_loadOut_0_bits_uop_robIdx_flag(lsq_io_loadOut_0_bits_uop_robIdx_flag),
    .io_loadOut_0_bits_uop_robIdx_value(lsq_io_loadOut_0_bits_uop_robIdx_value),
    .io_ldRawDataOut_0_lqData(lsq_io_ldRawDataOut_0_lqData),
    .io_ldRawDataOut_0_uop_ctrl_fuOpType(lsq_io_ldRawDataOut_0_uop_ctrl_fuOpType),
    .io_ldRawDataOut_0_uop_ctrl_fpWen(lsq_io_ldRawDataOut_0_uop_ctrl_fpWen),
    .io_ldRawDataOut_0_addrOffset(lsq_io_ldRawDataOut_0_addrOffset),
    .io_replay_0_ready(lsq_io_replay_0_ready),
    .io_replay_0_valid(lsq_io_replay_0_valid),
    .io_replay_0_bits_uop_cf_foldpc(lsq_io_replay_0_bits_uop_cf_foldpc),
    .io_replay_0_bits_uop_cf_trigger_backendEn_1(lsq_io_replay_0_bits_uop_cf_trigger_backendEn_1),
    .io_replay_0_bits_uop_cf_trigger_backendHit_0(lsq_io_replay_0_bits_uop_cf_trigger_backendHit_0),
    .io_replay_0_bits_uop_cf_trigger_backendHit_1(lsq_io_replay_0_bits_uop_cf_trigger_backendHit_1),
    .io_replay_0_bits_uop_cf_trigger_backendHit_4(lsq_io_replay_0_bits_uop_cf_trigger_backendHit_4),
    .io_replay_0_bits_uop_cf_waitForRobIdx_flag(lsq_io_replay_0_bits_uop_cf_waitForRobIdx_flag),
    .io_replay_0_bits_uop_cf_waitForRobIdx_value(lsq_io_replay_0_bits_uop_cf_waitForRobIdx_value),
    .io_replay_0_bits_uop_cf_loadWaitBit(lsq_io_replay_0_bits_uop_cf_loadWaitBit),
    .io_replay_0_bits_uop_cf_loadWaitStrict(lsq_io_replay_0_bits_uop_cf_loadWaitStrict),
    .io_replay_0_bits_uop_cf_ftqPtr_flag(lsq_io_replay_0_bits_uop_cf_ftqPtr_flag),
    .io_replay_0_bits_uop_cf_ftqPtr_value(lsq_io_replay_0_bits_uop_cf_ftqPtr_value),
    .io_replay_0_bits_uop_cf_ftqOffset(lsq_io_replay_0_bits_uop_cf_ftqOffset),
    .io_replay_0_bits_uop_ctrl_fuType(lsq_io_replay_0_bits_uop_ctrl_fuType),
    .io_replay_0_bits_uop_ctrl_fuOpType(lsq_io_replay_0_bits_uop_ctrl_fuOpType),
    .io_replay_0_bits_uop_ctrl_rfWen(lsq_io_replay_0_bits_uop_ctrl_rfWen),
    .io_replay_0_bits_uop_ctrl_fpWen(lsq_io_replay_0_bits_uop_ctrl_fpWen),
    .io_replay_0_bits_uop_pdest(lsq_io_replay_0_bits_uop_pdest),
    .io_replay_0_bits_uop_robIdx_flag(lsq_io_replay_0_bits_uop_robIdx_flag),
    .io_replay_0_bits_uop_robIdx_value(lsq_io_replay_0_bits_uop_robIdx_value),
    .io_replay_0_bits_uop_lqIdx_flag(lsq_io_replay_0_bits_uop_lqIdx_flag),
    .io_replay_0_bits_uop_lqIdx_value(lsq_io_replay_0_bits_uop_lqIdx_value),
    .io_replay_0_bits_uop_sqIdx_flag(lsq_io_replay_0_bits_uop_sqIdx_flag),
    .io_replay_0_bits_uop_sqIdx_value(lsq_io_replay_0_bits_uop_sqIdx_value),
    .io_replay_0_bits_vaddr(lsq_io_replay_0_bits_vaddr),
    .io_replay_0_bits_isFirstIssue(lsq_io_replay_0_bits_isFirstIssue),
    .io_replay_0_bits_replayCarry_real_way_en(lsq_io_replay_0_bits_replayCarry_real_way_en),
    .io_replay_0_bits_replayCarry_valid(lsq_io_replay_0_bits_replayCarry_valid),
    .io_replay_0_bits_mshrid(lsq_io_replay_0_bits_mshrid),
    .io_replay_0_bits_forward_tlDchannel(lsq_io_replay_0_bits_forward_tlDchannel),
    .io_replay_0_bits_rarAllocated(lsq_io_replay_0_bits_rarAllocated),
    .io_replay_0_bits_rarIndex(lsq_io_replay_0_bits_rarIndex),
    .io_replay_0_bits_rawAllocated(lsq_io_replay_0_bits_rawAllocated),
    .io_replay_0_bits_rawIndex(lsq_io_replay_0_bits_rawIndex),
    .io_replay_1_ready(lsq_io_replay_1_ready),
    .io_replay_1_valid(lsq_io_replay_1_valid),
    .io_replay_1_bits_uop_cf_foldpc(lsq_io_replay_1_bits_uop_cf_foldpc),
    .io_replay_1_bits_uop_cf_trigger_backendEn_1(lsq_io_replay_1_bits_uop_cf_trigger_backendEn_1),
    .io_replay_1_bits_uop_cf_trigger_backendHit_0(lsq_io_replay_1_bits_uop_cf_trigger_backendHit_0),
    .io_replay_1_bits_uop_cf_trigger_backendHit_1(lsq_io_replay_1_bits_uop_cf_trigger_backendHit_1),
    .io_replay_1_bits_uop_cf_trigger_backendHit_4(lsq_io_replay_1_bits_uop_cf_trigger_backendHit_4),
    .io_replay_1_bits_uop_cf_waitForRobIdx_flag(lsq_io_replay_1_bits_uop_cf_waitForRobIdx_flag),
    .io_replay_1_bits_uop_cf_waitForRobIdx_value(lsq_io_replay_1_bits_uop_cf_waitForRobIdx_value),
    .io_replay_1_bits_uop_cf_loadWaitBit(lsq_io_replay_1_bits_uop_cf_loadWaitBit),
    .io_replay_1_bits_uop_cf_loadWaitStrict(lsq_io_replay_1_bits_uop_cf_loadWaitStrict),
    .io_replay_1_bits_uop_cf_ftqPtr_flag(lsq_io_replay_1_bits_uop_cf_ftqPtr_flag),
    .io_replay_1_bits_uop_cf_ftqPtr_value(lsq_io_replay_1_bits_uop_cf_ftqPtr_value),
    .io_replay_1_bits_uop_cf_ftqOffset(lsq_io_replay_1_bits_uop_cf_ftqOffset),
    .io_replay_1_bits_uop_ctrl_fuType(lsq_io_replay_1_bits_uop_ctrl_fuType),
    .io_replay_1_bits_uop_ctrl_fuOpType(lsq_io_replay_1_bits_uop_ctrl_fuOpType),
    .io_replay_1_bits_uop_ctrl_rfWen(lsq_io_replay_1_bits_uop_ctrl_rfWen),
    .io_replay_1_bits_uop_ctrl_fpWen(lsq_io_replay_1_bits_uop_ctrl_fpWen),
    .io_replay_1_bits_uop_pdest(lsq_io_replay_1_bits_uop_pdest),
    .io_replay_1_bits_uop_robIdx_flag(lsq_io_replay_1_bits_uop_robIdx_flag),
    .io_replay_1_bits_uop_robIdx_value(lsq_io_replay_1_bits_uop_robIdx_value),
    .io_replay_1_bits_uop_lqIdx_flag(lsq_io_replay_1_bits_uop_lqIdx_flag),
    .io_replay_1_bits_uop_lqIdx_value(lsq_io_replay_1_bits_uop_lqIdx_value),
    .io_replay_1_bits_uop_sqIdx_flag(lsq_io_replay_1_bits_uop_sqIdx_flag),
    .io_replay_1_bits_uop_sqIdx_value(lsq_io_replay_1_bits_uop_sqIdx_value),
    .io_replay_1_bits_vaddr(lsq_io_replay_1_bits_vaddr),
    .io_replay_1_bits_isFirstIssue(lsq_io_replay_1_bits_isFirstIssue),
    .io_replay_1_bits_replayCarry_real_way_en(lsq_io_replay_1_bits_replayCarry_real_way_en),
    .io_replay_1_bits_replayCarry_valid(lsq_io_replay_1_bits_replayCarry_valid),
    .io_replay_1_bits_mshrid(lsq_io_replay_1_bits_mshrid),
    .io_replay_1_bits_forward_tlDchannel(lsq_io_replay_1_bits_forward_tlDchannel),
    .io_replay_1_bits_rarAllocated(lsq_io_replay_1_bits_rarAllocated),
    .io_replay_1_bits_rarIndex(lsq_io_replay_1_bits_rarIndex),
    .io_replay_1_bits_rawAllocated(lsq_io_replay_1_bits_rawAllocated),
    .io_replay_1_bits_rawIndex(lsq_io_replay_1_bits_rawIndex),
    .io_sbuffer_0_ready(lsq_io_sbuffer_0_ready),
    .io_sbuffer_0_valid(lsq_io_sbuffer_0_valid),
    .io_sbuffer_0_bits_addr(lsq_io_sbuffer_0_bits_addr),
    .io_sbuffer_0_bits_data(lsq_io_sbuffer_0_bits_data),
    .io_sbuffer_0_bits_mask(lsq_io_sbuffer_0_bits_mask),
    .io_sbuffer_0_bits_vaddr(lsq_io_sbuffer_0_bits_vaddr),
    .io_sbuffer_0_bits_wline(lsq_io_sbuffer_0_bits_wline),
    .io_sbuffer_1_ready(lsq_io_sbuffer_1_ready),
    .io_sbuffer_1_valid(lsq_io_sbuffer_1_valid),
    .io_sbuffer_1_bits_addr(lsq_io_sbuffer_1_bits_addr),
    .io_sbuffer_1_bits_data(lsq_io_sbuffer_1_bits_data),
    .io_sbuffer_1_bits_mask(lsq_io_sbuffer_1_bits_mask),
    .io_sbuffer_1_bits_vaddr(lsq_io_sbuffer_1_bits_vaddr),
    .io_sbuffer_1_bits_wline(lsq_io_sbuffer_1_bits_wline),
    .io_forward_0_vaddr(lsq_io_forward_0_vaddr),
    .io_forward_0_paddr(lsq_io_forward_0_paddr),
    .io_forward_0_uop_cf_waitForRobIdx_flag(lsq_io_forward_0_uop_cf_waitForRobIdx_flag),
    .io_forward_0_uop_cf_waitForRobIdx_value(lsq_io_forward_0_uop_cf_waitForRobIdx_value),
    .io_forward_0_uop_sqIdx_flag(lsq_io_forward_0_uop_sqIdx_flag),
    .io_forward_0_uop_sqIdx_value(lsq_io_forward_0_uop_sqIdx_value),
    .io_forward_0_valid(lsq_io_forward_0_valid),
    .io_forward_0_forwardMask_0(lsq_io_forward_0_forwardMask_0),
    .io_forward_0_forwardMask_1(lsq_io_forward_0_forwardMask_1),
    .io_forward_0_forwardMask_2(lsq_io_forward_0_forwardMask_2),
    .io_forward_0_forwardMask_3(lsq_io_forward_0_forwardMask_3),
    .io_forward_0_forwardMask_4(lsq_io_forward_0_forwardMask_4),
    .io_forward_0_forwardMask_5(lsq_io_forward_0_forwardMask_5),
    .io_forward_0_forwardMask_6(lsq_io_forward_0_forwardMask_6),
    .io_forward_0_forwardMask_7(lsq_io_forward_0_forwardMask_7),
    .io_forward_0_forwardMask_8(lsq_io_forward_0_forwardMask_8),
    .io_forward_0_forwardMask_9(lsq_io_forward_0_forwardMask_9),
    .io_forward_0_forwardMask_10(lsq_io_forward_0_forwardMask_10),
    .io_forward_0_forwardMask_11(lsq_io_forward_0_forwardMask_11),
    .io_forward_0_forwardMask_12(lsq_io_forward_0_forwardMask_12),
    .io_forward_0_forwardMask_13(lsq_io_forward_0_forwardMask_13),
    .io_forward_0_forwardMask_14(lsq_io_forward_0_forwardMask_14),
    .io_forward_0_forwardMask_15(lsq_io_forward_0_forwardMask_15),
    .io_forward_0_forwardData_0(lsq_io_forward_0_forwardData_0),
    .io_forward_0_forwardData_1(lsq_io_forward_0_forwardData_1),
    .io_forward_0_forwardData_2(lsq_io_forward_0_forwardData_2),
    .io_forward_0_forwardData_3(lsq_io_forward_0_forwardData_3),
    .io_forward_0_forwardData_4(lsq_io_forward_0_forwardData_4),
    .io_forward_0_forwardData_5(lsq_io_forward_0_forwardData_5),
    .io_forward_0_forwardData_6(lsq_io_forward_0_forwardData_6),
    .io_forward_0_forwardData_7(lsq_io_forward_0_forwardData_7),
    .io_forward_0_forwardData_8(lsq_io_forward_0_forwardData_8),
    .io_forward_0_forwardData_9(lsq_io_forward_0_forwardData_9),
    .io_forward_0_forwardData_10(lsq_io_forward_0_forwardData_10),
    .io_forward_0_forwardData_11(lsq_io_forward_0_forwardData_11),
    .io_forward_0_forwardData_12(lsq_io_forward_0_forwardData_12),
    .io_forward_0_forwardData_13(lsq_io_forward_0_forwardData_13),
    .io_forward_0_forwardData_14(lsq_io_forward_0_forwardData_14),
    .io_forward_0_forwardData_15(lsq_io_forward_0_forwardData_15),
    .io_forward_0_sqIdx_flag(lsq_io_forward_0_sqIdx_flag),
    .io_forward_0_dataInvalid(lsq_io_forward_0_dataInvalid),
    .io_forward_0_matchInvalid(lsq_io_forward_0_matchInvalid),
    .io_forward_0_schedWait(lsq_io_forward_0_schedWait),
    .io_forward_0_sqIdxMask(lsq_io_forward_0_sqIdxMask),
    .io_forward_0_dataInvalidSqIdx_flag(lsq_io_forward_0_dataInvalidSqIdx_flag),
    .io_forward_0_dataInvalidSqIdx_value(lsq_io_forward_0_dataInvalidSqIdx_value),
    .io_forward_0_addrInvalidSqIdx_flag(lsq_io_forward_0_addrInvalidSqIdx_flag),
    .io_forward_0_addrInvalidSqIdx_value(lsq_io_forward_0_addrInvalidSqIdx_value),
    .io_forward_1_vaddr(lsq_io_forward_1_vaddr),
    .io_forward_1_paddr(lsq_io_forward_1_paddr),
    .io_forward_1_uop_cf_waitForRobIdx_flag(lsq_io_forward_1_uop_cf_waitForRobIdx_flag),
    .io_forward_1_uop_cf_waitForRobIdx_value(lsq_io_forward_1_uop_cf_waitForRobIdx_value),
    .io_forward_1_uop_sqIdx_flag(lsq_io_forward_1_uop_sqIdx_flag),
    .io_forward_1_uop_sqIdx_value(lsq_io_forward_1_uop_sqIdx_value),
    .io_forward_1_valid(lsq_io_forward_1_valid),
    .io_forward_1_forwardMask_0(lsq_io_forward_1_forwardMask_0),
    .io_forward_1_forwardMask_1(lsq_io_forward_1_forwardMask_1),
    .io_forward_1_forwardMask_2(lsq_io_forward_1_forwardMask_2),
    .io_forward_1_forwardMask_3(lsq_io_forward_1_forwardMask_3),
    .io_forward_1_forwardMask_4(lsq_io_forward_1_forwardMask_4),
    .io_forward_1_forwardMask_5(lsq_io_forward_1_forwardMask_5),
    .io_forward_1_forwardMask_6(lsq_io_forward_1_forwardMask_6),
    .io_forward_1_forwardMask_7(lsq_io_forward_1_forwardMask_7),
    .io_forward_1_forwardMask_8(lsq_io_forward_1_forwardMask_8),
    .io_forward_1_forwardMask_9(lsq_io_forward_1_forwardMask_9),
    .io_forward_1_forwardMask_10(lsq_io_forward_1_forwardMask_10),
    .io_forward_1_forwardMask_11(lsq_io_forward_1_forwardMask_11),
    .io_forward_1_forwardMask_12(lsq_io_forward_1_forwardMask_12),
    .io_forward_1_forwardMask_13(lsq_io_forward_1_forwardMask_13),
    .io_forward_1_forwardMask_14(lsq_io_forward_1_forwardMask_14),
    .io_forward_1_forwardMask_15(lsq_io_forward_1_forwardMask_15),
    .io_forward_1_forwardData_0(lsq_io_forward_1_forwardData_0),
    .io_forward_1_forwardData_1(lsq_io_forward_1_forwardData_1),
    .io_forward_1_forwardData_2(lsq_io_forward_1_forwardData_2),
    .io_forward_1_forwardData_3(lsq_io_forward_1_forwardData_3),
    .io_forward_1_forwardData_4(lsq_io_forward_1_forwardData_4),
    .io_forward_1_forwardData_5(lsq_io_forward_1_forwardData_5),
    .io_forward_1_forwardData_6(lsq_io_forward_1_forwardData_6),
    .io_forward_1_forwardData_7(lsq_io_forward_1_forwardData_7),
    .io_forward_1_forwardData_8(lsq_io_forward_1_forwardData_8),
    .io_forward_1_forwardData_9(lsq_io_forward_1_forwardData_9),
    .io_forward_1_forwardData_10(lsq_io_forward_1_forwardData_10),
    .io_forward_1_forwardData_11(lsq_io_forward_1_forwardData_11),
    .io_forward_1_forwardData_12(lsq_io_forward_1_forwardData_12),
    .io_forward_1_forwardData_13(lsq_io_forward_1_forwardData_13),
    .io_forward_1_forwardData_14(lsq_io_forward_1_forwardData_14),
    .io_forward_1_forwardData_15(lsq_io_forward_1_forwardData_15),
    .io_forward_1_sqIdx_flag(lsq_io_forward_1_sqIdx_flag),
    .io_forward_1_dataInvalid(lsq_io_forward_1_dataInvalid),
    .io_forward_1_matchInvalid(lsq_io_forward_1_matchInvalid),
    .io_forward_1_schedWait(lsq_io_forward_1_schedWait),
    .io_forward_1_sqIdxMask(lsq_io_forward_1_sqIdxMask),
    .io_forward_1_dataInvalidSqIdx_flag(lsq_io_forward_1_dataInvalidSqIdx_flag),
    .io_forward_1_dataInvalidSqIdx_value(lsq_io_forward_1_dataInvalidSqIdx_value),
    .io_forward_1_addrInvalidSqIdx_flag(lsq_io_forward_1_addrInvalidSqIdx_flag),
    .io_forward_1_addrInvalidSqIdx_value(lsq_io_forward_1_addrInvalidSqIdx_value),
    .io_rob_scommit(lsq_io_rob_scommit),
    .io_rob_pendingld(lsq_io_rob_pendingld),
    .io_rob_pendingst(lsq_io_rob_pendingst),
    .io_rob_commit(lsq_io_rob_commit),
    .io_rob_isMMIO_0(lsq_io_rob_isMMIO_0),
    .io_rob_isMMIO_1(lsq_io_rob_isMMIO_1),
    .io_rob_uop_0_robIdx_value(lsq_io_rob_uop_0_robIdx_value),
    .io_rob_uop_1_robIdx_value(lsq_io_rob_uop_1_robIdx_value),
    .io_rollback_valid(lsq_io_rollback_valid),
    .io_rollback_bits_robIdx_flag(lsq_io_rollback_bits_robIdx_flag),
    .io_rollback_bits_robIdx_value(lsq_io_rollback_bits_robIdx_value),
    .io_rollback_bits_ftqIdx_flag(lsq_io_rollback_bits_ftqIdx_flag),
    .io_rollback_bits_ftqIdx_value(lsq_io_rollback_bits_ftqIdx_value),
    .io_rollback_bits_ftqOffset(lsq_io_rollback_bits_ftqOffset),
    .io_rollback_bits_stFtqIdx_value(lsq_io_rollback_bits_stFtqIdx_value),
    .io_rollback_bits_stFtqOffset(lsq_io_rollback_bits_stFtqOffset),
    .io_correctTableUpdate_valid(lsq_io_correctTableUpdate_valid),
    .io_correctTableUpdate_bits_addr(lsq_io_correctTableUpdate_bits_addr),
    .io_release_valid(lsq_io_release_valid),
    .io_release_bits_paddr(lsq_io_release_bits_paddr),
    .io_refill_valid(lsq_io_refill_valid),
    .io_refill_bits_id(lsq_io_refill_bits_id),
    .io_uncacheOutstanding(lsq_io_uncacheOutstanding),
    .io_uncache_req_ready(lsq_io_uncache_req_ready),
    .io_uncache_req_valid(lsq_io_uncache_req_valid),
    .io_uncache_req_bits_cmd(lsq_io_uncache_req_bits_cmd),
    .io_uncache_req_bits_addr(lsq_io_uncache_req_bits_addr),
    .io_uncache_req_bits_data(lsq_io_uncache_req_bits_data),
    .io_uncache_req_bits_mask(lsq_io_uncache_req_bits_mask),
    .io_uncache_req_bits_atomic(lsq_io_uncache_req_bits_atomic),
    .io_uncache_resp_ready(lsq_io_uncache_resp_ready),
    .io_uncache_resp_valid(lsq_io_uncache_resp_valid),
    .io_uncache_resp_bits_data(lsq_io_uncache_resp_bits_data),
    .io_mmioStout_ready(lsq_io_mmioStout_ready),
    .io_mmioStout_valid(lsq_io_mmioStout_valid),
    .io_mmioStout_bits_uop_cf_trigger_backendEn_0(lsq_io_mmioStout_bits_uop_cf_trigger_backendEn_0),
    .io_mmioStout_bits_uop_robIdx_flag(lsq_io_mmioStout_bits_uop_robIdx_flag),
    .io_mmioStout_bits_uop_robIdx_value(lsq_io_mmioStout_bits_uop_robIdx_value),
    .io_sqEmpty(lsq_io_sqEmpty),
    .io_lqReplayFull(lsq_io_lqReplayFull),
    .io_sqCancelCnt(lsq_io_sqCancelCnt),
    .io_lqCancelCnt(lsq_io_lqCancelCnt),
    .io_lqDeq(lsq_io_lqDeq),
    .io_sqDeq(lsq_io_sqDeq),
    .io_exceptionAddr_isStore(lsq_io_exceptionAddr_isStore),
    .io_exceptionAddr_vaddr(lsq_io_exceptionAddr_vaddr),
    .io_trigger_0_hitLoadAddrTriggerHitVec_0(lsq_io_trigger_0_hitLoadAddrTriggerHitVec_0),
    .io_trigger_0_hitLoadAddrTriggerHitVec_1(lsq_io_trigger_0_hitLoadAddrTriggerHitVec_1),
    .io_trigger_0_hitLoadAddrTriggerHitVec_2(lsq_io_trigger_0_hitLoadAddrTriggerHitVec_2),
    .io_trigger_0_lqLoadAddrTriggerHitVec_0(lsq_io_trigger_0_lqLoadAddrTriggerHitVec_0),
    .io_trigger_0_lqLoadAddrTriggerHitVec_1(lsq_io_trigger_0_lqLoadAddrTriggerHitVec_1),
    .io_trigger_0_lqLoadAddrTriggerHitVec_2(lsq_io_trigger_0_lqLoadAddrTriggerHitVec_2),
    .io_trigger_1_hitLoadAddrTriggerHitVec_0(lsq_io_trigger_1_hitLoadAddrTriggerHitVec_0),
    .io_trigger_1_hitLoadAddrTriggerHitVec_1(lsq_io_trigger_1_hitLoadAddrTriggerHitVec_1),
    .io_trigger_1_hitLoadAddrTriggerHitVec_2(lsq_io_trigger_1_hitLoadAddrTriggerHitVec_2),
    .io_perf_0_value(lsq_io_perf_0_value),
    .io_perf_1_value(lsq_io_perf_1_value),
    .io_perf_2_value(lsq_io_perf_2_value),
    .io_perf_3_value(lsq_io_perf_3_value),
    .io_perf_4_value(lsq_io_perf_4_value),
    .io_perf_5_value(lsq_io_perf_5_value),
    .io_perf_6_value(lsq_io_perf_6_value),
    .io_perf_7_value(lsq_io_perf_7_value),
    .io_perf_8_value(lsq_io_perf_8_value),
    .io_perf_9_value(lsq_io_perf_9_value),
    .io_perf_10_value(lsq_io_perf_10_value),
    .io_perf_11_value(lsq_io_perf_11_value),
    .io_perf_12_value(lsq_io_perf_12_value),
    .io_perf_13_value(lsq_io_perf_13_value),
    .io_perf_14_value(lsq_io_perf_14_value),
    .io_perf_15_value(lsq_io_perf_15_value),
    .io_perf_16_value(lsq_io_perf_16_value),
    .io_perf_17_value(lsq_io_perf_17_value),
    .io_perf_18_value(lsq_io_perf_18_value),
    .io_perf_19_value(lsq_io_perf_19_value),
    .io_perf_20_value(lsq_io_perf_20_value),
    .io_perf_21_value(lsq_io_perf_21_value),
    .io_perf_22_value(lsq_io_perf_22_value),
    .io_perf_23_value(lsq_io_perf_23_value),
    .io_perf_24_value(lsq_io_perf_24_value),
    .io_perf_25_value(lsq_io_perf_25_value),
    .io_perf_26_value(lsq_io_perf_26_value),
    .io_perf_27_value(lsq_io_perf_27_value),
    .io_perf_28_value(lsq_io_perf_28_value),
    .io_perf_29_value(lsq_io_perf_29_value)
  );
  Sbuffer sbuffer ( // @[MemBlock.scala 232:23]
    .clock(sbuffer_clock),
    .reset(sbuffer_reset),
    .io_in_0_ready(sbuffer_io_in_0_ready),
    .io_in_0_valid(sbuffer_io_in_0_valid),
    .io_in_0_bits_addr(sbuffer_io_in_0_bits_addr),
    .io_in_0_bits_data(sbuffer_io_in_0_bits_data),
    .io_in_0_bits_mask(sbuffer_io_in_0_bits_mask),
    .io_in_0_bits_vaddr(sbuffer_io_in_0_bits_vaddr),
    .io_in_0_bits_wline(sbuffer_io_in_0_bits_wline),
    .io_in_1_ready(sbuffer_io_in_1_ready),
    .io_in_1_valid(sbuffer_io_in_1_valid),
    .io_in_1_bits_addr(sbuffer_io_in_1_bits_addr),
    .io_in_1_bits_data(sbuffer_io_in_1_bits_data),
    .io_in_1_bits_mask(sbuffer_io_in_1_bits_mask),
    .io_in_1_bits_vaddr(sbuffer_io_in_1_bits_vaddr),
    .io_in_1_bits_wline(sbuffer_io_in_1_bits_wline),
    .io_dcache_req_ready(sbuffer_io_dcache_req_ready),
    .io_dcache_req_valid(sbuffer_io_dcache_req_valid),
    .io_dcache_req_bits_vaddr(sbuffer_io_dcache_req_bits_vaddr),
    .io_dcache_req_bits_addr(sbuffer_io_dcache_req_bits_addr),
    .io_dcache_req_bits_data(sbuffer_io_dcache_req_bits_data),
    .io_dcache_req_bits_mask(sbuffer_io_dcache_req_bits_mask),
    .io_dcache_req_bits_id(sbuffer_io_dcache_req_bits_id),
    .io_dcache_main_pipe_hit_resp_valid(sbuffer_io_dcache_main_pipe_hit_resp_valid),
    .io_dcache_main_pipe_hit_resp_bits_id(sbuffer_io_dcache_main_pipe_hit_resp_bits_id),
    .io_dcache_refill_hit_resp_valid(sbuffer_io_dcache_refill_hit_resp_valid),
    .io_dcache_refill_hit_resp_bits_id(sbuffer_io_dcache_refill_hit_resp_bits_id),
    .io_dcache_replay_resp_valid(sbuffer_io_dcache_replay_resp_valid),
    .io_dcache_replay_resp_bits_id(sbuffer_io_dcache_replay_resp_bits_id),
    .io_forward_0_vaddr(sbuffer_io_forward_0_vaddr),
    .io_forward_0_paddr(sbuffer_io_forward_0_paddr),
    .io_forward_0_valid(sbuffer_io_forward_0_valid),
    .io_forward_0_forwardMask_0(sbuffer_io_forward_0_forwardMask_0),
    .io_forward_0_forwardMask_1(sbuffer_io_forward_0_forwardMask_1),
    .io_forward_0_forwardMask_2(sbuffer_io_forward_0_forwardMask_2),
    .io_forward_0_forwardMask_3(sbuffer_io_forward_0_forwardMask_3),
    .io_forward_0_forwardMask_4(sbuffer_io_forward_0_forwardMask_4),
    .io_forward_0_forwardMask_5(sbuffer_io_forward_0_forwardMask_5),
    .io_forward_0_forwardMask_6(sbuffer_io_forward_0_forwardMask_6),
    .io_forward_0_forwardMask_7(sbuffer_io_forward_0_forwardMask_7),
    .io_forward_0_forwardMask_8(sbuffer_io_forward_0_forwardMask_8),
    .io_forward_0_forwardMask_9(sbuffer_io_forward_0_forwardMask_9),
    .io_forward_0_forwardMask_10(sbuffer_io_forward_0_forwardMask_10),
    .io_forward_0_forwardMask_11(sbuffer_io_forward_0_forwardMask_11),
    .io_forward_0_forwardMask_12(sbuffer_io_forward_0_forwardMask_12),
    .io_forward_0_forwardMask_13(sbuffer_io_forward_0_forwardMask_13),
    .io_forward_0_forwardMask_14(sbuffer_io_forward_0_forwardMask_14),
    .io_forward_0_forwardMask_15(sbuffer_io_forward_0_forwardMask_15),
    .io_forward_0_forwardData_0(sbuffer_io_forward_0_forwardData_0),
    .io_forward_0_forwardData_1(sbuffer_io_forward_0_forwardData_1),
    .io_forward_0_forwardData_2(sbuffer_io_forward_0_forwardData_2),
    .io_forward_0_forwardData_3(sbuffer_io_forward_0_forwardData_3),
    .io_forward_0_forwardData_4(sbuffer_io_forward_0_forwardData_4),
    .io_forward_0_forwardData_5(sbuffer_io_forward_0_forwardData_5),
    .io_forward_0_forwardData_6(sbuffer_io_forward_0_forwardData_6),
    .io_forward_0_forwardData_7(sbuffer_io_forward_0_forwardData_7),
    .io_forward_0_forwardData_8(sbuffer_io_forward_0_forwardData_8),
    .io_forward_0_forwardData_9(sbuffer_io_forward_0_forwardData_9),
    .io_forward_0_forwardData_10(sbuffer_io_forward_0_forwardData_10),
    .io_forward_0_forwardData_11(sbuffer_io_forward_0_forwardData_11),
    .io_forward_0_forwardData_12(sbuffer_io_forward_0_forwardData_12),
    .io_forward_0_forwardData_13(sbuffer_io_forward_0_forwardData_13),
    .io_forward_0_forwardData_14(sbuffer_io_forward_0_forwardData_14),
    .io_forward_0_forwardData_15(sbuffer_io_forward_0_forwardData_15),
    .io_forward_0_matchInvalid(sbuffer_io_forward_0_matchInvalid),
    .io_forward_1_vaddr(sbuffer_io_forward_1_vaddr),
    .io_forward_1_paddr(sbuffer_io_forward_1_paddr),
    .io_forward_1_valid(sbuffer_io_forward_1_valid),
    .io_forward_1_forwardMask_0(sbuffer_io_forward_1_forwardMask_0),
    .io_forward_1_forwardMask_1(sbuffer_io_forward_1_forwardMask_1),
    .io_forward_1_forwardMask_2(sbuffer_io_forward_1_forwardMask_2),
    .io_forward_1_forwardMask_3(sbuffer_io_forward_1_forwardMask_3),
    .io_forward_1_forwardMask_4(sbuffer_io_forward_1_forwardMask_4),
    .io_forward_1_forwardMask_5(sbuffer_io_forward_1_forwardMask_5),
    .io_forward_1_forwardMask_6(sbuffer_io_forward_1_forwardMask_6),
    .io_forward_1_forwardMask_7(sbuffer_io_forward_1_forwardMask_7),
    .io_forward_1_forwardMask_8(sbuffer_io_forward_1_forwardMask_8),
    .io_forward_1_forwardMask_9(sbuffer_io_forward_1_forwardMask_9),
    .io_forward_1_forwardMask_10(sbuffer_io_forward_1_forwardMask_10),
    .io_forward_1_forwardMask_11(sbuffer_io_forward_1_forwardMask_11),
    .io_forward_1_forwardMask_12(sbuffer_io_forward_1_forwardMask_12),
    .io_forward_1_forwardMask_13(sbuffer_io_forward_1_forwardMask_13),
    .io_forward_1_forwardMask_14(sbuffer_io_forward_1_forwardMask_14),
    .io_forward_1_forwardMask_15(sbuffer_io_forward_1_forwardMask_15),
    .io_forward_1_forwardData_0(sbuffer_io_forward_1_forwardData_0),
    .io_forward_1_forwardData_1(sbuffer_io_forward_1_forwardData_1),
    .io_forward_1_forwardData_2(sbuffer_io_forward_1_forwardData_2),
    .io_forward_1_forwardData_3(sbuffer_io_forward_1_forwardData_3),
    .io_forward_1_forwardData_4(sbuffer_io_forward_1_forwardData_4),
    .io_forward_1_forwardData_5(sbuffer_io_forward_1_forwardData_5),
    .io_forward_1_forwardData_6(sbuffer_io_forward_1_forwardData_6),
    .io_forward_1_forwardData_7(sbuffer_io_forward_1_forwardData_7),
    .io_forward_1_forwardData_8(sbuffer_io_forward_1_forwardData_8),
    .io_forward_1_forwardData_9(sbuffer_io_forward_1_forwardData_9),
    .io_forward_1_forwardData_10(sbuffer_io_forward_1_forwardData_10),
    .io_forward_1_forwardData_11(sbuffer_io_forward_1_forwardData_11),
    .io_forward_1_forwardData_12(sbuffer_io_forward_1_forwardData_12),
    .io_forward_1_forwardData_13(sbuffer_io_forward_1_forwardData_13),
    .io_forward_1_forwardData_14(sbuffer_io_forward_1_forwardData_14),
    .io_forward_1_forwardData_15(sbuffer_io_forward_1_forwardData_15),
    .io_forward_1_matchInvalid(sbuffer_io_forward_1_matchInvalid),
    .io_sqempty(sbuffer_io_sqempty),
    .io_flush_valid(sbuffer_io_flush_valid),
    .io_flush_empty(sbuffer_io_flush_empty),
    .io_csrCtrl_sbuffer_threshold(sbuffer_io_csrCtrl_sbuffer_threshold),
    .io_perf_0_value(sbuffer_io_perf_0_value),
    .io_perf_1_value(sbuffer_io_perf_1_value),
    .io_perf_2_value(sbuffer_io_perf_2_value),
    .io_perf_3_value(sbuffer_io_perf_3_value),
    .io_perf_4_value(sbuffer_io_perf_4_value),
    .io_perf_5_value(sbuffer_io_perf_5_value),
    .io_perf_6_value(sbuffer_io_perf_6_value),
    .io_perf_7_value(sbuffer_io_perf_7_value),
    .io_perf_8_value(sbuffer_io_perf_8_value),
    .io_perf_9_value(sbuffer_io_perf_9_value),
    .io_perf_10_value(sbuffer_io_perf_10_value),
    .io_perf_11_value(sbuffer_io_perf_11_value),
    .io_perf_12_value(sbuffer_io_perf_12_value),
    .io_perf_13_value(sbuffer_io_perf_13_value),
    .io_perf_14_value(sbuffer_io_perf_14_value),
    .io_perf_15_value(sbuffer_io_perf_15_value),
    .io_perf_16_value(sbuffer_io_perf_16_value)
  );
  TLBNonBlock dtlb_ld_tlb_ld ( // @[MemBlock.scala 246:24]
    .clock(dtlb_ld_tlb_ld_clock),
    .reset(dtlb_ld_tlb_ld_reset),
    .io_sfence_valid(dtlb_ld_tlb_ld_io_sfence_valid),
    .io_sfence_bits_rs1(dtlb_ld_tlb_ld_io_sfence_bits_rs1),
    .io_sfence_bits_rs2(dtlb_ld_tlb_ld_io_sfence_bits_rs2),
    .io_sfence_bits_addr(dtlb_ld_tlb_ld_io_sfence_bits_addr),
    .io_sfence_bits_asid(dtlb_ld_tlb_ld_io_sfence_bits_asid),
    .io_csr_satp_mode(dtlb_ld_tlb_ld_io_csr_satp_mode),
    .io_csr_satp_asid(dtlb_ld_tlb_ld_io_csr_satp_asid),
    .io_csr_satp_changed(dtlb_ld_tlb_ld_io_csr_satp_changed),
    .io_csr_priv_mxr(dtlb_ld_tlb_ld_io_csr_priv_mxr),
    .io_csr_priv_sum(dtlb_ld_tlb_ld_io_csr_priv_sum),
    .io_csr_priv_dmode(dtlb_ld_tlb_ld_io_csr_priv_dmode),
    .io_requestor_0_req_ready(dtlb_ld_tlb_ld_io_requestor_0_req_ready),
    .io_requestor_0_req_valid(dtlb_ld_tlb_ld_io_requestor_0_req_valid),
    .io_requestor_0_req_bits_vaddr(dtlb_ld_tlb_ld_io_requestor_0_req_bits_vaddr),
    .io_requestor_0_req_bits_cmd(dtlb_ld_tlb_ld_io_requestor_0_req_bits_cmd),
    .io_requestor_0_req_bits_no_translate(dtlb_ld_tlb_ld_io_requestor_0_req_bits_no_translate),
    .io_requestor_0_req_kill(dtlb_ld_tlb_ld_io_requestor_0_req_kill),
    .io_requestor_0_resp_valid(dtlb_ld_tlb_ld_io_requestor_0_resp_valid),
    .io_requestor_0_resp_bits_paddr_0(dtlb_ld_tlb_ld_io_requestor_0_resp_bits_paddr_0),
    .io_requestor_0_resp_bits_paddr_1(dtlb_ld_tlb_ld_io_requestor_0_resp_bits_paddr_1),
    .io_requestor_0_resp_bits_miss(dtlb_ld_tlb_ld_io_requestor_0_resp_bits_miss),
    .io_requestor_0_resp_bits_excp_0_pf_ld(dtlb_ld_tlb_ld_io_requestor_0_resp_bits_excp_0_pf_ld),
    .io_requestor_0_resp_bits_excp_0_pf_st(dtlb_ld_tlb_ld_io_requestor_0_resp_bits_excp_0_pf_st),
    .io_requestor_0_resp_bits_excp_0_af_ld(dtlb_ld_tlb_ld_io_requestor_0_resp_bits_excp_0_af_ld),
    .io_requestor_0_resp_bits_excp_0_af_st(dtlb_ld_tlb_ld_io_requestor_0_resp_bits_excp_0_af_st),
    .io_requestor_0_resp_bits_static_pm_valid(dtlb_ld_tlb_ld_io_requestor_0_resp_bits_static_pm_valid),
    .io_requestor_0_resp_bits_static_pm_bits(dtlb_ld_tlb_ld_io_requestor_0_resp_bits_static_pm_bits),
    .io_requestor_1_req_ready(dtlb_ld_tlb_ld_io_requestor_1_req_ready),
    .io_requestor_1_req_valid(dtlb_ld_tlb_ld_io_requestor_1_req_valid),
    .io_requestor_1_req_bits_vaddr(dtlb_ld_tlb_ld_io_requestor_1_req_bits_vaddr),
    .io_requestor_1_req_bits_cmd(dtlb_ld_tlb_ld_io_requestor_1_req_bits_cmd),
    .io_requestor_1_req_bits_no_translate(dtlb_ld_tlb_ld_io_requestor_1_req_bits_no_translate),
    .io_requestor_1_req_kill(dtlb_ld_tlb_ld_io_requestor_1_req_kill),
    .io_requestor_1_resp_valid(dtlb_ld_tlb_ld_io_requestor_1_resp_valid),
    .io_requestor_1_resp_bits_paddr_0(dtlb_ld_tlb_ld_io_requestor_1_resp_bits_paddr_0),
    .io_requestor_1_resp_bits_paddr_1(dtlb_ld_tlb_ld_io_requestor_1_resp_bits_paddr_1),
    .io_requestor_1_resp_bits_miss(dtlb_ld_tlb_ld_io_requestor_1_resp_bits_miss),
    .io_requestor_1_resp_bits_excp_0_pf_ld(dtlb_ld_tlb_ld_io_requestor_1_resp_bits_excp_0_pf_ld),
    .io_requestor_1_resp_bits_excp_0_af_ld(dtlb_ld_tlb_ld_io_requestor_1_resp_bits_excp_0_af_ld),
    .io_requestor_1_resp_bits_static_pm_valid(dtlb_ld_tlb_ld_io_requestor_1_resp_bits_static_pm_valid),
    .io_requestor_1_resp_bits_static_pm_bits(dtlb_ld_tlb_ld_io_requestor_1_resp_bits_static_pm_bits),
    .io_ptw_req_0_valid(dtlb_ld_tlb_ld_io_ptw_req_0_valid),
    .io_ptw_req_0_bits_vpn(dtlb_ld_tlb_ld_io_ptw_req_0_bits_vpn),
    .io_ptw_req_1_valid(dtlb_ld_tlb_ld_io_ptw_req_1_valid),
    .io_ptw_req_1_bits_vpn(dtlb_ld_tlb_ld_io_ptw_req_1_bits_vpn),
    .io_ptw_resp_ready(dtlb_ld_tlb_ld_io_ptw_resp_ready),
    .io_ptw_resp_valid(dtlb_ld_tlb_ld_io_ptw_resp_valid),
    .io_ptw_resp_bits_entry_tag(dtlb_ld_tlb_ld_io_ptw_resp_bits_entry_tag),
    .io_ptw_resp_bits_entry_asid(dtlb_ld_tlb_ld_io_ptw_resp_bits_entry_asid),
    .io_ptw_resp_bits_entry_ppn(dtlb_ld_tlb_ld_io_ptw_resp_bits_entry_ppn),
    .io_ptw_resp_bits_entry_perm_d(dtlb_ld_tlb_ld_io_ptw_resp_bits_entry_perm_d),
    .io_ptw_resp_bits_entry_perm_a(dtlb_ld_tlb_ld_io_ptw_resp_bits_entry_perm_a),
    .io_ptw_resp_bits_entry_perm_g(dtlb_ld_tlb_ld_io_ptw_resp_bits_entry_perm_g),
    .io_ptw_resp_bits_entry_perm_u(dtlb_ld_tlb_ld_io_ptw_resp_bits_entry_perm_u),
    .io_ptw_resp_bits_entry_perm_x(dtlb_ld_tlb_ld_io_ptw_resp_bits_entry_perm_x),
    .io_ptw_resp_bits_entry_perm_w(dtlb_ld_tlb_ld_io_ptw_resp_bits_entry_perm_w),
    .io_ptw_resp_bits_entry_perm_r(dtlb_ld_tlb_ld_io_ptw_resp_bits_entry_perm_r),
    .io_ptw_resp_bits_entry_level(dtlb_ld_tlb_ld_io_ptw_resp_bits_entry_level),
    .io_ptw_resp_bits_pf(dtlb_ld_tlb_ld_io_ptw_resp_bits_pf),
    .io_ptw_resp_bits_af(dtlb_ld_tlb_ld_io_ptw_resp_bits_af),
    .io_ptw_replenish_c(dtlb_ld_tlb_ld_io_ptw_replenish_c),
    .io_ptw_replenish_atomic(dtlb_ld_tlb_ld_io_ptw_replenish_atomic),
    .io_ptw_replenish_x(dtlb_ld_tlb_ld_io_ptw_replenish_x),
    .io_ptw_replenish_w(dtlb_ld_tlb_ld_io_ptw_replenish_w),
    .io_ptw_replenish_r(dtlb_ld_tlb_ld_io_ptw_replenish_r),
    .io_pmp_0_valid(dtlb_ld_tlb_ld_io_pmp_0_valid),
    .io_pmp_0_bits_addr(dtlb_ld_tlb_ld_io_pmp_0_bits_addr),
    .io_pmp_0_bits_cmd(dtlb_ld_tlb_ld_io_pmp_0_bits_cmd),
    .io_pmp_1_valid(dtlb_ld_tlb_ld_io_pmp_1_valid),
    .io_pmp_1_bits_addr(dtlb_ld_tlb_ld_io_pmp_1_bits_addr),
    .io_pmp_1_bits_cmd(dtlb_ld_tlb_ld_io_pmp_1_bits_cmd)
  );
  TLBNonBlock_1 dtlb_st_tlb_st ( // @[MemBlock.scala 250:24]
    .clock(dtlb_st_tlb_st_clock),
    .reset(dtlb_st_tlb_st_reset),
    .io_sfence_valid(dtlb_st_tlb_st_io_sfence_valid),
    .io_sfence_bits_rs1(dtlb_st_tlb_st_io_sfence_bits_rs1),
    .io_sfence_bits_rs2(dtlb_st_tlb_st_io_sfence_bits_rs2),
    .io_sfence_bits_addr(dtlb_st_tlb_st_io_sfence_bits_addr),
    .io_sfence_bits_asid(dtlb_st_tlb_st_io_sfence_bits_asid),
    .io_csr_satp_mode(dtlb_st_tlb_st_io_csr_satp_mode),
    .io_csr_satp_asid(dtlb_st_tlb_st_io_csr_satp_asid),
    .io_csr_satp_changed(dtlb_st_tlb_st_io_csr_satp_changed),
    .io_csr_priv_sum(dtlb_st_tlb_st_io_csr_priv_sum),
    .io_csr_priv_dmode(dtlb_st_tlb_st_io_csr_priv_dmode),
    .io_requestor_0_req_ready(dtlb_st_tlb_st_io_requestor_0_req_ready),
    .io_requestor_0_req_valid(dtlb_st_tlb_st_io_requestor_0_req_valid),
    .io_requestor_0_req_bits_vaddr(dtlb_st_tlb_st_io_requestor_0_req_bits_vaddr),
    .io_requestor_0_resp_valid(dtlb_st_tlb_st_io_requestor_0_resp_valid),
    .io_requestor_0_resp_bits_paddr_0(dtlb_st_tlb_st_io_requestor_0_resp_bits_paddr_0),
    .io_requestor_0_resp_bits_miss(dtlb_st_tlb_st_io_requestor_0_resp_bits_miss),
    .io_requestor_0_resp_bits_excp_0_pf_st(dtlb_st_tlb_st_io_requestor_0_resp_bits_excp_0_pf_st),
    .io_requestor_0_resp_bits_excp_0_af_st(dtlb_st_tlb_st_io_requestor_0_resp_bits_excp_0_af_st),
    .io_requestor_0_resp_bits_static_pm_valid(dtlb_st_tlb_st_io_requestor_0_resp_bits_static_pm_valid),
    .io_requestor_0_resp_bits_static_pm_bits(dtlb_st_tlb_st_io_requestor_0_resp_bits_static_pm_bits),
    .io_requestor_1_req_ready(dtlb_st_tlb_st_io_requestor_1_req_ready),
    .io_requestor_1_req_valid(dtlb_st_tlb_st_io_requestor_1_req_valid),
    .io_requestor_1_req_bits_vaddr(dtlb_st_tlb_st_io_requestor_1_req_bits_vaddr),
    .io_requestor_1_resp_valid(dtlb_st_tlb_st_io_requestor_1_resp_valid),
    .io_requestor_1_resp_bits_paddr_0(dtlb_st_tlb_st_io_requestor_1_resp_bits_paddr_0),
    .io_requestor_1_resp_bits_miss(dtlb_st_tlb_st_io_requestor_1_resp_bits_miss),
    .io_requestor_1_resp_bits_excp_0_pf_st(dtlb_st_tlb_st_io_requestor_1_resp_bits_excp_0_pf_st),
    .io_requestor_1_resp_bits_excp_0_af_st(dtlb_st_tlb_st_io_requestor_1_resp_bits_excp_0_af_st),
    .io_requestor_1_resp_bits_static_pm_valid(dtlb_st_tlb_st_io_requestor_1_resp_bits_static_pm_valid),
    .io_requestor_1_resp_bits_static_pm_bits(dtlb_st_tlb_st_io_requestor_1_resp_bits_static_pm_bits),
    .io_ptw_req_0_valid(dtlb_st_tlb_st_io_ptw_req_0_valid),
    .io_ptw_req_0_bits_vpn(dtlb_st_tlb_st_io_ptw_req_0_bits_vpn),
    .io_ptw_req_1_valid(dtlb_st_tlb_st_io_ptw_req_1_valid),
    .io_ptw_req_1_bits_vpn(dtlb_st_tlb_st_io_ptw_req_1_bits_vpn),
    .io_ptw_resp_ready(dtlb_st_tlb_st_io_ptw_resp_ready),
    .io_ptw_resp_valid(dtlb_st_tlb_st_io_ptw_resp_valid),
    .io_ptw_resp_bits_entry_tag(dtlb_st_tlb_st_io_ptw_resp_bits_entry_tag),
    .io_ptw_resp_bits_entry_asid(dtlb_st_tlb_st_io_ptw_resp_bits_entry_asid),
    .io_ptw_resp_bits_entry_ppn(dtlb_st_tlb_st_io_ptw_resp_bits_entry_ppn),
    .io_ptw_resp_bits_entry_perm_d(dtlb_st_tlb_st_io_ptw_resp_bits_entry_perm_d),
    .io_ptw_resp_bits_entry_perm_a(dtlb_st_tlb_st_io_ptw_resp_bits_entry_perm_a),
    .io_ptw_resp_bits_entry_perm_g(dtlb_st_tlb_st_io_ptw_resp_bits_entry_perm_g),
    .io_ptw_resp_bits_entry_perm_u(dtlb_st_tlb_st_io_ptw_resp_bits_entry_perm_u),
    .io_ptw_resp_bits_entry_perm_x(dtlb_st_tlb_st_io_ptw_resp_bits_entry_perm_x),
    .io_ptw_resp_bits_entry_perm_w(dtlb_st_tlb_st_io_ptw_resp_bits_entry_perm_w),
    .io_ptw_resp_bits_entry_perm_r(dtlb_st_tlb_st_io_ptw_resp_bits_entry_perm_r),
    .io_ptw_resp_bits_entry_level(dtlb_st_tlb_st_io_ptw_resp_bits_entry_level),
    .io_ptw_resp_bits_pf(dtlb_st_tlb_st_io_ptw_resp_bits_pf),
    .io_ptw_resp_bits_af(dtlb_st_tlb_st_io_ptw_resp_bits_af),
    .io_ptw_replenish_c(dtlb_st_tlb_st_io_ptw_replenish_c),
    .io_ptw_replenish_atomic(dtlb_st_tlb_st_io_ptw_replenish_atomic),
    .io_ptw_replenish_x(dtlb_st_tlb_st_io_ptw_replenish_x),
    .io_ptw_replenish_w(dtlb_st_tlb_st_io_ptw_replenish_w),
    .io_ptw_replenish_r(dtlb_st_tlb_st_io_ptw_replenish_r),
    .io_pmp_0_valid(dtlb_st_tlb_st_io_pmp_0_valid),
    .io_pmp_0_bits_addr(dtlb_st_tlb_st_io_pmp_0_bits_addr),
    .io_pmp_1_valid(dtlb_st_tlb_st_io_pmp_1_valid),
    .io_pmp_1_bits_addr(dtlb_st_tlb_st_io_pmp_1_bits_addr)
  );
  TLBNonBlock_2 dtlb_prefetch_tlb_prefetch ( // @[MemBlock.scala 254:30]
    .clock(dtlb_prefetch_tlb_prefetch_clock),
    .io_sfence_valid(dtlb_prefetch_tlb_prefetch_io_sfence_valid),
    .io_sfence_bits_rs1(dtlb_prefetch_tlb_prefetch_io_sfence_bits_rs1),
    .io_sfence_bits_rs2(dtlb_prefetch_tlb_prefetch_io_sfence_bits_rs2),
    .io_sfence_bits_addr(dtlb_prefetch_tlb_prefetch_io_sfence_bits_addr),
    .io_sfence_bits_asid(dtlb_prefetch_tlb_prefetch_io_sfence_bits_asid),
    .io_csr_satp_mode(dtlb_prefetch_tlb_prefetch_io_csr_satp_mode),
    .io_csr_satp_asid(dtlb_prefetch_tlb_prefetch_io_csr_satp_asid),
    .io_csr_satp_changed(dtlb_prefetch_tlb_prefetch_io_csr_satp_changed),
    .io_csr_priv_dmode(dtlb_prefetch_tlb_prefetch_io_csr_priv_dmode),
    .io_requestor_0_resp_valid(dtlb_prefetch_tlb_prefetch_io_requestor_0_resp_valid),
    .io_ptw_resp_ready(dtlb_prefetch_tlb_prefetch_io_ptw_resp_ready),
    .io_ptw_resp_valid(dtlb_prefetch_tlb_prefetch_io_ptw_resp_valid),
    .io_ptw_resp_bits_entry_tag(dtlb_prefetch_tlb_prefetch_io_ptw_resp_bits_entry_tag),
    .io_ptw_resp_bits_entry_asid(dtlb_prefetch_tlb_prefetch_io_ptw_resp_bits_entry_asid),
    .io_ptw_resp_bits_entry_ppn(dtlb_prefetch_tlb_prefetch_io_ptw_resp_bits_entry_ppn),
    .io_ptw_resp_bits_entry_level(dtlb_prefetch_tlb_prefetch_io_ptw_resp_bits_entry_level),
    .io_pmp_0_valid(dtlb_prefetch_tlb_prefetch_io_pmp_0_valid),
    .io_pmp_0_bits_addr(dtlb_prefetch_tlb_prefetch_io_pmp_0_bits_addr)
  );
  PMP_2 pmp ( // @[MemBlock.scala 311:19]
    .clock(pmp_clock),
    .reset(pmp_reset),
    .io_distribute_csr_wvalid(pmp_io_distribute_csr_wvalid),
    .io_distribute_csr_waddr(pmp_io_distribute_csr_waddr),
    .io_distribute_csr_wdata(pmp_io_distribute_csr_wdata),
    .io_pmp_0_cfg_l(pmp_io_pmp_0_cfg_l),
    .io_pmp_0_cfg_a(pmp_io_pmp_0_cfg_a),
    .io_pmp_0_cfg_x(pmp_io_pmp_0_cfg_x),
    .io_pmp_0_cfg_w(pmp_io_pmp_0_cfg_w),
    .io_pmp_0_cfg_r(pmp_io_pmp_0_cfg_r),
    .io_pmp_0_addr(pmp_io_pmp_0_addr),
    .io_pmp_0_mask(pmp_io_pmp_0_mask),
    .io_pmp_1_cfg_l(pmp_io_pmp_1_cfg_l),
    .io_pmp_1_cfg_a(pmp_io_pmp_1_cfg_a),
    .io_pmp_1_cfg_x(pmp_io_pmp_1_cfg_x),
    .io_pmp_1_cfg_w(pmp_io_pmp_1_cfg_w),
    .io_pmp_1_cfg_r(pmp_io_pmp_1_cfg_r),
    .io_pmp_1_addr(pmp_io_pmp_1_addr),
    .io_pmp_1_mask(pmp_io_pmp_1_mask),
    .io_pmp_2_cfg_l(pmp_io_pmp_2_cfg_l),
    .io_pmp_2_cfg_a(pmp_io_pmp_2_cfg_a),
    .io_pmp_2_cfg_x(pmp_io_pmp_2_cfg_x),
    .io_pmp_2_cfg_w(pmp_io_pmp_2_cfg_w),
    .io_pmp_2_cfg_r(pmp_io_pmp_2_cfg_r),
    .io_pmp_2_addr(pmp_io_pmp_2_addr),
    .io_pmp_2_mask(pmp_io_pmp_2_mask),
    .io_pmp_3_cfg_l(pmp_io_pmp_3_cfg_l),
    .io_pmp_3_cfg_a(pmp_io_pmp_3_cfg_a),
    .io_pmp_3_cfg_x(pmp_io_pmp_3_cfg_x),
    .io_pmp_3_cfg_w(pmp_io_pmp_3_cfg_w),
    .io_pmp_3_cfg_r(pmp_io_pmp_3_cfg_r),
    .io_pmp_3_addr(pmp_io_pmp_3_addr),
    .io_pmp_3_mask(pmp_io_pmp_3_mask),
    .io_pmp_4_cfg_l(pmp_io_pmp_4_cfg_l),
    .io_pmp_4_cfg_a(pmp_io_pmp_4_cfg_a),
    .io_pmp_4_cfg_x(pmp_io_pmp_4_cfg_x),
    .io_pmp_4_cfg_w(pmp_io_pmp_4_cfg_w),
    .io_pmp_4_cfg_r(pmp_io_pmp_4_cfg_r),
    .io_pmp_4_addr(pmp_io_pmp_4_addr),
    .io_pmp_4_mask(pmp_io_pmp_4_mask),
    .io_pmp_5_cfg_l(pmp_io_pmp_5_cfg_l),
    .io_pmp_5_cfg_a(pmp_io_pmp_5_cfg_a),
    .io_pmp_5_cfg_x(pmp_io_pmp_5_cfg_x),
    .io_pmp_5_cfg_w(pmp_io_pmp_5_cfg_w),
    .io_pmp_5_cfg_r(pmp_io_pmp_5_cfg_r),
    .io_pmp_5_addr(pmp_io_pmp_5_addr),
    .io_pmp_5_mask(pmp_io_pmp_5_mask),
    .io_pmp_6_cfg_l(pmp_io_pmp_6_cfg_l),
    .io_pmp_6_cfg_a(pmp_io_pmp_6_cfg_a),
    .io_pmp_6_cfg_x(pmp_io_pmp_6_cfg_x),
    .io_pmp_6_cfg_w(pmp_io_pmp_6_cfg_w),
    .io_pmp_6_cfg_r(pmp_io_pmp_6_cfg_r),
    .io_pmp_6_addr(pmp_io_pmp_6_addr),
    .io_pmp_6_mask(pmp_io_pmp_6_mask),
    .io_pmp_7_cfg_l(pmp_io_pmp_7_cfg_l),
    .io_pmp_7_cfg_a(pmp_io_pmp_7_cfg_a),
    .io_pmp_7_cfg_x(pmp_io_pmp_7_cfg_x),
    .io_pmp_7_cfg_w(pmp_io_pmp_7_cfg_w),
    .io_pmp_7_cfg_r(pmp_io_pmp_7_cfg_r),
    .io_pmp_7_addr(pmp_io_pmp_7_addr),
    .io_pmp_7_mask(pmp_io_pmp_7_mask),
    .io_pmp_8_cfg_l(pmp_io_pmp_8_cfg_l),
    .io_pmp_8_cfg_a(pmp_io_pmp_8_cfg_a),
    .io_pmp_8_cfg_x(pmp_io_pmp_8_cfg_x),
    .io_pmp_8_cfg_w(pmp_io_pmp_8_cfg_w),
    .io_pmp_8_cfg_r(pmp_io_pmp_8_cfg_r),
    .io_pmp_8_addr(pmp_io_pmp_8_addr),
    .io_pmp_8_mask(pmp_io_pmp_8_mask),
    .io_pmp_9_cfg_l(pmp_io_pmp_9_cfg_l),
    .io_pmp_9_cfg_a(pmp_io_pmp_9_cfg_a),
    .io_pmp_9_cfg_x(pmp_io_pmp_9_cfg_x),
    .io_pmp_9_cfg_w(pmp_io_pmp_9_cfg_w),
    .io_pmp_9_cfg_r(pmp_io_pmp_9_cfg_r),
    .io_pmp_9_addr(pmp_io_pmp_9_addr),
    .io_pmp_9_mask(pmp_io_pmp_9_mask),
    .io_pmp_10_cfg_l(pmp_io_pmp_10_cfg_l),
    .io_pmp_10_cfg_a(pmp_io_pmp_10_cfg_a),
    .io_pmp_10_cfg_x(pmp_io_pmp_10_cfg_x),
    .io_pmp_10_cfg_w(pmp_io_pmp_10_cfg_w),
    .io_pmp_10_cfg_r(pmp_io_pmp_10_cfg_r),
    .io_pmp_10_addr(pmp_io_pmp_10_addr),
    .io_pmp_10_mask(pmp_io_pmp_10_mask),
    .io_pmp_11_cfg_l(pmp_io_pmp_11_cfg_l),
    .io_pmp_11_cfg_a(pmp_io_pmp_11_cfg_a),
    .io_pmp_11_cfg_x(pmp_io_pmp_11_cfg_x),
    .io_pmp_11_cfg_w(pmp_io_pmp_11_cfg_w),
    .io_pmp_11_cfg_r(pmp_io_pmp_11_cfg_r),
    .io_pmp_11_addr(pmp_io_pmp_11_addr),
    .io_pmp_11_mask(pmp_io_pmp_11_mask),
    .io_pmp_12_cfg_l(pmp_io_pmp_12_cfg_l),
    .io_pmp_12_cfg_a(pmp_io_pmp_12_cfg_a),
    .io_pmp_12_cfg_x(pmp_io_pmp_12_cfg_x),
    .io_pmp_12_cfg_w(pmp_io_pmp_12_cfg_w),
    .io_pmp_12_cfg_r(pmp_io_pmp_12_cfg_r),
    .io_pmp_12_addr(pmp_io_pmp_12_addr),
    .io_pmp_12_mask(pmp_io_pmp_12_mask),
    .io_pmp_13_cfg_l(pmp_io_pmp_13_cfg_l),
    .io_pmp_13_cfg_a(pmp_io_pmp_13_cfg_a),
    .io_pmp_13_cfg_x(pmp_io_pmp_13_cfg_x),
    .io_pmp_13_cfg_w(pmp_io_pmp_13_cfg_w),
    .io_pmp_13_cfg_r(pmp_io_pmp_13_cfg_r),
    .io_pmp_13_addr(pmp_io_pmp_13_addr),
    .io_pmp_13_mask(pmp_io_pmp_13_mask),
    .io_pmp_14_cfg_l(pmp_io_pmp_14_cfg_l),
    .io_pmp_14_cfg_a(pmp_io_pmp_14_cfg_a),
    .io_pmp_14_cfg_x(pmp_io_pmp_14_cfg_x),
    .io_pmp_14_cfg_w(pmp_io_pmp_14_cfg_w),
    .io_pmp_14_cfg_r(pmp_io_pmp_14_cfg_r),
    .io_pmp_14_addr(pmp_io_pmp_14_addr),
    .io_pmp_14_mask(pmp_io_pmp_14_mask),
    .io_pmp_15_cfg_l(pmp_io_pmp_15_cfg_l),
    .io_pmp_15_cfg_a(pmp_io_pmp_15_cfg_a),
    .io_pmp_15_cfg_x(pmp_io_pmp_15_cfg_x),
    .io_pmp_15_cfg_w(pmp_io_pmp_15_cfg_w),
    .io_pmp_15_cfg_r(pmp_io_pmp_15_cfg_r),
    .io_pmp_15_addr(pmp_io_pmp_15_addr),
    .io_pmp_15_mask(pmp_io_pmp_15_mask),
    .io_pma_0_cfg_c(pmp_io_pma_0_cfg_c),
    .io_pma_0_cfg_atomic(pmp_io_pma_0_cfg_atomic),
    .io_pma_0_cfg_a(pmp_io_pma_0_cfg_a),
    .io_pma_0_cfg_x(pmp_io_pma_0_cfg_x),
    .io_pma_0_cfg_w(pmp_io_pma_0_cfg_w),
    .io_pma_0_cfg_r(pmp_io_pma_0_cfg_r),
    .io_pma_0_addr(pmp_io_pma_0_addr),
    .io_pma_0_mask(pmp_io_pma_0_mask),
    .io_pma_1_cfg_c(pmp_io_pma_1_cfg_c),
    .io_pma_1_cfg_atomic(pmp_io_pma_1_cfg_atomic),
    .io_pma_1_cfg_a(pmp_io_pma_1_cfg_a),
    .io_pma_1_cfg_x(pmp_io_pma_1_cfg_x),
    .io_pma_1_cfg_w(pmp_io_pma_1_cfg_w),
    .io_pma_1_cfg_r(pmp_io_pma_1_cfg_r),
    .io_pma_1_addr(pmp_io_pma_1_addr),
    .io_pma_1_mask(pmp_io_pma_1_mask),
    .io_pma_2_cfg_c(pmp_io_pma_2_cfg_c),
    .io_pma_2_cfg_atomic(pmp_io_pma_2_cfg_atomic),
    .io_pma_2_cfg_a(pmp_io_pma_2_cfg_a),
    .io_pma_2_cfg_x(pmp_io_pma_2_cfg_x),
    .io_pma_2_cfg_w(pmp_io_pma_2_cfg_w),
    .io_pma_2_cfg_r(pmp_io_pma_2_cfg_r),
    .io_pma_2_addr(pmp_io_pma_2_addr),
    .io_pma_2_mask(pmp_io_pma_2_mask),
    .io_pma_3_cfg_c(pmp_io_pma_3_cfg_c),
    .io_pma_3_cfg_atomic(pmp_io_pma_3_cfg_atomic),
    .io_pma_3_cfg_a(pmp_io_pma_3_cfg_a),
    .io_pma_3_cfg_x(pmp_io_pma_3_cfg_x),
    .io_pma_3_cfg_w(pmp_io_pma_3_cfg_w),
    .io_pma_3_cfg_r(pmp_io_pma_3_cfg_r),
    .io_pma_3_addr(pmp_io_pma_3_addr),
    .io_pma_3_mask(pmp_io_pma_3_mask),
    .io_pma_4_cfg_c(pmp_io_pma_4_cfg_c),
    .io_pma_4_cfg_atomic(pmp_io_pma_4_cfg_atomic),
    .io_pma_4_cfg_a(pmp_io_pma_4_cfg_a),
    .io_pma_4_cfg_x(pmp_io_pma_4_cfg_x),
    .io_pma_4_cfg_w(pmp_io_pma_4_cfg_w),
    .io_pma_4_cfg_r(pmp_io_pma_4_cfg_r),
    .io_pma_4_addr(pmp_io_pma_4_addr),
    .io_pma_4_mask(pmp_io_pma_4_mask),
    .io_pma_5_cfg_c(pmp_io_pma_5_cfg_c),
    .io_pma_5_cfg_atomic(pmp_io_pma_5_cfg_atomic),
    .io_pma_5_cfg_a(pmp_io_pma_5_cfg_a),
    .io_pma_5_cfg_x(pmp_io_pma_5_cfg_x),
    .io_pma_5_cfg_w(pmp_io_pma_5_cfg_w),
    .io_pma_5_cfg_r(pmp_io_pma_5_cfg_r),
    .io_pma_5_addr(pmp_io_pma_5_addr),
    .io_pma_5_mask(pmp_io_pma_5_mask),
    .io_pma_6_cfg_c(pmp_io_pma_6_cfg_c),
    .io_pma_6_cfg_atomic(pmp_io_pma_6_cfg_atomic),
    .io_pma_6_cfg_a(pmp_io_pma_6_cfg_a),
    .io_pma_6_cfg_x(pmp_io_pma_6_cfg_x),
    .io_pma_6_cfg_w(pmp_io_pma_6_cfg_w),
    .io_pma_6_cfg_r(pmp_io_pma_6_cfg_r),
    .io_pma_6_addr(pmp_io_pma_6_addr),
    .io_pma_6_mask(pmp_io_pma_6_mask),
    .io_pma_7_cfg_c(pmp_io_pma_7_cfg_c),
    .io_pma_7_cfg_atomic(pmp_io_pma_7_cfg_atomic),
    .io_pma_7_cfg_a(pmp_io_pma_7_cfg_a),
    .io_pma_7_cfg_x(pmp_io_pma_7_cfg_x),
    .io_pma_7_cfg_w(pmp_io_pma_7_cfg_w),
    .io_pma_7_cfg_r(pmp_io_pma_7_cfg_r),
    .io_pma_7_addr(pmp_io_pma_7_addr),
    .io_pma_7_mask(pmp_io_pma_7_mask),
    .io_pma_8_cfg_c(pmp_io_pma_8_cfg_c),
    .io_pma_8_cfg_atomic(pmp_io_pma_8_cfg_atomic),
    .io_pma_8_cfg_a(pmp_io_pma_8_cfg_a),
    .io_pma_8_cfg_x(pmp_io_pma_8_cfg_x),
    .io_pma_8_cfg_w(pmp_io_pma_8_cfg_w),
    .io_pma_8_cfg_r(pmp_io_pma_8_cfg_r),
    .io_pma_8_addr(pmp_io_pma_8_addr),
    .io_pma_8_mask(pmp_io_pma_8_mask),
    .io_pma_9_cfg_c(pmp_io_pma_9_cfg_c),
    .io_pma_9_cfg_atomic(pmp_io_pma_9_cfg_atomic),
    .io_pma_9_cfg_a(pmp_io_pma_9_cfg_a),
    .io_pma_9_cfg_x(pmp_io_pma_9_cfg_x),
    .io_pma_9_cfg_w(pmp_io_pma_9_cfg_w),
    .io_pma_9_cfg_r(pmp_io_pma_9_cfg_r),
    .io_pma_9_addr(pmp_io_pma_9_addr),
    .io_pma_9_mask(pmp_io_pma_9_mask),
    .io_pma_10_cfg_c(pmp_io_pma_10_cfg_c),
    .io_pma_10_cfg_atomic(pmp_io_pma_10_cfg_atomic),
    .io_pma_10_cfg_a(pmp_io_pma_10_cfg_a),
    .io_pma_10_cfg_x(pmp_io_pma_10_cfg_x),
    .io_pma_10_cfg_w(pmp_io_pma_10_cfg_w),
    .io_pma_10_cfg_r(pmp_io_pma_10_cfg_r),
    .io_pma_10_addr(pmp_io_pma_10_addr),
    .io_pma_10_mask(pmp_io_pma_10_mask),
    .io_pma_11_cfg_c(pmp_io_pma_11_cfg_c),
    .io_pma_11_cfg_atomic(pmp_io_pma_11_cfg_atomic),
    .io_pma_11_cfg_a(pmp_io_pma_11_cfg_a),
    .io_pma_11_cfg_x(pmp_io_pma_11_cfg_x),
    .io_pma_11_cfg_w(pmp_io_pma_11_cfg_w),
    .io_pma_11_cfg_r(pmp_io_pma_11_cfg_r),
    .io_pma_11_addr(pmp_io_pma_11_addr),
    .io_pma_11_mask(pmp_io_pma_11_mask),
    .io_pma_12_cfg_c(pmp_io_pma_12_cfg_c),
    .io_pma_12_cfg_atomic(pmp_io_pma_12_cfg_atomic),
    .io_pma_12_cfg_a(pmp_io_pma_12_cfg_a),
    .io_pma_12_cfg_x(pmp_io_pma_12_cfg_x),
    .io_pma_12_cfg_w(pmp_io_pma_12_cfg_w),
    .io_pma_12_cfg_r(pmp_io_pma_12_cfg_r),
    .io_pma_12_addr(pmp_io_pma_12_addr),
    .io_pma_12_mask(pmp_io_pma_12_mask),
    .io_pma_13_cfg_c(pmp_io_pma_13_cfg_c),
    .io_pma_13_cfg_atomic(pmp_io_pma_13_cfg_atomic),
    .io_pma_13_cfg_a(pmp_io_pma_13_cfg_a),
    .io_pma_13_cfg_x(pmp_io_pma_13_cfg_x),
    .io_pma_13_cfg_w(pmp_io_pma_13_cfg_w),
    .io_pma_13_cfg_r(pmp_io_pma_13_cfg_r),
    .io_pma_13_addr(pmp_io_pma_13_addr),
    .io_pma_13_mask(pmp_io_pma_13_mask),
    .io_pma_14_cfg_c(pmp_io_pma_14_cfg_c),
    .io_pma_14_cfg_atomic(pmp_io_pma_14_cfg_atomic),
    .io_pma_14_cfg_a(pmp_io_pma_14_cfg_a),
    .io_pma_14_cfg_x(pmp_io_pma_14_cfg_x),
    .io_pma_14_cfg_w(pmp_io_pma_14_cfg_w),
    .io_pma_14_cfg_r(pmp_io_pma_14_cfg_r),
    .io_pma_14_addr(pmp_io_pma_14_addr),
    .io_pma_14_mask(pmp_io_pma_14_mask),
    .io_pma_15_cfg_c(pmp_io_pma_15_cfg_c),
    .io_pma_15_cfg_atomic(pmp_io_pma_15_cfg_atomic),
    .io_pma_15_cfg_a(pmp_io_pma_15_cfg_a),
    .io_pma_15_cfg_x(pmp_io_pma_15_cfg_x),
    .io_pma_15_cfg_w(pmp_io_pma_15_cfg_w),
    .io_pma_15_cfg_r(pmp_io_pma_15_cfg_r),
    .io_pma_15_addr(pmp_io_pma_15_addr),
    .io_pma_15_mask(pmp_io_pma_15_mask)
  );
  PMPChecker_8 PMPChecker ( // @[MemBlock.scala 314:91]
    .clock(PMPChecker_clock),
    .io_check_env_mode(PMPChecker_io_check_env_mode),
    .io_check_env_pmp_0_cfg_l(PMPChecker_io_check_env_pmp_0_cfg_l),
    .io_check_env_pmp_0_cfg_a(PMPChecker_io_check_env_pmp_0_cfg_a),
    .io_check_env_pmp_0_cfg_w(PMPChecker_io_check_env_pmp_0_cfg_w),
    .io_check_env_pmp_0_cfg_r(PMPChecker_io_check_env_pmp_0_cfg_r),
    .io_check_env_pmp_0_addr(PMPChecker_io_check_env_pmp_0_addr),
    .io_check_env_pmp_0_mask(PMPChecker_io_check_env_pmp_0_mask),
    .io_check_env_pmp_1_cfg_l(PMPChecker_io_check_env_pmp_1_cfg_l),
    .io_check_env_pmp_1_cfg_a(PMPChecker_io_check_env_pmp_1_cfg_a),
    .io_check_env_pmp_1_cfg_w(PMPChecker_io_check_env_pmp_1_cfg_w),
    .io_check_env_pmp_1_cfg_r(PMPChecker_io_check_env_pmp_1_cfg_r),
    .io_check_env_pmp_1_addr(PMPChecker_io_check_env_pmp_1_addr),
    .io_check_env_pmp_1_mask(PMPChecker_io_check_env_pmp_1_mask),
    .io_check_env_pmp_2_cfg_l(PMPChecker_io_check_env_pmp_2_cfg_l),
    .io_check_env_pmp_2_cfg_a(PMPChecker_io_check_env_pmp_2_cfg_a),
    .io_check_env_pmp_2_cfg_w(PMPChecker_io_check_env_pmp_2_cfg_w),
    .io_check_env_pmp_2_cfg_r(PMPChecker_io_check_env_pmp_2_cfg_r),
    .io_check_env_pmp_2_addr(PMPChecker_io_check_env_pmp_2_addr),
    .io_check_env_pmp_2_mask(PMPChecker_io_check_env_pmp_2_mask),
    .io_check_env_pmp_3_cfg_l(PMPChecker_io_check_env_pmp_3_cfg_l),
    .io_check_env_pmp_3_cfg_a(PMPChecker_io_check_env_pmp_3_cfg_a),
    .io_check_env_pmp_3_cfg_w(PMPChecker_io_check_env_pmp_3_cfg_w),
    .io_check_env_pmp_3_cfg_r(PMPChecker_io_check_env_pmp_3_cfg_r),
    .io_check_env_pmp_3_addr(PMPChecker_io_check_env_pmp_3_addr),
    .io_check_env_pmp_3_mask(PMPChecker_io_check_env_pmp_3_mask),
    .io_check_env_pmp_4_cfg_l(PMPChecker_io_check_env_pmp_4_cfg_l),
    .io_check_env_pmp_4_cfg_a(PMPChecker_io_check_env_pmp_4_cfg_a),
    .io_check_env_pmp_4_cfg_w(PMPChecker_io_check_env_pmp_4_cfg_w),
    .io_check_env_pmp_4_cfg_r(PMPChecker_io_check_env_pmp_4_cfg_r),
    .io_check_env_pmp_4_addr(PMPChecker_io_check_env_pmp_4_addr),
    .io_check_env_pmp_4_mask(PMPChecker_io_check_env_pmp_4_mask),
    .io_check_env_pmp_5_cfg_l(PMPChecker_io_check_env_pmp_5_cfg_l),
    .io_check_env_pmp_5_cfg_a(PMPChecker_io_check_env_pmp_5_cfg_a),
    .io_check_env_pmp_5_cfg_w(PMPChecker_io_check_env_pmp_5_cfg_w),
    .io_check_env_pmp_5_cfg_r(PMPChecker_io_check_env_pmp_5_cfg_r),
    .io_check_env_pmp_5_addr(PMPChecker_io_check_env_pmp_5_addr),
    .io_check_env_pmp_5_mask(PMPChecker_io_check_env_pmp_5_mask),
    .io_check_env_pmp_6_cfg_l(PMPChecker_io_check_env_pmp_6_cfg_l),
    .io_check_env_pmp_6_cfg_a(PMPChecker_io_check_env_pmp_6_cfg_a),
    .io_check_env_pmp_6_cfg_w(PMPChecker_io_check_env_pmp_6_cfg_w),
    .io_check_env_pmp_6_cfg_r(PMPChecker_io_check_env_pmp_6_cfg_r),
    .io_check_env_pmp_6_addr(PMPChecker_io_check_env_pmp_6_addr),
    .io_check_env_pmp_6_mask(PMPChecker_io_check_env_pmp_6_mask),
    .io_check_env_pmp_7_cfg_l(PMPChecker_io_check_env_pmp_7_cfg_l),
    .io_check_env_pmp_7_cfg_a(PMPChecker_io_check_env_pmp_7_cfg_a),
    .io_check_env_pmp_7_cfg_w(PMPChecker_io_check_env_pmp_7_cfg_w),
    .io_check_env_pmp_7_cfg_r(PMPChecker_io_check_env_pmp_7_cfg_r),
    .io_check_env_pmp_7_addr(PMPChecker_io_check_env_pmp_7_addr),
    .io_check_env_pmp_7_mask(PMPChecker_io_check_env_pmp_7_mask),
    .io_check_env_pmp_8_cfg_l(PMPChecker_io_check_env_pmp_8_cfg_l),
    .io_check_env_pmp_8_cfg_a(PMPChecker_io_check_env_pmp_8_cfg_a),
    .io_check_env_pmp_8_cfg_w(PMPChecker_io_check_env_pmp_8_cfg_w),
    .io_check_env_pmp_8_cfg_r(PMPChecker_io_check_env_pmp_8_cfg_r),
    .io_check_env_pmp_8_addr(PMPChecker_io_check_env_pmp_8_addr),
    .io_check_env_pmp_8_mask(PMPChecker_io_check_env_pmp_8_mask),
    .io_check_env_pmp_9_cfg_l(PMPChecker_io_check_env_pmp_9_cfg_l),
    .io_check_env_pmp_9_cfg_a(PMPChecker_io_check_env_pmp_9_cfg_a),
    .io_check_env_pmp_9_cfg_w(PMPChecker_io_check_env_pmp_9_cfg_w),
    .io_check_env_pmp_9_cfg_r(PMPChecker_io_check_env_pmp_9_cfg_r),
    .io_check_env_pmp_9_addr(PMPChecker_io_check_env_pmp_9_addr),
    .io_check_env_pmp_9_mask(PMPChecker_io_check_env_pmp_9_mask),
    .io_check_env_pmp_10_cfg_l(PMPChecker_io_check_env_pmp_10_cfg_l),
    .io_check_env_pmp_10_cfg_a(PMPChecker_io_check_env_pmp_10_cfg_a),
    .io_check_env_pmp_10_cfg_w(PMPChecker_io_check_env_pmp_10_cfg_w),
    .io_check_env_pmp_10_cfg_r(PMPChecker_io_check_env_pmp_10_cfg_r),
    .io_check_env_pmp_10_addr(PMPChecker_io_check_env_pmp_10_addr),
    .io_check_env_pmp_10_mask(PMPChecker_io_check_env_pmp_10_mask),
    .io_check_env_pmp_11_cfg_l(PMPChecker_io_check_env_pmp_11_cfg_l),
    .io_check_env_pmp_11_cfg_a(PMPChecker_io_check_env_pmp_11_cfg_a),
    .io_check_env_pmp_11_cfg_w(PMPChecker_io_check_env_pmp_11_cfg_w),
    .io_check_env_pmp_11_cfg_r(PMPChecker_io_check_env_pmp_11_cfg_r),
    .io_check_env_pmp_11_addr(PMPChecker_io_check_env_pmp_11_addr),
    .io_check_env_pmp_11_mask(PMPChecker_io_check_env_pmp_11_mask),
    .io_check_env_pmp_12_cfg_l(PMPChecker_io_check_env_pmp_12_cfg_l),
    .io_check_env_pmp_12_cfg_a(PMPChecker_io_check_env_pmp_12_cfg_a),
    .io_check_env_pmp_12_cfg_w(PMPChecker_io_check_env_pmp_12_cfg_w),
    .io_check_env_pmp_12_cfg_r(PMPChecker_io_check_env_pmp_12_cfg_r),
    .io_check_env_pmp_12_addr(PMPChecker_io_check_env_pmp_12_addr),
    .io_check_env_pmp_12_mask(PMPChecker_io_check_env_pmp_12_mask),
    .io_check_env_pmp_13_cfg_l(PMPChecker_io_check_env_pmp_13_cfg_l),
    .io_check_env_pmp_13_cfg_a(PMPChecker_io_check_env_pmp_13_cfg_a),
    .io_check_env_pmp_13_cfg_w(PMPChecker_io_check_env_pmp_13_cfg_w),
    .io_check_env_pmp_13_cfg_r(PMPChecker_io_check_env_pmp_13_cfg_r),
    .io_check_env_pmp_13_addr(PMPChecker_io_check_env_pmp_13_addr),
    .io_check_env_pmp_13_mask(PMPChecker_io_check_env_pmp_13_mask),
    .io_check_env_pmp_14_cfg_l(PMPChecker_io_check_env_pmp_14_cfg_l),
    .io_check_env_pmp_14_cfg_a(PMPChecker_io_check_env_pmp_14_cfg_a),
    .io_check_env_pmp_14_cfg_w(PMPChecker_io_check_env_pmp_14_cfg_w),
    .io_check_env_pmp_14_cfg_r(PMPChecker_io_check_env_pmp_14_cfg_r),
    .io_check_env_pmp_14_addr(PMPChecker_io_check_env_pmp_14_addr),
    .io_check_env_pmp_14_mask(PMPChecker_io_check_env_pmp_14_mask),
    .io_check_env_pmp_15_cfg_l(PMPChecker_io_check_env_pmp_15_cfg_l),
    .io_check_env_pmp_15_cfg_a(PMPChecker_io_check_env_pmp_15_cfg_a),
    .io_check_env_pmp_15_cfg_w(PMPChecker_io_check_env_pmp_15_cfg_w),
    .io_check_env_pmp_15_cfg_r(PMPChecker_io_check_env_pmp_15_cfg_r),
    .io_check_env_pmp_15_addr(PMPChecker_io_check_env_pmp_15_addr),
    .io_check_env_pmp_15_mask(PMPChecker_io_check_env_pmp_15_mask),
    .io_check_env_pma_0_cfg_c(PMPChecker_io_check_env_pma_0_cfg_c),
    .io_check_env_pma_0_cfg_atomic(PMPChecker_io_check_env_pma_0_cfg_atomic),
    .io_check_env_pma_0_cfg_a(PMPChecker_io_check_env_pma_0_cfg_a),
    .io_check_env_pma_0_cfg_w(PMPChecker_io_check_env_pma_0_cfg_w),
    .io_check_env_pma_0_cfg_r(PMPChecker_io_check_env_pma_0_cfg_r),
    .io_check_env_pma_0_addr(PMPChecker_io_check_env_pma_0_addr),
    .io_check_env_pma_0_mask(PMPChecker_io_check_env_pma_0_mask),
    .io_check_env_pma_1_cfg_c(PMPChecker_io_check_env_pma_1_cfg_c),
    .io_check_env_pma_1_cfg_atomic(PMPChecker_io_check_env_pma_1_cfg_atomic),
    .io_check_env_pma_1_cfg_a(PMPChecker_io_check_env_pma_1_cfg_a),
    .io_check_env_pma_1_cfg_w(PMPChecker_io_check_env_pma_1_cfg_w),
    .io_check_env_pma_1_cfg_r(PMPChecker_io_check_env_pma_1_cfg_r),
    .io_check_env_pma_1_addr(PMPChecker_io_check_env_pma_1_addr),
    .io_check_env_pma_1_mask(PMPChecker_io_check_env_pma_1_mask),
    .io_check_env_pma_2_cfg_c(PMPChecker_io_check_env_pma_2_cfg_c),
    .io_check_env_pma_2_cfg_atomic(PMPChecker_io_check_env_pma_2_cfg_atomic),
    .io_check_env_pma_2_cfg_a(PMPChecker_io_check_env_pma_2_cfg_a),
    .io_check_env_pma_2_cfg_w(PMPChecker_io_check_env_pma_2_cfg_w),
    .io_check_env_pma_2_cfg_r(PMPChecker_io_check_env_pma_2_cfg_r),
    .io_check_env_pma_2_addr(PMPChecker_io_check_env_pma_2_addr),
    .io_check_env_pma_2_mask(PMPChecker_io_check_env_pma_2_mask),
    .io_check_env_pma_3_cfg_c(PMPChecker_io_check_env_pma_3_cfg_c),
    .io_check_env_pma_3_cfg_atomic(PMPChecker_io_check_env_pma_3_cfg_atomic),
    .io_check_env_pma_3_cfg_a(PMPChecker_io_check_env_pma_3_cfg_a),
    .io_check_env_pma_3_cfg_w(PMPChecker_io_check_env_pma_3_cfg_w),
    .io_check_env_pma_3_cfg_r(PMPChecker_io_check_env_pma_3_cfg_r),
    .io_check_env_pma_3_addr(PMPChecker_io_check_env_pma_3_addr),
    .io_check_env_pma_3_mask(PMPChecker_io_check_env_pma_3_mask),
    .io_check_env_pma_4_cfg_c(PMPChecker_io_check_env_pma_4_cfg_c),
    .io_check_env_pma_4_cfg_atomic(PMPChecker_io_check_env_pma_4_cfg_atomic),
    .io_check_env_pma_4_cfg_a(PMPChecker_io_check_env_pma_4_cfg_a),
    .io_check_env_pma_4_cfg_w(PMPChecker_io_check_env_pma_4_cfg_w),
    .io_check_env_pma_4_cfg_r(PMPChecker_io_check_env_pma_4_cfg_r),
    .io_check_env_pma_4_addr(PMPChecker_io_check_env_pma_4_addr),
    .io_check_env_pma_4_mask(PMPChecker_io_check_env_pma_4_mask),
    .io_check_env_pma_5_cfg_c(PMPChecker_io_check_env_pma_5_cfg_c),
    .io_check_env_pma_5_cfg_atomic(PMPChecker_io_check_env_pma_5_cfg_atomic),
    .io_check_env_pma_5_cfg_a(PMPChecker_io_check_env_pma_5_cfg_a),
    .io_check_env_pma_5_cfg_w(PMPChecker_io_check_env_pma_5_cfg_w),
    .io_check_env_pma_5_cfg_r(PMPChecker_io_check_env_pma_5_cfg_r),
    .io_check_env_pma_5_addr(PMPChecker_io_check_env_pma_5_addr),
    .io_check_env_pma_5_mask(PMPChecker_io_check_env_pma_5_mask),
    .io_check_env_pma_6_cfg_c(PMPChecker_io_check_env_pma_6_cfg_c),
    .io_check_env_pma_6_cfg_atomic(PMPChecker_io_check_env_pma_6_cfg_atomic),
    .io_check_env_pma_6_cfg_a(PMPChecker_io_check_env_pma_6_cfg_a),
    .io_check_env_pma_6_cfg_w(PMPChecker_io_check_env_pma_6_cfg_w),
    .io_check_env_pma_6_cfg_r(PMPChecker_io_check_env_pma_6_cfg_r),
    .io_check_env_pma_6_addr(PMPChecker_io_check_env_pma_6_addr),
    .io_check_env_pma_6_mask(PMPChecker_io_check_env_pma_6_mask),
    .io_check_env_pma_7_cfg_c(PMPChecker_io_check_env_pma_7_cfg_c),
    .io_check_env_pma_7_cfg_atomic(PMPChecker_io_check_env_pma_7_cfg_atomic),
    .io_check_env_pma_7_cfg_a(PMPChecker_io_check_env_pma_7_cfg_a),
    .io_check_env_pma_7_cfg_w(PMPChecker_io_check_env_pma_7_cfg_w),
    .io_check_env_pma_7_cfg_r(PMPChecker_io_check_env_pma_7_cfg_r),
    .io_check_env_pma_7_addr(PMPChecker_io_check_env_pma_7_addr),
    .io_check_env_pma_7_mask(PMPChecker_io_check_env_pma_7_mask),
    .io_check_env_pma_8_cfg_c(PMPChecker_io_check_env_pma_8_cfg_c),
    .io_check_env_pma_8_cfg_atomic(PMPChecker_io_check_env_pma_8_cfg_atomic),
    .io_check_env_pma_8_cfg_a(PMPChecker_io_check_env_pma_8_cfg_a),
    .io_check_env_pma_8_cfg_w(PMPChecker_io_check_env_pma_8_cfg_w),
    .io_check_env_pma_8_cfg_r(PMPChecker_io_check_env_pma_8_cfg_r),
    .io_check_env_pma_8_addr(PMPChecker_io_check_env_pma_8_addr),
    .io_check_env_pma_8_mask(PMPChecker_io_check_env_pma_8_mask),
    .io_check_env_pma_9_cfg_c(PMPChecker_io_check_env_pma_9_cfg_c),
    .io_check_env_pma_9_cfg_atomic(PMPChecker_io_check_env_pma_9_cfg_atomic),
    .io_check_env_pma_9_cfg_a(PMPChecker_io_check_env_pma_9_cfg_a),
    .io_check_env_pma_9_cfg_w(PMPChecker_io_check_env_pma_9_cfg_w),
    .io_check_env_pma_9_cfg_r(PMPChecker_io_check_env_pma_9_cfg_r),
    .io_check_env_pma_9_addr(PMPChecker_io_check_env_pma_9_addr),
    .io_check_env_pma_9_mask(PMPChecker_io_check_env_pma_9_mask),
    .io_check_env_pma_10_cfg_c(PMPChecker_io_check_env_pma_10_cfg_c),
    .io_check_env_pma_10_cfg_atomic(PMPChecker_io_check_env_pma_10_cfg_atomic),
    .io_check_env_pma_10_cfg_a(PMPChecker_io_check_env_pma_10_cfg_a),
    .io_check_env_pma_10_cfg_w(PMPChecker_io_check_env_pma_10_cfg_w),
    .io_check_env_pma_10_cfg_r(PMPChecker_io_check_env_pma_10_cfg_r),
    .io_check_env_pma_10_addr(PMPChecker_io_check_env_pma_10_addr),
    .io_check_env_pma_10_mask(PMPChecker_io_check_env_pma_10_mask),
    .io_check_env_pma_11_cfg_c(PMPChecker_io_check_env_pma_11_cfg_c),
    .io_check_env_pma_11_cfg_atomic(PMPChecker_io_check_env_pma_11_cfg_atomic),
    .io_check_env_pma_11_cfg_a(PMPChecker_io_check_env_pma_11_cfg_a),
    .io_check_env_pma_11_cfg_w(PMPChecker_io_check_env_pma_11_cfg_w),
    .io_check_env_pma_11_cfg_r(PMPChecker_io_check_env_pma_11_cfg_r),
    .io_check_env_pma_11_addr(PMPChecker_io_check_env_pma_11_addr),
    .io_check_env_pma_11_mask(PMPChecker_io_check_env_pma_11_mask),
    .io_check_env_pma_12_cfg_c(PMPChecker_io_check_env_pma_12_cfg_c),
    .io_check_env_pma_12_cfg_atomic(PMPChecker_io_check_env_pma_12_cfg_atomic),
    .io_check_env_pma_12_cfg_a(PMPChecker_io_check_env_pma_12_cfg_a),
    .io_check_env_pma_12_cfg_w(PMPChecker_io_check_env_pma_12_cfg_w),
    .io_check_env_pma_12_cfg_r(PMPChecker_io_check_env_pma_12_cfg_r),
    .io_check_env_pma_12_addr(PMPChecker_io_check_env_pma_12_addr),
    .io_check_env_pma_12_mask(PMPChecker_io_check_env_pma_12_mask),
    .io_check_env_pma_13_cfg_c(PMPChecker_io_check_env_pma_13_cfg_c),
    .io_check_env_pma_13_cfg_atomic(PMPChecker_io_check_env_pma_13_cfg_atomic),
    .io_check_env_pma_13_cfg_a(PMPChecker_io_check_env_pma_13_cfg_a),
    .io_check_env_pma_13_cfg_w(PMPChecker_io_check_env_pma_13_cfg_w),
    .io_check_env_pma_13_cfg_r(PMPChecker_io_check_env_pma_13_cfg_r),
    .io_check_env_pma_13_addr(PMPChecker_io_check_env_pma_13_addr),
    .io_check_env_pma_13_mask(PMPChecker_io_check_env_pma_13_mask),
    .io_check_env_pma_14_cfg_c(PMPChecker_io_check_env_pma_14_cfg_c),
    .io_check_env_pma_14_cfg_atomic(PMPChecker_io_check_env_pma_14_cfg_atomic),
    .io_check_env_pma_14_cfg_a(PMPChecker_io_check_env_pma_14_cfg_a),
    .io_check_env_pma_14_cfg_w(PMPChecker_io_check_env_pma_14_cfg_w),
    .io_check_env_pma_14_cfg_r(PMPChecker_io_check_env_pma_14_cfg_r),
    .io_check_env_pma_14_addr(PMPChecker_io_check_env_pma_14_addr),
    .io_check_env_pma_14_mask(PMPChecker_io_check_env_pma_14_mask),
    .io_check_env_pma_15_cfg_c(PMPChecker_io_check_env_pma_15_cfg_c),
    .io_check_env_pma_15_cfg_atomic(PMPChecker_io_check_env_pma_15_cfg_atomic),
    .io_check_env_pma_15_cfg_a(PMPChecker_io_check_env_pma_15_cfg_a),
    .io_check_env_pma_15_cfg_w(PMPChecker_io_check_env_pma_15_cfg_w),
    .io_check_env_pma_15_cfg_r(PMPChecker_io_check_env_pma_15_cfg_r),
    .io_check_env_pma_15_addr(PMPChecker_io_check_env_pma_15_addr),
    .io_check_env_pma_15_mask(PMPChecker_io_check_env_pma_15_mask),
    .io_req_valid(PMPChecker_io_req_valid),
    .io_req_bits_addr(PMPChecker_io_req_bits_addr),
    .io_req_bits_cmd(PMPChecker_io_req_bits_cmd),
    .io_resp_ld(PMPChecker_io_resp_ld),
    .io_resp_st(PMPChecker_io_resp_st),
    .io_resp_mmio(PMPChecker_io_resp_mmio),
    .io_resp_atomic(PMPChecker_io_resp_atomic)
  );
  PMPChecker_8 PMPChecker_1 ( // @[MemBlock.scala 314:91]
    .clock(PMPChecker_1_clock),
    .io_check_env_mode(PMPChecker_1_io_check_env_mode),
    .io_check_env_pmp_0_cfg_l(PMPChecker_1_io_check_env_pmp_0_cfg_l),
    .io_check_env_pmp_0_cfg_a(PMPChecker_1_io_check_env_pmp_0_cfg_a),
    .io_check_env_pmp_0_cfg_w(PMPChecker_1_io_check_env_pmp_0_cfg_w),
    .io_check_env_pmp_0_cfg_r(PMPChecker_1_io_check_env_pmp_0_cfg_r),
    .io_check_env_pmp_0_addr(PMPChecker_1_io_check_env_pmp_0_addr),
    .io_check_env_pmp_0_mask(PMPChecker_1_io_check_env_pmp_0_mask),
    .io_check_env_pmp_1_cfg_l(PMPChecker_1_io_check_env_pmp_1_cfg_l),
    .io_check_env_pmp_1_cfg_a(PMPChecker_1_io_check_env_pmp_1_cfg_a),
    .io_check_env_pmp_1_cfg_w(PMPChecker_1_io_check_env_pmp_1_cfg_w),
    .io_check_env_pmp_1_cfg_r(PMPChecker_1_io_check_env_pmp_1_cfg_r),
    .io_check_env_pmp_1_addr(PMPChecker_1_io_check_env_pmp_1_addr),
    .io_check_env_pmp_1_mask(PMPChecker_1_io_check_env_pmp_1_mask),
    .io_check_env_pmp_2_cfg_l(PMPChecker_1_io_check_env_pmp_2_cfg_l),
    .io_check_env_pmp_2_cfg_a(PMPChecker_1_io_check_env_pmp_2_cfg_a),
    .io_check_env_pmp_2_cfg_w(PMPChecker_1_io_check_env_pmp_2_cfg_w),
    .io_check_env_pmp_2_cfg_r(PMPChecker_1_io_check_env_pmp_2_cfg_r),
    .io_check_env_pmp_2_addr(PMPChecker_1_io_check_env_pmp_2_addr),
    .io_check_env_pmp_2_mask(PMPChecker_1_io_check_env_pmp_2_mask),
    .io_check_env_pmp_3_cfg_l(PMPChecker_1_io_check_env_pmp_3_cfg_l),
    .io_check_env_pmp_3_cfg_a(PMPChecker_1_io_check_env_pmp_3_cfg_a),
    .io_check_env_pmp_3_cfg_w(PMPChecker_1_io_check_env_pmp_3_cfg_w),
    .io_check_env_pmp_3_cfg_r(PMPChecker_1_io_check_env_pmp_3_cfg_r),
    .io_check_env_pmp_3_addr(PMPChecker_1_io_check_env_pmp_3_addr),
    .io_check_env_pmp_3_mask(PMPChecker_1_io_check_env_pmp_3_mask),
    .io_check_env_pmp_4_cfg_l(PMPChecker_1_io_check_env_pmp_4_cfg_l),
    .io_check_env_pmp_4_cfg_a(PMPChecker_1_io_check_env_pmp_4_cfg_a),
    .io_check_env_pmp_4_cfg_w(PMPChecker_1_io_check_env_pmp_4_cfg_w),
    .io_check_env_pmp_4_cfg_r(PMPChecker_1_io_check_env_pmp_4_cfg_r),
    .io_check_env_pmp_4_addr(PMPChecker_1_io_check_env_pmp_4_addr),
    .io_check_env_pmp_4_mask(PMPChecker_1_io_check_env_pmp_4_mask),
    .io_check_env_pmp_5_cfg_l(PMPChecker_1_io_check_env_pmp_5_cfg_l),
    .io_check_env_pmp_5_cfg_a(PMPChecker_1_io_check_env_pmp_5_cfg_a),
    .io_check_env_pmp_5_cfg_w(PMPChecker_1_io_check_env_pmp_5_cfg_w),
    .io_check_env_pmp_5_cfg_r(PMPChecker_1_io_check_env_pmp_5_cfg_r),
    .io_check_env_pmp_5_addr(PMPChecker_1_io_check_env_pmp_5_addr),
    .io_check_env_pmp_5_mask(PMPChecker_1_io_check_env_pmp_5_mask),
    .io_check_env_pmp_6_cfg_l(PMPChecker_1_io_check_env_pmp_6_cfg_l),
    .io_check_env_pmp_6_cfg_a(PMPChecker_1_io_check_env_pmp_6_cfg_a),
    .io_check_env_pmp_6_cfg_w(PMPChecker_1_io_check_env_pmp_6_cfg_w),
    .io_check_env_pmp_6_cfg_r(PMPChecker_1_io_check_env_pmp_6_cfg_r),
    .io_check_env_pmp_6_addr(PMPChecker_1_io_check_env_pmp_6_addr),
    .io_check_env_pmp_6_mask(PMPChecker_1_io_check_env_pmp_6_mask),
    .io_check_env_pmp_7_cfg_l(PMPChecker_1_io_check_env_pmp_7_cfg_l),
    .io_check_env_pmp_7_cfg_a(PMPChecker_1_io_check_env_pmp_7_cfg_a),
    .io_check_env_pmp_7_cfg_w(PMPChecker_1_io_check_env_pmp_7_cfg_w),
    .io_check_env_pmp_7_cfg_r(PMPChecker_1_io_check_env_pmp_7_cfg_r),
    .io_check_env_pmp_7_addr(PMPChecker_1_io_check_env_pmp_7_addr),
    .io_check_env_pmp_7_mask(PMPChecker_1_io_check_env_pmp_7_mask),
    .io_check_env_pmp_8_cfg_l(PMPChecker_1_io_check_env_pmp_8_cfg_l),
    .io_check_env_pmp_8_cfg_a(PMPChecker_1_io_check_env_pmp_8_cfg_a),
    .io_check_env_pmp_8_cfg_w(PMPChecker_1_io_check_env_pmp_8_cfg_w),
    .io_check_env_pmp_8_cfg_r(PMPChecker_1_io_check_env_pmp_8_cfg_r),
    .io_check_env_pmp_8_addr(PMPChecker_1_io_check_env_pmp_8_addr),
    .io_check_env_pmp_8_mask(PMPChecker_1_io_check_env_pmp_8_mask),
    .io_check_env_pmp_9_cfg_l(PMPChecker_1_io_check_env_pmp_9_cfg_l),
    .io_check_env_pmp_9_cfg_a(PMPChecker_1_io_check_env_pmp_9_cfg_a),
    .io_check_env_pmp_9_cfg_w(PMPChecker_1_io_check_env_pmp_9_cfg_w),
    .io_check_env_pmp_9_cfg_r(PMPChecker_1_io_check_env_pmp_9_cfg_r),
    .io_check_env_pmp_9_addr(PMPChecker_1_io_check_env_pmp_9_addr),
    .io_check_env_pmp_9_mask(PMPChecker_1_io_check_env_pmp_9_mask),
    .io_check_env_pmp_10_cfg_l(PMPChecker_1_io_check_env_pmp_10_cfg_l),
    .io_check_env_pmp_10_cfg_a(PMPChecker_1_io_check_env_pmp_10_cfg_a),
    .io_check_env_pmp_10_cfg_w(PMPChecker_1_io_check_env_pmp_10_cfg_w),
    .io_check_env_pmp_10_cfg_r(PMPChecker_1_io_check_env_pmp_10_cfg_r),
    .io_check_env_pmp_10_addr(PMPChecker_1_io_check_env_pmp_10_addr),
    .io_check_env_pmp_10_mask(PMPChecker_1_io_check_env_pmp_10_mask),
    .io_check_env_pmp_11_cfg_l(PMPChecker_1_io_check_env_pmp_11_cfg_l),
    .io_check_env_pmp_11_cfg_a(PMPChecker_1_io_check_env_pmp_11_cfg_a),
    .io_check_env_pmp_11_cfg_w(PMPChecker_1_io_check_env_pmp_11_cfg_w),
    .io_check_env_pmp_11_cfg_r(PMPChecker_1_io_check_env_pmp_11_cfg_r),
    .io_check_env_pmp_11_addr(PMPChecker_1_io_check_env_pmp_11_addr),
    .io_check_env_pmp_11_mask(PMPChecker_1_io_check_env_pmp_11_mask),
    .io_check_env_pmp_12_cfg_l(PMPChecker_1_io_check_env_pmp_12_cfg_l),
    .io_check_env_pmp_12_cfg_a(PMPChecker_1_io_check_env_pmp_12_cfg_a),
    .io_check_env_pmp_12_cfg_w(PMPChecker_1_io_check_env_pmp_12_cfg_w),
    .io_check_env_pmp_12_cfg_r(PMPChecker_1_io_check_env_pmp_12_cfg_r),
    .io_check_env_pmp_12_addr(PMPChecker_1_io_check_env_pmp_12_addr),
    .io_check_env_pmp_12_mask(PMPChecker_1_io_check_env_pmp_12_mask),
    .io_check_env_pmp_13_cfg_l(PMPChecker_1_io_check_env_pmp_13_cfg_l),
    .io_check_env_pmp_13_cfg_a(PMPChecker_1_io_check_env_pmp_13_cfg_a),
    .io_check_env_pmp_13_cfg_w(PMPChecker_1_io_check_env_pmp_13_cfg_w),
    .io_check_env_pmp_13_cfg_r(PMPChecker_1_io_check_env_pmp_13_cfg_r),
    .io_check_env_pmp_13_addr(PMPChecker_1_io_check_env_pmp_13_addr),
    .io_check_env_pmp_13_mask(PMPChecker_1_io_check_env_pmp_13_mask),
    .io_check_env_pmp_14_cfg_l(PMPChecker_1_io_check_env_pmp_14_cfg_l),
    .io_check_env_pmp_14_cfg_a(PMPChecker_1_io_check_env_pmp_14_cfg_a),
    .io_check_env_pmp_14_cfg_w(PMPChecker_1_io_check_env_pmp_14_cfg_w),
    .io_check_env_pmp_14_cfg_r(PMPChecker_1_io_check_env_pmp_14_cfg_r),
    .io_check_env_pmp_14_addr(PMPChecker_1_io_check_env_pmp_14_addr),
    .io_check_env_pmp_14_mask(PMPChecker_1_io_check_env_pmp_14_mask),
    .io_check_env_pmp_15_cfg_l(PMPChecker_1_io_check_env_pmp_15_cfg_l),
    .io_check_env_pmp_15_cfg_a(PMPChecker_1_io_check_env_pmp_15_cfg_a),
    .io_check_env_pmp_15_cfg_w(PMPChecker_1_io_check_env_pmp_15_cfg_w),
    .io_check_env_pmp_15_cfg_r(PMPChecker_1_io_check_env_pmp_15_cfg_r),
    .io_check_env_pmp_15_addr(PMPChecker_1_io_check_env_pmp_15_addr),
    .io_check_env_pmp_15_mask(PMPChecker_1_io_check_env_pmp_15_mask),
    .io_check_env_pma_0_cfg_c(PMPChecker_1_io_check_env_pma_0_cfg_c),
    .io_check_env_pma_0_cfg_atomic(PMPChecker_1_io_check_env_pma_0_cfg_atomic),
    .io_check_env_pma_0_cfg_a(PMPChecker_1_io_check_env_pma_0_cfg_a),
    .io_check_env_pma_0_cfg_w(PMPChecker_1_io_check_env_pma_0_cfg_w),
    .io_check_env_pma_0_cfg_r(PMPChecker_1_io_check_env_pma_0_cfg_r),
    .io_check_env_pma_0_addr(PMPChecker_1_io_check_env_pma_0_addr),
    .io_check_env_pma_0_mask(PMPChecker_1_io_check_env_pma_0_mask),
    .io_check_env_pma_1_cfg_c(PMPChecker_1_io_check_env_pma_1_cfg_c),
    .io_check_env_pma_1_cfg_atomic(PMPChecker_1_io_check_env_pma_1_cfg_atomic),
    .io_check_env_pma_1_cfg_a(PMPChecker_1_io_check_env_pma_1_cfg_a),
    .io_check_env_pma_1_cfg_w(PMPChecker_1_io_check_env_pma_1_cfg_w),
    .io_check_env_pma_1_cfg_r(PMPChecker_1_io_check_env_pma_1_cfg_r),
    .io_check_env_pma_1_addr(PMPChecker_1_io_check_env_pma_1_addr),
    .io_check_env_pma_1_mask(PMPChecker_1_io_check_env_pma_1_mask),
    .io_check_env_pma_2_cfg_c(PMPChecker_1_io_check_env_pma_2_cfg_c),
    .io_check_env_pma_2_cfg_atomic(PMPChecker_1_io_check_env_pma_2_cfg_atomic),
    .io_check_env_pma_2_cfg_a(PMPChecker_1_io_check_env_pma_2_cfg_a),
    .io_check_env_pma_2_cfg_w(PMPChecker_1_io_check_env_pma_2_cfg_w),
    .io_check_env_pma_2_cfg_r(PMPChecker_1_io_check_env_pma_2_cfg_r),
    .io_check_env_pma_2_addr(PMPChecker_1_io_check_env_pma_2_addr),
    .io_check_env_pma_2_mask(PMPChecker_1_io_check_env_pma_2_mask),
    .io_check_env_pma_3_cfg_c(PMPChecker_1_io_check_env_pma_3_cfg_c),
    .io_check_env_pma_3_cfg_atomic(PMPChecker_1_io_check_env_pma_3_cfg_atomic),
    .io_check_env_pma_3_cfg_a(PMPChecker_1_io_check_env_pma_3_cfg_a),
    .io_check_env_pma_3_cfg_w(PMPChecker_1_io_check_env_pma_3_cfg_w),
    .io_check_env_pma_3_cfg_r(PMPChecker_1_io_check_env_pma_3_cfg_r),
    .io_check_env_pma_3_addr(PMPChecker_1_io_check_env_pma_3_addr),
    .io_check_env_pma_3_mask(PMPChecker_1_io_check_env_pma_3_mask),
    .io_check_env_pma_4_cfg_c(PMPChecker_1_io_check_env_pma_4_cfg_c),
    .io_check_env_pma_4_cfg_atomic(PMPChecker_1_io_check_env_pma_4_cfg_atomic),
    .io_check_env_pma_4_cfg_a(PMPChecker_1_io_check_env_pma_4_cfg_a),
    .io_check_env_pma_4_cfg_w(PMPChecker_1_io_check_env_pma_4_cfg_w),
    .io_check_env_pma_4_cfg_r(PMPChecker_1_io_check_env_pma_4_cfg_r),
    .io_check_env_pma_4_addr(PMPChecker_1_io_check_env_pma_4_addr),
    .io_check_env_pma_4_mask(PMPChecker_1_io_check_env_pma_4_mask),
    .io_check_env_pma_5_cfg_c(PMPChecker_1_io_check_env_pma_5_cfg_c),
    .io_check_env_pma_5_cfg_atomic(PMPChecker_1_io_check_env_pma_5_cfg_atomic),
    .io_check_env_pma_5_cfg_a(PMPChecker_1_io_check_env_pma_5_cfg_a),
    .io_check_env_pma_5_cfg_w(PMPChecker_1_io_check_env_pma_5_cfg_w),
    .io_check_env_pma_5_cfg_r(PMPChecker_1_io_check_env_pma_5_cfg_r),
    .io_check_env_pma_5_addr(PMPChecker_1_io_check_env_pma_5_addr),
    .io_check_env_pma_5_mask(PMPChecker_1_io_check_env_pma_5_mask),
    .io_check_env_pma_6_cfg_c(PMPChecker_1_io_check_env_pma_6_cfg_c),
    .io_check_env_pma_6_cfg_atomic(PMPChecker_1_io_check_env_pma_6_cfg_atomic),
    .io_check_env_pma_6_cfg_a(PMPChecker_1_io_check_env_pma_6_cfg_a),
    .io_check_env_pma_6_cfg_w(PMPChecker_1_io_check_env_pma_6_cfg_w),
    .io_check_env_pma_6_cfg_r(PMPChecker_1_io_check_env_pma_6_cfg_r),
    .io_check_env_pma_6_addr(PMPChecker_1_io_check_env_pma_6_addr),
    .io_check_env_pma_6_mask(PMPChecker_1_io_check_env_pma_6_mask),
    .io_check_env_pma_7_cfg_c(PMPChecker_1_io_check_env_pma_7_cfg_c),
    .io_check_env_pma_7_cfg_atomic(PMPChecker_1_io_check_env_pma_7_cfg_atomic),
    .io_check_env_pma_7_cfg_a(PMPChecker_1_io_check_env_pma_7_cfg_a),
    .io_check_env_pma_7_cfg_w(PMPChecker_1_io_check_env_pma_7_cfg_w),
    .io_check_env_pma_7_cfg_r(PMPChecker_1_io_check_env_pma_7_cfg_r),
    .io_check_env_pma_7_addr(PMPChecker_1_io_check_env_pma_7_addr),
    .io_check_env_pma_7_mask(PMPChecker_1_io_check_env_pma_7_mask),
    .io_check_env_pma_8_cfg_c(PMPChecker_1_io_check_env_pma_8_cfg_c),
    .io_check_env_pma_8_cfg_atomic(PMPChecker_1_io_check_env_pma_8_cfg_atomic),
    .io_check_env_pma_8_cfg_a(PMPChecker_1_io_check_env_pma_8_cfg_a),
    .io_check_env_pma_8_cfg_w(PMPChecker_1_io_check_env_pma_8_cfg_w),
    .io_check_env_pma_8_cfg_r(PMPChecker_1_io_check_env_pma_8_cfg_r),
    .io_check_env_pma_8_addr(PMPChecker_1_io_check_env_pma_8_addr),
    .io_check_env_pma_8_mask(PMPChecker_1_io_check_env_pma_8_mask),
    .io_check_env_pma_9_cfg_c(PMPChecker_1_io_check_env_pma_9_cfg_c),
    .io_check_env_pma_9_cfg_atomic(PMPChecker_1_io_check_env_pma_9_cfg_atomic),
    .io_check_env_pma_9_cfg_a(PMPChecker_1_io_check_env_pma_9_cfg_a),
    .io_check_env_pma_9_cfg_w(PMPChecker_1_io_check_env_pma_9_cfg_w),
    .io_check_env_pma_9_cfg_r(PMPChecker_1_io_check_env_pma_9_cfg_r),
    .io_check_env_pma_9_addr(PMPChecker_1_io_check_env_pma_9_addr),
    .io_check_env_pma_9_mask(PMPChecker_1_io_check_env_pma_9_mask),
    .io_check_env_pma_10_cfg_c(PMPChecker_1_io_check_env_pma_10_cfg_c),
    .io_check_env_pma_10_cfg_atomic(PMPChecker_1_io_check_env_pma_10_cfg_atomic),
    .io_check_env_pma_10_cfg_a(PMPChecker_1_io_check_env_pma_10_cfg_a),
    .io_check_env_pma_10_cfg_w(PMPChecker_1_io_check_env_pma_10_cfg_w),
    .io_check_env_pma_10_cfg_r(PMPChecker_1_io_check_env_pma_10_cfg_r),
    .io_check_env_pma_10_addr(PMPChecker_1_io_check_env_pma_10_addr),
    .io_check_env_pma_10_mask(PMPChecker_1_io_check_env_pma_10_mask),
    .io_check_env_pma_11_cfg_c(PMPChecker_1_io_check_env_pma_11_cfg_c),
    .io_check_env_pma_11_cfg_atomic(PMPChecker_1_io_check_env_pma_11_cfg_atomic),
    .io_check_env_pma_11_cfg_a(PMPChecker_1_io_check_env_pma_11_cfg_a),
    .io_check_env_pma_11_cfg_w(PMPChecker_1_io_check_env_pma_11_cfg_w),
    .io_check_env_pma_11_cfg_r(PMPChecker_1_io_check_env_pma_11_cfg_r),
    .io_check_env_pma_11_addr(PMPChecker_1_io_check_env_pma_11_addr),
    .io_check_env_pma_11_mask(PMPChecker_1_io_check_env_pma_11_mask),
    .io_check_env_pma_12_cfg_c(PMPChecker_1_io_check_env_pma_12_cfg_c),
    .io_check_env_pma_12_cfg_atomic(PMPChecker_1_io_check_env_pma_12_cfg_atomic),
    .io_check_env_pma_12_cfg_a(PMPChecker_1_io_check_env_pma_12_cfg_a),
    .io_check_env_pma_12_cfg_w(PMPChecker_1_io_check_env_pma_12_cfg_w),
    .io_check_env_pma_12_cfg_r(PMPChecker_1_io_check_env_pma_12_cfg_r),
    .io_check_env_pma_12_addr(PMPChecker_1_io_check_env_pma_12_addr),
    .io_check_env_pma_12_mask(PMPChecker_1_io_check_env_pma_12_mask),
    .io_check_env_pma_13_cfg_c(PMPChecker_1_io_check_env_pma_13_cfg_c),
    .io_check_env_pma_13_cfg_atomic(PMPChecker_1_io_check_env_pma_13_cfg_atomic),
    .io_check_env_pma_13_cfg_a(PMPChecker_1_io_check_env_pma_13_cfg_a),
    .io_check_env_pma_13_cfg_w(PMPChecker_1_io_check_env_pma_13_cfg_w),
    .io_check_env_pma_13_cfg_r(PMPChecker_1_io_check_env_pma_13_cfg_r),
    .io_check_env_pma_13_addr(PMPChecker_1_io_check_env_pma_13_addr),
    .io_check_env_pma_13_mask(PMPChecker_1_io_check_env_pma_13_mask),
    .io_check_env_pma_14_cfg_c(PMPChecker_1_io_check_env_pma_14_cfg_c),
    .io_check_env_pma_14_cfg_atomic(PMPChecker_1_io_check_env_pma_14_cfg_atomic),
    .io_check_env_pma_14_cfg_a(PMPChecker_1_io_check_env_pma_14_cfg_a),
    .io_check_env_pma_14_cfg_w(PMPChecker_1_io_check_env_pma_14_cfg_w),
    .io_check_env_pma_14_cfg_r(PMPChecker_1_io_check_env_pma_14_cfg_r),
    .io_check_env_pma_14_addr(PMPChecker_1_io_check_env_pma_14_addr),
    .io_check_env_pma_14_mask(PMPChecker_1_io_check_env_pma_14_mask),
    .io_check_env_pma_15_cfg_c(PMPChecker_1_io_check_env_pma_15_cfg_c),
    .io_check_env_pma_15_cfg_atomic(PMPChecker_1_io_check_env_pma_15_cfg_atomic),
    .io_check_env_pma_15_cfg_a(PMPChecker_1_io_check_env_pma_15_cfg_a),
    .io_check_env_pma_15_cfg_w(PMPChecker_1_io_check_env_pma_15_cfg_w),
    .io_check_env_pma_15_cfg_r(PMPChecker_1_io_check_env_pma_15_cfg_r),
    .io_check_env_pma_15_addr(PMPChecker_1_io_check_env_pma_15_addr),
    .io_check_env_pma_15_mask(PMPChecker_1_io_check_env_pma_15_mask),
    .io_req_valid(PMPChecker_1_io_req_valid),
    .io_req_bits_addr(PMPChecker_1_io_req_bits_addr),
    .io_req_bits_cmd(PMPChecker_1_io_req_bits_cmd),
    .io_resp_ld(PMPChecker_1_io_resp_ld),
    .io_resp_st(PMPChecker_1_io_resp_st),
    .io_resp_mmio(PMPChecker_1_io_resp_mmio),
    .io_resp_atomic(PMPChecker_1_io_resp_atomic)
  );
  PMPChecker_8 PMPChecker_2 ( // @[MemBlock.scala 314:91]
    .clock(PMPChecker_2_clock),
    .io_check_env_mode(PMPChecker_2_io_check_env_mode),
    .io_check_env_pmp_0_cfg_l(PMPChecker_2_io_check_env_pmp_0_cfg_l),
    .io_check_env_pmp_0_cfg_a(PMPChecker_2_io_check_env_pmp_0_cfg_a),
    .io_check_env_pmp_0_cfg_w(PMPChecker_2_io_check_env_pmp_0_cfg_w),
    .io_check_env_pmp_0_cfg_r(PMPChecker_2_io_check_env_pmp_0_cfg_r),
    .io_check_env_pmp_0_addr(PMPChecker_2_io_check_env_pmp_0_addr),
    .io_check_env_pmp_0_mask(PMPChecker_2_io_check_env_pmp_0_mask),
    .io_check_env_pmp_1_cfg_l(PMPChecker_2_io_check_env_pmp_1_cfg_l),
    .io_check_env_pmp_1_cfg_a(PMPChecker_2_io_check_env_pmp_1_cfg_a),
    .io_check_env_pmp_1_cfg_w(PMPChecker_2_io_check_env_pmp_1_cfg_w),
    .io_check_env_pmp_1_cfg_r(PMPChecker_2_io_check_env_pmp_1_cfg_r),
    .io_check_env_pmp_1_addr(PMPChecker_2_io_check_env_pmp_1_addr),
    .io_check_env_pmp_1_mask(PMPChecker_2_io_check_env_pmp_1_mask),
    .io_check_env_pmp_2_cfg_l(PMPChecker_2_io_check_env_pmp_2_cfg_l),
    .io_check_env_pmp_2_cfg_a(PMPChecker_2_io_check_env_pmp_2_cfg_a),
    .io_check_env_pmp_2_cfg_w(PMPChecker_2_io_check_env_pmp_2_cfg_w),
    .io_check_env_pmp_2_cfg_r(PMPChecker_2_io_check_env_pmp_2_cfg_r),
    .io_check_env_pmp_2_addr(PMPChecker_2_io_check_env_pmp_2_addr),
    .io_check_env_pmp_2_mask(PMPChecker_2_io_check_env_pmp_2_mask),
    .io_check_env_pmp_3_cfg_l(PMPChecker_2_io_check_env_pmp_3_cfg_l),
    .io_check_env_pmp_3_cfg_a(PMPChecker_2_io_check_env_pmp_3_cfg_a),
    .io_check_env_pmp_3_cfg_w(PMPChecker_2_io_check_env_pmp_3_cfg_w),
    .io_check_env_pmp_3_cfg_r(PMPChecker_2_io_check_env_pmp_3_cfg_r),
    .io_check_env_pmp_3_addr(PMPChecker_2_io_check_env_pmp_3_addr),
    .io_check_env_pmp_3_mask(PMPChecker_2_io_check_env_pmp_3_mask),
    .io_check_env_pmp_4_cfg_l(PMPChecker_2_io_check_env_pmp_4_cfg_l),
    .io_check_env_pmp_4_cfg_a(PMPChecker_2_io_check_env_pmp_4_cfg_a),
    .io_check_env_pmp_4_cfg_w(PMPChecker_2_io_check_env_pmp_4_cfg_w),
    .io_check_env_pmp_4_cfg_r(PMPChecker_2_io_check_env_pmp_4_cfg_r),
    .io_check_env_pmp_4_addr(PMPChecker_2_io_check_env_pmp_4_addr),
    .io_check_env_pmp_4_mask(PMPChecker_2_io_check_env_pmp_4_mask),
    .io_check_env_pmp_5_cfg_l(PMPChecker_2_io_check_env_pmp_5_cfg_l),
    .io_check_env_pmp_5_cfg_a(PMPChecker_2_io_check_env_pmp_5_cfg_a),
    .io_check_env_pmp_5_cfg_w(PMPChecker_2_io_check_env_pmp_5_cfg_w),
    .io_check_env_pmp_5_cfg_r(PMPChecker_2_io_check_env_pmp_5_cfg_r),
    .io_check_env_pmp_5_addr(PMPChecker_2_io_check_env_pmp_5_addr),
    .io_check_env_pmp_5_mask(PMPChecker_2_io_check_env_pmp_5_mask),
    .io_check_env_pmp_6_cfg_l(PMPChecker_2_io_check_env_pmp_6_cfg_l),
    .io_check_env_pmp_6_cfg_a(PMPChecker_2_io_check_env_pmp_6_cfg_a),
    .io_check_env_pmp_6_cfg_w(PMPChecker_2_io_check_env_pmp_6_cfg_w),
    .io_check_env_pmp_6_cfg_r(PMPChecker_2_io_check_env_pmp_6_cfg_r),
    .io_check_env_pmp_6_addr(PMPChecker_2_io_check_env_pmp_6_addr),
    .io_check_env_pmp_6_mask(PMPChecker_2_io_check_env_pmp_6_mask),
    .io_check_env_pmp_7_cfg_l(PMPChecker_2_io_check_env_pmp_7_cfg_l),
    .io_check_env_pmp_7_cfg_a(PMPChecker_2_io_check_env_pmp_7_cfg_a),
    .io_check_env_pmp_7_cfg_w(PMPChecker_2_io_check_env_pmp_7_cfg_w),
    .io_check_env_pmp_7_cfg_r(PMPChecker_2_io_check_env_pmp_7_cfg_r),
    .io_check_env_pmp_7_addr(PMPChecker_2_io_check_env_pmp_7_addr),
    .io_check_env_pmp_7_mask(PMPChecker_2_io_check_env_pmp_7_mask),
    .io_check_env_pmp_8_cfg_l(PMPChecker_2_io_check_env_pmp_8_cfg_l),
    .io_check_env_pmp_8_cfg_a(PMPChecker_2_io_check_env_pmp_8_cfg_a),
    .io_check_env_pmp_8_cfg_w(PMPChecker_2_io_check_env_pmp_8_cfg_w),
    .io_check_env_pmp_8_cfg_r(PMPChecker_2_io_check_env_pmp_8_cfg_r),
    .io_check_env_pmp_8_addr(PMPChecker_2_io_check_env_pmp_8_addr),
    .io_check_env_pmp_8_mask(PMPChecker_2_io_check_env_pmp_8_mask),
    .io_check_env_pmp_9_cfg_l(PMPChecker_2_io_check_env_pmp_9_cfg_l),
    .io_check_env_pmp_9_cfg_a(PMPChecker_2_io_check_env_pmp_9_cfg_a),
    .io_check_env_pmp_9_cfg_w(PMPChecker_2_io_check_env_pmp_9_cfg_w),
    .io_check_env_pmp_9_cfg_r(PMPChecker_2_io_check_env_pmp_9_cfg_r),
    .io_check_env_pmp_9_addr(PMPChecker_2_io_check_env_pmp_9_addr),
    .io_check_env_pmp_9_mask(PMPChecker_2_io_check_env_pmp_9_mask),
    .io_check_env_pmp_10_cfg_l(PMPChecker_2_io_check_env_pmp_10_cfg_l),
    .io_check_env_pmp_10_cfg_a(PMPChecker_2_io_check_env_pmp_10_cfg_a),
    .io_check_env_pmp_10_cfg_w(PMPChecker_2_io_check_env_pmp_10_cfg_w),
    .io_check_env_pmp_10_cfg_r(PMPChecker_2_io_check_env_pmp_10_cfg_r),
    .io_check_env_pmp_10_addr(PMPChecker_2_io_check_env_pmp_10_addr),
    .io_check_env_pmp_10_mask(PMPChecker_2_io_check_env_pmp_10_mask),
    .io_check_env_pmp_11_cfg_l(PMPChecker_2_io_check_env_pmp_11_cfg_l),
    .io_check_env_pmp_11_cfg_a(PMPChecker_2_io_check_env_pmp_11_cfg_a),
    .io_check_env_pmp_11_cfg_w(PMPChecker_2_io_check_env_pmp_11_cfg_w),
    .io_check_env_pmp_11_cfg_r(PMPChecker_2_io_check_env_pmp_11_cfg_r),
    .io_check_env_pmp_11_addr(PMPChecker_2_io_check_env_pmp_11_addr),
    .io_check_env_pmp_11_mask(PMPChecker_2_io_check_env_pmp_11_mask),
    .io_check_env_pmp_12_cfg_l(PMPChecker_2_io_check_env_pmp_12_cfg_l),
    .io_check_env_pmp_12_cfg_a(PMPChecker_2_io_check_env_pmp_12_cfg_a),
    .io_check_env_pmp_12_cfg_w(PMPChecker_2_io_check_env_pmp_12_cfg_w),
    .io_check_env_pmp_12_cfg_r(PMPChecker_2_io_check_env_pmp_12_cfg_r),
    .io_check_env_pmp_12_addr(PMPChecker_2_io_check_env_pmp_12_addr),
    .io_check_env_pmp_12_mask(PMPChecker_2_io_check_env_pmp_12_mask),
    .io_check_env_pmp_13_cfg_l(PMPChecker_2_io_check_env_pmp_13_cfg_l),
    .io_check_env_pmp_13_cfg_a(PMPChecker_2_io_check_env_pmp_13_cfg_a),
    .io_check_env_pmp_13_cfg_w(PMPChecker_2_io_check_env_pmp_13_cfg_w),
    .io_check_env_pmp_13_cfg_r(PMPChecker_2_io_check_env_pmp_13_cfg_r),
    .io_check_env_pmp_13_addr(PMPChecker_2_io_check_env_pmp_13_addr),
    .io_check_env_pmp_13_mask(PMPChecker_2_io_check_env_pmp_13_mask),
    .io_check_env_pmp_14_cfg_l(PMPChecker_2_io_check_env_pmp_14_cfg_l),
    .io_check_env_pmp_14_cfg_a(PMPChecker_2_io_check_env_pmp_14_cfg_a),
    .io_check_env_pmp_14_cfg_w(PMPChecker_2_io_check_env_pmp_14_cfg_w),
    .io_check_env_pmp_14_cfg_r(PMPChecker_2_io_check_env_pmp_14_cfg_r),
    .io_check_env_pmp_14_addr(PMPChecker_2_io_check_env_pmp_14_addr),
    .io_check_env_pmp_14_mask(PMPChecker_2_io_check_env_pmp_14_mask),
    .io_check_env_pmp_15_cfg_l(PMPChecker_2_io_check_env_pmp_15_cfg_l),
    .io_check_env_pmp_15_cfg_a(PMPChecker_2_io_check_env_pmp_15_cfg_a),
    .io_check_env_pmp_15_cfg_w(PMPChecker_2_io_check_env_pmp_15_cfg_w),
    .io_check_env_pmp_15_cfg_r(PMPChecker_2_io_check_env_pmp_15_cfg_r),
    .io_check_env_pmp_15_addr(PMPChecker_2_io_check_env_pmp_15_addr),
    .io_check_env_pmp_15_mask(PMPChecker_2_io_check_env_pmp_15_mask),
    .io_check_env_pma_0_cfg_c(PMPChecker_2_io_check_env_pma_0_cfg_c),
    .io_check_env_pma_0_cfg_atomic(PMPChecker_2_io_check_env_pma_0_cfg_atomic),
    .io_check_env_pma_0_cfg_a(PMPChecker_2_io_check_env_pma_0_cfg_a),
    .io_check_env_pma_0_cfg_w(PMPChecker_2_io_check_env_pma_0_cfg_w),
    .io_check_env_pma_0_cfg_r(PMPChecker_2_io_check_env_pma_0_cfg_r),
    .io_check_env_pma_0_addr(PMPChecker_2_io_check_env_pma_0_addr),
    .io_check_env_pma_0_mask(PMPChecker_2_io_check_env_pma_0_mask),
    .io_check_env_pma_1_cfg_c(PMPChecker_2_io_check_env_pma_1_cfg_c),
    .io_check_env_pma_1_cfg_atomic(PMPChecker_2_io_check_env_pma_1_cfg_atomic),
    .io_check_env_pma_1_cfg_a(PMPChecker_2_io_check_env_pma_1_cfg_a),
    .io_check_env_pma_1_cfg_w(PMPChecker_2_io_check_env_pma_1_cfg_w),
    .io_check_env_pma_1_cfg_r(PMPChecker_2_io_check_env_pma_1_cfg_r),
    .io_check_env_pma_1_addr(PMPChecker_2_io_check_env_pma_1_addr),
    .io_check_env_pma_1_mask(PMPChecker_2_io_check_env_pma_1_mask),
    .io_check_env_pma_2_cfg_c(PMPChecker_2_io_check_env_pma_2_cfg_c),
    .io_check_env_pma_2_cfg_atomic(PMPChecker_2_io_check_env_pma_2_cfg_atomic),
    .io_check_env_pma_2_cfg_a(PMPChecker_2_io_check_env_pma_2_cfg_a),
    .io_check_env_pma_2_cfg_w(PMPChecker_2_io_check_env_pma_2_cfg_w),
    .io_check_env_pma_2_cfg_r(PMPChecker_2_io_check_env_pma_2_cfg_r),
    .io_check_env_pma_2_addr(PMPChecker_2_io_check_env_pma_2_addr),
    .io_check_env_pma_2_mask(PMPChecker_2_io_check_env_pma_2_mask),
    .io_check_env_pma_3_cfg_c(PMPChecker_2_io_check_env_pma_3_cfg_c),
    .io_check_env_pma_3_cfg_atomic(PMPChecker_2_io_check_env_pma_3_cfg_atomic),
    .io_check_env_pma_3_cfg_a(PMPChecker_2_io_check_env_pma_3_cfg_a),
    .io_check_env_pma_3_cfg_w(PMPChecker_2_io_check_env_pma_3_cfg_w),
    .io_check_env_pma_3_cfg_r(PMPChecker_2_io_check_env_pma_3_cfg_r),
    .io_check_env_pma_3_addr(PMPChecker_2_io_check_env_pma_3_addr),
    .io_check_env_pma_3_mask(PMPChecker_2_io_check_env_pma_3_mask),
    .io_check_env_pma_4_cfg_c(PMPChecker_2_io_check_env_pma_4_cfg_c),
    .io_check_env_pma_4_cfg_atomic(PMPChecker_2_io_check_env_pma_4_cfg_atomic),
    .io_check_env_pma_4_cfg_a(PMPChecker_2_io_check_env_pma_4_cfg_a),
    .io_check_env_pma_4_cfg_w(PMPChecker_2_io_check_env_pma_4_cfg_w),
    .io_check_env_pma_4_cfg_r(PMPChecker_2_io_check_env_pma_4_cfg_r),
    .io_check_env_pma_4_addr(PMPChecker_2_io_check_env_pma_4_addr),
    .io_check_env_pma_4_mask(PMPChecker_2_io_check_env_pma_4_mask),
    .io_check_env_pma_5_cfg_c(PMPChecker_2_io_check_env_pma_5_cfg_c),
    .io_check_env_pma_5_cfg_atomic(PMPChecker_2_io_check_env_pma_5_cfg_atomic),
    .io_check_env_pma_5_cfg_a(PMPChecker_2_io_check_env_pma_5_cfg_a),
    .io_check_env_pma_5_cfg_w(PMPChecker_2_io_check_env_pma_5_cfg_w),
    .io_check_env_pma_5_cfg_r(PMPChecker_2_io_check_env_pma_5_cfg_r),
    .io_check_env_pma_5_addr(PMPChecker_2_io_check_env_pma_5_addr),
    .io_check_env_pma_5_mask(PMPChecker_2_io_check_env_pma_5_mask),
    .io_check_env_pma_6_cfg_c(PMPChecker_2_io_check_env_pma_6_cfg_c),
    .io_check_env_pma_6_cfg_atomic(PMPChecker_2_io_check_env_pma_6_cfg_atomic),
    .io_check_env_pma_6_cfg_a(PMPChecker_2_io_check_env_pma_6_cfg_a),
    .io_check_env_pma_6_cfg_w(PMPChecker_2_io_check_env_pma_6_cfg_w),
    .io_check_env_pma_6_cfg_r(PMPChecker_2_io_check_env_pma_6_cfg_r),
    .io_check_env_pma_6_addr(PMPChecker_2_io_check_env_pma_6_addr),
    .io_check_env_pma_6_mask(PMPChecker_2_io_check_env_pma_6_mask),
    .io_check_env_pma_7_cfg_c(PMPChecker_2_io_check_env_pma_7_cfg_c),
    .io_check_env_pma_7_cfg_atomic(PMPChecker_2_io_check_env_pma_7_cfg_atomic),
    .io_check_env_pma_7_cfg_a(PMPChecker_2_io_check_env_pma_7_cfg_a),
    .io_check_env_pma_7_cfg_w(PMPChecker_2_io_check_env_pma_7_cfg_w),
    .io_check_env_pma_7_cfg_r(PMPChecker_2_io_check_env_pma_7_cfg_r),
    .io_check_env_pma_7_addr(PMPChecker_2_io_check_env_pma_7_addr),
    .io_check_env_pma_7_mask(PMPChecker_2_io_check_env_pma_7_mask),
    .io_check_env_pma_8_cfg_c(PMPChecker_2_io_check_env_pma_8_cfg_c),
    .io_check_env_pma_8_cfg_atomic(PMPChecker_2_io_check_env_pma_8_cfg_atomic),
    .io_check_env_pma_8_cfg_a(PMPChecker_2_io_check_env_pma_8_cfg_a),
    .io_check_env_pma_8_cfg_w(PMPChecker_2_io_check_env_pma_8_cfg_w),
    .io_check_env_pma_8_cfg_r(PMPChecker_2_io_check_env_pma_8_cfg_r),
    .io_check_env_pma_8_addr(PMPChecker_2_io_check_env_pma_8_addr),
    .io_check_env_pma_8_mask(PMPChecker_2_io_check_env_pma_8_mask),
    .io_check_env_pma_9_cfg_c(PMPChecker_2_io_check_env_pma_9_cfg_c),
    .io_check_env_pma_9_cfg_atomic(PMPChecker_2_io_check_env_pma_9_cfg_atomic),
    .io_check_env_pma_9_cfg_a(PMPChecker_2_io_check_env_pma_9_cfg_a),
    .io_check_env_pma_9_cfg_w(PMPChecker_2_io_check_env_pma_9_cfg_w),
    .io_check_env_pma_9_cfg_r(PMPChecker_2_io_check_env_pma_9_cfg_r),
    .io_check_env_pma_9_addr(PMPChecker_2_io_check_env_pma_9_addr),
    .io_check_env_pma_9_mask(PMPChecker_2_io_check_env_pma_9_mask),
    .io_check_env_pma_10_cfg_c(PMPChecker_2_io_check_env_pma_10_cfg_c),
    .io_check_env_pma_10_cfg_atomic(PMPChecker_2_io_check_env_pma_10_cfg_atomic),
    .io_check_env_pma_10_cfg_a(PMPChecker_2_io_check_env_pma_10_cfg_a),
    .io_check_env_pma_10_cfg_w(PMPChecker_2_io_check_env_pma_10_cfg_w),
    .io_check_env_pma_10_cfg_r(PMPChecker_2_io_check_env_pma_10_cfg_r),
    .io_check_env_pma_10_addr(PMPChecker_2_io_check_env_pma_10_addr),
    .io_check_env_pma_10_mask(PMPChecker_2_io_check_env_pma_10_mask),
    .io_check_env_pma_11_cfg_c(PMPChecker_2_io_check_env_pma_11_cfg_c),
    .io_check_env_pma_11_cfg_atomic(PMPChecker_2_io_check_env_pma_11_cfg_atomic),
    .io_check_env_pma_11_cfg_a(PMPChecker_2_io_check_env_pma_11_cfg_a),
    .io_check_env_pma_11_cfg_w(PMPChecker_2_io_check_env_pma_11_cfg_w),
    .io_check_env_pma_11_cfg_r(PMPChecker_2_io_check_env_pma_11_cfg_r),
    .io_check_env_pma_11_addr(PMPChecker_2_io_check_env_pma_11_addr),
    .io_check_env_pma_11_mask(PMPChecker_2_io_check_env_pma_11_mask),
    .io_check_env_pma_12_cfg_c(PMPChecker_2_io_check_env_pma_12_cfg_c),
    .io_check_env_pma_12_cfg_atomic(PMPChecker_2_io_check_env_pma_12_cfg_atomic),
    .io_check_env_pma_12_cfg_a(PMPChecker_2_io_check_env_pma_12_cfg_a),
    .io_check_env_pma_12_cfg_w(PMPChecker_2_io_check_env_pma_12_cfg_w),
    .io_check_env_pma_12_cfg_r(PMPChecker_2_io_check_env_pma_12_cfg_r),
    .io_check_env_pma_12_addr(PMPChecker_2_io_check_env_pma_12_addr),
    .io_check_env_pma_12_mask(PMPChecker_2_io_check_env_pma_12_mask),
    .io_check_env_pma_13_cfg_c(PMPChecker_2_io_check_env_pma_13_cfg_c),
    .io_check_env_pma_13_cfg_atomic(PMPChecker_2_io_check_env_pma_13_cfg_atomic),
    .io_check_env_pma_13_cfg_a(PMPChecker_2_io_check_env_pma_13_cfg_a),
    .io_check_env_pma_13_cfg_w(PMPChecker_2_io_check_env_pma_13_cfg_w),
    .io_check_env_pma_13_cfg_r(PMPChecker_2_io_check_env_pma_13_cfg_r),
    .io_check_env_pma_13_addr(PMPChecker_2_io_check_env_pma_13_addr),
    .io_check_env_pma_13_mask(PMPChecker_2_io_check_env_pma_13_mask),
    .io_check_env_pma_14_cfg_c(PMPChecker_2_io_check_env_pma_14_cfg_c),
    .io_check_env_pma_14_cfg_atomic(PMPChecker_2_io_check_env_pma_14_cfg_atomic),
    .io_check_env_pma_14_cfg_a(PMPChecker_2_io_check_env_pma_14_cfg_a),
    .io_check_env_pma_14_cfg_w(PMPChecker_2_io_check_env_pma_14_cfg_w),
    .io_check_env_pma_14_cfg_r(PMPChecker_2_io_check_env_pma_14_cfg_r),
    .io_check_env_pma_14_addr(PMPChecker_2_io_check_env_pma_14_addr),
    .io_check_env_pma_14_mask(PMPChecker_2_io_check_env_pma_14_mask),
    .io_check_env_pma_15_cfg_c(PMPChecker_2_io_check_env_pma_15_cfg_c),
    .io_check_env_pma_15_cfg_atomic(PMPChecker_2_io_check_env_pma_15_cfg_atomic),
    .io_check_env_pma_15_cfg_a(PMPChecker_2_io_check_env_pma_15_cfg_a),
    .io_check_env_pma_15_cfg_w(PMPChecker_2_io_check_env_pma_15_cfg_w),
    .io_check_env_pma_15_cfg_r(PMPChecker_2_io_check_env_pma_15_cfg_r),
    .io_check_env_pma_15_addr(PMPChecker_2_io_check_env_pma_15_addr),
    .io_check_env_pma_15_mask(PMPChecker_2_io_check_env_pma_15_mask),
    .io_req_valid(PMPChecker_2_io_req_valid),
    .io_req_bits_addr(PMPChecker_2_io_req_bits_addr),
    .io_req_bits_cmd(PMPChecker_2_io_req_bits_cmd),
    .io_resp_ld(PMPChecker_2_io_resp_ld),
    .io_resp_st(PMPChecker_2_io_resp_st),
    .io_resp_mmio(PMPChecker_2_io_resp_mmio),
    .io_resp_atomic(PMPChecker_2_io_resp_atomic)
  );
  PMPChecker_8 PMPChecker_3 ( // @[MemBlock.scala 314:91]
    .clock(PMPChecker_3_clock),
    .io_check_env_mode(PMPChecker_3_io_check_env_mode),
    .io_check_env_pmp_0_cfg_l(PMPChecker_3_io_check_env_pmp_0_cfg_l),
    .io_check_env_pmp_0_cfg_a(PMPChecker_3_io_check_env_pmp_0_cfg_a),
    .io_check_env_pmp_0_cfg_w(PMPChecker_3_io_check_env_pmp_0_cfg_w),
    .io_check_env_pmp_0_cfg_r(PMPChecker_3_io_check_env_pmp_0_cfg_r),
    .io_check_env_pmp_0_addr(PMPChecker_3_io_check_env_pmp_0_addr),
    .io_check_env_pmp_0_mask(PMPChecker_3_io_check_env_pmp_0_mask),
    .io_check_env_pmp_1_cfg_l(PMPChecker_3_io_check_env_pmp_1_cfg_l),
    .io_check_env_pmp_1_cfg_a(PMPChecker_3_io_check_env_pmp_1_cfg_a),
    .io_check_env_pmp_1_cfg_w(PMPChecker_3_io_check_env_pmp_1_cfg_w),
    .io_check_env_pmp_1_cfg_r(PMPChecker_3_io_check_env_pmp_1_cfg_r),
    .io_check_env_pmp_1_addr(PMPChecker_3_io_check_env_pmp_1_addr),
    .io_check_env_pmp_1_mask(PMPChecker_3_io_check_env_pmp_1_mask),
    .io_check_env_pmp_2_cfg_l(PMPChecker_3_io_check_env_pmp_2_cfg_l),
    .io_check_env_pmp_2_cfg_a(PMPChecker_3_io_check_env_pmp_2_cfg_a),
    .io_check_env_pmp_2_cfg_w(PMPChecker_3_io_check_env_pmp_2_cfg_w),
    .io_check_env_pmp_2_cfg_r(PMPChecker_3_io_check_env_pmp_2_cfg_r),
    .io_check_env_pmp_2_addr(PMPChecker_3_io_check_env_pmp_2_addr),
    .io_check_env_pmp_2_mask(PMPChecker_3_io_check_env_pmp_2_mask),
    .io_check_env_pmp_3_cfg_l(PMPChecker_3_io_check_env_pmp_3_cfg_l),
    .io_check_env_pmp_3_cfg_a(PMPChecker_3_io_check_env_pmp_3_cfg_a),
    .io_check_env_pmp_3_cfg_w(PMPChecker_3_io_check_env_pmp_3_cfg_w),
    .io_check_env_pmp_3_cfg_r(PMPChecker_3_io_check_env_pmp_3_cfg_r),
    .io_check_env_pmp_3_addr(PMPChecker_3_io_check_env_pmp_3_addr),
    .io_check_env_pmp_3_mask(PMPChecker_3_io_check_env_pmp_3_mask),
    .io_check_env_pmp_4_cfg_l(PMPChecker_3_io_check_env_pmp_4_cfg_l),
    .io_check_env_pmp_4_cfg_a(PMPChecker_3_io_check_env_pmp_4_cfg_a),
    .io_check_env_pmp_4_cfg_w(PMPChecker_3_io_check_env_pmp_4_cfg_w),
    .io_check_env_pmp_4_cfg_r(PMPChecker_3_io_check_env_pmp_4_cfg_r),
    .io_check_env_pmp_4_addr(PMPChecker_3_io_check_env_pmp_4_addr),
    .io_check_env_pmp_4_mask(PMPChecker_3_io_check_env_pmp_4_mask),
    .io_check_env_pmp_5_cfg_l(PMPChecker_3_io_check_env_pmp_5_cfg_l),
    .io_check_env_pmp_5_cfg_a(PMPChecker_3_io_check_env_pmp_5_cfg_a),
    .io_check_env_pmp_5_cfg_w(PMPChecker_3_io_check_env_pmp_5_cfg_w),
    .io_check_env_pmp_5_cfg_r(PMPChecker_3_io_check_env_pmp_5_cfg_r),
    .io_check_env_pmp_5_addr(PMPChecker_3_io_check_env_pmp_5_addr),
    .io_check_env_pmp_5_mask(PMPChecker_3_io_check_env_pmp_5_mask),
    .io_check_env_pmp_6_cfg_l(PMPChecker_3_io_check_env_pmp_6_cfg_l),
    .io_check_env_pmp_6_cfg_a(PMPChecker_3_io_check_env_pmp_6_cfg_a),
    .io_check_env_pmp_6_cfg_w(PMPChecker_3_io_check_env_pmp_6_cfg_w),
    .io_check_env_pmp_6_cfg_r(PMPChecker_3_io_check_env_pmp_6_cfg_r),
    .io_check_env_pmp_6_addr(PMPChecker_3_io_check_env_pmp_6_addr),
    .io_check_env_pmp_6_mask(PMPChecker_3_io_check_env_pmp_6_mask),
    .io_check_env_pmp_7_cfg_l(PMPChecker_3_io_check_env_pmp_7_cfg_l),
    .io_check_env_pmp_7_cfg_a(PMPChecker_3_io_check_env_pmp_7_cfg_a),
    .io_check_env_pmp_7_cfg_w(PMPChecker_3_io_check_env_pmp_7_cfg_w),
    .io_check_env_pmp_7_cfg_r(PMPChecker_3_io_check_env_pmp_7_cfg_r),
    .io_check_env_pmp_7_addr(PMPChecker_3_io_check_env_pmp_7_addr),
    .io_check_env_pmp_7_mask(PMPChecker_3_io_check_env_pmp_7_mask),
    .io_check_env_pmp_8_cfg_l(PMPChecker_3_io_check_env_pmp_8_cfg_l),
    .io_check_env_pmp_8_cfg_a(PMPChecker_3_io_check_env_pmp_8_cfg_a),
    .io_check_env_pmp_8_cfg_w(PMPChecker_3_io_check_env_pmp_8_cfg_w),
    .io_check_env_pmp_8_cfg_r(PMPChecker_3_io_check_env_pmp_8_cfg_r),
    .io_check_env_pmp_8_addr(PMPChecker_3_io_check_env_pmp_8_addr),
    .io_check_env_pmp_8_mask(PMPChecker_3_io_check_env_pmp_8_mask),
    .io_check_env_pmp_9_cfg_l(PMPChecker_3_io_check_env_pmp_9_cfg_l),
    .io_check_env_pmp_9_cfg_a(PMPChecker_3_io_check_env_pmp_9_cfg_a),
    .io_check_env_pmp_9_cfg_w(PMPChecker_3_io_check_env_pmp_9_cfg_w),
    .io_check_env_pmp_9_cfg_r(PMPChecker_3_io_check_env_pmp_9_cfg_r),
    .io_check_env_pmp_9_addr(PMPChecker_3_io_check_env_pmp_9_addr),
    .io_check_env_pmp_9_mask(PMPChecker_3_io_check_env_pmp_9_mask),
    .io_check_env_pmp_10_cfg_l(PMPChecker_3_io_check_env_pmp_10_cfg_l),
    .io_check_env_pmp_10_cfg_a(PMPChecker_3_io_check_env_pmp_10_cfg_a),
    .io_check_env_pmp_10_cfg_w(PMPChecker_3_io_check_env_pmp_10_cfg_w),
    .io_check_env_pmp_10_cfg_r(PMPChecker_3_io_check_env_pmp_10_cfg_r),
    .io_check_env_pmp_10_addr(PMPChecker_3_io_check_env_pmp_10_addr),
    .io_check_env_pmp_10_mask(PMPChecker_3_io_check_env_pmp_10_mask),
    .io_check_env_pmp_11_cfg_l(PMPChecker_3_io_check_env_pmp_11_cfg_l),
    .io_check_env_pmp_11_cfg_a(PMPChecker_3_io_check_env_pmp_11_cfg_a),
    .io_check_env_pmp_11_cfg_w(PMPChecker_3_io_check_env_pmp_11_cfg_w),
    .io_check_env_pmp_11_cfg_r(PMPChecker_3_io_check_env_pmp_11_cfg_r),
    .io_check_env_pmp_11_addr(PMPChecker_3_io_check_env_pmp_11_addr),
    .io_check_env_pmp_11_mask(PMPChecker_3_io_check_env_pmp_11_mask),
    .io_check_env_pmp_12_cfg_l(PMPChecker_3_io_check_env_pmp_12_cfg_l),
    .io_check_env_pmp_12_cfg_a(PMPChecker_3_io_check_env_pmp_12_cfg_a),
    .io_check_env_pmp_12_cfg_w(PMPChecker_3_io_check_env_pmp_12_cfg_w),
    .io_check_env_pmp_12_cfg_r(PMPChecker_3_io_check_env_pmp_12_cfg_r),
    .io_check_env_pmp_12_addr(PMPChecker_3_io_check_env_pmp_12_addr),
    .io_check_env_pmp_12_mask(PMPChecker_3_io_check_env_pmp_12_mask),
    .io_check_env_pmp_13_cfg_l(PMPChecker_3_io_check_env_pmp_13_cfg_l),
    .io_check_env_pmp_13_cfg_a(PMPChecker_3_io_check_env_pmp_13_cfg_a),
    .io_check_env_pmp_13_cfg_w(PMPChecker_3_io_check_env_pmp_13_cfg_w),
    .io_check_env_pmp_13_cfg_r(PMPChecker_3_io_check_env_pmp_13_cfg_r),
    .io_check_env_pmp_13_addr(PMPChecker_3_io_check_env_pmp_13_addr),
    .io_check_env_pmp_13_mask(PMPChecker_3_io_check_env_pmp_13_mask),
    .io_check_env_pmp_14_cfg_l(PMPChecker_3_io_check_env_pmp_14_cfg_l),
    .io_check_env_pmp_14_cfg_a(PMPChecker_3_io_check_env_pmp_14_cfg_a),
    .io_check_env_pmp_14_cfg_w(PMPChecker_3_io_check_env_pmp_14_cfg_w),
    .io_check_env_pmp_14_cfg_r(PMPChecker_3_io_check_env_pmp_14_cfg_r),
    .io_check_env_pmp_14_addr(PMPChecker_3_io_check_env_pmp_14_addr),
    .io_check_env_pmp_14_mask(PMPChecker_3_io_check_env_pmp_14_mask),
    .io_check_env_pmp_15_cfg_l(PMPChecker_3_io_check_env_pmp_15_cfg_l),
    .io_check_env_pmp_15_cfg_a(PMPChecker_3_io_check_env_pmp_15_cfg_a),
    .io_check_env_pmp_15_cfg_w(PMPChecker_3_io_check_env_pmp_15_cfg_w),
    .io_check_env_pmp_15_cfg_r(PMPChecker_3_io_check_env_pmp_15_cfg_r),
    .io_check_env_pmp_15_addr(PMPChecker_3_io_check_env_pmp_15_addr),
    .io_check_env_pmp_15_mask(PMPChecker_3_io_check_env_pmp_15_mask),
    .io_check_env_pma_0_cfg_c(PMPChecker_3_io_check_env_pma_0_cfg_c),
    .io_check_env_pma_0_cfg_atomic(PMPChecker_3_io_check_env_pma_0_cfg_atomic),
    .io_check_env_pma_0_cfg_a(PMPChecker_3_io_check_env_pma_0_cfg_a),
    .io_check_env_pma_0_cfg_w(PMPChecker_3_io_check_env_pma_0_cfg_w),
    .io_check_env_pma_0_cfg_r(PMPChecker_3_io_check_env_pma_0_cfg_r),
    .io_check_env_pma_0_addr(PMPChecker_3_io_check_env_pma_0_addr),
    .io_check_env_pma_0_mask(PMPChecker_3_io_check_env_pma_0_mask),
    .io_check_env_pma_1_cfg_c(PMPChecker_3_io_check_env_pma_1_cfg_c),
    .io_check_env_pma_1_cfg_atomic(PMPChecker_3_io_check_env_pma_1_cfg_atomic),
    .io_check_env_pma_1_cfg_a(PMPChecker_3_io_check_env_pma_1_cfg_a),
    .io_check_env_pma_1_cfg_w(PMPChecker_3_io_check_env_pma_1_cfg_w),
    .io_check_env_pma_1_cfg_r(PMPChecker_3_io_check_env_pma_1_cfg_r),
    .io_check_env_pma_1_addr(PMPChecker_3_io_check_env_pma_1_addr),
    .io_check_env_pma_1_mask(PMPChecker_3_io_check_env_pma_1_mask),
    .io_check_env_pma_2_cfg_c(PMPChecker_3_io_check_env_pma_2_cfg_c),
    .io_check_env_pma_2_cfg_atomic(PMPChecker_3_io_check_env_pma_2_cfg_atomic),
    .io_check_env_pma_2_cfg_a(PMPChecker_3_io_check_env_pma_2_cfg_a),
    .io_check_env_pma_2_cfg_w(PMPChecker_3_io_check_env_pma_2_cfg_w),
    .io_check_env_pma_2_cfg_r(PMPChecker_3_io_check_env_pma_2_cfg_r),
    .io_check_env_pma_2_addr(PMPChecker_3_io_check_env_pma_2_addr),
    .io_check_env_pma_2_mask(PMPChecker_3_io_check_env_pma_2_mask),
    .io_check_env_pma_3_cfg_c(PMPChecker_3_io_check_env_pma_3_cfg_c),
    .io_check_env_pma_3_cfg_atomic(PMPChecker_3_io_check_env_pma_3_cfg_atomic),
    .io_check_env_pma_3_cfg_a(PMPChecker_3_io_check_env_pma_3_cfg_a),
    .io_check_env_pma_3_cfg_w(PMPChecker_3_io_check_env_pma_3_cfg_w),
    .io_check_env_pma_3_cfg_r(PMPChecker_3_io_check_env_pma_3_cfg_r),
    .io_check_env_pma_3_addr(PMPChecker_3_io_check_env_pma_3_addr),
    .io_check_env_pma_3_mask(PMPChecker_3_io_check_env_pma_3_mask),
    .io_check_env_pma_4_cfg_c(PMPChecker_3_io_check_env_pma_4_cfg_c),
    .io_check_env_pma_4_cfg_atomic(PMPChecker_3_io_check_env_pma_4_cfg_atomic),
    .io_check_env_pma_4_cfg_a(PMPChecker_3_io_check_env_pma_4_cfg_a),
    .io_check_env_pma_4_cfg_w(PMPChecker_3_io_check_env_pma_4_cfg_w),
    .io_check_env_pma_4_cfg_r(PMPChecker_3_io_check_env_pma_4_cfg_r),
    .io_check_env_pma_4_addr(PMPChecker_3_io_check_env_pma_4_addr),
    .io_check_env_pma_4_mask(PMPChecker_3_io_check_env_pma_4_mask),
    .io_check_env_pma_5_cfg_c(PMPChecker_3_io_check_env_pma_5_cfg_c),
    .io_check_env_pma_5_cfg_atomic(PMPChecker_3_io_check_env_pma_5_cfg_atomic),
    .io_check_env_pma_5_cfg_a(PMPChecker_3_io_check_env_pma_5_cfg_a),
    .io_check_env_pma_5_cfg_w(PMPChecker_3_io_check_env_pma_5_cfg_w),
    .io_check_env_pma_5_cfg_r(PMPChecker_3_io_check_env_pma_5_cfg_r),
    .io_check_env_pma_5_addr(PMPChecker_3_io_check_env_pma_5_addr),
    .io_check_env_pma_5_mask(PMPChecker_3_io_check_env_pma_5_mask),
    .io_check_env_pma_6_cfg_c(PMPChecker_3_io_check_env_pma_6_cfg_c),
    .io_check_env_pma_6_cfg_atomic(PMPChecker_3_io_check_env_pma_6_cfg_atomic),
    .io_check_env_pma_6_cfg_a(PMPChecker_3_io_check_env_pma_6_cfg_a),
    .io_check_env_pma_6_cfg_w(PMPChecker_3_io_check_env_pma_6_cfg_w),
    .io_check_env_pma_6_cfg_r(PMPChecker_3_io_check_env_pma_6_cfg_r),
    .io_check_env_pma_6_addr(PMPChecker_3_io_check_env_pma_6_addr),
    .io_check_env_pma_6_mask(PMPChecker_3_io_check_env_pma_6_mask),
    .io_check_env_pma_7_cfg_c(PMPChecker_3_io_check_env_pma_7_cfg_c),
    .io_check_env_pma_7_cfg_atomic(PMPChecker_3_io_check_env_pma_7_cfg_atomic),
    .io_check_env_pma_7_cfg_a(PMPChecker_3_io_check_env_pma_7_cfg_a),
    .io_check_env_pma_7_cfg_w(PMPChecker_3_io_check_env_pma_7_cfg_w),
    .io_check_env_pma_7_cfg_r(PMPChecker_3_io_check_env_pma_7_cfg_r),
    .io_check_env_pma_7_addr(PMPChecker_3_io_check_env_pma_7_addr),
    .io_check_env_pma_7_mask(PMPChecker_3_io_check_env_pma_7_mask),
    .io_check_env_pma_8_cfg_c(PMPChecker_3_io_check_env_pma_8_cfg_c),
    .io_check_env_pma_8_cfg_atomic(PMPChecker_3_io_check_env_pma_8_cfg_atomic),
    .io_check_env_pma_8_cfg_a(PMPChecker_3_io_check_env_pma_8_cfg_a),
    .io_check_env_pma_8_cfg_w(PMPChecker_3_io_check_env_pma_8_cfg_w),
    .io_check_env_pma_8_cfg_r(PMPChecker_3_io_check_env_pma_8_cfg_r),
    .io_check_env_pma_8_addr(PMPChecker_3_io_check_env_pma_8_addr),
    .io_check_env_pma_8_mask(PMPChecker_3_io_check_env_pma_8_mask),
    .io_check_env_pma_9_cfg_c(PMPChecker_3_io_check_env_pma_9_cfg_c),
    .io_check_env_pma_9_cfg_atomic(PMPChecker_3_io_check_env_pma_9_cfg_atomic),
    .io_check_env_pma_9_cfg_a(PMPChecker_3_io_check_env_pma_9_cfg_a),
    .io_check_env_pma_9_cfg_w(PMPChecker_3_io_check_env_pma_9_cfg_w),
    .io_check_env_pma_9_cfg_r(PMPChecker_3_io_check_env_pma_9_cfg_r),
    .io_check_env_pma_9_addr(PMPChecker_3_io_check_env_pma_9_addr),
    .io_check_env_pma_9_mask(PMPChecker_3_io_check_env_pma_9_mask),
    .io_check_env_pma_10_cfg_c(PMPChecker_3_io_check_env_pma_10_cfg_c),
    .io_check_env_pma_10_cfg_atomic(PMPChecker_3_io_check_env_pma_10_cfg_atomic),
    .io_check_env_pma_10_cfg_a(PMPChecker_3_io_check_env_pma_10_cfg_a),
    .io_check_env_pma_10_cfg_w(PMPChecker_3_io_check_env_pma_10_cfg_w),
    .io_check_env_pma_10_cfg_r(PMPChecker_3_io_check_env_pma_10_cfg_r),
    .io_check_env_pma_10_addr(PMPChecker_3_io_check_env_pma_10_addr),
    .io_check_env_pma_10_mask(PMPChecker_3_io_check_env_pma_10_mask),
    .io_check_env_pma_11_cfg_c(PMPChecker_3_io_check_env_pma_11_cfg_c),
    .io_check_env_pma_11_cfg_atomic(PMPChecker_3_io_check_env_pma_11_cfg_atomic),
    .io_check_env_pma_11_cfg_a(PMPChecker_3_io_check_env_pma_11_cfg_a),
    .io_check_env_pma_11_cfg_w(PMPChecker_3_io_check_env_pma_11_cfg_w),
    .io_check_env_pma_11_cfg_r(PMPChecker_3_io_check_env_pma_11_cfg_r),
    .io_check_env_pma_11_addr(PMPChecker_3_io_check_env_pma_11_addr),
    .io_check_env_pma_11_mask(PMPChecker_3_io_check_env_pma_11_mask),
    .io_check_env_pma_12_cfg_c(PMPChecker_3_io_check_env_pma_12_cfg_c),
    .io_check_env_pma_12_cfg_atomic(PMPChecker_3_io_check_env_pma_12_cfg_atomic),
    .io_check_env_pma_12_cfg_a(PMPChecker_3_io_check_env_pma_12_cfg_a),
    .io_check_env_pma_12_cfg_w(PMPChecker_3_io_check_env_pma_12_cfg_w),
    .io_check_env_pma_12_cfg_r(PMPChecker_3_io_check_env_pma_12_cfg_r),
    .io_check_env_pma_12_addr(PMPChecker_3_io_check_env_pma_12_addr),
    .io_check_env_pma_12_mask(PMPChecker_3_io_check_env_pma_12_mask),
    .io_check_env_pma_13_cfg_c(PMPChecker_3_io_check_env_pma_13_cfg_c),
    .io_check_env_pma_13_cfg_atomic(PMPChecker_3_io_check_env_pma_13_cfg_atomic),
    .io_check_env_pma_13_cfg_a(PMPChecker_3_io_check_env_pma_13_cfg_a),
    .io_check_env_pma_13_cfg_w(PMPChecker_3_io_check_env_pma_13_cfg_w),
    .io_check_env_pma_13_cfg_r(PMPChecker_3_io_check_env_pma_13_cfg_r),
    .io_check_env_pma_13_addr(PMPChecker_3_io_check_env_pma_13_addr),
    .io_check_env_pma_13_mask(PMPChecker_3_io_check_env_pma_13_mask),
    .io_check_env_pma_14_cfg_c(PMPChecker_3_io_check_env_pma_14_cfg_c),
    .io_check_env_pma_14_cfg_atomic(PMPChecker_3_io_check_env_pma_14_cfg_atomic),
    .io_check_env_pma_14_cfg_a(PMPChecker_3_io_check_env_pma_14_cfg_a),
    .io_check_env_pma_14_cfg_w(PMPChecker_3_io_check_env_pma_14_cfg_w),
    .io_check_env_pma_14_cfg_r(PMPChecker_3_io_check_env_pma_14_cfg_r),
    .io_check_env_pma_14_addr(PMPChecker_3_io_check_env_pma_14_addr),
    .io_check_env_pma_14_mask(PMPChecker_3_io_check_env_pma_14_mask),
    .io_check_env_pma_15_cfg_c(PMPChecker_3_io_check_env_pma_15_cfg_c),
    .io_check_env_pma_15_cfg_atomic(PMPChecker_3_io_check_env_pma_15_cfg_atomic),
    .io_check_env_pma_15_cfg_a(PMPChecker_3_io_check_env_pma_15_cfg_a),
    .io_check_env_pma_15_cfg_w(PMPChecker_3_io_check_env_pma_15_cfg_w),
    .io_check_env_pma_15_cfg_r(PMPChecker_3_io_check_env_pma_15_cfg_r),
    .io_check_env_pma_15_addr(PMPChecker_3_io_check_env_pma_15_addr),
    .io_check_env_pma_15_mask(PMPChecker_3_io_check_env_pma_15_mask),
    .io_req_valid(PMPChecker_3_io_req_valid),
    .io_req_bits_addr(PMPChecker_3_io_req_bits_addr),
    .io_req_bits_cmd(PMPChecker_3_io_req_bits_cmd),
    .io_resp_ld(PMPChecker_3_io_resp_ld),
    .io_resp_st(PMPChecker_3_io_resp_st),
    .io_resp_mmio(PMPChecker_3_io_resp_mmio),
    .io_resp_atomic(PMPChecker_3_io_resp_atomic)
  );
  PMPChecker_8 PMPChecker_4 ( // @[MemBlock.scala 314:91]
    .clock(PMPChecker_4_clock),
    .io_check_env_mode(PMPChecker_4_io_check_env_mode),
    .io_check_env_pmp_0_cfg_l(PMPChecker_4_io_check_env_pmp_0_cfg_l),
    .io_check_env_pmp_0_cfg_a(PMPChecker_4_io_check_env_pmp_0_cfg_a),
    .io_check_env_pmp_0_cfg_w(PMPChecker_4_io_check_env_pmp_0_cfg_w),
    .io_check_env_pmp_0_cfg_r(PMPChecker_4_io_check_env_pmp_0_cfg_r),
    .io_check_env_pmp_0_addr(PMPChecker_4_io_check_env_pmp_0_addr),
    .io_check_env_pmp_0_mask(PMPChecker_4_io_check_env_pmp_0_mask),
    .io_check_env_pmp_1_cfg_l(PMPChecker_4_io_check_env_pmp_1_cfg_l),
    .io_check_env_pmp_1_cfg_a(PMPChecker_4_io_check_env_pmp_1_cfg_a),
    .io_check_env_pmp_1_cfg_w(PMPChecker_4_io_check_env_pmp_1_cfg_w),
    .io_check_env_pmp_1_cfg_r(PMPChecker_4_io_check_env_pmp_1_cfg_r),
    .io_check_env_pmp_1_addr(PMPChecker_4_io_check_env_pmp_1_addr),
    .io_check_env_pmp_1_mask(PMPChecker_4_io_check_env_pmp_1_mask),
    .io_check_env_pmp_2_cfg_l(PMPChecker_4_io_check_env_pmp_2_cfg_l),
    .io_check_env_pmp_2_cfg_a(PMPChecker_4_io_check_env_pmp_2_cfg_a),
    .io_check_env_pmp_2_cfg_w(PMPChecker_4_io_check_env_pmp_2_cfg_w),
    .io_check_env_pmp_2_cfg_r(PMPChecker_4_io_check_env_pmp_2_cfg_r),
    .io_check_env_pmp_2_addr(PMPChecker_4_io_check_env_pmp_2_addr),
    .io_check_env_pmp_2_mask(PMPChecker_4_io_check_env_pmp_2_mask),
    .io_check_env_pmp_3_cfg_l(PMPChecker_4_io_check_env_pmp_3_cfg_l),
    .io_check_env_pmp_3_cfg_a(PMPChecker_4_io_check_env_pmp_3_cfg_a),
    .io_check_env_pmp_3_cfg_w(PMPChecker_4_io_check_env_pmp_3_cfg_w),
    .io_check_env_pmp_3_cfg_r(PMPChecker_4_io_check_env_pmp_3_cfg_r),
    .io_check_env_pmp_3_addr(PMPChecker_4_io_check_env_pmp_3_addr),
    .io_check_env_pmp_3_mask(PMPChecker_4_io_check_env_pmp_3_mask),
    .io_check_env_pmp_4_cfg_l(PMPChecker_4_io_check_env_pmp_4_cfg_l),
    .io_check_env_pmp_4_cfg_a(PMPChecker_4_io_check_env_pmp_4_cfg_a),
    .io_check_env_pmp_4_cfg_w(PMPChecker_4_io_check_env_pmp_4_cfg_w),
    .io_check_env_pmp_4_cfg_r(PMPChecker_4_io_check_env_pmp_4_cfg_r),
    .io_check_env_pmp_4_addr(PMPChecker_4_io_check_env_pmp_4_addr),
    .io_check_env_pmp_4_mask(PMPChecker_4_io_check_env_pmp_4_mask),
    .io_check_env_pmp_5_cfg_l(PMPChecker_4_io_check_env_pmp_5_cfg_l),
    .io_check_env_pmp_5_cfg_a(PMPChecker_4_io_check_env_pmp_5_cfg_a),
    .io_check_env_pmp_5_cfg_w(PMPChecker_4_io_check_env_pmp_5_cfg_w),
    .io_check_env_pmp_5_cfg_r(PMPChecker_4_io_check_env_pmp_5_cfg_r),
    .io_check_env_pmp_5_addr(PMPChecker_4_io_check_env_pmp_5_addr),
    .io_check_env_pmp_5_mask(PMPChecker_4_io_check_env_pmp_5_mask),
    .io_check_env_pmp_6_cfg_l(PMPChecker_4_io_check_env_pmp_6_cfg_l),
    .io_check_env_pmp_6_cfg_a(PMPChecker_4_io_check_env_pmp_6_cfg_a),
    .io_check_env_pmp_6_cfg_w(PMPChecker_4_io_check_env_pmp_6_cfg_w),
    .io_check_env_pmp_6_cfg_r(PMPChecker_4_io_check_env_pmp_6_cfg_r),
    .io_check_env_pmp_6_addr(PMPChecker_4_io_check_env_pmp_6_addr),
    .io_check_env_pmp_6_mask(PMPChecker_4_io_check_env_pmp_6_mask),
    .io_check_env_pmp_7_cfg_l(PMPChecker_4_io_check_env_pmp_7_cfg_l),
    .io_check_env_pmp_7_cfg_a(PMPChecker_4_io_check_env_pmp_7_cfg_a),
    .io_check_env_pmp_7_cfg_w(PMPChecker_4_io_check_env_pmp_7_cfg_w),
    .io_check_env_pmp_7_cfg_r(PMPChecker_4_io_check_env_pmp_7_cfg_r),
    .io_check_env_pmp_7_addr(PMPChecker_4_io_check_env_pmp_7_addr),
    .io_check_env_pmp_7_mask(PMPChecker_4_io_check_env_pmp_7_mask),
    .io_check_env_pmp_8_cfg_l(PMPChecker_4_io_check_env_pmp_8_cfg_l),
    .io_check_env_pmp_8_cfg_a(PMPChecker_4_io_check_env_pmp_8_cfg_a),
    .io_check_env_pmp_8_cfg_w(PMPChecker_4_io_check_env_pmp_8_cfg_w),
    .io_check_env_pmp_8_cfg_r(PMPChecker_4_io_check_env_pmp_8_cfg_r),
    .io_check_env_pmp_8_addr(PMPChecker_4_io_check_env_pmp_8_addr),
    .io_check_env_pmp_8_mask(PMPChecker_4_io_check_env_pmp_8_mask),
    .io_check_env_pmp_9_cfg_l(PMPChecker_4_io_check_env_pmp_9_cfg_l),
    .io_check_env_pmp_9_cfg_a(PMPChecker_4_io_check_env_pmp_9_cfg_a),
    .io_check_env_pmp_9_cfg_w(PMPChecker_4_io_check_env_pmp_9_cfg_w),
    .io_check_env_pmp_9_cfg_r(PMPChecker_4_io_check_env_pmp_9_cfg_r),
    .io_check_env_pmp_9_addr(PMPChecker_4_io_check_env_pmp_9_addr),
    .io_check_env_pmp_9_mask(PMPChecker_4_io_check_env_pmp_9_mask),
    .io_check_env_pmp_10_cfg_l(PMPChecker_4_io_check_env_pmp_10_cfg_l),
    .io_check_env_pmp_10_cfg_a(PMPChecker_4_io_check_env_pmp_10_cfg_a),
    .io_check_env_pmp_10_cfg_w(PMPChecker_4_io_check_env_pmp_10_cfg_w),
    .io_check_env_pmp_10_cfg_r(PMPChecker_4_io_check_env_pmp_10_cfg_r),
    .io_check_env_pmp_10_addr(PMPChecker_4_io_check_env_pmp_10_addr),
    .io_check_env_pmp_10_mask(PMPChecker_4_io_check_env_pmp_10_mask),
    .io_check_env_pmp_11_cfg_l(PMPChecker_4_io_check_env_pmp_11_cfg_l),
    .io_check_env_pmp_11_cfg_a(PMPChecker_4_io_check_env_pmp_11_cfg_a),
    .io_check_env_pmp_11_cfg_w(PMPChecker_4_io_check_env_pmp_11_cfg_w),
    .io_check_env_pmp_11_cfg_r(PMPChecker_4_io_check_env_pmp_11_cfg_r),
    .io_check_env_pmp_11_addr(PMPChecker_4_io_check_env_pmp_11_addr),
    .io_check_env_pmp_11_mask(PMPChecker_4_io_check_env_pmp_11_mask),
    .io_check_env_pmp_12_cfg_l(PMPChecker_4_io_check_env_pmp_12_cfg_l),
    .io_check_env_pmp_12_cfg_a(PMPChecker_4_io_check_env_pmp_12_cfg_a),
    .io_check_env_pmp_12_cfg_w(PMPChecker_4_io_check_env_pmp_12_cfg_w),
    .io_check_env_pmp_12_cfg_r(PMPChecker_4_io_check_env_pmp_12_cfg_r),
    .io_check_env_pmp_12_addr(PMPChecker_4_io_check_env_pmp_12_addr),
    .io_check_env_pmp_12_mask(PMPChecker_4_io_check_env_pmp_12_mask),
    .io_check_env_pmp_13_cfg_l(PMPChecker_4_io_check_env_pmp_13_cfg_l),
    .io_check_env_pmp_13_cfg_a(PMPChecker_4_io_check_env_pmp_13_cfg_a),
    .io_check_env_pmp_13_cfg_w(PMPChecker_4_io_check_env_pmp_13_cfg_w),
    .io_check_env_pmp_13_cfg_r(PMPChecker_4_io_check_env_pmp_13_cfg_r),
    .io_check_env_pmp_13_addr(PMPChecker_4_io_check_env_pmp_13_addr),
    .io_check_env_pmp_13_mask(PMPChecker_4_io_check_env_pmp_13_mask),
    .io_check_env_pmp_14_cfg_l(PMPChecker_4_io_check_env_pmp_14_cfg_l),
    .io_check_env_pmp_14_cfg_a(PMPChecker_4_io_check_env_pmp_14_cfg_a),
    .io_check_env_pmp_14_cfg_w(PMPChecker_4_io_check_env_pmp_14_cfg_w),
    .io_check_env_pmp_14_cfg_r(PMPChecker_4_io_check_env_pmp_14_cfg_r),
    .io_check_env_pmp_14_addr(PMPChecker_4_io_check_env_pmp_14_addr),
    .io_check_env_pmp_14_mask(PMPChecker_4_io_check_env_pmp_14_mask),
    .io_check_env_pmp_15_cfg_l(PMPChecker_4_io_check_env_pmp_15_cfg_l),
    .io_check_env_pmp_15_cfg_a(PMPChecker_4_io_check_env_pmp_15_cfg_a),
    .io_check_env_pmp_15_cfg_w(PMPChecker_4_io_check_env_pmp_15_cfg_w),
    .io_check_env_pmp_15_cfg_r(PMPChecker_4_io_check_env_pmp_15_cfg_r),
    .io_check_env_pmp_15_addr(PMPChecker_4_io_check_env_pmp_15_addr),
    .io_check_env_pmp_15_mask(PMPChecker_4_io_check_env_pmp_15_mask),
    .io_check_env_pma_0_cfg_c(PMPChecker_4_io_check_env_pma_0_cfg_c),
    .io_check_env_pma_0_cfg_atomic(PMPChecker_4_io_check_env_pma_0_cfg_atomic),
    .io_check_env_pma_0_cfg_a(PMPChecker_4_io_check_env_pma_0_cfg_a),
    .io_check_env_pma_0_cfg_w(PMPChecker_4_io_check_env_pma_0_cfg_w),
    .io_check_env_pma_0_cfg_r(PMPChecker_4_io_check_env_pma_0_cfg_r),
    .io_check_env_pma_0_addr(PMPChecker_4_io_check_env_pma_0_addr),
    .io_check_env_pma_0_mask(PMPChecker_4_io_check_env_pma_0_mask),
    .io_check_env_pma_1_cfg_c(PMPChecker_4_io_check_env_pma_1_cfg_c),
    .io_check_env_pma_1_cfg_atomic(PMPChecker_4_io_check_env_pma_1_cfg_atomic),
    .io_check_env_pma_1_cfg_a(PMPChecker_4_io_check_env_pma_1_cfg_a),
    .io_check_env_pma_1_cfg_w(PMPChecker_4_io_check_env_pma_1_cfg_w),
    .io_check_env_pma_1_cfg_r(PMPChecker_4_io_check_env_pma_1_cfg_r),
    .io_check_env_pma_1_addr(PMPChecker_4_io_check_env_pma_1_addr),
    .io_check_env_pma_1_mask(PMPChecker_4_io_check_env_pma_1_mask),
    .io_check_env_pma_2_cfg_c(PMPChecker_4_io_check_env_pma_2_cfg_c),
    .io_check_env_pma_2_cfg_atomic(PMPChecker_4_io_check_env_pma_2_cfg_atomic),
    .io_check_env_pma_2_cfg_a(PMPChecker_4_io_check_env_pma_2_cfg_a),
    .io_check_env_pma_2_cfg_w(PMPChecker_4_io_check_env_pma_2_cfg_w),
    .io_check_env_pma_2_cfg_r(PMPChecker_4_io_check_env_pma_2_cfg_r),
    .io_check_env_pma_2_addr(PMPChecker_4_io_check_env_pma_2_addr),
    .io_check_env_pma_2_mask(PMPChecker_4_io_check_env_pma_2_mask),
    .io_check_env_pma_3_cfg_c(PMPChecker_4_io_check_env_pma_3_cfg_c),
    .io_check_env_pma_3_cfg_atomic(PMPChecker_4_io_check_env_pma_3_cfg_atomic),
    .io_check_env_pma_3_cfg_a(PMPChecker_4_io_check_env_pma_3_cfg_a),
    .io_check_env_pma_3_cfg_w(PMPChecker_4_io_check_env_pma_3_cfg_w),
    .io_check_env_pma_3_cfg_r(PMPChecker_4_io_check_env_pma_3_cfg_r),
    .io_check_env_pma_3_addr(PMPChecker_4_io_check_env_pma_3_addr),
    .io_check_env_pma_3_mask(PMPChecker_4_io_check_env_pma_3_mask),
    .io_check_env_pma_4_cfg_c(PMPChecker_4_io_check_env_pma_4_cfg_c),
    .io_check_env_pma_4_cfg_atomic(PMPChecker_4_io_check_env_pma_4_cfg_atomic),
    .io_check_env_pma_4_cfg_a(PMPChecker_4_io_check_env_pma_4_cfg_a),
    .io_check_env_pma_4_cfg_w(PMPChecker_4_io_check_env_pma_4_cfg_w),
    .io_check_env_pma_4_cfg_r(PMPChecker_4_io_check_env_pma_4_cfg_r),
    .io_check_env_pma_4_addr(PMPChecker_4_io_check_env_pma_4_addr),
    .io_check_env_pma_4_mask(PMPChecker_4_io_check_env_pma_4_mask),
    .io_check_env_pma_5_cfg_c(PMPChecker_4_io_check_env_pma_5_cfg_c),
    .io_check_env_pma_5_cfg_atomic(PMPChecker_4_io_check_env_pma_5_cfg_atomic),
    .io_check_env_pma_5_cfg_a(PMPChecker_4_io_check_env_pma_5_cfg_a),
    .io_check_env_pma_5_cfg_w(PMPChecker_4_io_check_env_pma_5_cfg_w),
    .io_check_env_pma_5_cfg_r(PMPChecker_4_io_check_env_pma_5_cfg_r),
    .io_check_env_pma_5_addr(PMPChecker_4_io_check_env_pma_5_addr),
    .io_check_env_pma_5_mask(PMPChecker_4_io_check_env_pma_5_mask),
    .io_check_env_pma_6_cfg_c(PMPChecker_4_io_check_env_pma_6_cfg_c),
    .io_check_env_pma_6_cfg_atomic(PMPChecker_4_io_check_env_pma_6_cfg_atomic),
    .io_check_env_pma_6_cfg_a(PMPChecker_4_io_check_env_pma_6_cfg_a),
    .io_check_env_pma_6_cfg_w(PMPChecker_4_io_check_env_pma_6_cfg_w),
    .io_check_env_pma_6_cfg_r(PMPChecker_4_io_check_env_pma_6_cfg_r),
    .io_check_env_pma_6_addr(PMPChecker_4_io_check_env_pma_6_addr),
    .io_check_env_pma_6_mask(PMPChecker_4_io_check_env_pma_6_mask),
    .io_check_env_pma_7_cfg_c(PMPChecker_4_io_check_env_pma_7_cfg_c),
    .io_check_env_pma_7_cfg_atomic(PMPChecker_4_io_check_env_pma_7_cfg_atomic),
    .io_check_env_pma_7_cfg_a(PMPChecker_4_io_check_env_pma_7_cfg_a),
    .io_check_env_pma_7_cfg_w(PMPChecker_4_io_check_env_pma_7_cfg_w),
    .io_check_env_pma_7_cfg_r(PMPChecker_4_io_check_env_pma_7_cfg_r),
    .io_check_env_pma_7_addr(PMPChecker_4_io_check_env_pma_7_addr),
    .io_check_env_pma_7_mask(PMPChecker_4_io_check_env_pma_7_mask),
    .io_check_env_pma_8_cfg_c(PMPChecker_4_io_check_env_pma_8_cfg_c),
    .io_check_env_pma_8_cfg_atomic(PMPChecker_4_io_check_env_pma_8_cfg_atomic),
    .io_check_env_pma_8_cfg_a(PMPChecker_4_io_check_env_pma_8_cfg_a),
    .io_check_env_pma_8_cfg_w(PMPChecker_4_io_check_env_pma_8_cfg_w),
    .io_check_env_pma_8_cfg_r(PMPChecker_4_io_check_env_pma_8_cfg_r),
    .io_check_env_pma_8_addr(PMPChecker_4_io_check_env_pma_8_addr),
    .io_check_env_pma_8_mask(PMPChecker_4_io_check_env_pma_8_mask),
    .io_check_env_pma_9_cfg_c(PMPChecker_4_io_check_env_pma_9_cfg_c),
    .io_check_env_pma_9_cfg_atomic(PMPChecker_4_io_check_env_pma_9_cfg_atomic),
    .io_check_env_pma_9_cfg_a(PMPChecker_4_io_check_env_pma_9_cfg_a),
    .io_check_env_pma_9_cfg_w(PMPChecker_4_io_check_env_pma_9_cfg_w),
    .io_check_env_pma_9_cfg_r(PMPChecker_4_io_check_env_pma_9_cfg_r),
    .io_check_env_pma_9_addr(PMPChecker_4_io_check_env_pma_9_addr),
    .io_check_env_pma_9_mask(PMPChecker_4_io_check_env_pma_9_mask),
    .io_check_env_pma_10_cfg_c(PMPChecker_4_io_check_env_pma_10_cfg_c),
    .io_check_env_pma_10_cfg_atomic(PMPChecker_4_io_check_env_pma_10_cfg_atomic),
    .io_check_env_pma_10_cfg_a(PMPChecker_4_io_check_env_pma_10_cfg_a),
    .io_check_env_pma_10_cfg_w(PMPChecker_4_io_check_env_pma_10_cfg_w),
    .io_check_env_pma_10_cfg_r(PMPChecker_4_io_check_env_pma_10_cfg_r),
    .io_check_env_pma_10_addr(PMPChecker_4_io_check_env_pma_10_addr),
    .io_check_env_pma_10_mask(PMPChecker_4_io_check_env_pma_10_mask),
    .io_check_env_pma_11_cfg_c(PMPChecker_4_io_check_env_pma_11_cfg_c),
    .io_check_env_pma_11_cfg_atomic(PMPChecker_4_io_check_env_pma_11_cfg_atomic),
    .io_check_env_pma_11_cfg_a(PMPChecker_4_io_check_env_pma_11_cfg_a),
    .io_check_env_pma_11_cfg_w(PMPChecker_4_io_check_env_pma_11_cfg_w),
    .io_check_env_pma_11_cfg_r(PMPChecker_4_io_check_env_pma_11_cfg_r),
    .io_check_env_pma_11_addr(PMPChecker_4_io_check_env_pma_11_addr),
    .io_check_env_pma_11_mask(PMPChecker_4_io_check_env_pma_11_mask),
    .io_check_env_pma_12_cfg_c(PMPChecker_4_io_check_env_pma_12_cfg_c),
    .io_check_env_pma_12_cfg_atomic(PMPChecker_4_io_check_env_pma_12_cfg_atomic),
    .io_check_env_pma_12_cfg_a(PMPChecker_4_io_check_env_pma_12_cfg_a),
    .io_check_env_pma_12_cfg_w(PMPChecker_4_io_check_env_pma_12_cfg_w),
    .io_check_env_pma_12_cfg_r(PMPChecker_4_io_check_env_pma_12_cfg_r),
    .io_check_env_pma_12_addr(PMPChecker_4_io_check_env_pma_12_addr),
    .io_check_env_pma_12_mask(PMPChecker_4_io_check_env_pma_12_mask),
    .io_check_env_pma_13_cfg_c(PMPChecker_4_io_check_env_pma_13_cfg_c),
    .io_check_env_pma_13_cfg_atomic(PMPChecker_4_io_check_env_pma_13_cfg_atomic),
    .io_check_env_pma_13_cfg_a(PMPChecker_4_io_check_env_pma_13_cfg_a),
    .io_check_env_pma_13_cfg_w(PMPChecker_4_io_check_env_pma_13_cfg_w),
    .io_check_env_pma_13_cfg_r(PMPChecker_4_io_check_env_pma_13_cfg_r),
    .io_check_env_pma_13_addr(PMPChecker_4_io_check_env_pma_13_addr),
    .io_check_env_pma_13_mask(PMPChecker_4_io_check_env_pma_13_mask),
    .io_check_env_pma_14_cfg_c(PMPChecker_4_io_check_env_pma_14_cfg_c),
    .io_check_env_pma_14_cfg_atomic(PMPChecker_4_io_check_env_pma_14_cfg_atomic),
    .io_check_env_pma_14_cfg_a(PMPChecker_4_io_check_env_pma_14_cfg_a),
    .io_check_env_pma_14_cfg_w(PMPChecker_4_io_check_env_pma_14_cfg_w),
    .io_check_env_pma_14_cfg_r(PMPChecker_4_io_check_env_pma_14_cfg_r),
    .io_check_env_pma_14_addr(PMPChecker_4_io_check_env_pma_14_addr),
    .io_check_env_pma_14_mask(PMPChecker_4_io_check_env_pma_14_mask),
    .io_check_env_pma_15_cfg_c(PMPChecker_4_io_check_env_pma_15_cfg_c),
    .io_check_env_pma_15_cfg_atomic(PMPChecker_4_io_check_env_pma_15_cfg_atomic),
    .io_check_env_pma_15_cfg_a(PMPChecker_4_io_check_env_pma_15_cfg_a),
    .io_check_env_pma_15_cfg_w(PMPChecker_4_io_check_env_pma_15_cfg_w),
    .io_check_env_pma_15_cfg_r(PMPChecker_4_io_check_env_pma_15_cfg_r),
    .io_check_env_pma_15_addr(PMPChecker_4_io_check_env_pma_15_addr),
    .io_check_env_pma_15_mask(PMPChecker_4_io_check_env_pma_15_mask),
    .io_req_valid(PMPChecker_4_io_req_valid),
    .io_req_bits_addr(PMPChecker_4_io_req_bits_addr),
    .io_req_bits_cmd(PMPChecker_4_io_req_bits_cmd),
    .io_resp_ld(PMPChecker_4_io_resp_ld),
    .io_resp_st(PMPChecker_4_io_resp_st),
    .io_resp_mmio(PMPChecker_4_io_resp_mmio),
    .io_resp_atomic(PMPChecker_4_io_resp_atomic)
  );
  PMPCheckerv2 pmp_check_ptw ( // @[MemBlock.scala 319:29]
    .clock(pmp_check_ptw_clock),
    .reset(pmp_check_ptw_reset),
    .io_check_env_mode(pmp_check_ptw_io_check_env_mode),
    .io_check_env_pmp_0_cfg_l(pmp_check_ptw_io_check_env_pmp_0_cfg_l),
    .io_check_env_pmp_0_cfg_a(pmp_check_ptw_io_check_env_pmp_0_cfg_a),
    .io_check_env_pmp_0_cfg_x(pmp_check_ptw_io_check_env_pmp_0_cfg_x),
    .io_check_env_pmp_0_cfg_w(pmp_check_ptw_io_check_env_pmp_0_cfg_w),
    .io_check_env_pmp_0_cfg_r(pmp_check_ptw_io_check_env_pmp_0_cfg_r),
    .io_check_env_pmp_0_addr(pmp_check_ptw_io_check_env_pmp_0_addr),
    .io_check_env_pmp_0_mask(pmp_check_ptw_io_check_env_pmp_0_mask),
    .io_check_env_pmp_1_cfg_l(pmp_check_ptw_io_check_env_pmp_1_cfg_l),
    .io_check_env_pmp_1_cfg_a(pmp_check_ptw_io_check_env_pmp_1_cfg_a),
    .io_check_env_pmp_1_cfg_x(pmp_check_ptw_io_check_env_pmp_1_cfg_x),
    .io_check_env_pmp_1_cfg_w(pmp_check_ptw_io_check_env_pmp_1_cfg_w),
    .io_check_env_pmp_1_cfg_r(pmp_check_ptw_io_check_env_pmp_1_cfg_r),
    .io_check_env_pmp_1_addr(pmp_check_ptw_io_check_env_pmp_1_addr),
    .io_check_env_pmp_1_mask(pmp_check_ptw_io_check_env_pmp_1_mask),
    .io_check_env_pmp_2_cfg_l(pmp_check_ptw_io_check_env_pmp_2_cfg_l),
    .io_check_env_pmp_2_cfg_a(pmp_check_ptw_io_check_env_pmp_2_cfg_a),
    .io_check_env_pmp_2_cfg_x(pmp_check_ptw_io_check_env_pmp_2_cfg_x),
    .io_check_env_pmp_2_cfg_w(pmp_check_ptw_io_check_env_pmp_2_cfg_w),
    .io_check_env_pmp_2_cfg_r(pmp_check_ptw_io_check_env_pmp_2_cfg_r),
    .io_check_env_pmp_2_addr(pmp_check_ptw_io_check_env_pmp_2_addr),
    .io_check_env_pmp_2_mask(pmp_check_ptw_io_check_env_pmp_2_mask),
    .io_check_env_pmp_3_cfg_l(pmp_check_ptw_io_check_env_pmp_3_cfg_l),
    .io_check_env_pmp_3_cfg_a(pmp_check_ptw_io_check_env_pmp_3_cfg_a),
    .io_check_env_pmp_3_cfg_x(pmp_check_ptw_io_check_env_pmp_3_cfg_x),
    .io_check_env_pmp_3_cfg_w(pmp_check_ptw_io_check_env_pmp_3_cfg_w),
    .io_check_env_pmp_3_cfg_r(pmp_check_ptw_io_check_env_pmp_3_cfg_r),
    .io_check_env_pmp_3_addr(pmp_check_ptw_io_check_env_pmp_3_addr),
    .io_check_env_pmp_3_mask(pmp_check_ptw_io_check_env_pmp_3_mask),
    .io_check_env_pmp_4_cfg_l(pmp_check_ptw_io_check_env_pmp_4_cfg_l),
    .io_check_env_pmp_4_cfg_a(pmp_check_ptw_io_check_env_pmp_4_cfg_a),
    .io_check_env_pmp_4_cfg_x(pmp_check_ptw_io_check_env_pmp_4_cfg_x),
    .io_check_env_pmp_4_cfg_w(pmp_check_ptw_io_check_env_pmp_4_cfg_w),
    .io_check_env_pmp_4_cfg_r(pmp_check_ptw_io_check_env_pmp_4_cfg_r),
    .io_check_env_pmp_4_addr(pmp_check_ptw_io_check_env_pmp_4_addr),
    .io_check_env_pmp_4_mask(pmp_check_ptw_io_check_env_pmp_4_mask),
    .io_check_env_pmp_5_cfg_l(pmp_check_ptw_io_check_env_pmp_5_cfg_l),
    .io_check_env_pmp_5_cfg_a(pmp_check_ptw_io_check_env_pmp_5_cfg_a),
    .io_check_env_pmp_5_cfg_x(pmp_check_ptw_io_check_env_pmp_5_cfg_x),
    .io_check_env_pmp_5_cfg_w(pmp_check_ptw_io_check_env_pmp_5_cfg_w),
    .io_check_env_pmp_5_cfg_r(pmp_check_ptw_io_check_env_pmp_5_cfg_r),
    .io_check_env_pmp_5_addr(pmp_check_ptw_io_check_env_pmp_5_addr),
    .io_check_env_pmp_5_mask(pmp_check_ptw_io_check_env_pmp_5_mask),
    .io_check_env_pmp_6_cfg_l(pmp_check_ptw_io_check_env_pmp_6_cfg_l),
    .io_check_env_pmp_6_cfg_a(pmp_check_ptw_io_check_env_pmp_6_cfg_a),
    .io_check_env_pmp_6_cfg_x(pmp_check_ptw_io_check_env_pmp_6_cfg_x),
    .io_check_env_pmp_6_cfg_w(pmp_check_ptw_io_check_env_pmp_6_cfg_w),
    .io_check_env_pmp_6_cfg_r(pmp_check_ptw_io_check_env_pmp_6_cfg_r),
    .io_check_env_pmp_6_addr(pmp_check_ptw_io_check_env_pmp_6_addr),
    .io_check_env_pmp_6_mask(pmp_check_ptw_io_check_env_pmp_6_mask),
    .io_check_env_pmp_7_cfg_l(pmp_check_ptw_io_check_env_pmp_7_cfg_l),
    .io_check_env_pmp_7_cfg_a(pmp_check_ptw_io_check_env_pmp_7_cfg_a),
    .io_check_env_pmp_7_cfg_x(pmp_check_ptw_io_check_env_pmp_7_cfg_x),
    .io_check_env_pmp_7_cfg_w(pmp_check_ptw_io_check_env_pmp_7_cfg_w),
    .io_check_env_pmp_7_cfg_r(pmp_check_ptw_io_check_env_pmp_7_cfg_r),
    .io_check_env_pmp_7_addr(pmp_check_ptw_io_check_env_pmp_7_addr),
    .io_check_env_pmp_7_mask(pmp_check_ptw_io_check_env_pmp_7_mask),
    .io_check_env_pmp_8_cfg_l(pmp_check_ptw_io_check_env_pmp_8_cfg_l),
    .io_check_env_pmp_8_cfg_a(pmp_check_ptw_io_check_env_pmp_8_cfg_a),
    .io_check_env_pmp_8_cfg_x(pmp_check_ptw_io_check_env_pmp_8_cfg_x),
    .io_check_env_pmp_8_cfg_w(pmp_check_ptw_io_check_env_pmp_8_cfg_w),
    .io_check_env_pmp_8_cfg_r(pmp_check_ptw_io_check_env_pmp_8_cfg_r),
    .io_check_env_pmp_8_addr(pmp_check_ptw_io_check_env_pmp_8_addr),
    .io_check_env_pmp_8_mask(pmp_check_ptw_io_check_env_pmp_8_mask),
    .io_check_env_pmp_9_cfg_l(pmp_check_ptw_io_check_env_pmp_9_cfg_l),
    .io_check_env_pmp_9_cfg_a(pmp_check_ptw_io_check_env_pmp_9_cfg_a),
    .io_check_env_pmp_9_cfg_x(pmp_check_ptw_io_check_env_pmp_9_cfg_x),
    .io_check_env_pmp_9_cfg_w(pmp_check_ptw_io_check_env_pmp_9_cfg_w),
    .io_check_env_pmp_9_cfg_r(pmp_check_ptw_io_check_env_pmp_9_cfg_r),
    .io_check_env_pmp_9_addr(pmp_check_ptw_io_check_env_pmp_9_addr),
    .io_check_env_pmp_9_mask(pmp_check_ptw_io_check_env_pmp_9_mask),
    .io_check_env_pmp_10_cfg_l(pmp_check_ptw_io_check_env_pmp_10_cfg_l),
    .io_check_env_pmp_10_cfg_a(pmp_check_ptw_io_check_env_pmp_10_cfg_a),
    .io_check_env_pmp_10_cfg_x(pmp_check_ptw_io_check_env_pmp_10_cfg_x),
    .io_check_env_pmp_10_cfg_w(pmp_check_ptw_io_check_env_pmp_10_cfg_w),
    .io_check_env_pmp_10_cfg_r(pmp_check_ptw_io_check_env_pmp_10_cfg_r),
    .io_check_env_pmp_10_addr(pmp_check_ptw_io_check_env_pmp_10_addr),
    .io_check_env_pmp_10_mask(pmp_check_ptw_io_check_env_pmp_10_mask),
    .io_check_env_pmp_11_cfg_l(pmp_check_ptw_io_check_env_pmp_11_cfg_l),
    .io_check_env_pmp_11_cfg_a(pmp_check_ptw_io_check_env_pmp_11_cfg_a),
    .io_check_env_pmp_11_cfg_x(pmp_check_ptw_io_check_env_pmp_11_cfg_x),
    .io_check_env_pmp_11_cfg_w(pmp_check_ptw_io_check_env_pmp_11_cfg_w),
    .io_check_env_pmp_11_cfg_r(pmp_check_ptw_io_check_env_pmp_11_cfg_r),
    .io_check_env_pmp_11_addr(pmp_check_ptw_io_check_env_pmp_11_addr),
    .io_check_env_pmp_11_mask(pmp_check_ptw_io_check_env_pmp_11_mask),
    .io_check_env_pmp_12_cfg_l(pmp_check_ptw_io_check_env_pmp_12_cfg_l),
    .io_check_env_pmp_12_cfg_a(pmp_check_ptw_io_check_env_pmp_12_cfg_a),
    .io_check_env_pmp_12_cfg_x(pmp_check_ptw_io_check_env_pmp_12_cfg_x),
    .io_check_env_pmp_12_cfg_w(pmp_check_ptw_io_check_env_pmp_12_cfg_w),
    .io_check_env_pmp_12_cfg_r(pmp_check_ptw_io_check_env_pmp_12_cfg_r),
    .io_check_env_pmp_12_addr(pmp_check_ptw_io_check_env_pmp_12_addr),
    .io_check_env_pmp_12_mask(pmp_check_ptw_io_check_env_pmp_12_mask),
    .io_check_env_pmp_13_cfg_l(pmp_check_ptw_io_check_env_pmp_13_cfg_l),
    .io_check_env_pmp_13_cfg_a(pmp_check_ptw_io_check_env_pmp_13_cfg_a),
    .io_check_env_pmp_13_cfg_x(pmp_check_ptw_io_check_env_pmp_13_cfg_x),
    .io_check_env_pmp_13_cfg_w(pmp_check_ptw_io_check_env_pmp_13_cfg_w),
    .io_check_env_pmp_13_cfg_r(pmp_check_ptw_io_check_env_pmp_13_cfg_r),
    .io_check_env_pmp_13_addr(pmp_check_ptw_io_check_env_pmp_13_addr),
    .io_check_env_pmp_13_mask(pmp_check_ptw_io_check_env_pmp_13_mask),
    .io_check_env_pmp_14_cfg_l(pmp_check_ptw_io_check_env_pmp_14_cfg_l),
    .io_check_env_pmp_14_cfg_a(pmp_check_ptw_io_check_env_pmp_14_cfg_a),
    .io_check_env_pmp_14_cfg_x(pmp_check_ptw_io_check_env_pmp_14_cfg_x),
    .io_check_env_pmp_14_cfg_w(pmp_check_ptw_io_check_env_pmp_14_cfg_w),
    .io_check_env_pmp_14_cfg_r(pmp_check_ptw_io_check_env_pmp_14_cfg_r),
    .io_check_env_pmp_14_addr(pmp_check_ptw_io_check_env_pmp_14_addr),
    .io_check_env_pmp_14_mask(pmp_check_ptw_io_check_env_pmp_14_mask),
    .io_check_env_pmp_15_cfg_l(pmp_check_ptw_io_check_env_pmp_15_cfg_l),
    .io_check_env_pmp_15_cfg_a(pmp_check_ptw_io_check_env_pmp_15_cfg_a),
    .io_check_env_pmp_15_cfg_x(pmp_check_ptw_io_check_env_pmp_15_cfg_x),
    .io_check_env_pmp_15_cfg_w(pmp_check_ptw_io_check_env_pmp_15_cfg_w),
    .io_check_env_pmp_15_cfg_r(pmp_check_ptw_io_check_env_pmp_15_cfg_r),
    .io_check_env_pmp_15_addr(pmp_check_ptw_io_check_env_pmp_15_addr),
    .io_check_env_pmp_15_mask(pmp_check_ptw_io_check_env_pmp_15_mask),
    .io_check_env_pma_0_cfg_c(pmp_check_ptw_io_check_env_pma_0_cfg_c),
    .io_check_env_pma_0_cfg_atomic(pmp_check_ptw_io_check_env_pma_0_cfg_atomic),
    .io_check_env_pma_0_cfg_a(pmp_check_ptw_io_check_env_pma_0_cfg_a),
    .io_check_env_pma_0_cfg_x(pmp_check_ptw_io_check_env_pma_0_cfg_x),
    .io_check_env_pma_0_cfg_w(pmp_check_ptw_io_check_env_pma_0_cfg_w),
    .io_check_env_pma_0_cfg_r(pmp_check_ptw_io_check_env_pma_0_cfg_r),
    .io_check_env_pma_0_addr(pmp_check_ptw_io_check_env_pma_0_addr),
    .io_check_env_pma_0_mask(pmp_check_ptw_io_check_env_pma_0_mask),
    .io_check_env_pma_1_cfg_c(pmp_check_ptw_io_check_env_pma_1_cfg_c),
    .io_check_env_pma_1_cfg_atomic(pmp_check_ptw_io_check_env_pma_1_cfg_atomic),
    .io_check_env_pma_1_cfg_a(pmp_check_ptw_io_check_env_pma_1_cfg_a),
    .io_check_env_pma_1_cfg_x(pmp_check_ptw_io_check_env_pma_1_cfg_x),
    .io_check_env_pma_1_cfg_w(pmp_check_ptw_io_check_env_pma_1_cfg_w),
    .io_check_env_pma_1_cfg_r(pmp_check_ptw_io_check_env_pma_1_cfg_r),
    .io_check_env_pma_1_addr(pmp_check_ptw_io_check_env_pma_1_addr),
    .io_check_env_pma_1_mask(pmp_check_ptw_io_check_env_pma_1_mask),
    .io_check_env_pma_2_cfg_c(pmp_check_ptw_io_check_env_pma_2_cfg_c),
    .io_check_env_pma_2_cfg_atomic(pmp_check_ptw_io_check_env_pma_2_cfg_atomic),
    .io_check_env_pma_2_cfg_a(pmp_check_ptw_io_check_env_pma_2_cfg_a),
    .io_check_env_pma_2_cfg_x(pmp_check_ptw_io_check_env_pma_2_cfg_x),
    .io_check_env_pma_2_cfg_w(pmp_check_ptw_io_check_env_pma_2_cfg_w),
    .io_check_env_pma_2_cfg_r(pmp_check_ptw_io_check_env_pma_2_cfg_r),
    .io_check_env_pma_2_addr(pmp_check_ptw_io_check_env_pma_2_addr),
    .io_check_env_pma_2_mask(pmp_check_ptw_io_check_env_pma_2_mask),
    .io_check_env_pma_3_cfg_c(pmp_check_ptw_io_check_env_pma_3_cfg_c),
    .io_check_env_pma_3_cfg_atomic(pmp_check_ptw_io_check_env_pma_3_cfg_atomic),
    .io_check_env_pma_3_cfg_a(pmp_check_ptw_io_check_env_pma_3_cfg_a),
    .io_check_env_pma_3_cfg_x(pmp_check_ptw_io_check_env_pma_3_cfg_x),
    .io_check_env_pma_3_cfg_w(pmp_check_ptw_io_check_env_pma_3_cfg_w),
    .io_check_env_pma_3_cfg_r(pmp_check_ptw_io_check_env_pma_3_cfg_r),
    .io_check_env_pma_3_addr(pmp_check_ptw_io_check_env_pma_3_addr),
    .io_check_env_pma_3_mask(pmp_check_ptw_io_check_env_pma_3_mask),
    .io_check_env_pma_4_cfg_c(pmp_check_ptw_io_check_env_pma_4_cfg_c),
    .io_check_env_pma_4_cfg_atomic(pmp_check_ptw_io_check_env_pma_4_cfg_atomic),
    .io_check_env_pma_4_cfg_a(pmp_check_ptw_io_check_env_pma_4_cfg_a),
    .io_check_env_pma_4_cfg_x(pmp_check_ptw_io_check_env_pma_4_cfg_x),
    .io_check_env_pma_4_cfg_w(pmp_check_ptw_io_check_env_pma_4_cfg_w),
    .io_check_env_pma_4_cfg_r(pmp_check_ptw_io_check_env_pma_4_cfg_r),
    .io_check_env_pma_4_addr(pmp_check_ptw_io_check_env_pma_4_addr),
    .io_check_env_pma_4_mask(pmp_check_ptw_io_check_env_pma_4_mask),
    .io_check_env_pma_5_cfg_c(pmp_check_ptw_io_check_env_pma_5_cfg_c),
    .io_check_env_pma_5_cfg_atomic(pmp_check_ptw_io_check_env_pma_5_cfg_atomic),
    .io_check_env_pma_5_cfg_a(pmp_check_ptw_io_check_env_pma_5_cfg_a),
    .io_check_env_pma_5_cfg_x(pmp_check_ptw_io_check_env_pma_5_cfg_x),
    .io_check_env_pma_5_cfg_w(pmp_check_ptw_io_check_env_pma_5_cfg_w),
    .io_check_env_pma_5_cfg_r(pmp_check_ptw_io_check_env_pma_5_cfg_r),
    .io_check_env_pma_5_addr(pmp_check_ptw_io_check_env_pma_5_addr),
    .io_check_env_pma_5_mask(pmp_check_ptw_io_check_env_pma_5_mask),
    .io_check_env_pma_6_cfg_c(pmp_check_ptw_io_check_env_pma_6_cfg_c),
    .io_check_env_pma_6_cfg_atomic(pmp_check_ptw_io_check_env_pma_6_cfg_atomic),
    .io_check_env_pma_6_cfg_a(pmp_check_ptw_io_check_env_pma_6_cfg_a),
    .io_check_env_pma_6_cfg_x(pmp_check_ptw_io_check_env_pma_6_cfg_x),
    .io_check_env_pma_6_cfg_w(pmp_check_ptw_io_check_env_pma_6_cfg_w),
    .io_check_env_pma_6_cfg_r(pmp_check_ptw_io_check_env_pma_6_cfg_r),
    .io_check_env_pma_6_addr(pmp_check_ptw_io_check_env_pma_6_addr),
    .io_check_env_pma_6_mask(pmp_check_ptw_io_check_env_pma_6_mask),
    .io_check_env_pma_7_cfg_c(pmp_check_ptw_io_check_env_pma_7_cfg_c),
    .io_check_env_pma_7_cfg_atomic(pmp_check_ptw_io_check_env_pma_7_cfg_atomic),
    .io_check_env_pma_7_cfg_a(pmp_check_ptw_io_check_env_pma_7_cfg_a),
    .io_check_env_pma_7_cfg_x(pmp_check_ptw_io_check_env_pma_7_cfg_x),
    .io_check_env_pma_7_cfg_w(pmp_check_ptw_io_check_env_pma_7_cfg_w),
    .io_check_env_pma_7_cfg_r(pmp_check_ptw_io_check_env_pma_7_cfg_r),
    .io_check_env_pma_7_addr(pmp_check_ptw_io_check_env_pma_7_addr),
    .io_check_env_pma_7_mask(pmp_check_ptw_io_check_env_pma_7_mask),
    .io_check_env_pma_8_cfg_c(pmp_check_ptw_io_check_env_pma_8_cfg_c),
    .io_check_env_pma_8_cfg_atomic(pmp_check_ptw_io_check_env_pma_8_cfg_atomic),
    .io_check_env_pma_8_cfg_a(pmp_check_ptw_io_check_env_pma_8_cfg_a),
    .io_check_env_pma_8_cfg_x(pmp_check_ptw_io_check_env_pma_8_cfg_x),
    .io_check_env_pma_8_cfg_w(pmp_check_ptw_io_check_env_pma_8_cfg_w),
    .io_check_env_pma_8_cfg_r(pmp_check_ptw_io_check_env_pma_8_cfg_r),
    .io_check_env_pma_8_addr(pmp_check_ptw_io_check_env_pma_8_addr),
    .io_check_env_pma_8_mask(pmp_check_ptw_io_check_env_pma_8_mask),
    .io_check_env_pma_9_cfg_c(pmp_check_ptw_io_check_env_pma_9_cfg_c),
    .io_check_env_pma_9_cfg_atomic(pmp_check_ptw_io_check_env_pma_9_cfg_atomic),
    .io_check_env_pma_9_cfg_a(pmp_check_ptw_io_check_env_pma_9_cfg_a),
    .io_check_env_pma_9_cfg_x(pmp_check_ptw_io_check_env_pma_9_cfg_x),
    .io_check_env_pma_9_cfg_w(pmp_check_ptw_io_check_env_pma_9_cfg_w),
    .io_check_env_pma_9_cfg_r(pmp_check_ptw_io_check_env_pma_9_cfg_r),
    .io_check_env_pma_9_addr(pmp_check_ptw_io_check_env_pma_9_addr),
    .io_check_env_pma_9_mask(pmp_check_ptw_io_check_env_pma_9_mask),
    .io_check_env_pma_10_cfg_c(pmp_check_ptw_io_check_env_pma_10_cfg_c),
    .io_check_env_pma_10_cfg_atomic(pmp_check_ptw_io_check_env_pma_10_cfg_atomic),
    .io_check_env_pma_10_cfg_a(pmp_check_ptw_io_check_env_pma_10_cfg_a),
    .io_check_env_pma_10_cfg_x(pmp_check_ptw_io_check_env_pma_10_cfg_x),
    .io_check_env_pma_10_cfg_w(pmp_check_ptw_io_check_env_pma_10_cfg_w),
    .io_check_env_pma_10_cfg_r(pmp_check_ptw_io_check_env_pma_10_cfg_r),
    .io_check_env_pma_10_addr(pmp_check_ptw_io_check_env_pma_10_addr),
    .io_check_env_pma_10_mask(pmp_check_ptw_io_check_env_pma_10_mask),
    .io_check_env_pma_11_cfg_c(pmp_check_ptw_io_check_env_pma_11_cfg_c),
    .io_check_env_pma_11_cfg_atomic(pmp_check_ptw_io_check_env_pma_11_cfg_atomic),
    .io_check_env_pma_11_cfg_a(pmp_check_ptw_io_check_env_pma_11_cfg_a),
    .io_check_env_pma_11_cfg_x(pmp_check_ptw_io_check_env_pma_11_cfg_x),
    .io_check_env_pma_11_cfg_w(pmp_check_ptw_io_check_env_pma_11_cfg_w),
    .io_check_env_pma_11_cfg_r(pmp_check_ptw_io_check_env_pma_11_cfg_r),
    .io_check_env_pma_11_addr(pmp_check_ptw_io_check_env_pma_11_addr),
    .io_check_env_pma_11_mask(pmp_check_ptw_io_check_env_pma_11_mask),
    .io_check_env_pma_12_cfg_c(pmp_check_ptw_io_check_env_pma_12_cfg_c),
    .io_check_env_pma_12_cfg_atomic(pmp_check_ptw_io_check_env_pma_12_cfg_atomic),
    .io_check_env_pma_12_cfg_a(pmp_check_ptw_io_check_env_pma_12_cfg_a),
    .io_check_env_pma_12_cfg_x(pmp_check_ptw_io_check_env_pma_12_cfg_x),
    .io_check_env_pma_12_cfg_w(pmp_check_ptw_io_check_env_pma_12_cfg_w),
    .io_check_env_pma_12_cfg_r(pmp_check_ptw_io_check_env_pma_12_cfg_r),
    .io_check_env_pma_12_addr(pmp_check_ptw_io_check_env_pma_12_addr),
    .io_check_env_pma_12_mask(pmp_check_ptw_io_check_env_pma_12_mask),
    .io_check_env_pma_13_cfg_c(pmp_check_ptw_io_check_env_pma_13_cfg_c),
    .io_check_env_pma_13_cfg_atomic(pmp_check_ptw_io_check_env_pma_13_cfg_atomic),
    .io_check_env_pma_13_cfg_a(pmp_check_ptw_io_check_env_pma_13_cfg_a),
    .io_check_env_pma_13_cfg_x(pmp_check_ptw_io_check_env_pma_13_cfg_x),
    .io_check_env_pma_13_cfg_w(pmp_check_ptw_io_check_env_pma_13_cfg_w),
    .io_check_env_pma_13_cfg_r(pmp_check_ptw_io_check_env_pma_13_cfg_r),
    .io_check_env_pma_13_addr(pmp_check_ptw_io_check_env_pma_13_addr),
    .io_check_env_pma_13_mask(pmp_check_ptw_io_check_env_pma_13_mask),
    .io_check_env_pma_14_cfg_c(pmp_check_ptw_io_check_env_pma_14_cfg_c),
    .io_check_env_pma_14_cfg_atomic(pmp_check_ptw_io_check_env_pma_14_cfg_atomic),
    .io_check_env_pma_14_cfg_a(pmp_check_ptw_io_check_env_pma_14_cfg_a),
    .io_check_env_pma_14_cfg_x(pmp_check_ptw_io_check_env_pma_14_cfg_x),
    .io_check_env_pma_14_cfg_w(pmp_check_ptw_io_check_env_pma_14_cfg_w),
    .io_check_env_pma_14_cfg_r(pmp_check_ptw_io_check_env_pma_14_cfg_r),
    .io_check_env_pma_14_addr(pmp_check_ptw_io_check_env_pma_14_addr),
    .io_check_env_pma_14_mask(pmp_check_ptw_io_check_env_pma_14_mask),
    .io_check_env_pma_15_cfg_c(pmp_check_ptw_io_check_env_pma_15_cfg_c),
    .io_check_env_pma_15_cfg_atomic(pmp_check_ptw_io_check_env_pma_15_cfg_atomic),
    .io_check_env_pma_15_cfg_a(pmp_check_ptw_io_check_env_pma_15_cfg_a),
    .io_check_env_pma_15_cfg_x(pmp_check_ptw_io_check_env_pma_15_cfg_x),
    .io_check_env_pma_15_cfg_w(pmp_check_ptw_io_check_env_pma_15_cfg_w),
    .io_check_env_pma_15_cfg_r(pmp_check_ptw_io_check_env_pma_15_cfg_r),
    .io_check_env_pma_15_addr(pmp_check_ptw_io_check_env_pma_15_addr),
    .io_check_env_pma_15_mask(pmp_check_ptw_io_check_env_pma_15_mask),
    .io_req_valid(pmp_check_ptw_io_req_valid),
    .io_req_bits_addr(pmp_check_ptw_io_req_bits_addr),
    .io_resp_c(pmp_check_ptw_io_resp_c),
    .io_resp_atomic(pmp_check_ptw_io_resp_atomic),
    .io_resp_x(pmp_check_ptw_io_resp_x),
    .io_resp_w(pmp_check_ptw_io_resp_w),
    .io_resp_r(pmp_check_ptw_io_resp_r)
  );
  PipelineRegModule_27 pipelineReg ( // @[MemCommon.scala 396:29]
    .clock(pipelineReg_clock),
    .reset(pipelineReg_reset),
    .io_in_ready(pipelineReg_io_in_ready),
    .io_in_valid(pipelineReg_io_in_valid),
    .io_in_bits_cmd(pipelineReg_io_in_bits_cmd),
    .io_in_bits_addr(pipelineReg_io_in_bits_addr),
    .io_in_bits_data(pipelineReg_io_in_bits_data),
    .io_in_bits_mask(pipelineReg_io_in_bits_mask),
    .io_in_bits_atomic(pipelineReg_io_in_bits_atomic),
    .io_out_ready(pipelineReg_io_out_ready),
    .io_out_valid(pipelineReg_io_out_valid),
    .io_out_bits_cmd(pipelineReg_io_out_bits_cmd),
    .io_out_bits_addr(pipelineReg_io_out_bits_addr),
    .io_out_bits_data(pipelineReg_io_out_bits_data),
    .io_out_bits_mask(pipelineReg_io_out_bits_mask),
    .io_out_bits_atomic(pipelineReg_io_out_bits_atomic)
  );
  PipelineRegModule_28 pipelineReg_1 ( // @[MemCommon.scala 396:29]
    .clock(pipelineReg_1_clock),
    .reset(pipelineReg_1_reset),
    .io_in_ready(pipelineReg_1_io_in_ready),
    .io_in_valid(pipelineReg_1_io_in_valid),
    .io_in_bits_data(pipelineReg_1_io_in_bits_data),
    .io_out_valid(pipelineReg_1_io_out_valid),
    .io_out_bits_data(pipelineReg_1_io_out_bits_data)
  );
  DelayN_246 delay ( // @[Hold.scala 97:23]
    .clock(delay_clock),
    .io_in(delay_io_in),
    .io_out(delay_io_out)
  );
  PFEvent pfevent ( // @[MemBlock.scala 687:23]
    .clock(pfevent_clock),
    .reset(pfevent_reset),
    .io_distribute_csr_wvalid(pfevent_io_distribute_csr_wvalid),
    .io_distribute_csr_waddr(pfevent_io_distribute_csr_waddr),
    .io_distribute_csr_wdata(pfevent_io_distribute_csr_wdata),
    .io_hpmevent_0(pfevent_io_hpmevent_0),
    .io_hpmevent_1(pfevent_io_hpmevent_1),
    .io_hpmevent_2(pfevent_io_hpmevent_2),
    .io_hpmevent_3(pfevent_io_hpmevent_3),
    .io_hpmevent_4(pfevent_io_hpmevent_4),
    .io_hpmevent_5(pfevent_io_hpmevent_5),
    .io_hpmevent_6(pfevent_io_hpmevent_6),
    .io_hpmevent_7(pfevent_io_hpmevent_7),
    .io_hpmevent_8(pfevent_io_hpmevent_8),
    .io_hpmevent_9(pfevent_io_hpmevent_9),
    .io_hpmevent_10(pfevent_io_hpmevent_10),
    .io_hpmevent_11(pfevent_io_hpmevent_11),
    .io_hpmevent_12(pfevent_io_hpmevent_12),
    .io_hpmevent_13(pfevent_io_hpmevent_13),
    .io_hpmevent_14(pfevent_io_hpmevent_14),
    .io_hpmevent_15(pfevent_io_hpmevent_15),
    .io_hpmevent_16(pfevent_io_hpmevent_16),
    .io_hpmevent_17(pfevent_io_hpmevent_17),
    .io_hpmevent_18(pfevent_io_hpmevent_18),
    .io_hpmevent_19(pfevent_io_hpmevent_19),
    .io_hpmevent_20(pfevent_io_hpmevent_20),
    .io_hpmevent_21(pfevent_io_hpmevent_21),
    .io_hpmevent_22(pfevent_io_hpmevent_22),
    .io_hpmevent_23(pfevent_io_hpmevent_23)
  );
  HPerfMonitor_2 hpm ( // @[PerfCounterUtils.scala 255:21]
    .clock(hpm_clock),
    .io_hpm_event_0(hpm_io_hpm_event_0),
    .io_hpm_event_1(hpm_io_hpm_event_1),
    .io_hpm_event_2(hpm_io_hpm_event_2),
    .io_hpm_event_3(hpm_io_hpm_event_3),
    .io_hpm_event_4(hpm_io_hpm_event_4),
    .io_hpm_event_5(hpm_io_hpm_event_5),
    .io_hpm_event_6(hpm_io_hpm_event_6),
    .io_hpm_event_7(hpm_io_hpm_event_7),
    .io_events_sets_0_value(hpm_io_events_sets_0_value),
    .io_events_sets_1_value(hpm_io_events_sets_1_value),
    .io_events_sets_2_value(hpm_io_events_sets_2_value),
    .io_events_sets_3_value(hpm_io_events_sets_3_value),
    .io_events_sets_4_value(hpm_io_events_sets_4_value),
    .io_events_sets_5_value(hpm_io_events_sets_5_value),
    .io_events_sets_6_value(hpm_io_events_sets_6_value),
    .io_events_sets_7_value(hpm_io_events_sets_7_value),
    .io_events_sets_8_value(hpm_io_events_sets_8_value),
    .io_events_sets_9_value(hpm_io_events_sets_9_value),
    .io_events_sets_10_value(hpm_io_events_sets_10_value),
    .io_events_sets_11_value(hpm_io_events_sets_11_value),
    .io_events_sets_12_value(hpm_io_events_sets_12_value),
    .io_events_sets_13_value(hpm_io_events_sets_13_value),
    .io_events_sets_14_value(hpm_io_events_sets_14_value),
    .io_events_sets_15_value(hpm_io_events_sets_15_value),
    .io_events_sets_16_value(hpm_io_events_sets_16_value),
    .io_events_sets_17_value(hpm_io_events_sets_17_value),
    .io_events_sets_18_value(hpm_io_events_sets_18_value),
    .io_events_sets_19_value(hpm_io_events_sets_19_value),
    .io_events_sets_20_value(hpm_io_events_sets_20_value),
    .io_events_sets_21_value(hpm_io_events_sets_21_value),
    .io_events_sets_22_value(hpm_io_events_sets_22_value),
    .io_events_sets_23_value(hpm_io_events_sets_23_value),
    .io_events_sets_24_value(hpm_io_events_sets_24_value),
    .io_events_sets_25_value(hpm_io_events_sets_25_value),
    .io_events_sets_26_value(hpm_io_events_sets_26_value),
    .io_events_sets_27_value(hpm_io_events_sets_27_value),
    .io_events_sets_28_value(hpm_io_events_sets_28_value),
    .io_events_sets_29_value(hpm_io_events_sets_29_value),
    .io_events_sets_30_value(hpm_io_events_sets_30_value),
    .io_events_sets_31_value(hpm_io_events_sets_31_value),
    .io_events_sets_32_value(hpm_io_events_sets_32_value),
    .io_events_sets_33_value(hpm_io_events_sets_33_value),
    .io_events_sets_34_value(hpm_io_events_sets_34_value),
    .io_events_sets_35_value(hpm_io_events_sets_35_value),
    .io_events_sets_36_value(hpm_io_events_sets_36_value),
    .io_events_sets_37_value(hpm_io_events_sets_37_value),
    .io_events_sets_38_value(hpm_io_events_sets_38_value),
    .io_events_sets_39_value(hpm_io_events_sets_39_value),
    .io_events_sets_40_value(hpm_io_events_sets_40_value),
    .io_events_sets_41_value(hpm_io_events_sets_41_value),
    .io_events_sets_42_value(hpm_io_events_sets_42_value),
    .io_events_sets_43_value(hpm_io_events_sets_43_value),
    .io_events_sets_44_value(hpm_io_events_sets_44_value),
    .io_events_sets_45_value(hpm_io_events_sets_45_value),
    .io_events_sets_46_value(hpm_io_events_sets_46_value),
    .io_events_sets_47_value(hpm_io_events_sets_47_value),
    .io_events_sets_48_value(hpm_io_events_sets_48_value),
    .io_events_sets_49_value(hpm_io_events_sets_49_value),
    .io_events_sets_50_value(hpm_io_events_sets_50_value),
    .io_events_sets_51_value(hpm_io_events_sets_51_value),
    .io_events_sets_52_value(hpm_io_events_sets_52_value),
    .io_events_sets_53_value(hpm_io_events_sets_53_value),
    .io_events_sets_54_value(hpm_io_events_sets_54_value),
    .io_events_sets_55_value(hpm_io_events_sets_55_value),
    .io_events_sets_56_value(hpm_io_events_sets_56_value),
    .io_events_sets_57_value(hpm_io_events_sets_57_value),
    .io_events_sets_58_value(hpm_io_events_sets_58_value),
    .io_events_sets_59_value(hpm_io_events_sets_59_value),
    .io_events_sets_60_value(hpm_io_events_sets_60_value),
    .io_events_sets_61_value(hpm_io_events_sets_61_value),
    .io_events_sets_62_value(hpm_io_events_sets_62_value),
    .io_events_sets_63_value(hpm_io_events_sets_63_value),
    .io_events_sets_64_value(hpm_io_events_sets_64_value),
    .io_events_sets_65_value(hpm_io_events_sets_65_value),
    .io_events_sets_66_value(hpm_io_events_sets_66_value),
    .io_events_sets_67_value(hpm_io_events_sets_67_value),
    .io_events_sets_68_value(hpm_io_events_sets_68_value),
    .io_events_sets_69_value(hpm_io_events_sets_69_value),
    .io_events_sets_70_value(hpm_io_events_sets_70_value),
    .io_events_sets_71_value(hpm_io_events_sets_71_value),
    .io_events_sets_72_value(hpm_io_events_sets_72_value),
    .io_events_sets_73_value(hpm_io_events_sets_73_value),
    .io_events_sets_74_value(hpm_io_events_sets_74_value),
    .io_events_sets_75_value(hpm_io_events_sets_75_value),
    .io_events_sets_76_value(hpm_io_events_sets_76_value),
    .io_events_sets_77_value(hpm_io_events_sets_77_value),
    .io_events_sets_78_value(hpm_io_events_sets_78_value),
    .io_events_sets_79_value(hpm_io_events_sets_79_value),
    .io_events_sets_80_value(hpm_io_events_sets_80_value),
    .io_events_sets_81_value(hpm_io_events_sets_81_value),
    .io_events_sets_82_value(hpm_io_events_sets_82_value),
    .io_events_sets_83_value(hpm_io_events_sets_83_value),
    .io_events_sets_84_value(hpm_io_events_sets_84_value),
    .io_events_sets_85_value(hpm_io_events_sets_85_value),
    .io_events_sets_86_value(hpm_io_events_sets_86_value),
    .io_events_sets_87_value(hpm_io_events_sets_87_value),
    .io_events_sets_88_value(hpm_io_events_sets_88_value),
    .io_events_sets_89_value(hpm_io_events_sets_89_value),
    .io_events_sets_90_value(hpm_io_events_sets_90_value),
    .io_events_sets_91_value(hpm_io_events_sets_91_value),
    .io_events_sets_92_value(hpm_io_events_sets_92_value),
    .io_events_sets_93_value(hpm_io_events_sets_93_value),
    .io_events_sets_94_value(hpm_io_events_sets_94_value),
    .io_events_sets_95_value(hpm_io_events_sets_95_value),
    .io_events_sets_96_value(hpm_io_events_sets_96_value),
    .io_events_sets_97_value(hpm_io_events_sets_97_value),
    .io_events_sets_98_value(hpm_io_events_sets_98_value),
    .io_events_sets_99_value(hpm_io_events_sets_99_value),
    .io_events_sets_100_value(hpm_io_events_sets_100_value),
    .io_events_sets_101_value(hpm_io_events_sets_101_value),
    .io_events_sets_102_value(hpm_io_events_sets_102_value),
    .io_events_sets_103_value(hpm_io_events_sets_103_value),
    .io_events_sets_104_value(hpm_io_events_sets_104_value),
    .io_events_sets_105_value(hpm_io_events_sets_105_value),
    .io_events_sets_106_value(hpm_io_events_sets_106_value),
    .io_events_sets_107_value(hpm_io_events_sets_107_value),
    .io_events_sets_108_value(hpm_io_events_sets_108_value),
    .io_perf_0_value(hpm_io_perf_0_value),
    .io_perf_1_value(hpm_io_perf_1_value),
    .io_perf_2_value(hpm_io_perf_2_value),
    .io_perf_3_value(hpm_io_perf_3_value),
    .io_perf_4_value(hpm_io_perf_4_value),
    .io_perf_5_value(hpm_io_perf_5_value),
    .io_perf_6_value(hpm_io_perf_6_value),
    .io_perf_7_value(hpm_io_perf_7_value)
  );
  assign auto_uncache_client_out_a_valid = uncache_auto_client_out_a_valid; // @[LazyModule.scala 311:12]
  assign auto_uncache_client_out_a_bits_opcode = uncache_auto_client_out_a_bits_opcode; // @[LazyModule.scala 311:12]
  assign auto_uncache_client_out_a_bits_size = uncache_auto_client_out_a_bits_size; // @[LazyModule.scala 311:12]
  assign auto_uncache_client_out_a_bits_source = uncache_auto_client_out_a_bits_source; // @[LazyModule.scala 311:12]
  assign auto_uncache_client_out_a_bits_address = uncache_auto_client_out_a_bits_address; // @[LazyModule.scala 311:12]
  assign auto_uncache_client_out_a_bits_mask = uncache_auto_client_out_a_bits_mask; // @[LazyModule.scala 311:12]
  assign auto_uncache_client_out_a_bits_data = uncache_auto_client_out_a_bits_data; // @[LazyModule.scala 311:12]
  assign auto_uncache_client_out_d_ready = uncache_auto_client_out_d_ready; // @[LazyModule.scala 311:12]
  assign auto_dcache_client_out_a_valid = dcache_auto_client_out_a_valid; // @[LazyModule.scala 311:12]
  assign auto_dcache_client_out_a_bits_opcode = dcache_auto_client_out_a_bits_opcode; // @[LazyModule.scala 311:12]
  assign auto_dcache_client_out_a_bits_param = dcache_auto_client_out_a_bits_param; // @[LazyModule.scala 311:12]
  assign auto_dcache_client_out_a_bits_size = dcache_auto_client_out_a_bits_size; // @[LazyModule.scala 311:12]
  assign auto_dcache_client_out_a_bits_source = dcache_auto_client_out_a_bits_source; // @[LazyModule.scala 311:12]
  assign auto_dcache_client_out_a_bits_address = dcache_auto_client_out_a_bits_address; // @[LazyModule.scala 311:12]
  assign auto_dcache_client_out_a_bits_mask = dcache_auto_client_out_a_bits_mask; // @[LazyModule.scala 311:12]
  assign auto_dcache_client_out_bready = dcache_auto_client_out_bready; // @[LazyModule.scala 311:12]
  assign auto_dcache_client_out_c_valid = dcache_auto_client_out_c_valid; // @[LazyModule.scala 311:12]
  assign auto_dcache_client_out_c_bits_opcode = dcache_auto_client_out_c_bits_opcode; // @[LazyModule.scala 311:12]
  assign auto_dcache_client_out_c_bits_param = dcache_auto_client_out_c_bits_param; // @[LazyModule.scala 311:12]
  assign auto_dcache_client_out_c_bits_size = dcache_auto_client_out_c_bits_size; // @[LazyModule.scala 311:12]
  assign auto_dcache_client_out_c_bits_source = dcache_auto_client_out_c_bits_source; // @[LazyModule.scala 311:12]
  assign auto_dcache_client_out_c_bits_address = dcache_auto_client_out_c_bits_address; // @[LazyModule.scala 311:12]
  assign auto_dcache_client_out_c_bits_echo_blockisdirty = dcache_auto_client_out_c_bits_echo_blockisdirty; // @[LazyModule.scala 311:12]
  assign auto_dcache_client_out_c_bits_data = dcache_auto_client_out_c_bits_data; // @[LazyModule.scala 311:12]
  assign auto_dcache_client_out_d_ready = dcache_auto_client_out_d_ready; // @[LazyModule.scala 311:12]
  assign auto_dcache_client_out_e_valid = dcache_auto_client_out_e_valid; // @[LazyModule.scala 311:12]
  assign auto_dcache_client_out_e_bits_sink = dcache_auto_client_out_e_bits_sink; // @[LazyModule.scala 311:12]
  assign io_issue_0_ready = LoadUnit_0_io_loadIn_ready; // @[MemBlock.scala 344:28]
  assign io_issue_1_ready = LoadUnit_1_io_loadIn_ready; // @[MemBlock.scala 344:28]
  assign io_issue_2_ready = st_atomics_0 ? atomicsUnit_io_in_ready : 1'h1; // @[MemBlock.scala 460:25 602:63 603:34]
  assign io_issue_3_ready = st_atomics_1 ? atomicsUnit_io_in_ready : 1'h1; // @[MemBlock.scala 460:25 602:63 603:34]
  assign io_issue_4_ready = stdExeUnits_0_io_fromInt_ready; // @[MemBlock.scala 451:31]
  assign io_issue_5_ready = stdExeUnits_1_io_fromInt_ready; // @[MemBlock.scala 451:31]
  assign io_rsfeedback_0_feedbackSlow_valid = _T_43 ? atomicsUnit_io_feedbackSlow_valid :
    StoreUnit_0_io_feedbackSlow_valid; // @[MemBlock.scala 456:25 652:73 653:33]
  assign io_rsfeedback_0_feedbackSlow_bits_rsIdx = _T_43 ? atomicsUnit_io_feedbackSlow_bits_rsIdx :
    StoreUnit_0_io_feedbackSlow_bits_rsIdx; // @[MemBlock.scala 456:25 652:73 653:33]
  assign io_rsfeedback_0_feedbackSlow_bits_hit = _T_43 | StoreUnit_0_io_feedbackSlow_bits_hit; // @[MemBlock.scala 456:25 652:73 653:33]
  assign io_rsfeedback_1_feedbackSlow_valid = _T_44 ? atomicsUnit_io_feedbackSlow_valid :
    StoreUnit_1_io_feedbackSlow_valid; // @[MemBlock.scala 456:25 652:73 653:33]
  assign io_rsfeedback_1_feedbackSlow_bits_rsIdx = _T_44 ? atomicsUnit_io_feedbackSlow_bits_rsIdx :
    StoreUnit_1_io_feedbackSlow_bits_rsIdx; // @[MemBlock.scala 456:25 652:73 653:33]
  assign io_rsfeedback_1_feedbackSlow_bits_hit = _T_44 | StoreUnit_1_io_feedbackSlow_bits_hit; // @[MemBlock.scala 456:25 652:73 653:33]
  assign io_writeback_0_valid = atomicsUnit_io_out_valid | LoadUnit_0_io_loadOut_valid; // @[MemBlock.scala 184:46]
  assign io_writeback_0_bits_uop_cf_exceptionVec_4 = atomicsUnit_io_out_valid ? 1'h0 :
    loadWritebackOverride_uop_cf_exceptionVec_4; // @[MemBlock.scala 185:18 188:33 189:39]
  assign io_writeback_0_bits_uop_cf_exceptionVec_5 = atomicsUnit_io_out_valid ? 1'h0 :
    loadWritebackOverride_uop_cf_exceptionVec_5; // @[MemBlock.scala 185:18 188:33 189:39]
  assign io_writeback_0_bits_uop_cf_exceptionVec_13 = atomicsUnit_io_out_valid ? 1'h0 :
    loadWritebackOverride_uop_cf_exceptionVec_13; // @[MemBlock.scala 185:18 188:33 189:39]
  assign io_writeback_0_bits_uop_cf_trigger_backendEn_1 = atomicsUnit_io_out_valid ?
    atomicsUnit_io_out_bits_uop_cf_trigger_backendEn_1 : LoadUnit_0_io_loadOut_bits_uop_cf_trigger_backendEn_1; // @[MemBlock.scala 182:35]
  assign io_writeback_0_bits_uop_cf_trigger_backendHit_0 = atomicsUnit_io_out_valid ? 1'h0 : _GEN_200; // @[MemBlock.scala 521:35 529:54]
  assign io_writeback_0_bits_uop_cf_trigger_backendHit_1 = atomicsUnit_io_out_valid ? 1'h0 : _GEN_201; // @[MemBlock.scala 521:35 529:54]
  assign io_writeback_0_bits_uop_cf_trigger_backendHit_2 = atomicsUnit_io_out_valid ? 1'h0 : _GEN_188; // @[MemBlock.scala 521:35 529:54]
  assign io_writeback_0_bits_uop_cf_trigger_backendHit_3 = atomicsUnit_io_out_valid ? 1'h0 : _GEN_189; // @[MemBlock.scala 521:35 529:54]
  assign io_writeback_0_bits_uop_cf_trigger_backendHit_4 = atomicsUnit_io_out_valid ? 1'h0 :
    loadWritebackOverride_uop_cf_trigger_backendHit_4; // @[MemBlock.scala 193:16 521:35 529:54]
  assign io_writeback_0_bits_uop_cf_trigger_backendHit_5 = atomicsUnit_io_out_valid ? 1'h0 : _GEN_190; // @[MemBlock.scala 521:35 529:54]
  assign io_writeback_0_bits_uop_ctrl_rfWen = atomicsUnit_io_out_valid ? atomicsUnit_io_out_bits_uop_ctrl_rfWen :
    LoadUnit_0_io_loadOut_bits_uop_ctrl_rfWen; // @[MemBlock.scala 182:35]
  assign io_writeback_0_bits_uop_ctrl_fpWen = atomicsUnit_io_out_valid ? atomicsUnit_io_out_bits_uop_ctrl_fpWen :
    LoadUnit_0_io_loadOut_bits_uop_ctrl_fpWen; // @[MemBlock.scala 182:35]
  assign io_writeback_0_bits_uop_ctrl_flushPipe = atomicsUnit_io_out_valid ? 1'h0 :
    LoadUnit_0_io_loadOut_bits_uop_ctrl_flushPipe; // @[MemBlock.scala 182:35]
  assign io_writeback_0_bits_uop_ctrl_replayInst = atomicsUnit_io_out_valid ? 1'h0 :
    LoadUnit_0_io_loadOut_bits_uop_ctrl_replayInst; // @[MemBlock.scala 182:35]
  assign io_writeback_0_bits_uop_pdest = atomicsUnit_io_out_valid ? atomicsUnit_io_out_bits_uop_pdest :
    LoadUnit_0_io_loadOut_bits_uop_pdest; // @[MemBlock.scala 182:35]
  assign io_writeback_0_bits_uop_robIdx_flag = atomicsUnit_io_out_valid ? atomicsUnit_io_out_bits_uop_robIdx_flag :
    LoadUnit_0_io_loadOut_bits_uop_robIdx_flag; // @[MemBlock.scala 182:35]
  assign io_writeback_0_bits_uop_robIdx_value = atomicsUnit_io_out_valid ? atomicsUnit_io_out_bits_uop_robIdx_value :
    LoadUnit_0_io_loadOut_bits_uop_robIdx_value; // @[MemBlock.scala 182:35]
  assign io_writeback_0_bits_data = atomicsUnit_io_out_valid ? atomicsUnit_io_out_bits_data :
    LoadUnit_0_io_loadOut_bits_data; // @[MemBlock.scala 182:35]
  assign io_writeback_0_bits_debug_isMMIO = atomicsUnit_io_out_valid ? atomicsUnit_io_out_bits_debug_isMMIO :
    LoadUnit_0_io_loadOut_bits_debug_isMMIO; // @[MemBlock.scala 182:35]
  assign io_writeback_1_valid = LoadUnit_1_io_loadOut_valid; // @[MemBlock.scala 193:16]
  assign io_writeback_1_bits_uop_cf_exceptionVec_4 = LoadUnit_1_io_loadOut_bits_uop_cf_exceptionVec_4; // @[MemBlock.scala 193:16]
  assign io_writeback_1_bits_uop_cf_exceptionVec_5 = LoadUnit_1_io_loadOut_bits_uop_cf_exceptionVec_5; // @[MemBlock.scala 193:16]
  assign io_writeback_1_bits_uop_cf_exceptionVec_13 = LoadUnit_1_io_loadOut_bits_uop_cf_exceptionVec_13; // @[MemBlock.scala 193:16]
  assign io_writeback_1_bits_uop_cf_trigger_backendEn_1 = LoadUnit_1_io_loadOut_bits_uop_cf_trigger_backendEn_1; // @[MemBlock.scala 193:16]
  assign io_writeback_1_bits_uop_cf_trigger_backendHit_0 = atomicsUnit_io_out_valid ? 1'h0 : _GEN_208; // @[MemBlock.scala 521:35 529:54]
  assign io_writeback_1_bits_uop_cf_trigger_backendHit_1 = atomicsUnit_io_out_valid ? 1'h0 : _GEN_209; // @[MemBlock.scala 521:35 529:54]
  assign io_writeback_1_bits_uop_cf_trigger_backendHit_2 = atomicsUnit_io_out_valid ? 1'h0 : _GEN_191; // @[MemBlock.scala 521:35 529:54]
  assign io_writeback_1_bits_uop_cf_trigger_backendHit_3 = atomicsUnit_io_out_valid ? 1'h0 : _GEN_192; // @[MemBlock.scala 521:35 529:54]
  assign io_writeback_1_bits_uop_cf_trigger_backendHit_4 = atomicsUnit_io_out_valid ? 1'h0 :
    LoadUnit_1_io_loadOut_bits_uop_cf_trigger_backendHit_4; // @[MemBlock.scala 193:16 521:35 529:54]
  assign io_writeback_1_bits_uop_cf_trigger_backendHit_5 = atomicsUnit_io_out_valid ? 1'h0 : _GEN_193; // @[MemBlock.scala 521:35 529:54]
  assign io_writeback_1_bits_uop_ctrl_rfWen = LoadUnit_1_io_loadOut_bits_uop_ctrl_rfWen; // @[MemBlock.scala 193:16]
  assign io_writeback_1_bits_uop_ctrl_fpWen = LoadUnit_1_io_loadOut_bits_uop_ctrl_fpWen; // @[MemBlock.scala 193:16]
  assign io_writeback_1_bits_uop_ctrl_flushPipe = LoadUnit_1_io_loadOut_bits_uop_ctrl_flushPipe; // @[MemBlock.scala 193:16]
  assign io_writeback_1_bits_uop_ctrl_replayInst = LoadUnit_1_io_loadOut_bits_uop_ctrl_replayInst; // @[MemBlock.scala 193:16]
  assign io_writeback_1_bits_uop_pdest = LoadUnit_1_io_loadOut_bits_uop_pdest; // @[MemBlock.scala 193:16]
  assign io_writeback_1_bits_uop_robIdx_flag = LoadUnit_1_io_loadOut_bits_uop_robIdx_flag; // @[MemBlock.scala 193:16]
  assign io_writeback_1_bits_uop_robIdx_value = LoadUnit_1_io_loadOut_bits_uop_robIdx_value; // @[MemBlock.scala 193:16]
  assign io_writeback_1_bits_data = LoadUnit_1_io_loadOut_bits_data; // @[MemBlock.scala 193:16]
  assign io_writeback_1_bits_debug_isMMIO = LoadUnit_1_io_loadOut_bits_debug_isMMIO; // @[MemBlock.scala 193:16]
  assign io_writeback_2_valid = atomicsUnit_io_out_valid | _GEN_210; // @[MemBlock.scala 521:35 523:20]
  assign io_writeback_2_bits_uop_cf_exceptionVec_4 = atomicsUnit_io_out_valid &
    atomicsUnit_io_out_bits_uop_cf_exceptionVec_4; // @[MemBlock.scala 521:35 524:20]
  assign io_writeback_2_bits_uop_cf_exceptionVec_5 = atomicsUnit_io_out_valid &
    atomicsUnit_io_out_bits_uop_cf_exceptionVec_5; // @[MemBlock.scala 521:35 524:20]
  assign io_writeback_2_bits_uop_cf_exceptionVec_6 = atomicsUnit_io_out_valid ?
    atomicsUnit_io_out_bits_uop_cf_exceptionVec_6 : _GEN_220; // @[MemBlock.scala 521:35 524:20]
  assign io_writeback_2_bits_uop_cf_exceptionVec_7 = atomicsUnit_io_out_valid ?
    atomicsUnit_io_out_bits_uop_cf_exceptionVec_7 : _GEN_221; // @[MemBlock.scala 521:35 524:20]
  assign io_writeback_2_bits_uop_cf_exceptionVec_13 = atomicsUnit_io_out_valid &
    atomicsUnit_io_out_bits_uop_cf_exceptionVec_13; // @[MemBlock.scala 521:35 524:20]
  assign io_writeback_2_bits_uop_cf_exceptionVec_15 = atomicsUnit_io_out_valid ?
    atomicsUnit_io_out_bits_uop_cf_exceptionVec_15 : _GEN_229; // @[MemBlock.scala 521:35 524:20]
  assign io_writeback_2_bits_uop_cf_trigger_backendEn_0 = atomicsUnit_io_out_valid ?
    atomicsUnit_io_out_bits_uop_cf_trigger_backendEn_0 : _GEN_234; // @[MemBlock.scala 521:35 524:20]
  assign io_writeback_2_bits_uop_cf_trigger_backendHit_0 = atomicsUnit_io_out_valid ?
    atomicsUnit_io_out_bits_uop_cf_trigger_backendHit_0 : _GEN_236; // @[MemBlock.scala 521:35 524:20]
  assign io_writeback_2_bits_uop_cf_trigger_backendHit_1 = atomicsUnit_io_out_valid ?
    atomicsUnit_io_out_bits_uop_cf_trigger_backendHit_1 : _GEN_237; // @[MemBlock.scala 521:35 524:20]
  assign io_writeback_2_bits_uop_cf_trigger_backendHit_2 = atomicsUnit_io_out_valid &
    atomicsUnit_io_out_bits_uop_cf_trigger_backendHit_2; // @[MemBlock.scala 521:35 524:20]
  assign io_writeback_2_bits_uop_cf_trigger_backendHit_3 = atomicsUnit_io_out_valid &
    atomicsUnit_io_out_bits_uop_cf_trigger_backendHit_3; // @[MemBlock.scala 521:35 524:20]
  assign io_writeback_2_bits_uop_cf_trigger_backendHit_4 = atomicsUnit_io_out_valid ?
    atomicsUnit_io_out_bits_uop_cf_trigger_backendHit_4 : _GEN_240; // @[MemBlock.scala 521:35 524:20]
  assign io_writeback_2_bits_uop_cf_trigger_backendHit_5 = atomicsUnit_io_out_valid &
    atomicsUnit_io_out_bits_uop_cf_trigger_backendHit_5; // @[MemBlock.scala 521:35 524:20]
  assign io_writeback_2_bits_uop_robIdx_flag = atomicsUnit_io_out_valid ? atomicsUnit_io_out_bits_uop_robIdx_flag :
    _GEN_302; // @[MemBlock.scala 521:35 524:20]
  assign io_writeback_2_bits_uop_robIdx_value = atomicsUnit_io_out_valid ? atomicsUnit_io_out_bits_uop_robIdx_value :
    _GEN_303; // @[MemBlock.scala 521:35 524:20]
  assign io_writeback_2_bits_debug_isMMIO = atomicsUnit_io_out_valid ? atomicsUnit_io_out_bits_debug_isMMIO : _GEN_397; // @[MemBlock.scala 521:35 524:20]
  assign io_writeback_2_bits_debug_vaddr = atomicsUnit_io_out_valid ? 39'h0 : _GEN_400; // @[MemBlock.scala 521:35 524:20]
  assign io_writeback_3_valid = StoreUnit_1_io_stout_valid; // @[MemBlock.scala 193:{41,41}]
  assign io_writeback_3_bits_uop_cf_exceptionVec_6 = StoreUnit_1_io_stout_bits_uop_cf_exceptionVec_6; // @[MemBlock.scala 193:{41,41}]
  assign io_writeback_3_bits_uop_cf_exceptionVec_7 = StoreUnit_1_io_stout_bits_uop_cf_exceptionVec_7; // @[MemBlock.scala 193:{41,41}]
  assign io_writeback_3_bits_uop_cf_exceptionVec_15 = StoreUnit_1_io_stout_bits_uop_cf_exceptionVec_15; // @[MemBlock.scala 193:{41,41}]
  assign io_writeback_3_bits_uop_cf_trigger_backendEn_0 = StoreUnit_1_io_stout_bits_uop_cf_trigger_backendEn_0; // @[MemBlock.scala 193:{41,41}]
  assign io_writeback_3_bits_uop_cf_trigger_backendHit_0 = io_writeback_3_valid & hit_3_0; // @[MemBlock.scala 193:16 489:26 498:68]
  assign io_writeback_3_bits_uop_cf_trigger_backendHit_1 = io_writeback_3_valid & hit_3_1; // @[MemBlock.scala 193:16 489:26 498:68]
  assign io_writeback_3_bits_uop_cf_trigger_backendHit_4 = io_writeback_3_valid & _GEN_204; // @[MemBlock.scala 193:16 489:26]
  assign io_writeback_3_bits_uop_robIdx_flag = StoreUnit_1_io_stout_bits_uop_robIdx_flag; // @[MemBlock.scala 193:{41,41}]
  assign io_writeback_3_bits_uop_robIdx_value = StoreUnit_1_io_stout_bits_uop_robIdx_value; // @[MemBlock.scala 193:{41,41}]
  assign io_writeback_3_bits_debug_isMMIO = StoreUnit_1_io_stout_bits_debug_isMMIO; // @[MemBlock.scala 193:{41,41}]
  assign io_writeback_3_bits_debug_vaddr = StoreUnit_1_io_stout_bits_debug_vaddr; // @[MemBlock.scala 193:{41,41}]
  assign io_writeback_4_valid = stdExeUnits_0_io_out_valid; // @[MemBlock.scala 193:{80,80}]
  assign io_writeback_4_bits_uop_robIdx_flag = stdExeUnits_0_io_out_bits_uop_robIdx_flag; // @[MemBlock.scala 193:{80,80}]
  assign io_writeback_4_bits_uop_robIdx_value = stdExeUnits_0_io_out_bits_uop_robIdx_value; // @[MemBlock.scala 193:{80,80}]
  assign io_writeback_5_valid = stdExeUnits_1_io_out_valid; // @[MemBlock.scala 193:{80,80}]
  assign io_writeback_5_bits_uop_robIdx_flag = stdExeUnits_1_io_out_bits_uop_robIdx_flag; // @[MemBlock.scala 193:{80,80}]
  assign io_writeback_5_bits_uop_robIdx_value = stdExeUnits_1_io_out_bits_uop_robIdx_value; // @[MemBlock.scala 193:{80,80}]
  assign io_stIn_0_valid = StoreUnit_0_io_issue_valid; // @[MemBlock.scala 481:22]
  assign io_stIn_0_bits_uop_cf_storeSetHit = StoreUnit_0_io_issue_bits_uop_cf_storeSetHit; // @[MemBlock.scala 482:21]
  assign io_stIn_0_bits_uop_cf_ssid = StoreUnit_0_io_issue_bits_uop_cf_ssid; // @[MemBlock.scala 482:21]
  assign io_stIn_0_bits_uop_robIdx_value = StoreUnit_0_io_issue_bits_uop_robIdx_value; // @[MemBlock.scala 482:21]
  assign io_stIn_1_valid = StoreUnit_1_io_issue_valid; // @[MemBlock.scala 481:22]
  assign io_stIn_1_bits_uop_cf_storeSetHit = StoreUnit_1_io_issue_bits_uop_cf_storeSetHit; // @[MemBlock.scala 482:21]
  assign io_stIn_1_bits_uop_cf_ssid = StoreUnit_1_io_issue_bits_uop_cf_ssid; // @[MemBlock.scala 482:21]
  assign io_stIn_1_bits_uop_robIdx_value = StoreUnit_1_io_issue_bits_uop_robIdx_value; // @[MemBlock.scala 482:21]
  assign io_memoryViolation_valid = lsq_io_rollback_valid; // @[MemBlock.scala 543:25]
  assign io_memoryViolation_bits_robIdx_flag = lsq_io_rollback_bits_robIdx_flag; // @[MemBlock.scala 543:25]
  assign io_memoryViolation_bits_robIdx_value = lsq_io_rollback_bits_robIdx_value; // @[MemBlock.scala 543:25]
  assign io_memoryViolation_bits_ftqIdx_flag = lsq_io_rollback_bits_ftqIdx_flag; // @[MemBlock.scala 543:25]
  assign io_memoryViolation_bits_ftqIdx_value = lsq_io_rollback_bits_ftqIdx_value; // @[MemBlock.scala 543:25]
  assign io_memoryViolation_bits_ftqOffset = lsq_io_rollback_bits_ftqOffset; // @[MemBlock.scala 543:25]
  assign io_memoryViolation_bits_stFtqIdx_value = lsq_io_rollback_bits_stFtqIdx_value; // @[MemBlock.scala 543:25]
  assign io_memoryViolation_bits_stFtqOffset = lsq_io_rollback_bits_stFtqOffset; // @[MemBlock.scala 543:25]
  assign io_ptw_req_0_valid = dtlb_ld_0_ptw_req_0_valid & ~(ptw_resp_v & vector_hit & _io_ptw_req_0_valid_T_7); // @[MemBlock.scala 291:38]
  assign io_ptw_req_0_bits_vpn = dtlb_ld_tlb_ld_io_ptw_req_0_bits_vpn; // @[MemBlock.scala 245:{24,24}]
  assign io_ptw_req_1_valid = dtlb_ld_0_ptw_req_1_valid & ~(ptw_resp_v & vector_hit & _io_ptw_req_1_valid_T_7); // @[MemBlock.scala 291:38]
  assign io_ptw_req_1_bits_vpn = dtlb_ld_tlb_ld_io_ptw_req_1_bits_vpn; // @[MemBlock.scala 245:{24,24}]
  assign io_ptw_req_2_valid = dtlb_st_0_ptw_req_0_valid & ~(ptw_resp_v & vector_hit_2 & _io_ptw_req_2_valid_T_7); // @[MemBlock.scala 291:38]
  assign io_ptw_req_2_bits_vpn = dtlb_st_tlb_st_io_ptw_req_0_bits_vpn; // @[MemBlock.scala 249:{24,24}]
  assign io_ptw_req_3_valid = dtlb_st_0_ptw_req_1_valid & ~(ptw_resp_v & vector_hit_2 & _io_ptw_req_3_valid_T_7); // @[MemBlock.scala 291:38]
  assign io_ptw_req_3_bits_vpn = dtlb_st_tlb_st_io_ptw_req_1_bits_vpn; // @[MemBlock.scala 249:{24,24}]
  assign io_fenceToSbuffer_sbIsEmpty = io_fenceToSbuffer_sbIsEmpty_REG; // @[MemBlock.scala 567:31]
  assign io_lsqio_exceptionAddr_vaddr = io_lsqio_exceptionAddr_vaddr_REG; // @[MemBlock.scala 668:32]
  assign io_lsqio_rob_isMMIO_0 = lsq_io_rob_isMMIO_0; // @[MemBlock.scala 539:25]
  assign io_lsqio_rob_isMMIO_1 = lsq_io_rob_isMMIO_1; // @[MemBlock.scala 539:25]
  assign io_lsqio_rob_uop_0_robIdx_value = lsq_io_rob_uop_0_robIdx_value; // @[MemBlock.scala 539:25]
  assign io_lsqio_rob_uop_1_robIdx_value = lsq_io_rob_uop_1_robIdx_value; // @[MemBlock.scala 539:25]
  assign io_csrUpdate_wvalid = io_csrUpdate_REG_wvalid; // @[MemBlock.scala 132:16]
  assign io_csrUpdate_waddr = io_csrUpdate_REG_waddr; // @[MemBlock.scala 132:16]
  assign io_csrUpdate_wdata = io_csrUpdate_REG_wdata; // @[MemBlock.scala 132:16]
  assign io_error_paddr = io_error_REG_1_paddr; // @[MemBlock.scala 133:12]
  assign io_error_report_to_beu = ~csrCtrl_delay_io_out_cache_error_enable ? 1'h0 : io_error_REG_1_report_to_beu; // @[MemBlock.scala 133:12 134:36 135:28]
  assign io_lqCancelCnt = lsq_io_lqCancelCnt; // @[MemBlock.scala 550:22]
  assign io_sqCancelCnt = lsq_io_sqCancelCnt; // @[MemBlock.scala 551:22]
  assign io_sqDeq = lsq_io_sqDeq; // @[MemBlock.scala 553:16]
  assign io_lqDeq = lsq_io_lqDeq; // @[MemBlock.scala 552:16]
  assign io_perf_0_value = io_perf_0_value_REG_1; // @[PerfCounterUtils.scala 188:17]
  assign io_perf_1_value = io_perf_1_value_REG_1; // @[PerfCounterUtils.scala 188:17]
  assign io_perf_2_value = io_perf_2_value_REG_1; // @[PerfCounterUtils.scala 188:17]
  assign io_perf_3_value = io_perf_3_value_REG_1; // @[PerfCounterUtils.scala 188:17]
  assign io_perf_4_value = io_perf_4_value_REG_1; // @[PerfCounterUtils.scala 188:17]
  assign io_perf_5_value = io_perf_5_value_REG_1; // @[PerfCounterUtils.scala 188:17]
  assign io_perf_6_value = io_perf_6_value_REG_1; // @[PerfCounterUtils.scala 188:17]
  assign io_perf_7_value = io_perf_7_value_REG_1; // @[PerfCounterUtils.scala 188:17]
  assign dcache_clock = clock;
  assign dcache_reset = reset;
  assign dcache_auto_client_out_a_ready = auto_dcache_client_out_a_ready; // @[LazyModule.scala 311:12]
  assign dcache_auto_client_out_bvalid = auto_dcache_client_out_bvalid; // @[LazyModule.scala 311:12]
  assign dcache_auto_client_out_bparam = auto_dcache_client_out_bparam; // @[LazyModule.scala 311:12]
  assign dcache_auto_client_out_baddress = auto_dcache_client_out_baddress; // @[LazyModule.scala 311:12]
  assign dcache_auto_client_out_bdata = auto_dcache_client_out_bdata; // @[LazyModule.scala 311:12]
  assign dcache_auto_client_out_c_ready = auto_dcache_client_out_c_ready; // @[LazyModule.scala 311:12]
  assign dcache_auto_client_out_d_valid = auto_dcache_client_out_d_valid; // @[LazyModule.scala 311:12]
  assign dcache_auto_client_out_d_bits_opcode = auto_dcache_client_out_d_bits_opcode; // @[LazyModule.scala 311:12]
  assign dcache_auto_client_out_d_bits_param = auto_dcache_client_out_d_bits_param; // @[LazyModule.scala 311:12]
  assign dcache_auto_client_out_d_bits_size = auto_dcache_client_out_d_bits_size; // @[LazyModule.scala 311:12]
  assign dcache_auto_client_out_d_bits_source = auto_dcache_client_out_d_bits_source; // @[LazyModule.scala 311:12]
  assign dcache_auto_client_out_d_bits_sink = auto_dcache_client_out_d_bits_sink; // @[LazyModule.scala 311:12]
  assign dcache_auto_client_out_d_bits_denied = auto_dcache_client_out_d_bits_denied; // @[LazyModule.scala 311:12]
  assign dcache_auto_client_out_d_bits_echo_blockisdirty = auto_dcache_client_out_d_bits_echo_blockisdirty; // @[LazyModule.scala 311:12]
  assign dcache_auto_client_out_d_bits_data = auto_dcache_client_out_d_bits_data; // @[LazyModule.scala 311:12]
  assign dcache_auto_client_out_d_bits_corrupt = auto_dcache_client_out_d_bits_corrupt; // @[LazyModule.scala 311:12]
  assign dcache_auto_client_out_e_ready = auto_dcache_client_out_e_ready; // @[LazyModule.scala 311:12]
  assign dcache_io_lsu_load_0_req_valid = LoadUnit_0_io_dcache_req_valid; // @[MemBlock.scala 348:28]
  assign dcache_io_lsu_load_0_req_bits_cmd = LoadUnit_0_io_dcache_req_bits_cmd; // @[MemBlock.scala 348:28]
  assign dcache_io_lsu_load_0_req_bits_addr = LoadUnit_0_io_dcache_req_bits_addr; // @[MemBlock.scala 348:28]
  assign dcache_io_lsu_load_0_req_bits_instrtype = LoadUnit_0_io_dcache_req_bits_instrtype; // @[MemBlock.scala 348:28]
  assign dcache_io_lsu_load_0_req_bits_replayCarry_real_way_en = LoadUnit_0_io_dcache_req_bits_replayCarry_real_way_en; // @[MemBlock.scala 348:28]
  assign dcache_io_lsu_load_0_req_bits_replayCarry_valid = LoadUnit_0_io_dcache_req_bits_replayCarry_valid; // @[MemBlock.scala 348:28]
  assign dcache_io_lsu_load_0_s1_kill = LoadUnit_0_io_dcache_s1_kill; // @[MemBlock.scala 348:28]
  assign dcache_io_lsu_load_0_s2_kill = LoadUnit_0_io_dcache_s2_kill; // @[MemBlock.scala 348:28]
  assign dcache_io_lsu_load_0_s1_paddr_dup_lsu = LoadUnit_0_io_dcache_s1_paddr_dup_lsu; // @[MemBlock.scala 348:28]
  assign dcache_io_lsu_load_0_s1_paddr_dup_dcache = LoadUnit_0_io_dcache_s1_paddr_dup_dcache; // @[MemBlock.scala 348:28]
  assign dcache_io_lsu_load_1_req_valid = LoadUnit_1_io_dcache_req_valid; // @[MemBlock.scala 348:28]
  assign dcache_io_lsu_load_1_req_bits_cmd = LoadUnit_1_io_dcache_req_bits_cmd; // @[MemBlock.scala 348:28]
  assign dcache_io_lsu_load_1_req_bits_addr = LoadUnit_1_io_dcache_req_bits_addr; // @[MemBlock.scala 348:28]
  assign dcache_io_lsu_load_1_req_bits_instrtype = LoadUnit_1_io_dcache_req_bits_instrtype; // @[MemBlock.scala 348:28]
  assign dcache_io_lsu_load_1_req_bits_replayCarry_real_way_en = LoadUnit_1_io_dcache_req_bits_replayCarry_real_way_en; // @[MemBlock.scala 348:28]
  assign dcache_io_lsu_load_1_req_bits_replayCarry_valid = LoadUnit_1_io_dcache_req_bits_replayCarry_valid; // @[MemBlock.scala 348:28]
  assign dcache_io_lsu_load_1_s1_kill = LoadUnit_1_io_dcache_s1_kill; // @[MemBlock.scala 348:28]
  assign dcache_io_lsu_load_1_s2_kill = LoadUnit_1_io_dcache_s2_kill; // @[MemBlock.scala 348:28]
  assign dcache_io_lsu_load_1_s1_paddr_dup_lsu = LoadUnit_1_io_dcache_s1_paddr_dup_lsu; // @[MemBlock.scala 348:28]
  assign dcache_io_lsu_load_1_s1_paddr_dup_dcache = LoadUnit_1_io_dcache_s1_paddr_dup_dcache; // @[MemBlock.scala 348:28]
  assign dcache_io_lsu_store_req_valid = sbuffer_io_dcache_req_valid; // @[MemBlock.scala 561:25]
  assign dcache_io_lsu_store_req_bits_vaddr = sbuffer_io_dcache_req_bits_vaddr; // @[MemBlock.scala 561:25]
  assign dcache_io_lsu_store_req_bits_addr = sbuffer_io_dcache_req_bits_addr; // @[MemBlock.scala 561:25]
  assign dcache_io_lsu_store_req_bits_data = sbuffer_io_dcache_req_bits_data; // @[MemBlock.scala 561:25]
  assign dcache_io_lsu_store_req_bits_mask = sbuffer_io_dcache_req_bits_mask; // @[MemBlock.scala 561:25]
  assign dcache_io_lsu_store_req_bits_id = sbuffer_io_dcache_req_bits_id; // @[MemBlock.scala 561:25]
  assign dcache_io_lsu_atomics_req_valid = atomicsUnit_io_dcache_req_valid; // @[MemBlock.scala 632:25]
  assign dcache_io_lsu_atomics_req_bits_cmd = atomicsUnit_io_dcache_req_bits_cmd; // @[MemBlock.scala 632:25]
  assign dcache_io_lsu_atomics_req_bits_vaddr = atomicsUnit_io_dcache_req_bits_vaddr; // @[MemBlock.scala 632:25]
  assign dcache_io_lsu_atomics_req_bits_addr = atomicsUnit_io_dcache_req_bits_addr; // @[MemBlock.scala 632:25]
  assign dcache_io_lsu_atomics_req_bits_word_idx = atomicsUnit_io_dcache_req_bits_word_idx; // @[MemBlock.scala 632:25]
  assign dcache_io_lsu_atomics_req_bits_amo_data = atomicsUnit_io_dcache_req_bits_amo_data; // @[MemBlock.scala 632:25]
  assign dcache_io_lsu_atomics_req_bits_amo_mask = atomicsUnit_io_dcache_req_bits_amo_mask; // @[MemBlock.scala 632:25]
  assign dcache_io_lsu_forward_mshr_0_valid = LoadUnit_0_io_forward_mshr_valid; // @[MemBlock.scala 355:34]
  assign dcache_io_lsu_forward_mshr_0_mshrid = LoadUnit_0_io_forward_mshr_mshrid; // @[MemBlock.scala 355:34]
  assign dcache_io_lsu_forward_mshr_0_paddr = LoadUnit_0_io_forward_mshr_paddr; // @[MemBlock.scala 355:34]
  assign dcache_io_lsu_forward_mshr_1_valid = LoadUnit_1_io_forward_mshr_valid; // @[MemBlock.scala 355:34]
  assign dcache_io_lsu_forward_mshr_1_mshrid = LoadUnit_1_io_forward_mshr_mshrid; // @[MemBlock.scala 355:34]
  assign dcache_io_lsu_forward_mshr_1_paddr = LoadUnit_1_io_forward_mshr_paddr; // @[MemBlock.scala 355:34]
  assign dcache_io_csr_distribute_csr_wvalid = csrCtrl_delay_io_out_distribute_csr_wvalid; // @[MemBlock.scala 130:32]
  assign dcache_io_csr_distribute_csr_waddr = csrCtrl_delay_io_out_distribute_csr_waddr; // @[MemBlock.scala 130:32]
  assign dcache_io_csr_distribute_csr_wdata = csrCtrl_delay_io_out_distribute_csr_wdata; // @[MemBlock.scala 130:32]
  assign uncache_clock = clock;
  assign uncache_reset = reset;
  assign uncache_auto_client_out_a_ready = auto_uncache_client_out_a_ready; // @[LazyModule.scala 311:12]
  assign uncache_auto_client_out_d_valid = auto_uncache_client_out_d_valid; // @[LazyModule.scala 311:12]
  assign uncache_auto_client_out_d_bits_opcode = auto_uncache_client_out_d_bits_opcode; // @[LazyModule.scala 311:12]
  assign uncache_auto_client_out_d_bits_data = auto_uncache_client_out_d_bits_data; // @[LazyModule.scala 311:12]
  assign uncache_io_hartId = io_hartId; // @[MemBlock.scala 535:21]
  assign uncache_io_enableOutstanding = io_csrCtrl_uncache_write_outstanding_enable; // @[MemBlock.scala 534:32]
  assign uncache_io_lsq_req_valid = pipelineReg_io_out_valid; // @[MemCommon.scala 399:11]
  assign uncache_io_lsq_req_bits_cmd = pipelineReg_io_out_bits_cmd; // @[MemCommon.scala 399:11]
  assign uncache_io_lsq_req_bits_addr = pipelineReg_io_out_bits_addr; // @[MemCommon.scala 399:11]
  assign uncache_io_lsq_req_bits_data = pipelineReg_io_out_bits_data; // @[MemCommon.scala 399:11]
  assign uncache_io_lsq_req_bits_mask = pipelineReg_io_out_bits_mask; // @[MemCommon.scala 399:11]
  assign uncache_io_lsq_req_bits_atomic = pipelineReg_io_out_bits_atomic; // @[MemCommon.scala 399:11]
  assign csrCtrl_delay_clock = clock;
  assign csrCtrl_delay_io_in_icache_parity_enable = io_csrCtrl_icache_parity_enable; // @[Hold.scala 98:17]
  assign csrCtrl_delay_io_in_lvpred_disable = io_csrCtrl_lvpred_disable; // @[Hold.scala 98:17]
  assign csrCtrl_delay_io_in_no_spec_load = io_csrCtrl_no_spec_load; // @[Hold.scala 98:17]
  assign csrCtrl_delay_io_in_storeset_wait_store = io_csrCtrl_storeset_wait_store; // @[Hold.scala 98:17]
  assign csrCtrl_delay_io_in_lvpred_timeout = io_csrCtrl_lvpred_timeout; // @[Hold.scala 98:17]
  assign csrCtrl_delay_io_in_bp_ctrl_ubtb_enable = io_csrCtrl_bp_ctrl_ubtb_enable; // @[Hold.scala 98:17]
  assign csrCtrl_delay_io_in_bp_ctrl_btb_enable = io_csrCtrl_bp_ctrl_btb_enable; // @[Hold.scala 98:17]
  assign csrCtrl_delay_io_in_bp_ctrl_tage_enable = io_csrCtrl_bp_ctrl_tage_enable; // @[Hold.scala 98:17]
  assign csrCtrl_delay_io_in_bp_ctrl_sc_enable = io_csrCtrl_bp_ctrl_sc_enable; // @[Hold.scala 98:17]
  assign csrCtrl_delay_io_in_bp_ctrl_ras_enable = io_csrCtrl_bp_ctrl_ras_enable; // @[Hold.scala 98:17]
  assign csrCtrl_delay_io_in_sbuffer_threshold = io_csrCtrl_sbuffer_threshold; // @[Hold.scala 98:17]
  assign csrCtrl_delay_io_in_ldld_vio_check_enable = io_csrCtrl_ldld_vio_check_enable; // @[Hold.scala 98:17]
  assign csrCtrl_delay_io_in_cache_error_enable = io_csrCtrl_cache_error_enable; // @[Hold.scala 98:17]
  assign csrCtrl_delay_io_in_uncache_write_outstanding_enable = io_csrCtrl_uncache_write_outstanding_enable; // @[Hold.scala 98:17]
  assign csrCtrl_delay_io_in_fusion_enable = io_csrCtrl_fusion_enable; // @[Hold.scala 98:17]
  assign csrCtrl_delay_io_in_wfi_enable = io_csrCtrl_wfi_enable; // @[Hold.scala 98:17]
  assign csrCtrl_delay_io_in_svinval_enable = io_csrCtrl_svinval_enable; // @[Hold.scala 98:17]
  assign csrCtrl_delay_io_in_distribute_csr_wvalid = io_csrCtrl_distribute_csr_wvalid; // @[Hold.scala 98:17]
  assign csrCtrl_delay_io_in_distribute_csr_waddr = io_csrCtrl_distribute_csr_waddr; // @[Hold.scala 98:17]
  assign csrCtrl_delay_io_in_distribute_csr_wdata = io_csrCtrl_distribute_csr_wdata; // @[Hold.scala 98:17]
  assign csrCtrl_delay_io_in_singlestep = io_csrCtrl_singlestep; // @[Hold.scala 98:17]
  assign csrCtrl_delay_io_in_frontend_trigger_t_valid = io_csrCtrl_frontend_trigger_t_valid; // @[Hold.scala 98:17]
  assign csrCtrl_delay_io_in_frontend_trigger_t_bits_addr = io_csrCtrl_frontend_trigger_t_bits_addr; // @[Hold.scala 98:17]
  assign csrCtrl_delay_io_in_frontend_trigger_t_bits_tdata_matchType =
    io_csrCtrl_frontend_trigger_t_bits_tdata_matchType; // @[Hold.scala 98:17]
  assign csrCtrl_delay_io_in_frontend_trigger_t_bits_tdata_select = io_csrCtrl_frontend_trigger_t_bits_tdata_select; // @[Hold.scala 98:17]
  assign csrCtrl_delay_io_in_frontend_trigger_t_bits_tdata_timing = io_csrCtrl_frontend_trigger_t_bits_tdata_timing; // @[Hold.scala 98:17]
  assign csrCtrl_delay_io_in_frontend_trigger_t_bits_tdata_chain = io_csrCtrl_frontend_trigger_t_bits_tdata_chain; // @[Hold.scala 98:17]
  assign csrCtrl_delay_io_in_frontend_trigger_t_bits_tdata_tdata2 = io_csrCtrl_frontend_trigger_t_bits_tdata_tdata2; // @[Hold.scala 98:17]
  assign csrCtrl_delay_io_in_mem_trigger_t_valid = io_csrCtrl_mem_trigger_t_valid; // @[Hold.scala 98:17]
  assign csrCtrl_delay_io_in_mem_trigger_t_bits_addr = io_csrCtrl_mem_trigger_t_bits_addr; // @[Hold.scala 98:17]
  assign csrCtrl_delay_io_in_mem_trigger_t_bits_tdata_matchType = io_csrCtrl_mem_trigger_t_bits_tdata_matchType; // @[Hold.scala 98:17]
  assign csrCtrl_delay_io_in_mem_trigger_t_bits_tdata_select = io_csrCtrl_mem_trigger_t_bits_tdata_select; // @[Hold.scala 98:17]
  assign csrCtrl_delay_io_in_mem_trigger_t_bits_tdata_chain = io_csrCtrl_mem_trigger_t_bits_tdata_chain; // @[Hold.scala 98:17]
  assign csrCtrl_delay_io_in_mem_trigger_t_bits_tdata_tdata2 = io_csrCtrl_mem_trigger_t_bits_tdata_tdata2; // @[Hold.scala 98:17]
  assign csrCtrl_delay_io_in_trigger_enable_0 = io_csrCtrl_trigger_enable_0; // @[Hold.scala 98:17]
  assign csrCtrl_delay_io_in_trigger_enable_1 = io_csrCtrl_trigger_enable_1; // @[Hold.scala 98:17]
  assign csrCtrl_delay_io_in_trigger_enable_2 = io_csrCtrl_trigger_enable_2; // @[Hold.scala 98:17]
  assign csrCtrl_delay_io_in_trigger_enable_3 = io_csrCtrl_trigger_enable_3; // @[Hold.scala 98:17]
  assign csrCtrl_delay_io_in_trigger_enable_4 = io_csrCtrl_trigger_enable_4; // @[Hold.scala 98:17]
  assign csrCtrl_delay_io_in_trigger_enable_5 = io_csrCtrl_trigger_enable_5; // @[Hold.scala 98:17]
  assign csrCtrl_delay_io_in_trigger_enable_6 = io_csrCtrl_trigger_enable_6; // @[Hold.scala 98:17]
  assign csrCtrl_delay_io_in_trigger_enable_7 = io_csrCtrl_trigger_enable_7; // @[Hold.scala 98:17]
  assign csrCtrl_delay_io_in_trigger_enable_8 = io_csrCtrl_trigger_enable_8; // @[Hold.scala 98:17]
  assign csrCtrl_delay_io_in_trigger_enable_9 = io_csrCtrl_trigger_enable_9; // @[Hold.scala 98:17]
  assign LoadUnit_0_clock = clock;
  assign LoadUnit_0_reset = reset;
  assign LoadUnit_0_io_loadIn_valid = io_issue_0_valid; // @[MemBlock.scala 344:28]
  assign LoadUnit_0_io_loadIn_bits_uop_cf_foldpc = io_issue_0_bits_uop_cf_foldpc; // @[MemBlock.scala 344:28]
  assign LoadUnit_0_io_loadIn_bits_uop_cf_trigger_backendEn_1 = io_issue_0_bits_uop_cf_trigger_backendEn_1; // @[MemBlock.scala 344:28]
  assign LoadUnit_0_io_loadIn_bits_uop_cf_waitForRobIdx_flag = io_issue_0_bits_uop_cf_waitForRobIdx_flag; // @[MemBlock.scala 344:28]
  assign LoadUnit_0_io_loadIn_bits_uop_cf_waitForRobIdx_value = io_issue_0_bits_uop_cf_waitForRobIdx_value; // @[MemBlock.scala 344:28]
  assign LoadUnit_0_io_loadIn_bits_uop_cf_loadWaitBit = io_issue_0_bits_uop_cf_loadWaitBit; // @[MemBlock.scala 344:28]
  assign LoadUnit_0_io_loadIn_bits_uop_cf_loadWaitStrict = io_issue_0_bits_uop_cf_loadWaitStrict; // @[MemBlock.scala 344:28]
  assign LoadUnit_0_io_loadIn_bits_uop_cf_ftqPtr_flag = io_issue_0_bits_uop_cf_ftqPtr_flag; // @[MemBlock.scala 344:28]
  assign LoadUnit_0_io_loadIn_bits_uop_cf_ftqPtr_value = io_issue_0_bits_uop_cf_ftqPtr_value; // @[MemBlock.scala 344:28]
  assign LoadUnit_0_io_loadIn_bits_uop_cf_ftqOffset = io_issue_0_bits_uop_cf_ftqOffset; // @[MemBlock.scala 344:28]
  assign LoadUnit_0_io_loadIn_bits_uop_ctrl_fuType = io_issue_0_bits_uop_ctrl_fuType; // @[MemBlock.scala 344:28]
  assign LoadUnit_0_io_loadIn_bits_uop_ctrl_fuOpType = io_issue_0_bits_uop_ctrl_fuOpType; // @[MemBlock.scala 344:28]
  assign LoadUnit_0_io_loadIn_bits_uop_ctrl_rfWen = io_issue_0_bits_uop_ctrl_rfWen; // @[MemBlock.scala 344:28]
  assign LoadUnit_0_io_loadIn_bits_uop_ctrl_fpWen = io_issue_0_bits_uop_ctrl_fpWen; // @[MemBlock.scala 344:28]
  assign LoadUnit_0_io_loadIn_bits_uop_ctrl_imm = io_issue_0_bits_uop_ctrl_imm; // @[MemBlock.scala 344:28]
  assign LoadUnit_0_io_loadIn_bits_uop_pdest = io_issue_0_bits_uop_pdest; // @[MemBlock.scala 344:28]
  assign LoadUnit_0_io_loadIn_bits_uop_robIdx_flag = io_issue_0_bits_uop_robIdx_flag; // @[MemBlock.scala 344:28]
  assign LoadUnit_0_io_loadIn_bits_uop_robIdx_value = io_issue_0_bits_uop_robIdx_value; // @[MemBlock.scala 344:28]
  assign LoadUnit_0_io_loadIn_bits_uop_lqIdx_flag = io_issue_0_bits_uop_lqIdx_flag; // @[MemBlock.scala 344:28]
  assign LoadUnit_0_io_loadIn_bits_uop_lqIdx_value = io_issue_0_bits_uop_lqIdx_value; // @[MemBlock.scala 344:28]
  assign LoadUnit_0_io_loadIn_bits_uop_sqIdx_flag = io_issue_0_bits_uop_sqIdx_flag; // @[MemBlock.scala 344:28]
  assign LoadUnit_0_io_loadIn_bits_uop_sqIdx_value = io_issue_0_bits_uop_sqIdx_value; // @[MemBlock.scala 344:28]
  assign LoadUnit_0_io_loadIn_bits_src_0 = io_issue_0_bits_src_0; // @[MemBlock.scala 344:28]
  assign LoadUnit_0_io_VecloadIn_valid = vlflowqueue_io_loadPipeOut_0_valid; // @[MemBlock.scala 346:31]
  assign LoadUnit_0_io_VecloadIn_bits_vaddr = vlflowqueue_io_loadPipeOut_0_bits_vaddr; // @[MemBlock.scala 346:31]
  assign LoadUnit_0_io_redirect_valid = redirect_next_valid_REG; // @[BitUtils.scala 26:20 28:18]
  assign LoadUnit_0_io_redirect_bits_robIdx_flag = redirect_next_bits_rrobIdx_flag; // @[BitUtils.scala 26:20 33:15]
  assign LoadUnit_0_io_redirect_bits_robIdx_value = redirect_next_bits_rrobIdx_value; // @[BitUtils.scala 26:20 33:15]
  assign LoadUnit_0_io_redirect_bits_level = redirect_next_bits_rlevel; // @[BitUtils.scala 26:20 33:15]
  assign LoadUnit_0_io_dcache_req_ready = dcache_io_lsu_load_0_req_ready; // @[MemBlock.scala 348:28]
  assign LoadUnit_0_io_dcache_resp_bits_data_delayed = dcache_io_lsu_load_0_resp_bits_data_delayed; // @[MemBlock.scala 348:28]
  assign LoadUnit_0_io_dcache_resp_bits_miss = dcache_io_lsu_load_0_resp_bits_miss; // @[MemBlock.scala 348:28]
  assign LoadUnit_0_io_dcache_resp_bits_replay = dcache_io_lsu_load_0_resp_bits_replay; // @[MemBlock.scala 348:28]
  assign LoadUnit_0_io_dcache_resp_bits_replayCarry_real_way_en = dcache_io_lsu_load_0_resp_bits_replayCarry_real_way_en
    ; // @[MemBlock.scala 348:28]
  assign LoadUnit_0_io_dcache_resp_bits_replayCarry_valid = dcache_io_lsu_load_0_resp_bits_replayCarry_valid; // @[MemBlock.scala 348:28]
  assign LoadUnit_0_io_dcache_resp_bits_tag_error = dcache_io_lsu_load_0_resp_bits_tag_error; // @[MemBlock.scala 348:28]
  assign LoadUnit_0_io_dcache_resp_bits_mshr_id = dcache_io_lsu_load_0_resp_bits_mshr_id; // @[MemBlock.scala 348:28]
  assign LoadUnit_0_io_dcache_resp_bits_error_delayed = dcache_io_lsu_load_0_resp_bits_error_delayed; // @[MemBlock.scala 348:28]
  assign LoadUnit_0_io_dcache_s1_bank_conflict = dcache_io_lsu_load_0_s1_bank_conflict; // @[MemBlock.scala 348:28]
  assign LoadUnit_0_io_sbuffer_forwardMask_0 = sbuffer_io_forward_0_forwardMask_0; // @[MemBlock.scala 351:29]
  assign LoadUnit_0_io_sbuffer_forwardMask_1 = sbuffer_io_forward_0_forwardMask_1; // @[MemBlock.scala 351:29]
  assign LoadUnit_0_io_sbuffer_forwardMask_2 = sbuffer_io_forward_0_forwardMask_2; // @[MemBlock.scala 351:29]
  assign LoadUnit_0_io_sbuffer_forwardMask_3 = sbuffer_io_forward_0_forwardMask_3; // @[MemBlock.scala 351:29]
  assign LoadUnit_0_io_sbuffer_forwardMask_4 = sbuffer_io_forward_0_forwardMask_4; // @[MemBlock.scala 351:29]
  assign LoadUnit_0_io_sbuffer_forwardMask_5 = sbuffer_io_forward_0_forwardMask_5; // @[MemBlock.scala 351:29]
  assign LoadUnit_0_io_sbuffer_forwardMask_6 = sbuffer_io_forward_0_forwardMask_6; // @[MemBlock.scala 351:29]
  assign LoadUnit_0_io_sbuffer_forwardMask_7 = sbuffer_io_forward_0_forwardMask_7; // @[MemBlock.scala 351:29]
  assign LoadUnit_0_io_sbuffer_forwardMask_8 = sbuffer_io_forward_0_forwardMask_8; // @[MemBlock.scala 351:29]
  assign LoadUnit_0_io_sbuffer_forwardMask_9 = sbuffer_io_forward_0_forwardMask_9; // @[MemBlock.scala 351:29]
  assign LoadUnit_0_io_sbuffer_forwardMask_10 = sbuffer_io_forward_0_forwardMask_10; // @[MemBlock.scala 351:29]
  assign LoadUnit_0_io_sbuffer_forwardMask_11 = sbuffer_io_forward_0_forwardMask_11; // @[MemBlock.scala 351:29]
  assign LoadUnit_0_io_sbuffer_forwardMask_12 = sbuffer_io_forward_0_forwardMask_12; // @[MemBlock.scala 351:29]
  assign LoadUnit_0_io_sbuffer_forwardMask_13 = sbuffer_io_forward_0_forwardMask_13; // @[MemBlock.scala 351:29]
  assign LoadUnit_0_io_sbuffer_forwardMask_14 = sbuffer_io_forward_0_forwardMask_14; // @[MemBlock.scala 351:29]
  assign LoadUnit_0_io_sbuffer_forwardMask_15 = sbuffer_io_forward_0_forwardMask_15; // @[MemBlock.scala 351:29]
  assign LoadUnit_0_io_sbuffer_forwardData_0 = sbuffer_io_forward_0_forwardData_0; // @[MemBlock.scala 351:29]
  assign LoadUnit_0_io_sbuffer_forwardData_1 = sbuffer_io_forward_0_forwardData_1; // @[MemBlock.scala 351:29]
  assign LoadUnit_0_io_sbuffer_forwardData_2 = sbuffer_io_forward_0_forwardData_2; // @[MemBlock.scala 351:29]
  assign LoadUnit_0_io_sbuffer_forwardData_3 = sbuffer_io_forward_0_forwardData_3; // @[MemBlock.scala 351:29]
  assign LoadUnit_0_io_sbuffer_forwardData_4 = sbuffer_io_forward_0_forwardData_4; // @[MemBlock.scala 351:29]
  assign LoadUnit_0_io_sbuffer_forwardData_5 = sbuffer_io_forward_0_forwardData_5; // @[MemBlock.scala 351:29]
  assign LoadUnit_0_io_sbuffer_forwardData_6 = sbuffer_io_forward_0_forwardData_6; // @[MemBlock.scala 351:29]
  assign LoadUnit_0_io_sbuffer_forwardData_7 = sbuffer_io_forward_0_forwardData_7; // @[MemBlock.scala 351:29]
  assign LoadUnit_0_io_sbuffer_forwardData_8 = sbuffer_io_forward_0_forwardData_8; // @[MemBlock.scala 351:29]
  assign LoadUnit_0_io_sbuffer_forwardData_9 = sbuffer_io_forward_0_forwardData_9; // @[MemBlock.scala 351:29]
  assign LoadUnit_0_io_sbuffer_forwardData_10 = sbuffer_io_forward_0_forwardData_10; // @[MemBlock.scala 351:29]
  assign LoadUnit_0_io_sbuffer_forwardData_11 = sbuffer_io_forward_0_forwardData_11; // @[MemBlock.scala 351:29]
  assign LoadUnit_0_io_sbuffer_forwardData_12 = sbuffer_io_forward_0_forwardData_12; // @[MemBlock.scala 351:29]
  assign LoadUnit_0_io_sbuffer_forwardData_13 = sbuffer_io_forward_0_forwardData_13; // @[MemBlock.scala 351:29]
  assign LoadUnit_0_io_sbuffer_forwardData_14 = sbuffer_io_forward_0_forwardData_14; // @[MemBlock.scala 351:29]
  assign LoadUnit_0_io_sbuffer_forwardData_15 = sbuffer_io_forward_0_forwardData_15; // @[MemBlock.scala 351:29]
  assign LoadUnit_0_io_sbuffer_matchInvalid = sbuffer_io_forward_0_matchInvalid; // @[MemBlock.scala 351:29]
  assign LoadUnit_0_io_lsq_loadOut_valid = lsq_io_loadOut_0_valid; // @[MemBlock.scala 400:23]
  assign LoadUnit_0_io_lsq_loadOut_bits_uop_cf_exceptionVec_4 = lsq_io_loadOut_0_bits_uop_cf_exceptionVec_4; // @[MemBlock.scala 400:23]
  assign LoadUnit_0_io_lsq_loadOut_bits_uop_cf_exceptionVec_5 = lsq_io_loadOut_0_bits_uop_cf_exceptionVec_5; // @[MemBlock.scala 400:23]
  assign LoadUnit_0_io_lsq_loadOut_bits_uop_cf_exceptionVec_13 = lsq_io_loadOut_0_bits_uop_cf_exceptionVec_13; // @[MemBlock.scala 400:23]
  assign LoadUnit_0_io_lsq_loadOut_bits_uop_cf_trigger_backendEn_1 = lsq_io_loadOut_0_bits_uop_cf_trigger_backendEn_1; // @[MemBlock.scala 400:23]
  assign LoadUnit_0_io_lsq_loadOut_bits_uop_cf_trigger_backendHit_0 = lsq_io_loadOut_0_bits_uop_cf_trigger_backendHit_0; // @[MemBlock.scala 400:23]
  assign LoadUnit_0_io_lsq_loadOut_bits_uop_cf_trigger_backendHit_1 = lsq_io_loadOut_0_bits_uop_cf_trigger_backendHit_1; // @[MemBlock.scala 400:23]
  assign LoadUnit_0_io_lsq_loadOut_bits_uop_cf_trigger_backendHit_4 = lsq_io_loadOut_0_bits_uop_cf_trigger_backendHit_4; // @[MemBlock.scala 400:23]
  assign LoadUnit_0_io_lsq_loadOut_bits_uop_ctrl_rfWen = lsq_io_loadOut_0_bits_uop_ctrl_rfWen; // @[MemBlock.scala 400:23]
  assign LoadUnit_0_io_lsq_loadOut_bits_uop_ctrl_fpWen = lsq_io_loadOut_0_bits_uop_ctrl_fpWen; // @[MemBlock.scala 400:23]
  assign LoadUnit_0_io_lsq_loadOut_bits_uop_ctrl_flushPipe = lsq_io_loadOut_0_bits_uop_ctrl_flushPipe; // @[MemBlock.scala 400:23]
  assign LoadUnit_0_io_lsq_loadOut_bits_uop_ctrl_replayInst = lsq_io_loadOut_0_bits_uop_ctrl_replayInst; // @[MemBlock.scala 400:23]
  assign LoadUnit_0_io_lsq_loadOut_bits_uop_pdest = lsq_io_loadOut_0_bits_uop_pdest; // @[MemBlock.scala 400:23]
  assign LoadUnit_0_io_lsq_loadOut_bits_uop_robIdx_flag = lsq_io_loadOut_0_bits_uop_robIdx_flag; // @[MemBlock.scala 400:23]
  assign LoadUnit_0_io_lsq_loadOut_bits_uop_robIdx_value = lsq_io_loadOut_0_bits_uop_robIdx_value; // @[MemBlock.scala 400:23]
  assign LoadUnit_0_io_lsq_loadOut_bits_debug_isMMIO = 1'h1; // @[MemBlock.scala 400:23]
  assign LoadUnit_0_io_lsq_ldRawData_lqData = lsq_io_ldRawDataOut_0_lqData; // @[MemBlock.scala 401:28]
  assign LoadUnit_0_io_lsq_ldRawData_uop_ctrl_fuOpType = lsq_io_ldRawDataOut_0_uop_ctrl_fuOpType; // @[MemBlock.scala 401:28]
  assign LoadUnit_0_io_lsq_ldRawData_uop_ctrl_fpWen = lsq_io_ldRawDataOut_0_uop_ctrl_fpWen; // @[MemBlock.scala 401:28]
  assign LoadUnit_0_io_lsq_ldRawData_addrOffset = lsq_io_ldRawDataOut_0_addrOffset; // @[MemBlock.scala 401:28]
  assign LoadUnit_0_io_lsq_forward_forwardMask_0 = lsq_io_forward_0_forwardMask_0; // @[MemBlock.scala 350:33]
  assign LoadUnit_0_io_lsq_forward_forwardMask_1 = lsq_io_forward_0_forwardMask_1; // @[MemBlock.scala 350:33]
  assign LoadUnit_0_io_lsq_forward_forwardMask_2 = lsq_io_forward_0_forwardMask_2; // @[MemBlock.scala 350:33]
  assign LoadUnit_0_io_lsq_forward_forwardMask_3 = lsq_io_forward_0_forwardMask_3; // @[MemBlock.scala 350:33]
  assign LoadUnit_0_io_lsq_forward_forwardMask_4 = lsq_io_forward_0_forwardMask_4; // @[MemBlock.scala 350:33]
  assign LoadUnit_0_io_lsq_forward_forwardMask_5 = lsq_io_forward_0_forwardMask_5; // @[MemBlock.scala 350:33]
  assign LoadUnit_0_io_lsq_forward_forwardMask_6 = lsq_io_forward_0_forwardMask_6; // @[MemBlock.scala 350:33]
  assign LoadUnit_0_io_lsq_forward_forwardMask_7 = lsq_io_forward_0_forwardMask_7; // @[MemBlock.scala 350:33]
  assign LoadUnit_0_io_lsq_forward_forwardMask_8 = lsq_io_forward_0_forwardMask_8; // @[MemBlock.scala 350:33]
  assign LoadUnit_0_io_lsq_forward_forwardMask_9 = lsq_io_forward_0_forwardMask_9; // @[MemBlock.scala 350:33]
  assign LoadUnit_0_io_lsq_forward_forwardMask_10 = lsq_io_forward_0_forwardMask_10; // @[MemBlock.scala 350:33]
  assign LoadUnit_0_io_lsq_forward_forwardMask_11 = lsq_io_forward_0_forwardMask_11; // @[MemBlock.scala 350:33]
  assign LoadUnit_0_io_lsq_forward_forwardMask_12 = lsq_io_forward_0_forwardMask_12; // @[MemBlock.scala 350:33]
  assign LoadUnit_0_io_lsq_forward_forwardMask_13 = lsq_io_forward_0_forwardMask_13; // @[MemBlock.scala 350:33]
  assign LoadUnit_0_io_lsq_forward_forwardMask_14 = lsq_io_forward_0_forwardMask_14; // @[MemBlock.scala 350:33]
  assign LoadUnit_0_io_lsq_forward_forwardMask_15 = lsq_io_forward_0_forwardMask_15; // @[MemBlock.scala 350:33]
  assign LoadUnit_0_io_lsq_forward_forwardData_0 = lsq_io_forward_0_forwardData_0; // @[MemBlock.scala 350:33]
  assign LoadUnit_0_io_lsq_forward_forwardData_1 = lsq_io_forward_0_forwardData_1; // @[MemBlock.scala 350:33]
  assign LoadUnit_0_io_lsq_forward_forwardData_2 = lsq_io_forward_0_forwardData_2; // @[MemBlock.scala 350:33]
  assign LoadUnit_0_io_lsq_forward_forwardData_3 = lsq_io_forward_0_forwardData_3; // @[MemBlock.scala 350:33]
  assign LoadUnit_0_io_lsq_forward_forwardData_4 = lsq_io_forward_0_forwardData_4; // @[MemBlock.scala 350:33]
  assign LoadUnit_0_io_lsq_forward_forwardData_5 = lsq_io_forward_0_forwardData_5; // @[MemBlock.scala 350:33]
  assign LoadUnit_0_io_lsq_forward_forwardData_6 = lsq_io_forward_0_forwardData_6; // @[MemBlock.scala 350:33]
  assign LoadUnit_0_io_lsq_forward_forwardData_7 = lsq_io_forward_0_forwardData_7; // @[MemBlock.scala 350:33]
  assign LoadUnit_0_io_lsq_forward_forwardData_8 = lsq_io_forward_0_forwardData_8; // @[MemBlock.scala 350:33]
  assign LoadUnit_0_io_lsq_forward_forwardData_9 = lsq_io_forward_0_forwardData_9; // @[MemBlock.scala 350:33]
  assign LoadUnit_0_io_lsq_forward_forwardData_10 = lsq_io_forward_0_forwardData_10; // @[MemBlock.scala 350:33]
  assign LoadUnit_0_io_lsq_forward_forwardData_11 = lsq_io_forward_0_forwardData_11; // @[MemBlock.scala 350:33]
  assign LoadUnit_0_io_lsq_forward_forwardData_12 = lsq_io_forward_0_forwardData_12; // @[MemBlock.scala 350:33]
  assign LoadUnit_0_io_lsq_forward_forwardData_13 = lsq_io_forward_0_forwardData_13; // @[MemBlock.scala 350:33]
  assign LoadUnit_0_io_lsq_forward_forwardData_14 = lsq_io_forward_0_forwardData_14; // @[MemBlock.scala 350:33]
  assign LoadUnit_0_io_lsq_forward_forwardData_15 = lsq_io_forward_0_forwardData_15; // @[MemBlock.scala 350:33]
  assign LoadUnit_0_io_lsq_forward_dataInvalid = lsq_io_forward_0_dataInvalid; // @[MemBlock.scala 350:33]
  assign LoadUnit_0_io_lsq_forward_matchInvalid = lsq_io_forward_0_matchInvalid; // @[MemBlock.scala 350:33]
  assign LoadUnit_0_io_lsq_forward_schedWait = lsq_io_forward_0_schedWait; // @[MemBlock.scala 350:33]
  assign LoadUnit_0_io_lsq_forward_dataInvalidSqIdx_flag = lsq_io_forward_0_dataInvalidSqIdx_flag; // @[MemBlock.scala 350:33]
  assign LoadUnit_0_io_lsq_forward_dataInvalidSqIdx_value = lsq_io_forward_0_dataInvalidSqIdx_value; // @[MemBlock.scala 350:33]
  assign LoadUnit_0_io_lsq_forward_addrInvalidSqIdx_flag = lsq_io_forward_0_addrInvalidSqIdx_flag; // @[MemBlock.scala 350:33]
  assign LoadUnit_0_io_lsq_forward_addrInvalidSqIdx_value = lsq_io_forward_0_addrInvalidSqIdx_value; // @[MemBlock.scala 350:33]
  assign LoadUnit_0_io_lsq_storeLoadViolationQuery_resp_bits_index =
    lsq_io_ldu_s2_storeLoadViolationQuery_0_resp_bits_index; // @[MemBlock.scala 358:49]
  assign LoadUnit_0_io_lsq_storeLoadViolationQuery_resp_bits_canAccept =
    lsq_io_ldu_s2_storeLoadViolationQuery_0_resp_bits_canAccept; // @[MemBlock.scala 358:49]
  assign LoadUnit_0_io_lsq_storeLoadViolationQuery_resp_bits_allocated =
    lsq_io_ldu_s2_storeLoadViolationQuery_0_resp_bits_allocated; // @[MemBlock.scala 358:49]
  assign LoadUnit_0_io_lsq_loadLoadViolationQuery_resp_valid = lsq_io_ldu_s2_loadLoadViolationQuery_0_resp_valid; // @[MemBlock.scala 357:48]
  assign LoadUnit_0_io_lsq_loadLoadViolationQuery_resp_bits_index =
    lsq_io_ldu_s2_loadLoadViolationQuery_0_resp_bits_index; // @[MemBlock.scala 357:48]
  assign LoadUnit_0_io_lsq_loadLoadViolationQuery_resp_bits_canAccept =
    lsq_io_ldu_s2_loadLoadViolationQuery_0_resp_bits_canAccept; // @[MemBlock.scala 357:48]
  assign LoadUnit_0_io_lsq_loadLoadViolationQuery_resp_bits_allocated =
    lsq_io_ldu_s2_loadLoadViolationQuery_0_resp_bits_allocated; // @[MemBlock.scala 357:48]
  assign LoadUnit_0_io_lsq_loadLoadViolationQuery_resp_bits_replayFromFetch =
    lsq_io_ldu_s2_loadLoadViolationQuery_0_resp_bits_replayFromFetch; // @[MemBlock.scala 357:48]
  assign LoadUnit_0_io_lsq_trigger_lqLoadAddrTriggerHitVec_0 = lsq_io_trigger_0_lqLoadAddrTriggerHitVec_0; // @[MemBlock.scala 402:23]
  assign LoadUnit_0_io_lsq_trigger_lqLoadAddrTriggerHitVec_1 = lsq_io_trigger_0_lqLoadAddrTriggerHitVec_1; // @[MemBlock.scala 402:23]
  assign LoadUnit_0_io_lsq_trigger_lqLoadAddrTriggerHitVec_2 = lsq_io_trigger_0_lqLoadAddrTriggerHitVec_2; // @[MemBlock.scala 402:23]
  assign LoadUnit_0_io_tlDchannel_valid = dcache_io_lsu_forward_D_0_valid; // @[MemBlock.scala 354:32]
  assign LoadUnit_0_io_tlDchannel_data = dcache_io_lsu_forward_D_0_data; // @[MemBlock.scala 354:32]
  assign LoadUnit_0_io_tlDchannel_mshrid = dcache_io_lsu_forward_D_0_mshrid; // @[MemBlock.scala 354:32]
  assign LoadUnit_0_io_tlDchannel_last = dcache_io_lsu_forward_D_0_last; // @[MemBlock.scala 354:32]
  assign LoadUnit_0_io_forward_mshr_forward_mshr = dcache_io_lsu_forward_mshr_0_forward_mshr; // @[MemBlock.scala 355:34]
  assign LoadUnit_0_io_forward_mshr_forwardData_0 = dcache_io_lsu_forward_mshr_0_forwardData_0; // @[MemBlock.scala 355:34]
  assign LoadUnit_0_io_forward_mshr_forwardData_1 = dcache_io_lsu_forward_mshr_0_forwardData_1; // @[MemBlock.scala 355:34]
  assign LoadUnit_0_io_forward_mshr_forwardData_2 = dcache_io_lsu_forward_mshr_0_forwardData_2; // @[MemBlock.scala 355:34]
  assign LoadUnit_0_io_forward_mshr_forwardData_3 = dcache_io_lsu_forward_mshr_0_forwardData_3; // @[MemBlock.scala 355:34]
  assign LoadUnit_0_io_forward_mshr_forwardData_4 = dcache_io_lsu_forward_mshr_0_forwardData_4; // @[MemBlock.scala 355:34]
  assign LoadUnit_0_io_forward_mshr_forwardData_5 = dcache_io_lsu_forward_mshr_0_forwardData_5; // @[MemBlock.scala 355:34]
  assign LoadUnit_0_io_forward_mshr_forwardData_6 = dcache_io_lsu_forward_mshr_0_forwardData_6; // @[MemBlock.scala 355:34]
  assign LoadUnit_0_io_forward_mshr_forwardData_7 = dcache_io_lsu_forward_mshr_0_forwardData_7; // @[MemBlock.scala 355:34]
  assign LoadUnit_0_io_forward_mshr_forwardData_8 = dcache_io_lsu_forward_mshr_0_forwardData_8; // @[MemBlock.scala 355:34]
  assign LoadUnit_0_io_forward_mshr_forwardData_9 = dcache_io_lsu_forward_mshr_0_forwardData_9; // @[MemBlock.scala 355:34]
  assign LoadUnit_0_io_forward_mshr_forwardData_10 = dcache_io_lsu_forward_mshr_0_forwardData_10; // @[MemBlock.scala 355:34]
  assign LoadUnit_0_io_forward_mshr_forwardData_11 = dcache_io_lsu_forward_mshr_0_forwardData_11; // @[MemBlock.scala 355:34]
  assign LoadUnit_0_io_forward_mshr_forwardData_12 = dcache_io_lsu_forward_mshr_0_forwardData_12; // @[MemBlock.scala 355:34]
  assign LoadUnit_0_io_forward_mshr_forwardData_13 = dcache_io_lsu_forward_mshr_0_forwardData_13; // @[MemBlock.scala 355:34]
  assign LoadUnit_0_io_forward_mshr_forwardData_14 = dcache_io_lsu_forward_mshr_0_forwardData_14; // @[MemBlock.scala 355:34]
  assign LoadUnit_0_io_forward_mshr_forwardData_15 = dcache_io_lsu_forward_mshr_0_forwardData_15; // @[MemBlock.scala 355:34]
  assign LoadUnit_0_io_forward_mshr_forward_result_valid = dcache_io_lsu_forward_mshr_0_forward_result_valid; // @[MemBlock.scala 355:34]
  assign LoadUnit_0_io_trigger_0_tdata2 = tdata_2_tdata2; // @[MemBlock.scala 416:41]
  assign LoadUnit_0_io_trigger_0_matchType = tdata_2_matchType; // @[MemBlock.scala 417:44]
  assign LoadUnit_0_io_trigger_0_tEnable = tEnable_2; // @[MemBlock.scala 418:42]
  assign LoadUnit_0_io_trigger_1_tdata2 = tdata_3_tdata2; // @[MemBlock.scala 416:41]
  assign LoadUnit_0_io_trigger_1_matchType = tdata_3_matchType; // @[MemBlock.scala 417:44]
  assign LoadUnit_0_io_trigger_1_tEnable = tEnable_3; // @[MemBlock.scala 418:42]
  assign LoadUnit_0_io_trigger_2_tdata2 = tdata_5_tdata2; // @[MemBlock.scala 416:41]
  assign LoadUnit_0_io_trigger_2_matchType = tdata_5_matchType; // @[MemBlock.scala 417:44]
  assign LoadUnit_0_io_trigger_2_tEnable = tEnable_5; // @[MemBlock.scala 418:42]
  assign LoadUnit_0_io_tlb_resp_bits_paddr_0 = dtlb_ld_tlb_ld_io_requestor_0_resp_bits_paddr_0; // @[MemBlock.scala 245:{24,24}]
  assign LoadUnit_0_io_tlb_resp_bits_paddr_1 = dtlb_ld_tlb_ld_io_requestor_0_resp_bits_paddr_1; // @[MemBlock.scala 245:{24,24}]
  assign LoadUnit_0_io_tlb_resp_bits_miss = dtlb_ld_tlb_ld_io_requestor_0_resp_bits_miss; // @[MemBlock.scala 245:{24,24}]
  assign LoadUnit_0_io_tlb_resp_bits_excp_0_pf_ld = dtlb_ld_tlb_ld_io_requestor_0_resp_bits_excp_0_pf_ld; // @[MemBlock.scala 245:{24,24}]
  assign LoadUnit_0_io_tlb_resp_bits_excp_0_af_ld = dtlb_ld_tlb_ld_io_requestor_0_resp_bits_excp_0_af_ld; // @[MemBlock.scala 245:{24,24}]
  assign LoadUnit_0_io_tlb_resp_bits_static_pm_valid = dtlb_ld_tlb_ld_io_requestor_0_resp_bits_static_pm_valid; // @[MemBlock.scala 245:{24,24}]
  assign LoadUnit_0_io_tlb_resp_bits_static_pm_bits = dtlb_ld_tlb_ld_io_requestor_0_resp_bits_static_pm_bits; // @[MemBlock.scala 245:{24,24}]
  assign LoadUnit_0_io_pmp_ld = PMPChecker_io_resp_ld; // @[MemBlock.scala 314:{26,26}]
  assign LoadUnit_0_io_pmp_mmio = PMPChecker_io_resp_mmio; // @[MemBlock.scala 314:{26,26}]
  assign LoadUnit_0_io_fastpathIn_data = LoadUnit_0_io_fastpathOut_valid ? LoadUnit_0_io_fastpathOut_data :
    LoadUnit_1_io_fastpathOut_data; // @[ParallelMux.scala 90:77]
  assign LoadUnit_0_io_fastpathIn_valid = |_LoadUnit_0_io_fastpathIn_valid_T; // @[MemBlock.scala 391:70]
  assign LoadUnit_0_io_loadFastMatch = LoadUnit_0_io_fastpathOut_valid ? fastMatchVec_0 : fastMatchVec_1; // @[ParallelMux.scala 90:77]
  assign LoadUnit_0_io_loadFastImm = io_loadFastImm_0; // @[MemBlock.scala 395:33]
  assign LoadUnit_0_io_csrCtrl_ldld_vio_check_enable = csrCtrl_delay_io_out_ldld_vio_check_enable; // @[MemBlock.scala 359:35]
  assign LoadUnit_0_io_csrCtrl_cache_error_enable = csrCtrl_delay_io_out_cache_error_enable; // @[MemBlock.scala 359:35]
  assign LoadUnit_0_io_correctTableQuery_resp_strict = correctTable_io_issue_0_resp_strict; // @[MemBlock.scala 367:39]
  assign LoadUnit_0_io_reExecuteQuery_0_valid = StoreUnit_0_io_reExecuteQuery_valid; // @[MemBlock.scala 371:41]
  assign LoadUnit_0_io_reExecuteQuery_0_bits_robIdx_flag = StoreUnit_0_io_reExecuteQuery_bits_robIdx_flag; // @[MemBlock.scala 371:41]
  assign LoadUnit_0_io_reExecuteQuery_0_bits_robIdx_value = StoreUnit_0_io_reExecuteQuery_bits_robIdx_value; // @[MemBlock.scala 371:41]
  assign LoadUnit_0_io_reExecuteQuery_0_bits_paddr = StoreUnit_0_io_reExecuteQuery_bits_paddr; // @[MemBlock.scala 371:41]
  assign LoadUnit_0_io_reExecuteQuery_0_bits_mask = StoreUnit_0_io_reExecuteQuery_bits_mask; // @[MemBlock.scala 371:41]
  assign LoadUnit_0_io_reExecuteQuery_1_valid = StoreUnit_1_io_reExecuteQuery_valid; // @[MemBlock.scala 371:41]
  assign LoadUnit_0_io_reExecuteQuery_1_bits_robIdx_flag = StoreUnit_1_io_reExecuteQuery_bits_robIdx_flag; // @[MemBlock.scala 371:41]
  assign LoadUnit_0_io_reExecuteQuery_1_bits_robIdx_value = StoreUnit_1_io_reExecuteQuery_bits_robIdx_value; // @[MemBlock.scala 371:41]
  assign LoadUnit_0_io_reExecuteQuery_1_bits_paddr = StoreUnit_1_io_reExecuteQuery_bits_paddr; // @[MemBlock.scala 371:41]
  assign LoadUnit_0_io_reExecuteQuery_1_bits_mask = StoreUnit_1_io_reExecuteQuery_bits_mask; // @[MemBlock.scala 371:41]
  assign LoadUnit_0_io_replay_valid = lsq_io_replay_0_valid; // @[MemBlock.scala 396:28]
  assign LoadUnit_0_io_replay_bits_uop_cf_foldpc = lsq_io_replay_0_bits_uop_cf_foldpc; // @[MemBlock.scala 396:28]
  assign LoadUnit_0_io_replay_bits_uop_cf_trigger_backendEn_1 = lsq_io_replay_0_bits_uop_cf_trigger_backendEn_1; // @[MemBlock.scala 396:28]
  assign LoadUnit_0_io_replay_bits_uop_cf_trigger_backendHit_0 = lsq_io_replay_0_bits_uop_cf_trigger_backendHit_0; // @[MemBlock.scala 396:28]
  assign LoadUnit_0_io_replay_bits_uop_cf_trigger_backendHit_1 = lsq_io_replay_0_bits_uop_cf_trigger_backendHit_1; // @[MemBlock.scala 396:28]
  assign LoadUnit_0_io_replay_bits_uop_cf_trigger_backendHit_4 = lsq_io_replay_0_bits_uop_cf_trigger_backendHit_4; // @[MemBlock.scala 396:28]
  assign LoadUnit_0_io_replay_bits_uop_cf_waitForRobIdx_flag = lsq_io_replay_0_bits_uop_cf_waitForRobIdx_flag; // @[MemBlock.scala 396:28]
  assign LoadUnit_0_io_replay_bits_uop_cf_waitForRobIdx_value = lsq_io_replay_0_bits_uop_cf_waitForRobIdx_value; // @[MemBlock.scala 396:28]
  assign LoadUnit_0_io_replay_bits_uop_cf_loadWaitBit = lsq_io_replay_0_bits_uop_cf_loadWaitBit; // @[MemBlock.scala 396:28]
  assign LoadUnit_0_io_replay_bits_uop_cf_loadWaitStrict = lsq_io_replay_0_bits_uop_cf_loadWaitStrict; // @[MemBlock.scala 396:28]
  assign LoadUnit_0_io_replay_bits_uop_cf_ftqPtr_flag = lsq_io_replay_0_bits_uop_cf_ftqPtr_flag; // @[MemBlock.scala 396:28]
  assign LoadUnit_0_io_replay_bits_uop_cf_ftqPtr_value = lsq_io_replay_0_bits_uop_cf_ftqPtr_value; // @[MemBlock.scala 396:28]
  assign LoadUnit_0_io_replay_bits_uop_cf_ftqOffset = lsq_io_replay_0_bits_uop_cf_ftqOffset; // @[MemBlock.scala 396:28]
  assign LoadUnit_0_io_replay_bits_uop_ctrl_fuType = lsq_io_replay_0_bits_uop_ctrl_fuType; // @[MemBlock.scala 396:28]
  assign LoadUnit_0_io_replay_bits_uop_ctrl_fuOpType = lsq_io_replay_0_bits_uop_ctrl_fuOpType; // @[MemBlock.scala 396:28]
  assign LoadUnit_0_io_replay_bits_uop_ctrl_rfWen = lsq_io_replay_0_bits_uop_ctrl_rfWen; // @[MemBlock.scala 396:28]
  assign LoadUnit_0_io_replay_bits_uop_ctrl_fpWen = lsq_io_replay_0_bits_uop_ctrl_fpWen; // @[MemBlock.scala 396:28]
  assign LoadUnit_0_io_replay_bits_uop_pdest = lsq_io_replay_0_bits_uop_pdest; // @[MemBlock.scala 396:28]
  assign LoadUnit_0_io_replay_bits_uop_robIdx_flag = lsq_io_replay_0_bits_uop_robIdx_flag; // @[MemBlock.scala 396:28]
  assign LoadUnit_0_io_replay_bits_uop_robIdx_value = lsq_io_replay_0_bits_uop_robIdx_value; // @[MemBlock.scala 396:28]
  assign LoadUnit_0_io_replay_bits_uop_lqIdx_flag = lsq_io_replay_0_bits_uop_lqIdx_flag; // @[MemBlock.scala 396:28]
  assign LoadUnit_0_io_replay_bits_uop_lqIdx_value = lsq_io_replay_0_bits_uop_lqIdx_value; // @[MemBlock.scala 396:28]
  assign LoadUnit_0_io_replay_bits_uop_sqIdx_flag = lsq_io_replay_0_bits_uop_sqIdx_flag; // @[MemBlock.scala 396:28]
  assign LoadUnit_0_io_replay_bits_uop_sqIdx_value = lsq_io_replay_0_bits_uop_sqIdx_value; // @[MemBlock.scala 396:28]
  assign LoadUnit_0_io_replay_bits_vaddr = lsq_io_replay_0_bits_vaddr; // @[MemBlock.scala 396:28]
  assign LoadUnit_0_io_replay_bits_isFirstIssue = lsq_io_replay_0_bits_isFirstIssue; // @[MemBlock.scala 396:28]
  assign LoadUnit_0_io_replay_bits_replayCarry_real_way_en = lsq_io_replay_0_bits_replayCarry_real_way_en; // @[MemBlock.scala 396:28]
  assign LoadUnit_0_io_replay_bits_replayCarry_valid = lsq_io_replay_0_bits_replayCarry_valid; // @[MemBlock.scala 396:28]
  assign LoadUnit_0_io_replay_bits_mshrid = lsq_io_replay_0_bits_mshrid; // @[MemBlock.scala 396:28]
  assign LoadUnit_0_io_replay_bits_forward_tlDchannel = lsq_io_replay_0_bits_forward_tlDchannel; // @[MemBlock.scala 396:28]
  assign LoadUnit_0_io_replay_bits_rarAllocated = lsq_io_replay_0_bits_rarAllocated; // @[MemBlock.scala 396:28]
  assign LoadUnit_0_io_replay_bits_rarIndex = lsq_io_replay_0_bits_rarIndex; // @[MemBlock.scala 396:28]
  assign LoadUnit_0_io_replay_bits_rawAllocated = lsq_io_replay_0_bits_rawAllocated; // @[MemBlock.scala 396:28]
  assign LoadUnit_0_io_replay_bits_rawIndex = lsq_io_replay_0_bits_rawIndex; // @[MemBlock.scala 396:28]
  assign LoadUnit_0_io_lqReplayFull = lsq_io_lqReplayFull; // @[MemBlock.scala 373:34]
  assign LoadUnit_1_clock = clock;
  assign LoadUnit_1_reset = reset;
  assign LoadUnit_1_io_loadIn_valid = io_issue_1_valid; // @[MemBlock.scala 344:28]
  assign LoadUnit_1_io_loadIn_bits_uop_cf_foldpc = io_issue_1_bits_uop_cf_foldpc; // @[MemBlock.scala 344:28]
  assign LoadUnit_1_io_loadIn_bits_uop_cf_trigger_backendEn_1 = io_issue_1_bits_uop_cf_trigger_backendEn_1; // @[MemBlock.scala 344:28]
  assign LoadUnit_1_io_loadIn_bits_uop_cf_waitForRobIdx_flag = io_issue_1_bits_uop_cf_waitForRobIdx_flag; // @[MemBlock.scala 344:28]
  assign LoadUnit_1_io_loadIn_bits_uop_cf_waitForRobIdx_value = io_issue_1_bits_uop_cf_waitForRobIdx_value; // @[MemBlock.scala 344:28]
  assign LoadUnit_1_io_loadIn_bits_uop_cf_loadWaitBit = io_issue_1_bits_uop_cf_loadWaitBit; // @[MemBlock.scala 344:28]
  assign LoadUnit_1_io_loadIn_bits_uop_cf_loadWaitStrict = io_issue_1_bits_uop_cf_loadWaitStrict; // @[MemBlock.scala 344:28]
  assign LoadUnit_1_io_loadIn_bits_uop_cf_ftqPtr_flag = io_issue_1_bits_uop_cf_ftqPtr_flag; // @[MemBlock.scala 344:28]
  assign LoadUnit_1_io_loadIn_bits_uop_cf_ftqPtr_value = io_issue_1_bits_uop_cf_ftqPtr_value; // @[MemBlock.scala 344:28]
  assign LoadUnit_1_io_loadIn_bits_uop_cf_ftqOffset = io_issue_1_bits_uop_cf_ftqOffset; // @[MemBlock.scala 344:28]
  assign LoadUnit_1_io_loadIn_bits_uop_ctrl_fuType = io_issue_1_bits_uop_ctrl_fuType; // @[MemBlock.scala 344:28]
  assign LoadUnit_1_io_loadIn_bits_uop_ctrl_fuOpType = io_issue_1_bits_uop_ctrl_fuOpType; // @[MemBlock.scala 344:28]
  assign LoadUnit_1_io_loadIn_bits_uop_ctrl_rfWen = io_issue_1_bits_uop_ctrl_rfWen; // @[MemBlock.scala 344:28]
  assign LoadUnit_1_io_loadIn_bits_uop_ctrl_fpWen = io_issue_1_bits_uop_ctrl_fpWen; // @[MemBlock.scala 344:28]
  assign LoadUnit_1_io_loadIn_bits_uop_ctrl_imm = io_issue_1_bits_uop_ctrl_imm; // @[MemBlock.scala 344:28]
  assign LoadUnit_1_io_loadIn_bits_uop_pdest = io_issue_1_bits_uop_pdest; // @[MemBlock.scala 344:28]
  assign LoadUnit_1_io_loadIn_bits_uop_robIdx_flag = io_issue_1_bits_uop_robIdx_flag; // @[MemBlock.scala 344:28]
  assign LoadUnit_1_io_loadIn_bits_uop_robIdx_value = io_issue_1_bits_uop_robIdx_value; // @[MemBlock.scala 344:28]
  assign LoadUnit_1_io_loadIn_bits_uop_lqIdx_flag = io_issue_1_bits_uop_lqIdx_flag; // @[MemBlock.scala 344:28]
  assign LoadUnit_1_io_loadIn_bits_uop_lqIdx_value = io_issue_1_bits_uop_lqIdx_value; // @[MemBlock.scala 344:28]
  assign LoadUnit_1_io_loadIn_bits_uop_sqIdx_flag = io_issue_1_bits_uop_sqIdx_flag; // @[MemBlock.scala 344:28]
  assign LoadUnit_1_io_loadIn_bits_uop_sqIdx_value = io_issue_1_bits_uop_sqIdx_value; // @[MemBlock.scala 344:28]
  assign LoadUnit_1_io_loadIn_bits_src_0 = io_issue_1_bits_src_0; // @[MemBlock.scala 344:28]
  assign LoadUnit_1_io_VecloadIn_valid = vlflowqueue_io_loadPipeOut_1_valid; // @[MemBlock.scala 346:31]
  assign LoadUnit_1_io_VecloadIn_bits_vaddr = vlflowqueue_io_loadPipeOut_1_bits_vaddr; // @[MemBlock.scala 346:31]
  assign LoadUnit_1_io_redirect_valid = redirect_next_valid_REG; // @[BitUtils.scala 26:20 28:18]
  assign LoadUnit_1_io_redirect_bits_robIdx_flag = redirect_next_bits_rrobIdx_flag; // @[BitUtils.scala 26:20 33:15]
  assign LoadUnit_1_io_redirect_bits_robIdx_value = redirect_next_bits_rrobIdx_value; // @[BitUtils.scala 26:20 33:15]
  assign LoadUnit_1_io_redirect_bits_level = redirect_next_bits_rlevel; // @[BitUtils.scala 26:20 33:15]
  assign LoadUnit_1_io_dcache_req_ready = dcache_io_lsu_load_1_req_ready; // @[MemBlock.scala 348:28]
  assign LoadUnit_1_io_dcache_resp_bits_data_delayed = dcache_io_lsu_load_1_resp_bits_data_delayed; // @[MemBlock.scala 348:28]
  assign LoadUnit_1_io_dcache_resp_bits_miss = dcache_io_lsu_load_1_resp_bits_miss; // @[MemBlock.scala 348:28]
  assign LoadUnit_1_io_dcache_resp_bits_replay = dcache_io_lsu_load_1_resp_bits_replay; // @[MemBlock.scala 348:28]
  assign LoadUnit_1_io_dcache_resp_bits_replayCarry_real_way_en = dcache_io_lsu_load_1_resp_bits_replayCarry_real_way_en
    ; // @[MemBlock.scala 348:28]
  assign LoadUnit_1_io_dcache_resp_bits_replayCarry_valid = dcache_io_lsu_load_1_resp_bits_replayCarry_valid; // @[MemBlock.scala 348:28]
  assign LoadUnit_1_io_dcache_resp_bits_tag_error = dcache_io_lsu_load_1_resp_bits_tag_error; // @[MemBlock.scala 348:28]
  assign LoadUnit_1_io_dcache_resp_bits_mshr_id = dcache_io_lsu_load_1_resp_bits_mshr_id; // @[MemBlock.scala 348:28]
  assign LoadUnit_1_io_dcache_resp_bits_error_delayed = dcache_io_lsu_load_1_resp_bits_error_delayed; // @[MemBlock.scala 348:28]
  assign LoadUnit_1_io_dcache_s1_bank_conflict = dcache_io_lsu_load_1_s1_bank_conflict; // @[MemBlock.scala 348:28]
  assign LoadUnit_1_io_sbuffer_forwardMask_0 = sbuffer_io_forward_1_forwardMask_0; // @[MemBlock.scala 351:29]
  assign LoadUnit_1_io_sbuffer_forwardMask_1 = sbuffer_io_forward_1_forwardMask_1; // @[MemBlock.scala 351:29]
  assign LoadUnit_1_io_sbuffer_forwardMask_2 = sbuffer_io_forward_1_forwardMask_2; // @[MemBlock.scala 351:29]
  assign LoadUnit_1_io_sbuffer_forwardMask_3 = sbuffer_io_forward_1_forwardMask_3; // @[MemBlock.scala 351:29]
  assign LoadUnit_1_io_sbuffer_forwardMask_4 = sbuffer_io_forward_1_forwardMask_4; // @[MemBlock.scala 351:29]
  assign LoadUnit_1_io_sbuffer_forwardMask_5 = sbuffer_io_forward_1_forwardMask_5; // @[MemBlock.scala 351:29]
  assign LoadUnit_1_io_sbuffer_forwardMask_6 = sbuffer_io_forward_1_forwardMask_6; // @[MemBlock.scala 351:29]
  assign LoadUnit_1_io_sbuffer_forwardMask_7 = sbuffer_io_forward_1_forwardMask_7; // @[MemBlock.scala 351:29]
  assign LoadUnit_1_io_sbuffer_forwardMask_8 = sbuffer_io_forward_1_forwardMask_8; // @[MemBlock.scala 351:29]
  assign LoadUnit_1_io_sbuffer_forwardMask_9 = sbuffer_io_forward_1_forwardMask_9; // @[MemBlock.scala 351:29]
  assign LoadUnit_1_io_sbuffer_forwardMask_10 = sbuffer_io_forward_1_forwardMask_10; // @[MemBlock.scala 351:29]
  assign LoadUnit_1_io_sbuffer_forwardMask_11 = sbuffer_io_forward_1_forwardMask_11; // @[MemBlock.scala 351:29]
  assign LoadUnit_1_io_sbuffer_forwardMask_12 = sbuffer_io_forward_1_forwardMask_12; // @[MemBlock.scala 351:29]
  assign LoadUnit_1_io_sbuffer_forwardMask_13 = sbuffer_io_forward_1_forwardMask_13; // @[MemBlock.scala 351:29]
  assign LoadUnit_1_io_sbuffer_forwardMask_14 = sbuffer_io_forward_1_forwardMask_14; // @[MemBlock.scala 351:29]
  assign LoadUnit_1_io_sbuffer_forwardMask_15 = sbuffer_io_forward_1_forwardMask_15; // @[MemBlock.scala 351:29]
  assign LoadUnit_1_io_sbuffer_forwardData_0 = sbuffer_io_forward_1_forwardData_0; // @[MemBlock.scala 351:29]
  assign LoadUnit_1_io_sbuffer_forwardData_1 = sbuffer_io_forward_1_forwardData_1; // @[MemBlock.scala 351:29]
  assign LoadUnit_1_io_sbuffer_forwardData_2 = sbuffer_io_forward_1_forwardData_2; // @[MemBlock.scala 351:29]
  assign LoadUnit_1_io_sbuffer_forwardData_3 = sbuffer_io_forward_1_forwardData_3; // @[MemBlock.scala 351:29]
  assign LoadUnit_1_io_sbuffer_forwardData_4 = sbuffer_io_forward_1_forwardData_4; // @[MemBlock.scala 351:29]
  assign LoadUnit_1_io_sbuffer_forwardData_5 = sbuffer_io_forward_1_forwardData_5; // @[MemBlock.scala 351:29]
  assign LoadUnit_1_io_sbuffer_forwardData_6 = sbuffer_io_forward_1_forwardData_6; // @[MemBlock.scala 351:29]
  assign LoadUnit_1_io_sbuffer_forwardData_7 = sbuffer_io_forward_1_forwardData_7; // @[MemBlock.scala 351:29]
  assign LoadUnit_1_io_sbuffer_forwardData_8 = sbuffer_io_forward_1_forwardData_8; // @[MemBlock.scala 351:29]
  assign LoadUnit_1_io_sbuffer_forwardData_9 = sbuffer_io_forward_1_forwardData_9; // @[MemBlock.scala 351:29]
  assign LoadUnit_1_io_sbuffer_forwardData_10 = sbuffer_io_forward_1_forwardData_10; // @[MemBlock.scala 351:29]
  assign LoadUnit_1_io_sbuffer_forwardData_11 = sbuffer_io_forward_1_forwardData_11; // @[MemBlock.scala 351:29]
  assign LoadUnit_1_io_sbuffer_forwardData_12 = sbuffer_io_forward_1_forwardData_12; // @[MemBlock.scala 351:29]
  assign LoadUnit_1_io_sbuffer_forwardData_13 = sbuffer_io_forward_1_forwardData_13; // @[MemBlock.scala 351:29]
  assign LoadUnit_1_io_sbuffer_forwardData_14 = sbuffer_io_forward_1_forwardData_14; // @[MemBlock.scala 351:29]
  assign LoadUnit_1_io_sbuffer_forwardData_15 = sbuffer_io_forward_1_forwardData_15; // @[MemBlock.scala 351:29]
  assign LoadUnit_1_io_sbuffer_matchInvalid = sbuffer_io_forward_1_matchInvalid; // @[MemBlock.scala 351:29]
  assign LoadUnit_1_io_lsq_loadOut_valid = 1'h0; // @[MemBlock.scala 400:23]
  assign LoadUnit_1_io_lsq_loadOut_bits_uop_cf_exceptionVec_4 = 1'h0; // @[MemBlock.scala 400:23]
  assign LoadUnit_1_io_lsq_loadOut_bits_uop_cf_exceptionVec_5 = 1'h0; // @[MemBlock.scala 400:23]
  assign LoadUnit_1_io_lsq_loadOut_bits_uop_cf_exceptionVec_13 = 1'h0; // @[MemBlock.scala 400:23]
  assign LoadUnit_1_io_lsq_loadOut_bits_uop_cf_trigger_backendEn_1 = 1'h0; // @[MemBlock.scala 400:23]
  assign LoadUnit_1_io_lsq_loadOut_bits_uop_cf_trigger_backendHit_0 = 1'h0; // @[MemBlock.scala 400:23]
  assign LoadUnit_1_io_lsq_loadOut_bits_uop_cf_trigger_backendHit_1 = 1'h0; // @[MemBlock.scala 400:23]
  assign LoadUnit_1_io_lsq_loadOut_bits_uop_cf_trigger_backendHit_4 = 1'h0; // @[MemBlock.scala 400:23]
  assign LoadUnit_1_io_lsq_loadOut_bits_uop_ctrl_rfWen = 1'h0; // @[MemBlock.scala 400:23]
  assign LoadUnit_1_io_lsq_loadOut_bits_uop_ctrl_fpWen = 1'h0; // @[MemBlock.scala 400:23]
  assign LoadUnit_1_io_lsq_loadOut_bits_uop_ctrl_flushPipe = 1'h0; // @[MemBlock.scala 400:23]
  assign LoadUnit_1_io_lsq_loadOut_bits_uop_ctrl_replayInst = 1'h0; // @[MemBlock.scala 400:23]
  assign LoadUnit_1_io_lsq_loadOut_bits_uop_pdest = 6'h0; // @[MemBlock.scala 400:23]
  assign LoadUnit_1_io_lsq_loadOut_bits_uop_robIdx_flag = 1'h0; // @[MemBlock.scala 400:23]
  assign LoadUnit_1_io_lsq_loadOut_bits_uop_robIdx_value = 5'h0; // @[MemBlock.scala 400:23]
  assign LoadUnit_1_io_lsq_loadOut_bits_debug_isMMIO = 1'h0; // @[MemBlock.scala 400:23]
  assign LoadUnit_1_io_lsq_ldRawData_lqData = 64'h0; // @[MemBlock.scala 401:28]
  assign LoadUnit_1_io_lsq_ldRawData_uop_ctrl_fuOpType = 7'h0; // @[MemBlock.scala 401:28]
  assign LoadUnit_1_io_lsq_ldRawData_uop_ctrl_fpWen = 1'h0; // @[MemBlock.scala 401:28]
  assign LoadUnit_1_io_lsq_ldRawData_addrOffset = 3'h0; // @[MemBlock.scala 401:28]
  assign LoadUnit_1_io_lsq_forward_forwardMask_0 = lsq_io_forward_1_forwardMask_0; // @[MemBlock.scala 350:33]
  assign LoadUnit_1_io_lsq_forward_forwardMask_1 = lsq_io_forward_1_forwardMask_1; // @[MemBlock.scala 350:33]
  assign LoadUnit_1_io_lsq_forward_forwardMask_2 = lsq_io_forward_1_forwardMask_2; // @[MemBlock.scala 350:33]
  assign LoadUnit_1_io_lsq_forward_forwardMask_3 = lsq_io_forward_1_forwardMask_3; // @[MemBlock.scala 350:33]
  assign LoadUnit_1_io_lsq_forward_forwardMask_4 = lsq_io_forward_1_forwardMask_4; // @[MemBlock.scala 350:33]
  assign LoadUnit_1_io_lsq_forward_forwardMask_5 = lsq_io_forward_1_forwardMask_5; // @[MemBlock.scala 350:33]
  assign LoadUnit_1_io_lsq_forward_forwardMask_6 = lsq_io_forward_1_forwardMask_6; // @[MemBlock.scala 350:33]
  assign LoadUnit_1_io_lsq_forward_forwardMask_7 = lsq_io_forward_1_forwardMask_7; // @[MemBlock.scala 350:33]
  assign LoadUnit_1_io_lsq_forward_forwardMask_8 = lsq_io_forward_1_forwardMask_8; // @[MemBlock.scala 350:33]
  assign LoadUnit_1_io_lsq_forward_forwardMask_9 = lsq_io_forward_1_forwardMask_9; // @[MemBlock.scala 350:33]
  assign LoadUnit_1_io_lsq_forward_forwardMask_10 = lsq_io_forward_1_forwardMask_10; // @[MemBlock.scala 350:33]
  assign LoadUnit_1_io_lsq_forward_forwardMask_11 = lsq_io_forward_1_forwardMask_11; // @[MemBlock.scala 350:33]
  assign LoadUnit_1_io_lsq_forward_forwardMask_12 = lsq_io_forward_1_forwardMask_12; // @[MemBlock.scala 350:33]
  assign LoadUnit_1_io_lsq_forward_forwardMask_13 = lsq_io_forward_1_forwardMask_13; // @[MemBlock.scala 350:33]
  assign LoadUnit_1_io_lsq_forward_forwardMask_14 = lsq_io_forward_1_forwardMask_14; // @[MemBlock.scala 350:33]
  assign LoadUnit_1_io_lsq_forward_forwardMask_15 = lsq_io_forward_1_forwardMask_15; // @[MemBlock.scala 350:33]
  assign LoadUnit_1_io_lsq_forward_forwardData_0 = lsq_io_forward_1_forwardData_0; // @[MemBlock.scala 350:33]
  assign LoadUnit_1_io_lsq_forward_forwardData_1 = lsq_io_forward_1_forwardData_1; // @[MemBlock.scala 350:33]
  assign LoadUnit_1_io_lsq_forward_forwardData_2 = lsq_io_forward_1_forwardData_2; // @[MemBlock.scala 350:33]
  assign LoadUnit_1_io_lsq_forward_forwardData_3 = lsq_io_forward_1_forwardData_3; // @[MemBlock.scala 350:33]
  assign LoadUnit_1_io_lsq_forward_forwardData_4 = lsq_io_forward_1_forwardData_4; // @[MemBlock.scala 350:33]
  assign LoadUnit_1_io_lsq_forward_forwardData_5 = lsq_io_forward_1_forwardData_5; // @[MemBlock.scala 350:33]
  assign LoadUnit_1_io_lsq_forward_forwardData_6 = lsq_io_forward_1_forwardData_6; // @[MemBlock.scala 350:33]
  assign LoadUnit_1_io_lsq_forward_forwardData_7 = lsq_io_forward_1_forwardData_7; // @[MemBlock.scala 350:33]
  assign LoadUnit_1_io_lsq_forward_forwardData_8 = lsq_io_forward_1_forwardData_8; // @[MemBlock.scala 350:33]
  assign LoadUnit_1_io_lsq_forward_forwardData_9 = lsq_io_forward_1_forwardData_9; // @[MemBlock.scala 350:33]
  assign LoadUnit_1_io_lsq_forward_forwardData_10 = lsq_io_forward_1_forwardData_10; // @[MemBlock.scala 350:33]
  assign LoadUnit_1_io_lsq_forward_forwardData_11 = lsq_io_forward_1_forwardData_11; // @[MemBlock.scala 350:33]
  assign LoadUnit_1_io_lsq_forward_forwardData_12 = lsq_io_forward_1_forwardData_12; // @[MemBlock.scala 350:33]
  assign LoadUnit_1_io_lsq_forward_forwardData_13 = lsq_io_forward_1_forwardData_13; // @[MemBlock.scala 350:33]
  assign LoadUnit_1_io_lsq_forward_forwardData_14 = lsq_io_forward_1_forwardData_14; // @[MemBlock.scala 350:33]
  assign LoadUnit_1_io_lsq_forward_forwardData_15 = lsq_io_forward_1_forwardData_15; // @[MemBlock.scala 350:33]
  assign LoadUnit_1_io_lsq_forward_dataInvalid = lsq_io_forward_1_dataInvalid; // @[MemBlock.scala 350:33]
  assign LoadUnit_1_io_lsq_forward_matchInvalid = lsq_io_forward_1_matchInvalid; // @[MemBlock.scala 350:33]
  assign LoadUnit_1_io_lsq_forward_schedWait = lsq_io_forward_1_schedWait; // @[MemBlock.scala 350:33]
  assign LoadUnit_1_io_lsq_forward_dataInvalidSqIdx_flag = lsq_io_forward_1_dataInvalidSqIdx_flag; // @[MemBlock.scala 350:33]
  assign LoadUnit_1_io_lsq_forward_dataInvalidSqIdx_value = lsq_io_forward_1_dataInvalidSqIdx_value; // @[MemBlock.scala 350:33]
  assign LoadUnit_1_io_lsq_forward_addrInvalidSqIdx_flag = lsq_io_forward_1_addrInvalidSqIdx_flag; // @[MemBlock.scala 350:33]
  assign LoadUnit_1_io_lsq_forward_addrInvalidSqIdx_value = lsq_io_forward_1_addrInvalidSqIdx_value; // @[MemBlock.scala 350:33]
  assign LoadUnit_1_io_lsq_storeLoadViolationQuery_resp_bits_index =
    lsq_io_ldu_s2_storeLoadViolationQuery_1_resp_bits_index; // @[MemBlock.scala 358:49]
  assign LoadUnit_1_io_lsq_storeLoadViolationQuery_resp_bits_canAccept =
    lsq_io_ldu_s2_storeLoadViolationQuery_1_resp_bits_canAccept; // @[MemBlock.scala 358:49]
  assign LoadUnit_1_io_lsq_storeLoadViolationQuery_resp_bits_allocated =
    lsq_io_ldu_s2_storeLoadViolationQuery_1_resp_bits_allocated; // @[MemBlock.scala 358:49]
  assign LoadUnit_1_io_lsq_loadLoadViolationQuery_resp_valid = lsq_io_ldu_s2_loadLoadViolationQuery_1_resp_valid; // @[MemBlock.scala 357:48]
  assign LoadUnit_1_io_lsq_loadLoadViolationQuery_resp_bits_index =
    lsq_io_ldu_s2_loadLoadViolationQuery_1_resp_bits_index; // @[MemBlock.scala 357:48]
  assign LoadUnit_1_io_lsq_loadLoadViolationQuery_resp_bits_canAccept =
    lsq_io_ldu_s2_loadLoadViolationQuery_1_resp_bits_canAccept; // @[MemBlock.scala 357:48]
  assign LoadUnit_1_io_lsq_loadLoadViolationQuery_resp_bits_allocated =
    lsq_io_ldu_s2_loadLoadViolationQuery_1_resp_bits_allocated; // @[MemBlock.scala 357:48]
  assign LoadUnit_1_io_lsq_loadLoadViolationQuery_resp_bits_replayFromFetch =
    lsq_io_ldu_s2_loadLoadViolationQuery_1_resp_bits_replayFromFetch; // @[MemBlock.scala 357:48]
  assign LoadUnit_1_io_lsq_trigger_lqLoadAddrTriggerHitVec_0 = 1'h0; // @[MemBlock.scala 402:23]
  assign LoadUnit_1_io_lsq_trigger_lqLoadAddrTriggerHitVec_1 = 1'h0; // @[MemBlock.scala 402:23]
  assign LoadUnit_1_io_lsq_trigger_lqLoadAddrTriggerHitVec_2 = 1'h0; // @[MemBlock.scala 402:23]
  assign LoadUnit_1_io_tlDchannel_valid = dcache_io_lsu_forward_D_1_valid; // @[MemBlock.scala 354:32]
  assign LoadUnit_1_io_tlDchannel_data = dcache_io_lsu_forward_D_1_data; // @[MemBlock.scala 354:32]
  assign LoadUnit_1_io_tlDchannel_mshrid = dcache_io_lsu_forward_D_1_mshrid; // @[MemBlock.scala 354:32]
  assign LoadUnit_1_io_tlDchannel_last = dcache_io_lsu_forward_D_1_last; // @[MemBlock.scala 354:32]
  assign LoadUnit_1_io_forward_mshr_forward_mshr = dcache_io_lsu_forward_mshr_1_forward_mshr; // @[MemBlock.scala 355:34]
  assign LoadUnit_1_io_forward_mshr_forwardData_0 = dcache_io_lsu_forward_mshr_1_forwardData_0; // @[MemBlock.scala 355:34]
  assign LoadUnit_1_io_forward_mshr_forwardData_1 = dcache_io_lsu_forward_mshr_1_forwardData_1; // @[MemBlock.scala 355:34]
  assign LoadUnit_1_io_forward_mshr_forwardData_2 = dcache_io_lsu_forward_mshr_1_forwardData_2; // @[MemBlock.scala 355:34]
  assign LoadUnit_1_io_forward_mshr_forwardData_3 = dcache_io_lsu_forward_mshr_1_forwardData_3; // @[MemBlock.scala 355:34]
  assign LoadUnit_1_io_forward_mshr_forwardData_4 = dcache_io_lsu_forward_mshr_1_forwardData_4; // @[MemBlock.scala 355:34]
  assign LoadUnit_1_io_forward_mshr_forwardData_5 = dcache_io_lsu_forward_mshr_1_forwardData_5; // @[MemBlock.scala 355:34]
  assign LoadUnit_1_io_forward_mshr_forwardData_6 = dcache_io_lsu_forward_mshr_1_forwardData_6; // @[MemBlock.scala 355:34]
  assign LoadUnit_1_io_forward_mshr_forwardData_7 = dcache_io_lsu_forward_mshr_1_forwardData_7; // @[MemBlock.scala 355:34]
  assign LoadUnit_1_io_forward_mshr_forwardData_8 = dcache_io_lsu_forward_mshr_1_forwardData_8; // @[MemBlock.scala 355:34]
  assign LoadUnit_1_io_forward_mshr_forwardData_9 = dcache_io_lsu_forward_mshr_1_forwardData_9; // @[MemBlock.scala 355:34]
  assign LoadUnit_1_io_forward_mshr_forwardData_10 = dcache_io_lsu_forward_mshr_1_forwardData_10; // @[MemBlock.scala 355:34]
  assign LoadUnit_1_io_forward_mshr_forwardData_11 = dcache_io_lsu_forward_mshr_1_forwardData_11; // @[MemBlock.scala 355:34]
  assign LoadUnit_1_io_forward_mshr_forwardData_12 = dcache_io_lsu_forward_mshr_1_forwardData_12; // @[MemBlock.scala 355:34]
  assign LoadUnit_1_io_forward_mshr_forwardData_13 = dcache_io_lsu_forward_mshr_1_forwardData_13; // @[MemBlock.scala 355:34]
  assign LoadUnit_1_io_forward_mshr_forwardData_14 = dcache_io_lsu_forward_mshr_1_forwardData_14; // @[MemBlock.scala 355:34]
  assign LoadUnit_1_io_forward_mshr_forwardData_15 = dcache_io_lsu_forward_mshr_1_forwardData_15; // @[MemBlock.scala 355:34]
  assign LoadUnit_1_io_forward_mshr_forward_result_valid = dcache_io_lsu_forward_mshr_1_forward_result_valid; // @[MemBlock.scala 355:34]
  assign LoadUnit_1_io_trigger_0_tdata2 = tdata_2_tdata2; // @[MemBlock.scala 416:41]
  assign LoadUnit_1_io_trigger_0_matchType = tdata_2_matchType; // @[MemBlock.scala 417:44]
  assign LoadUnit_1_io_trigger_0_tEnable = tEnable_2; // @[MemBlock.scala 418:42]
  assign LoadUnit_1_io_trigger_1_tdata2 = tdata_3_tdata2; // @[MemBlock.scala 416:41]
  assign LoadUnit_1_io_trigger_1_matchType = tdata_3_matchType; // @[MemBlock.scala 417:44]
  assign LoadUnit_1_io_trigger_1_tEnable = tEnable_3; // @[MemBlock.scala 418:42]
  assign LoadUnit_1_io_trigger_2_tdata2 = tdata_5_tdata2; // @[MemBlock.scala 416:41]
  assign LoadUnit_1_io_trigger_2_matchType = tdata_5_matchType; // @[MemBlock.scala 417:44]
  assign LoadUnit_1_io_trigger_2_tEnable = tEnable_5; // @[MemBlock.scala 418:42]
  assign LoadUnit_1_io_tlb_resp_bits_paddr_0 = dtlb_ld_tlb_ld_io_requestor_1_resp_bits_paddr_0; // @[MemBlock.scala 245:{24,24}]
  assign LoadUnit_1_io_tlb_resp_bits_paddr_1 = dtlb_ld_tlb_ld_io_requestor_1_resp_bits_paddr_1; // @[MemBlock.scala 245:{24,24}]
  assign LoadUnit_1_io_tlb_resp_bits_miss = dtlb_ld_tlb_ld_io_requestor_1_resp_bits_miss; // @[MemBlock.scala 245:{24,24}]
  assign LoadUnit_1_io_tlb_resp_bits_excp_0_pf_ld = dtlb_ld_tlb_ld_io_requestor_1_resp_bits_excp_0_pf_ld; // @[MemBlock.scala 245:{24,24}]
  assign LoadUnit_1_io_tlb_resp_bits_excp_0_af_ld = dtlb_ld_tlb_ld_io_requestor_1_resp_bits_excp_0_af_ld; // @[MemBlock.scala 245:{24,24}]
  assign LoadUnit_1_io_tlb_resp_bits_static_pm_valid = dtlb_ld_tlb_ld_io_requestor_1_resp_bits_static_pm_valid; // @[MemBlock.scala 245:{24,24}]
  assign LoadUnit_1_io_tlb_resp_bits_static_pm_bits = dtlb_ld_tlb_ld_io_requestor_1_resp_bits_static_pm_bits; // @[MemBlock.scala 245:{24,24}]
  assign LoadUnit_1_io_pmp_ld = PMPChecker_1_io_resp_ld; // @[MemBlock.scala 314:{26,26}]
  assign LoadUnit_1_io_pmp_mmio = PMPChecker_1_io_resp_mmio; // @[MemBlock.scala 314:{26,26}]
  assign LoadUnit_1_io_fastpathIn_data = LoadUnit_1_io_fastpathOut_valid ? LoadUnit_1_io_fastpathOut_data :
    LoadUnit_0_io_fastpathOut_data; // @[ParallelMux.scala 90:77]
  assign LoadUnit_1_io_fastpathIn_valid = |_LoadUnit_1_io_fastpathIn_valid_T; // @[MemBlock.scala 391:70]
  assign LoadUnit_1_io_loadFastMatch = LoadUnit_1_io_fastpathOut_valid ? fastMatchVec_0_1 : fastMatchVec_1_1; // @[ParallelMux.scala 90:77]
  assign LoadUnit_1_io_loadFastImm = io_loadFastImm_1; // @[MemBlock.scala 395:33]
  assign LoadUnit_1_io_csrCtrl_ldld_vio_check_enable = csrCtrl_delay_io_out_ldld_vio_check_enable; // @[MemBlock.scala 359:35]
  assign LoadUnit_1_io_csrCtrl_cache_error_enable = csrCtrl_delay_io_out_cache_error_enable; // @[MemBlock.scala 359:35]
  assign LoadUnit_1_io_correctTableQuery_resp_strict = correctTable_io_issue_1_resp_strict; // @[MemBlock.scala 367:39]
  assign LoadUnit_1_io_reExecuteQuery_0_valid = StoreUnit_0_io_reExecuteQuery_valid; // @[MemBlock.scala 371:41]
  assign LoadUnit_1_io_reExecuteQuery_0_bits_robIdx_flag = StoreUnit_0_io_reExecuteQuery_bits_robIdx_flag; // @[MemBlock.scala 371:41]
  assign LoadUnit_1_io_reExecuteQuery_0_bits_robIdx_value = StoreUnit_0_io_reExecuteQuery_bits_robIdx_value; // @[MemBlock.scala 371:41]
  assign LoadUnit_1_io_reExecuteQuery_0_bits_paddr = StoreUnit_0_io_reExecuteQuery_bits_paddr; // @[MemBlock.scala 371:41]
  assign LoadUnit_1_io_reExecuteQuery_0_bits_mask = StoreUnit_0_io_reExecuteQuery_bits_mask; // @[MemBlock.scala 371:41]
  assign LoadUnit_1_io_reExecuteQuery_1_valid = StoreUnit_1_io_reExecuteQuery_valid; // @[MemBlock.scala 371:41]
  assign LoadUnit_1_io_reExecuteQuery_1_bits_robIdx_flag = StoreUnit_1_io_reExecuteQuery_bits_robIdx_flag; // @[MemBlock.scala 371:41]
  assign LoadUnit_1_io_reExecuteQuery_1_bits_robIdx_value = StoreUnit_1_io_reExecuteQuery_bits_robIdx_value; // @[MemBlock.scala 371:41]
  assign LoadUnit_1_io_reExecuteQuery_1_bits_paddr = StoreUnit_1_io_reExecuteQuery_bits_paddr; // @[MemBlock.scala 371:41]
  assign LoadUnit_1_io_reExecuteQuery_1_bits_mask = StoreUnit_1_io_reExecuteQuery_bits_mask; // @[MemBlock.scala 371:41]
  assign LoadUnit_1_io_replay_valid = lsq_io_replay_1_valid; // @[MemBlock.scala 396:28]
  assign LoadUnit_1_io_replay_bits_uop_cf_foldpc = lsq_io_replay_1_bits_uop_cf_foldpc; // @[MemBlock.scala 396:28]
  assign LoadUnit_1_io_replay_bits_uop_cf_trigger_backendEn_1 = lsq_io_replay_1_bits_uop_cf_trigger_backendEn_1; // @[MemBlock.scala 396:28]
  assign LoadUnit_1_io_replay_bits_uop_cf_trigger_backendHit_0 = lsq_io_replay_1_bits_uop_cf_trigger_backendHit_0; // @[MemBlock.scala 396:28]
  assign LoadUnit_1_io_replay_bits_uop_cf_trigger_backendHit_1 = lsq_io_replay_1_bits_uop_cf_trigger_backendHit_1; // @[MemBlock.scala 396:28]
  assign LoadUnit_1_io_replay_bits_uop_cf_trigger_backendHit_4 = lsq_io_replay_1_bits_uop_cf_trigger_backendHit_4; // @[MemBlock.scala 396:28]
  assign LoadUnit_1_io_replay_bits_uop_cf_waitForRobIdx_flag = lsq_io_replay_1_bits_uop_cf_waitForRobIdx_flag; // @[MemBlock.scala 396:28]
  assign LoadUnit_1_io_replay_bits_uop_cf_waitForRobIdx_value = lsq_io_replay_1_bits_uop_cf_waitForRobIdx_value; // @[MemBlock.scala 396:28]
  assign LoadUnit_1_io_replay_bits_uop_cf_loadWaitBit = lsq_io_replay_1_bits_uop_cf_loadWaitBit; // @[MemBlock.scala 396:28]
  assign LoadUnit_1_io_replay_bits_uop_cf_loadWaitStrict = lsq_io_replay_1_bits_uop_cf_loadWaitStrict; // @[MemBlock.scala 396:28]
  assign LoadUnit_1_io_replay_bits_uop_cf_ftqPtr_flag = lsq_io_replay_1_bits_uop_cf_ftqPtr_flag; // @[MemBlock.scala 396:28]
  assign LoadUnit_1_io_replay_bits_uop_cf_ftqPtr_value = lsq_io_replay_1_bits_uop_cf_ftqPtr_value; // @[MemBlock.scala 396:28]
  assign LoadUnit_1_io_replay_bits_uop_cf_ftqOffset = lsq_io_replay_1_bits_uop_cf_ftqOffset; // @[MemBlock.scala 396:28]
  assign LoadUnit_1_io_replay_bits_uop_ctrl_fuType = lsq_io_replay_1_bits_uop_ctrl_fuType; // @[MemBlock.scala 396:28]
  assign LoadUnit_1_io_replay_bits_uop_ctrl_fuOpType = lsq_io_replay_1_bits_uop_ctrl_fuOpType; // @[MemBlock.scala 396:28]
  assign LoadUnit_1_io_replay_bits_uop_ctrl_rfWen = lsq_io_replay_1_bits_uop_ctrl_rfWen; // @[MemBlock.scala 396:28]
  assign LoadUnit_1_io_replay_bits_uop_ctrl_fpWen = lsq_io_replay_1_bits_uop_ctrl_fpWen; // @[MemBlock.scala 396:28]
  assign LoadUnit_1_io_replay_bits_uop_pdest = lsq_io_replay_1_bits_uop_pdest; // @[MemBlock.scala 396:28]
  assign LoadUnit_1_io_replay_bits_uop_robIdx_flag = lsq_io_replay_1_bits_uop_robIdx_flag; // @[MemBlock.scala 396:28]
  assign LoadUnit_1_io_replay_bits_uop_robIdx_value = lsq_io_replay_1_bits_uop_robIdx_value; // @[MemBlock.scala 396:28]
  assign LoadUnit_1_io_replay_bits_uop_lqIdx_flag = lsq_io_replay_1_bits_uop_lqIdx_flag; // @[MemBlock.scala 396:28]
  assign LoadUnit_1_io_replay_bits_uop_lqIdx_value = lsq_io_replay_1_bits_uop_lqIdx_value; // @[MemBlock.scala 396:28]
  assign LoadUnit_1_io_replay_bits_uop_sqIdx_flag = lsq_io_replay_1_bits_uop_sqIdx_flag; // @[MemBlock.scala 396:28]
  assign LoadUnit_1_io_replay_bits_uop_sqIdx_value = lsq_io_replay_1_bits_uop_sqIdx_value; // @[MemBlock.scala 396:28]
  assign LoadUnit_1_io_replay_bits_vaddr = lsq_io_replay_1_bits_vaddr; // @[MemBlock.scala 396:28]
  assign LoadUnit_1_io_replay_bits_isFirstIssue = lsq_io_replay_1_bits_isFirstIssue; // @[MemBlock.scala 396:28]
  assign LoadUnit_1_io_replay_bits_replayCarry_real_way_en = lsq_io_replay_1_bits_replayCarry_real_way_en; // @[MemBlock.scala 396:28]
  assign LoadUnit_1_io_replay_bits_replayCarry_valid = lsq_io_replay_1_bits_replayCarry_valid; // @[MemBlock.scala 396:28]
  assign LoadUnit_1_io_replay_bits_mshrid = lsq_io_replay_1_bits_mshrid; // @[MemBlock.scala 396:28]
  assign LoadUnit_1_io_replay_bits_forward_tlDchannel = lsq_io_replay_1_bits_forward_tlDchannel; // @[MemBlock.scala 396:28]
  assign LoadUnit_1_io_replay_bits_rarAllocated = lsq_io_replay_1_bits_rarAllocated; // @[MemBlock.scala 396:28]
  assign LoadUnit_1_io_replay_bits_rarIndex = lsq_io_replay_1_bits_rarIndex; // @[MemBlock.scala 396:28]
  assign LoadUnit_1_io_replay_bits_rawAllocated = lsq_io_replay_1_bits_rawAllocated; // @[MemBlock.scala 396:28]
  assign LoadUnit_1_io_replay_bits_rawIndex = lsq_io_replay_1_bits_rawIndex; // @[MemBlock.scala 396:28]
  assign LoadUnit_1_io_lqReplayFull = lsq_io_lqReplayFull; // @[MemBlock.scala 373:34]
  assign StoreUnit_0_clock = clock;
  assign StoreUnit_0_reset = reset;
  assign StoreUnit_0_io_stin_valid = st_atomics_0 ? 1'h0 : io_issue_2_valid; // @[MemBlock.scala 460:25 602:63 604:33]
  assign StoreUnit_0_io_stin_bits_uop_cf_trigger_backendEn_0 = io_issue_2_bits_uop_cf_trigger_backendEn_0; // @[MemBlock.scala 460:25]
  assign StoreUnit_0_io_stin_bits_uop_cf_storeSetHit = io_issue_2_bits_uop_cf_storeSetHit; // @[MemBlock.scala 460:25]
  assign StoreUnit_0_io_stin_bits_uop_cf_ssid = io_issue_2_bits_uop_cf_ssid; // @[MemBlock.scala 460:25]
  assign StoreUnit_0_io_stin_bits_uop_cf_ftqPtr_value = io_issue_2_bits_uop_cf_ftqPtr_value; // @[MemBlock.scala 460:25]
  assign StoreUnit_0_io_stin_bits_uop_cf_ftqOffset = io_issue_2_bits_uop_cf_ftqOffset; // @[MemBlock.scala 460:25]
  assign StoreUnit_0_io_stin_bits_uop_ctrl_fuOpType = io_issue_2_bits_uop_ctrl_fuOpType; // @[MemBlock.scala 460:25]
  assign StoreUnit_0_io_stin_bits_uop_ctrl_imm = io_issue_2_bits_uop_ctrl_imm; // @[MemBlock.scala 460:25]
  assign StoreUnit_0_io_stin_bits_uop_robIdx_flag = io_issue_2_bits_uop_robIdx_flag; // @[MemBlock.scala 460:25]
  assign StoreUnit_0_io_stin_bits_uop_robIdx_value = io_issue_2_bits_uop_robIdx_value; // @[MemBlock.scala 460:25]
  assign StoreUnit_0_io_stin_bits_uop_sqIdx_flag = io_issue_2_bits_uop_sqIdx_flag; // @[MemBlock.scala 460:25]
  assign StoreUnit_0_io_stin_bits_uop_sqIdx_value = io_issue_2_bits_uop_sqIdx_value; // @[MemBlock.scala 460:25]
  assign StoreUnit_0_io_stin_bits_src_0 = io_issue_2_bits_src_0; // @[MemBlock.scala 460:25]
  assign StoreUnit_0_io_redirect_valid = redirect_next_valid_REG; // @[BitUtils.scala 26:20 28:18]
  assign StoreUnit_0_io_redirect_bits_robIdx_flag = redirect_next_bits_rrobIdx_flag; // @[BitUtils.scala 26:20 33:15]
  assign StoreUnit_0_io_redirect_bits_robIdx_value = redirect_next_bits_rrobIdx_value; // @[BitUtils.scala 26:20 33:15]
  assign StoreUnit_0_io_redirect_bits_level = redirect_next_bits_rlevel; // @[BitUtils.scala 26:20 33:15]
  assign StoreUnit_0_io_tlb_resp_bits_paddr_0 = dtlb_st_tlb_st_io_requestor_0_resp_bits_paddr_0; // @[MemBlock.scala 249:{24,24}]
  assign StoreUnit_0_io_tlb_resp_bits_miss = dtlb_st_tlb_st_io_requestor_0_resp_bits_miss; // @[MemBlock.scala 249:{24,24}]
  assign StoreUnit_0_io_tlb_resp_bits_excp_0_pf_st = dtlb_st_tlb_st_io_requestor_0_resp_bits_excp_0_pf_st; // @[MemBlock.scala 249:{24,24}]
  assign StoreUnit_0_io_tlb_resp_bits_excp_0_af_st = dtlb_st_tlb_st_io_requestor_0_resp_bits_excp_0_af_st; // @[MemBlock.scala 249:{24,24}]
  assign StoreUnit_0_io_tlb_resp_bits_static_pm_valid = dtlb_st_tlb_st_io_requestor_0_resp_bits_static_pm_valid; // @[MemBlock.scala 249:{24,24}]
  assign StoreUnit_0_io_tlb_resp_bits_static_pm_bits = dtlb_st_tlb_st_io_requestor_0_resp_bits_static_pm_bits; // @[MemBlock.scala 249:{24,24}]
  assign StoreUnit_0_io_pmp_st = PMPChecker_2_io_resp_st; // @[MemBlock.scala 314:{26,26}]
  assign StoreUnit_0_io_pmp_mmio = PMPChecker_2_io_resp_mmio; // @[MemBlock.scala 314:{26,26}]
  assign StoreUnit_0_io_pmp_atomic = PMPChecker_2_io_resp_atomic; // @[MemBlock.scala 314:{26,26}]
  assign StoreUnit_0_io_rsIdx = io_rsfeedback_0_rsIdx; // @[MemBlock.scala 457:25]
  assign StoreUnit_1_clock = clock;
  assign StoreUnit_1_reset = reset;
  assign StoreUnit_1_io_stin_valid = st_atomics_1 ? 1'h0 : io_issue_3_valid; // @[MemBlock.scala 460:25 602:63 604:33]
  assign StoreUnit_1_io_stin_bits_uop_cf_trigger_backendEn_0 = io_issue_3_bits_uop_cf_trigger_backendEn_0; // @[MemBlock.scala 460:25]
  assign StoreUnit_1_io_stin_bits_uop_cf_storeSetHit = io_issue_3_bits_uop_cf_storeSetHit; // @[MemBlock.scala 460:25]
  assign StoreUnit_1_io_stin_bits_uop_cf_ssid = io_issue_3_bits_uop_cf_ssid; // @[MemBlock.scala 460:25]
  assign StoreUnit_1_io_stin_bits_uop_cf_ftqPtr_value = io_issue_3_bits_uop_cf_ftqPtr_value; // @[MemBlock.scala 460:25]
  assign StoreUnit_1_io_stin_bits_uop_cf_ftqOffset = io_issue_3_bits_uop_cf_ftqOffset; // @[MemBlock.scala 460:25]
  assign StoreUnit_1_io_stin_bits_uop_ctrl_fuOpType = io_issue_3_bits_uop_ctrl_fuOpType; // @[MemBlock.scala 460:25]
  assign StoreUnit_1_io_stin_bits_uop_ctrl_imm = io_issue_3_bits_uop_ctrl_imm; // @[MemBlock.scala 460:25]
  assign StoreUnit_1_io_stin_bits_uop_robIdx_flag = io_issue_3_bits_uop_robIdx_flag; // @[MemBlock.scala 460:25]
  assign StoreUnit_1_io_stin_bits_uop_robIdx_value = io_issue_3_bits_uop_robIdx_value; // @[MemBlock.scala 460:25]
  assign StoreUnit_1_io_stin_bits_uop_sqIdx_flag = io_issue_3_bits_uop_sqIdx_flag; // @[MemBlock.scala 460:25]
  assign StoreUnit_1_io_stin_bits_uop_sqIdx_value = io_issue_3_bits_uop_sqIdx_value; // @[MemBlock.scala 460:25]
  assign StoreUnit_1_io_stin_bits_src_0 = io_issue_3_bits_src_0; // @[MemBlock.scala 460:25]
  assign StoreUnit_1_io_redirect_valid = redirect_next_valid_REG; // @[BitUtils.scala 26:20 28:18]
  assign StoreUnit_1_io_redirect_bits_robIdx_flag = redirect_next_bits_rrobIdx_flag; // @[BitUtils.scala 26:20 33:15]
  assign StoreUnit_1_io_redirect_bits_robIdx_value = redirect_next_bits_rrobIdx_value; // @[BitUtils.scala 26:20 33:15]
  assign StoreUnit_1_io_redirect_bits_level = redirect_next_bits_rlevel; // @[BitUtils.scala 26:20 33:15]
  assign StoreUnit_1_io_tlb_resp_bits_paddr_0 = dtlb_st_tlb_st_io_requestor_1_resp_bits_paddr_0; // @[MemBlock.scala 249:{24,24}]
  assign StoreUnit_1_io_tlb_resp_bits_miss = dtlb_st_tlb_st_io_requestor_1_resp_bits_miss; // @[MemBlock.scala 249:{24,24}]
  assign StoreUnit_1_io_tlb_resp_bits_excp_0_pf_st = dtlb_st_tlb_st_io_requestor_1_resp_bits_excp_0_pf_st; // @[MemBlock.scala 249:{24,24}]
  assign StoreUnit_1_io_tlb_resp_bits_excp_0_af_st = dtlb_st_tlb_st_io_requestor_1_resp_bits_excp_0_af_st; // @[MemBlock.scala 249:{24,24}]
  assign StoreUnit_1_io_tlb_resp_bits_static_pm_valid = dtlb_st_tlb_st_io_requestor_1_resp_bits_static_pm_valid; // @[MemBlock.scala 249:{24,24}]
  assign StoreUnit_1_io_tlb_resp_bits_static_pm_bits = dtlb_st_tlb_st_io_requestor_1_resp_bits_static_pm_bits; // @[MemBlock.scala 249:{24,24}]
  assign StoreUnit_1_io_pmp_st = PMPChecker_3_io_resp_st; // @[MemBlock.scala 314:{26,26}]
  assign StoreUnit_1_io_pmp_mmio = PMPChecker_3_io_resp_mmio; // @[MemBlock.scala 314:{26,26}]
  assign StoreUnit_1_io_pmp_atomic = PMPChecker_3_io_resp_atomic; // @[MemBlock.scala 314:{26,26}]
  assign StoreUnit_1_io_rsIdx = io_rsfeedback_1_rsIdx; // @[MemBlock.scala 457:25]
  assign stdExeUnits_0_io_fromInt_valid = io_issue_4_valid; // @[MemBlock.scala 451:31]
  assign stdExeUnits_0_io_fromInt_bits_uop_ctrl_fuType = io_issue_4_bits_uop_ctrl_fuType; // @[MemBlock.scala 451:31]
  assign stdExeUnits_0_io_fromInt_bits_uop_ctrl_fuOpType = io_issue_4_bits_uop_ctrl_fuOpType; // @[MemBlock.scala 451:31]
  assign stdExeUnits_0_io_fromInt_bits_uop_robIdx_flag = io_issue_4_bits_uop_robIdx_flag; // @[MemBlock.scala 451:31]
  assign stdExeUnits_0_io_fromInt_bits_uop_robIdx_value = io_issue_4_bits_uop_robIdx_value; // @[MemBlock.scala 451:31]
  assign stdExeUnits_0_io_fromInt_bits_uop_sqIdx_flag = io_issue_4_bits_uop_sqIdx_flag; // @[MemBlock.scala 451:31]
  assign stdExeUnits_0_io_fromInt_bits_uop_sqIdx_value = io_issue_4_bits_uop_sqIdx_value; // @[MemBlock.scala 451:31]
  assign stdExeUnits_0_io_fromInt_bits_src_0 = io_issue_4_bits_src_0; // @[MemBlock.scala 451:31]
  assign stdExeUnits_1_io_fromInt_valid = io_issue_5_valid; // @[MemBlock.scala 451:31]
  assign stdExeUnits_1_io_fromInt_bits_uop_ctrl_fuType = io_issue_5_bits_uop_ctrl_fuType; // @[MemBlock.scala 451:31]
  assign stdExeUnits_1_io_fromInt_bits_uop_ctrl_fuOpType = io_issue_5_bits_uop_ctrl_fuOpType; // @[MemBlock.scala 451:31]
  assign stdExeUnits_1_io_fromInt_bits_uop_robIdx_flag = io_issue_5_bits_uop_robIdx_flag; // @[MemBlock.scala 451:31]
  assign stdExeUnits_1_io_fromInt_bits_uop_robIdx_value = io_issue_5_bits_uop_robIdx_value; // @[MemBlock.scala 451:31]
  assign stdExeUnits_1_io_fromInt_bits_uop_sqIdx_flag = io_issue_5_bits_uop_sqIdx_flag; // @[MemBlock.scala 451:31]
  assign stdExeUnits_1_io_fromInt_bits_uop_sqIdx_value = io_issue_5_bits_uop_sqIdx_value; // @[MemBlock.scala 451:31]
  assign stdExeUnits_1_io_fromInt_bits_src_0 = io_issue_5_bits_src_0; // @[MemBlock.scala 451:31]
  assign correctTable_clock = clock;
  assign correctTable_io_issue_0_req_addr = LoadUnit_0_io_correctTableQuery_req_addr; // @[MemBlock.scala 367:39]
  assign correctTable_io_issue_1_req_addr = LoadUnit_1_io_correctTableQuery_req_addr; // @[MemBlock.scala 367:39]
  assign correctTable_io_update_0_valid = LoadUnit_0_io_correctTableUpdate_valid; // @[MemBlock.scala 368:40]
  assign correctTable_io_update_0_bits_addr = LoadUnit_0_io_correctTableUpdate_bits_addr; // @[MemBlock.scala 368:40]
  assign correctTable_io_update_0_bits_strict = LoadUnit_0_io_correctTableUpdate_bits_strict; // @[MemBlock.scala 368:40]
  assign correctTable_io_update_0_bits_violation = LoadUnit_0_io_correctTableUpdate_bits_violation; // @[MemBlock.scala 368:40]
  assign correctTable_io_update_1_valid = LoadUnit_1_io_correctTableUpdate_valid; // @[MemBlock.scala 368:40]
  assign correctTable_io_update_1_bits_addr = LoadUnit_1_io_correctTableUpdate_bits_addr; // @[MemBlock.scala 368:40]
  assign correctTable_io_update_1_bits_strict = LoadUnit_1_io_correctTableUpdate_bits_strict; // @[MemBlock.scala 368:40]
  assign correctTable_io_update_1_bits_violation = LoadUnit_1_io_correctTableUpdate_bits_violation; // @[MemBlock.scala 368:40]
  assign correctTable_io_update_2_valid = lsq_io_correctTableUpdate_valid; // @[MemBlock.scala 542:29]
  assign correctTable_io_update_2_bits_addr = lsq_io_correctTableUpdate_bits_addr; // @[MemBlock.scala 542:29]
  assign atomicsUnit_clock = clock;
  assign atomicsUnit_reset = reset;
  assign atomicsUnit_io_hartId = io_hartId; // @[MemBlock.scala 240:25]
  assign atomicsUnit_io_in_valid = st_atomics_0 | st_atomics_1; // @[MemBlock.scala 615:50]
  assign atomicsUnit_io_in_bits_uop_cf_trigger_backendEn_0 = st_atomics_0 & io_issue_2_bits_uop_cf_trigger_backendEn_0
     | st_atomics_1 & io_issue_3_bits_uop_cf_trigger_backendEn_0; // @[Mux.scala 27:73]
  assign atomicsUnit_io_in_bits_uop_cf_trigger_backendEn_1 = st_atomics_0 & io_issue_2_bits_uop_cf_trigger_backendEn_1
     | st_atomics_1 & io_issue_3_bits_uop_cf_trigger_backendEn_1; // @[Mux.scala 27:73]
  assign atomicsUnit_io_in_bits_uop_ctrl_fuOpType = _atomicsUnit_io_in_bits_T_162 | _atomicsUnit_io_in_bits_T_163; // @[Mux.scala 27:73]
  assign atomicsUnit_io_in_bits_uop_ctrl_rfWen = st_atomics_0 & io_issue_2_bits_uop_ctrl_rfWen | st_atomics_1 &
    io_issue_3_bits_uop_ctrl_rfWen; // @[Mux.scala 27:73]
  assign atomicsUnit_io_in_bits_uop_ctrl_fpWen = st_atomics_0 & io_issue_2_bits_uop_ctrl_fpWen | st_atomics_1 &
    io_issue_3_bits_uop_ctrl_fpWen; // @[Mux.scala 27:73]
  assign atomicsUnit_io_in_bits_uop_pdest = _atomicsUnit_io_in_bits_T_63 | _atomicsUnit_io_in_bits_T_64; // @[Mux.scala 27:73]
  assign atomicsUnit_io_in_bits_uop_robIdx_flag = st_atomics_0 & io_issue_2_bits_uop_robIdx_flag | st_atomics_1 &
    io_issue_3_bits_uop_robIdx_flag; // @[Mux.scala 27:73]
  assign atomicsUnit_io_in_bits_uop_robIdx_value = _atomicsUnit_io_in_bits_T_54 | _atomicsUnit_io_in_bits_T_55; // @[Mux.scala 27:73]
  assign atomicsUnit_io_in_bits_src_0 = _atomicsUnit_io_in_bits_T | _atomicsUnit_io_in_bits_T_1; // @[Mux.scala 27:73]
  assign atomicsUnit_io_storeDataIn_valid = st_data_atomics_0 | st_data_atomics_1; // @[MemBlock.scala 618:64]
  assign atomicsUnit_io_storeDataIn_bits_data = _atomicsUnit_io_storeDataIn_bits_T_243 |
    _atomicsUnit_io_storeDataIn_bits_T_244; // @[Mux.scala 27:73]
  assign atomicsUnit_io_dcache_req_ready = dcache_io_lsu_atomics_req_ready; // @[MemBlock.scala 632:25]
  assign atomicsUnit_io_dcache_resp_valid = dcache_io_lsu_atomics_resp_valid; // @[MemBlock.scala 632:25]
  assign atomicsUnit_io_dcache_resp_bits_data = dcache_io_lsu_atomics_resp_bits_data; // @[MemBlock.scala 632:25]
  assign atomicsUnit_io_dcache_resp_bits_miss = dcache_io_lsu_atomics_resp_bits_miss; // @[MemBlock.scala 632:25]
  assign atomicsUnit_io_dcache_resp_bits_replay = dcache_io_lsu_atomics_resp_bits_replay; // @[MemBlock.scala 632:25]
  assign atomicsUnit_io_dcache_resp_bits_error = dcache_io_lsu_atomics_resp_bits_error; // @[MemBlock.scala 632:25]
  assign atomicsUnit_io_dcache_resp_bits_id = dcache_io_lsu_atomics_resp_bits_id; // @[MemBlock.scala 632:25]
  assign atomicsUnit_io_dcache_block_lr = dcache_io_lsu_atomics_block_lr; // @[MemBlock.scala 632:25]
  assign atomicsUnit_io_dtlb_resp_valid = state != 2'h0 & dtlb_ld_0_requestor_0_resp_valid; // @[MemBlock.scala 639:29 643:25 627:34]
  assign atomicsUnit_io_dtlb_resp_bits_paddr_0 = dtlb_ld_tlb_ld_io_requestor_0_resp_bits_paddr_0; // @[MemBlock.scala 245:{24,24}]
  assign atomicsUnit_io_dtlb_resp_bits_miss = dtlb_ld_tlb_ld_io_requestor_0_resp_bits_miss; // @[MemBlock.scala 245:{24,24}]
  assign atomicsUnit_io_dtlb_resp_bits_excp_0_pf_ld = dtlb_ld_tlb_ld_io_requestor_0_resp_bits_excp_0_pf_ld; // @[MemBlock.scala 245:{24,24}]
  assign atomicsUnit_io_dtlb_resp_bits_excp_0_pf_st = dtlb_ld_tlb_ld_io_requestor_0_resp_bits_excp_0_pf_st; // @[MemBlock.scala 245:{24,24}]
  assign atomicsUnit_io_dtlb_resp_bits_excp_0_af_ld = dtlb_ld_tlb_ld_io_requestor_0_resp_bits_excp_0_af_ld; // @[MemBlock.scala 245:{24,24}]
  assign atomicsUnit_io_dtlb_resp_bits_excp_0_af_st = dtlb_ld_tlb_ld_io_requestor_0_resp_bits_excp_0_af_st; // @[MemBlock.scala 245:{24,24}]
  assign atomicsUnit_io_dtlb_resp_bits_static_pm_valid = dtlb_ld_tlb_ld_io_requestor_0_resp_bits_static_pm_valid; // @[MemBlock.scala 245:{24,24}]
  assign atomicsUnit_io_dtlb_resp_bits_static_pm_bits = dtlb_ld_tlb_ld_io_requestor_0_resp_bits_static_pm_bits; // @[MemBlock.scala 245:{24,24}]
  assign atomicsUnit_io_pmpResp_ld = PMPChecker_io_resp_ld; // @[MemBlock.scala 314:{26,26}]
  assign atomicsUnit_io_pmpResp_st = PMPChecker_io_resp_st; // @[MemBlock.scala 314:{26,26}]
  assign atomicsUnit_io_pmpResp_mmio = PMPChecker_io_resp_mmio; // @[MemBlock.scala 314:{26,26}]
  assign atomicsUnit_io_rsIdx = _atomicsUnit_io_rsIdx_T | _atomicsUnit_io_rsIdx_T_1; // @[Mux.scala 27:73]
  assign atomicsUnit_io_flush_sbuffer_empty = sbuffer_io_flush_empty & uncache_io_flush_empty; // @[MemBlock.scala 566:42]
  assign atomicsUnit_io_redirect_valid = redirect_next_valid_REG; // @[BitUtils.scala 26:20 28:18]
  assign atomicsUnit_io_csrCtrl_cache_error_enable = csrCtrl_delay_io_out_cache_error_enable; // @[MemBlock.scala 635:26]
  assign atomicsUnit_io_csrCtrl_mem_trigger_t_valid = csrCtrl_delay_io_out_mem_trigger_t_valid; // @[MemBlock.scala 635:26]
  assign atomicsUnit_io_csrCtrl_mem_trigger_t_bits_addr = csrCtrl_delay_io_out_mem_trigger_t_bits_addr; // @[MemBlock.scala 635:26]
  assign atomicsUnit_io_csrCtrl_mem_trigger_t_bits_tdata_matchType =
    csrCtrl_delay_io_out_mem_trigger_t_bits_tdata_matchType; // @[MemBlock.scala 635:26]
  assign atomicsUnit_io_csrCtrl_mem_trigger_t_bits_tdata_select = csrCtrl_delay_io_out_mem_trigger_t_bits_tdata_select; // @[MemBlock.scala 635:26]
  assign atomicsUnit_io_csrCtrl_mem_trigger_t_bits_tdata_chain = csrCtrl_delay_io_out_mem_trigger_t_bits_tdata_chain; // @[MemBlock.scala 635:26]
  assign atomicsUnit_io_csrCtrl_mem_trigger_t_bits_tdata_tdata2 = csrCtrl_delay_io_out_mem_trigger_t_bits_tdata_tdata2; // @[MemBlock.scala 635:26]
  assign atomicsUnit_io_csrCtrl_trigger_enable_2 = csrCtrl_delay_io_out_trigger_enable_2; // @[MemBlock.scala 635:26]
  assign atomicsUnit_io_csrCtrl_trigger_enable_3 = csrCtrl_delay_io_out_trigger_enable_3; // @[MemBlock.scala 635:26]
  assign atomicsUnit_io_csrCtrl_trigger_enable_4 = csrCtrl_delay_io_out_trigger_enable_4; // @[MemBlock.scala 635:26]
  assign atomicsUnit_io_csrCtrl_trigger_enable_5 = csrCtrl_delay_io_out_trigger_enable_5; // @[MemBlock.scala 635:26]
  assign atomicsUnit_io_csrCtrl_trigger_enable_7 = csrCtrl_delay_io_out_trigger_enable_7; // @[MemBlock.scala 635:26]
  assign atomicsUnit_io_csrCtrl_trigger_enable_9 = csrCtrl_delay_io_out_trigger_enable_9; // @[MemBlock.scala 635:26]
  assign vlflowqueue_clock = clock;
  assign vlflowqueue_reset = reset;
  assign vlflowqueue_io_loadRegIn_0_valid = vlExcSignal_io_vecloadRegIn_0_valid; // @[MemBlock.scala 577:28]
  assign vlflowqueue_io_loadRegIn_0_bits_uop_robIdx_value = vlExcSignal_io_vecloadRegIn_0_bits_uop_robIdx_value; // @[MemBlock.scala 577:28]
  assign vlflowqueue_io_loadRegIn_0_bits_baseaddr = vlExcSignal_io_vecloadRegIn_0_bits_baseaddr; // @[MemBlock.scala 577:28]
  assign vlflowqueue_io_loadRegIn_1_valid = vlExcSignal_io_vecloadRegIn_1_valid; // @[MemBlock.scala 577:28]
  assign vlflowqueue_io_loadRegIn_1_bits_uop_robIdx_value = vlExcSignal_io_vecloadRegIn_1_bits_uop_robIdx_value; // @[MemBlock.scala 577:28]
  assign vlflowqueue_io_loadRegIn_1_bits_baseaddr = vlExcSignal_io_vecloadRegIn_1_bits_baseaddr; // @[MemBlock.scala 577:28]
  assign vlflowqueue_io_loadPipeOut_0_ready = LoadUnit_0_io_VecloadIn_ready; // @[MemBlock.scala 346:31]
  assign vlflowqueue_io_loadPipeOut_1_ready = LoadUnit_1_io_VecloadIn_ready; // @[MemBlock.scala 346:31]
  assign vlExcSignal_clock = clock;
  assign vlExcSignal_reset = reset;
  assign lsq_clock = clock;
  assign lsq_reset = reset;
  assign lsq_io_brqRedirect_valid = redirect_next_valid_REG; // @[BitUtils.scala 26:20 28:18]
  assign lsq_io_brqRedirect_bits_robIdx_flag = redirect_next_bits_rrobIdx_flag; // @[BitUtils.scala 26:20 33:15]
  assign lsq_io_brqRedirect_bits_robIdx_value = redirect_next_bits_rrobIdx_value; // @[BitUtils.scala 26:20 33:15]
  assign lsq_io_brqRedirect_bits_level = redirect_next_bits_rlevel; // @[BitUtils.scala 26:20 33:15]
  assign lsq_io_enq_needAlloc_0 = io_enqLsq_needAlloc_0; // @[MemBlock.scala 540:25]
  assign lsq_io_enq_needAlloc_1 = io_enqLsq_needAlloc_1; // @[MemBlock.scala 540:25]
  assign lsq_io_enq_needAlloc_2 = io_enqLsq_needAlloc_2; // @[MemBlock.scala 540:25]
  assign lsq_io_enq_needAlloc_3 = io_enqLsq_needAlloc_3; // @[MemBlock.scala 540:25]
  assign lsq_io_enq_req_0_valid = io_enqLsq_req_0_valid; // @[MemBlock.scala 540:25]
  assign lsq_io_enq_req_0_bits_cf_trigger_backendEn_0 = io_enqLsq_req_0_bits_cf_trigger_backendEn_0; // @[MemBlock.scala 540:25]
  assign lsq_io_enq_req_0_bits_cf_trigger_backendEn_1 = io_enqLsq_req_0_bits_cf_trigger_backendEn_1; // @[MemBlock.scala 540:25]
  assign lsq_io_enq_req_0_bits_ctrl_fuOpType = io_enqLsq_req_0_bits_ctrl_fuOpType; // @[MemBlock.scala 540:25]
  assign lsq_io_enq_req_0_bits_ctrl_rfWen = io_enqLsq_req_0_bits_ctrl_rfWen; // @[MemBlock.scala 540:25]
  assign lsq_io_enq_req_0_bits_ctrl_fpWen = io_enqLsq_req_0_bits_ctrl_fpWen; // @[MemBlock.scala 540:25]
  assign lsq_io_enq_req_0_bits_ctrl_flushPipe = io_enqLsq_req_0_bits_ctrl_flushPipe; // @[MemBlock.scala 540:25]
  assign lsq_io_enq_req_0_bits_ctrl_replayInst = io_enqLsq_req_0_bits_ctrl_replayInst; // @[MemBlock.scala 540:25]
  assign lsq_io_enq_req_0_bits_pdest = io_enqLsq_req_0_bits_pdest; // @[MemBlock.scala 540:25]
  assign lsq_io_enq_req_0_bits_robIdx_flag = io_enqLsq_req_0_bits_robIdx_flag; // @[MemBlock.scala 540:25]
  assign lsq_io_enq_req_0_bits_robIdx_value = io_enqLsq_req_0_bits_robIdx_value; // @[MemBlock.scala 540:25]
  assign lsq_io_enq_req_0_bits_lqIdx_value = io_enqLsq_req_0_bits_lqIdx_value; // @[MemBlock.scala 540:25]
  assign lsq_io_enq_req_0_bits_sqIdx_value = io_enqLsq_req_0_bits_sqIdx_value; // @[MemBlock.scala 540:25]
  assign lsq_io_enq_req_1_valid = io_enqLsq_req_1_valid; // @[MemBlock.scala 540:25]
  assign lsq_io_enq_req_1_bits_cf_trigger_backendEn_0 = io_enqLsq_req_1_bits_cf_trigger_backendEn_0; // @[MemBlock.scala 540:25]
  assign lsq_io_enq_req_1_bits_cf_trigger_backendEn_1 = io_enqLsq_req_1_bits_cf_trigger_backendEn_1; // @[MemBlock.scala 540:25]
  assign lsq_io_enq_req_1_bits_ctrl_fuOpType = io_enqLsq_req_1_bits_ctrl_fuOpType; // @[MemBlock.scala 540:25]
  assign lsq_io_enq_req_1_bits_ctrl_rfWen = io_enqLsq_req_1_bits_ctrl_rfWen; // @[MemBlock.scala 540:25]
  assign lsq_io_enq_req_1_bits_ctrl_fpWen = io_enqLsq_req_1_bits_ctrl_fpWen; // @[MemBlock.scala 540:25]
  assign lsq_io_enq_req_1_bits_ctrl_flushPipe = io_enqLsq_req_1_bits_ctrl_flushPipe; // @[MemBlock.scala 540:25]
  assign lsq_io_enq_req_1_bits_ctrl_replayInst = io_enqLsq_req_1_bits_ctrl_replayInst; // @[MemBlock.scala 540:25]
  assign lsq_io_enq_req_1_bits_pdest = io_enqLsq_req_1_bits_pdest; // @[MemBlock.scala 540:25]
  assign lsq_io_enq_req_1_bits_robIdx_flag = io_enqLsq_req_1_bits_robIdx_flag; // @[MemBlock.scala 540:25]
  assign lsq_io_enq_req_1_bits_robIdx_value = io_enqLsq_req_1_bits_robIdx_value; // @[MemBlock.scala 540:25]
  assign lsq_io_enq_req_1_bits_lqIdx_value = io_enqLsq_req_1_bits_lqIdx_value; // @[MemBlock.scala 540:25]
  assign lsq_io_enq_req_1_bits_sqIdx_value = io_enqLsq_req_1_bits_sqIdx_value; // @[MemBlock.scala 540:25]
  assign lsq_io_enq_req_2_valid = io_enqLsq_req_2_valid; // @[MemBlock.scala 540:25]
  assign lsq_io_enq_req_2_bits_cf_trigger_backendEn_0 = io_enqLsq_req_2_bits_cf_trigger_backendEn_0; // @[MemBlock.scala 540:25]
  assign lsq_io_enq_req_2_bits_cf_trigger_backendEn_1 = io_enqLsq_req_2_bits_cf_trigger_backendEn_1; // @[MemBlock.scala 540:25]
  assign lsq_io_enq_req_2_bits_ctrl_fuOpType = io_enqLsq_req_2_bits_ctrl_fuOpType; // @[MemBlock.scala 540:25]
  assign lsq_io_enq_req_2_bits_ctrl_rfWen = io_enqLsq_req_2_bits_ctrl_rfWen; // @[MemBlock.scala 540:25]
  assign lsq_io_enq_req_2_bits_ctrl_fpWen = io_enqLsq_req_2_bits_ctrl_fpWen; // @[MemBlock.scala 540:25]
  assign lsq_io_enq_req_2_bits_ctrl_flushPipe = io_enqLsq_req_2_bits_ctrl_flushPipe; // @[MemBlock.scala 540:25]
  assign lsq_io_enq_req_2_bits_ctrl_replayInst = io_enqLsq_req_2_bits_ctrl_replayInst; // @[MemBlock.scala 540:25]
  assign lsq_io_enq_req_2_bits_pdest = io_enqLsq_req_2_bits_pdest; // @[MemBlock.scala 540:25]
  assign lsq_io_enq_req_2_bits_robIdx_flag = io_enqLsq_req_2_bits_robIdx_flag; // @[MemBlock.scala 540:25]
  assign lsq_io_enq_req_2_bits_robIdx_value = io_enqLsq_req_2_bits_robIdx_value; // @[MemBlock.scala 540:25]
  assign lsq_io_enq_req_2_bits_lqIdx_value = io_enqLsq_req_2_bits_lqIdx_value; // @[MemBlock.scala 540:25]
  assign lsq_io_enq_req_2_bits_sqIdx_value = io_enqLsq_req_2_bits_sqIdx_value; // @[MemBlock.scala 540:25]
  assign lsq_io_enq_req_3_valid = io_enqLsq_req_3_valid; // @[MemBlock.scala 540:25]
  assign lsq_io_enq_req_3_bits_cf_trigger_backendEn_0 = io_enqLsq_req_3_bits_cf_trigger_backendEn_0; // @[MemBlock.scala 540:25]
  assign lsq_io_enq_req_3_bits_cf_trigger_backendEn_1 = io_enqLsq_req_3_bits_cf_trigger_backendEn_1; // @[MemBlock.scala 540:25]
  assign lsq_io_enq_req_3_bits_ctrl_fuOpType = io_enqLsq_req_3_bits_ctrl_fuOpType; // @[MemBlock.scala 540:25]
  assign lsq_io_enq_req_3_bits_ctrl_rfWen = io_enqLsq_req_3_bits_ctrl_rfWen; // @[MemBlock.scala 540:25]
  assign lsq_io_enq_req_3_bits_ctrl_fpWen = io_enqLsq_req_3_bits_ctrl_fpWen; // @[MemBlock.scala 540:25]
  assign lsq_io_enq_req_3_bits_ctrl_flushPipe = io_enqLsq_req_3_bits_ctrl_flushPipe; // @[MemBlock.scala 540:25]
  assign lsq_io_enq_req_3_bits_ctrl_replayInst = io_enqLsq_req_3_bits_ctrl_replayInst; // @[MemBlock.scala 540:25]
  assign lsq_io_enq_req_3_bits_pdest = io_enqLsq_req_3_bits_pdest; // @[MemBlock.scala 540:25]
  assign lsq_io_enq_req_3_bits_robIdx_flag = io_enqLsq_req_3_bits_robIdx_flag; // @[MemBlock.scala 540:25]
  assign lsq_io_enq_req_3_bits_robIdx_value = io_enqLsq_req_3_bits_robIdx_value; // @[MemBlock.scala 540:25]
  assign lsq_io_enq_req_3_bits_lqIdx_value = io_enqLsq_req_3_bits_lqIdx_value; // @[MemBlock.scala 540:25]
  assign lsq_io_enq_req_3_bits_sqIdx_value = io_enqLsq_req_3_bits_sqIdx_value; // @[MemBlock.scala 540:25]
  assign lsq_io_ldu_s2_storeLoadViolationQuery_0_req_valid = LoadUnit_0_io_lsq_storeLoadViolationQuery_req_valid; // @[MemBlock.scala 358:49]
  assign lsq_io_ldu_s2_storeLoadViolationQuery_0_req_bits_uop_cf_foldpc =
    LoadUnit_0_io_lsq_storeLoadViolationQuery_req_bits_uop_cf_foldpc; // @[MemBlock.scala 358:49]
  assign lsq_io_ldu_s2_storeLoadViolationQuery_0_req_bits_uop_cf_ftqPtr_flag =
    LoadUnit_0_io_lsq_storeLoadViolationQuery_req_bits_uop_cf_ftqPtr_flag; // @[MemBlock.scala 358:49]
  assign lsq_io_ldu_s2_storeLoadViolationQuery_0_req_bits_uop_cf_ftqPtr_value =
    LoadUnit_0_io_lsq_storeLoadViolationQuery_req_bits_uop_cf_ftqPtr_value; // @[MemBlock.scala 358:49]
  assign lsq_io_ldu_s2_storeLoadViolationQuery_0_req_bits_uop_cf_ftqOffset =
    LoadUnit_0_io_lsq_storeLoadViolationQuery_req_bits_uop_cf_ftqOffset; // @[MemBlock.scala 358:49]
  assign lsq_io_ldu_s2_storeLoadViolationQuery_0_req_bits_uop_robIdx_flag =
    LoadUnit_0_io_lsq_storeLoadViolationQuery_req_bits_uop_robIdx_flag; // @[MemBlock.scala 358:49]
  assign lsq_io_ldu_s2_storeLoadViolationQuery_0_req_bits_uop_robIdx_value =
    LoadUnit_0_io_lsq_storeLoadViolationQuery_req_bits_uop_robIdx_value; // @[MemBlock.scala 358:49]
  assign lsq_io_ldu_s2_storeLoadViolationQuery_0_req_bits_uop_sqIdx_flag =
    LoadUnit_0_io_lsq_storeLoadViolationQuery_req_bits_uop_sqIdx_flag; // @[MemBlock.scala 358:49]
  assign lsq_io_ldu_s2_storeLoadViolationQuery_0_req_bits_uop_sqIdx_value =
    LoadUnit_0_io_lsq_storeLoadViolationQuery_req_bits_uop_sqIdx_value; // @[MemBlock.scala 358:49]
  assign lsq_io_ldu_s2_storeLoadViolationQuery_0_req_bits_index =
    LoadUnit_0_io_lsq_storeLoadViolationQuery_req_bits_index; // @[MemBlock.scala 358:49]
  assign lsq_io_ldu_s2_storeLoadViolationQuery_0_req_bits_allocated =
    LoadUnit_0_io_lsq_storeLoadViolationQuery_req_bits_allocated; // @[MemBlock.scala 358:49]
  assign lsq_io_ldu_s2_storeLoadViolationQuery_0_req_bits_datavalid =
    LoadUnit_0_io_lsq_storeLoadViolationQuery_req_bits_datavalid; // @[MemBlock.scala 358:49]
  assign lsq_io_ldu_s2_storeLoadViolationQuery_0_req_bits_mask = LoadUnit_0_io_lsq_storeLoadViolationQuery_req_bits_mask
    ; // @[MemBlock.scala 358:49]
  assign lsq_io_ldu_s2_storeLoadViolationQuery_0_req_bits_paddr =
    LoadUnit_0_io_lsq_storeLoadViolationQuery_req_bits_paddr; // @[MemBlock.scala 358:49]
  assign lsq_io_ldu_s2_storeLoadViolationQuery_1_req_valid = LoadUnit_1_io_lsq_storeLoadViolationQuery_req_valid; // @[MemBlock.scala 358:49]
  assign lsq_io_ldu_s2_storeLoadViolationQuery_1_req_bits_uop_cf_foldpc =
    LoadUnit_1_io_lsq_storeLoadViolationQuery_req_bits_uop_cf_foldpc; // @[MemBlock.scala 358:49]
  assign lsq_io_ldu_s2_storeLoadViolationQuery_1_req_bits_uop_cf_ftqPtr_flag =
    LoadUnit_1_io_lsq_storeLoadViolationQuery_req_bits_uop_cf_ftqPtr_flag; // @[MemBlock.scala 358:49]
  assign lsq_io_ldu_s2_storeLoadViolationQuery_1_req_bits_uop_cf_ftqPtr_value =
    LoadUnit_1_io_lsq_storeLoadViolationQuery_req_bits_uop_cf_ftqPtr_value; // @[MemBlock.scala 358:49]
  assign lsq_io_ldu_s2_storeLoadViolationQuery_1_req_bits_uop_cf_ftqOffset =
    LoadUnit_1_io_lsq_storeLoadViolationQuery_req_bits_uop_cf_ftqOffset; // @[MemBlock.scala 358:49]
  assign lsq_io_ldu_s2_storeLoadViolationQuery_1_req_bits_uop_robIdx_flag =
    LoadUnit_1_io_lsq_storeLoadViolationQuery_req_bits_uop_robIdx_flag; // @[MemBlock.scala 358:49]
  assign lsq_io_ldu_s2_storeLoadViolationQuery_1_req_bits_uop_robIdx_value =
    LoadUnit_1_io_lsq_storeLoadViolationQuery_req_bits_uop_robIdx_value; // @[MemBlock.scala 358:49]
  assign lsq_io_ldu_s2_storeLoadViolationQuery_1_req_bits_uop_sqIdx_flag =
    LoadUnit_1_io_lsq_storeLoadViolationQuery_req_bits_uop_sqIdx_flag; // @[MemBlock.scala 358:49]
  assign lsq_io_ldu_s2_storeLoadViolationQuery_1_req_bits_uop_sqIdx_value =
    LoadUnit_1_io_lsq_storeLoadViolationQuery_req_bits_uop_sqIdx_value; // @[MemBlock.scala 358:49]
  assign lsq_io_ldu_s2_storeLoadViolationQuery_1_req_bits_index =
    LoadUnit_1_io_lsq_storeLoadViolationQuery_req_bits_index; // @[MemBlock.scala 358:49]
  assign lsq_io_ldu_s2_storeLoadViolationQuery_1_req_bits_allocated =
    LoadUnit_1_io_lsq_storeLoadViolationQuery_req_bits_allocated; // @[MemBlock.scala 358:49]
  assign lsq_io_ldu_s2_storeLoadViolationQuery_1_req_bits_datavalid =
    LoadUnit_1_io_lsq_storeLoadViolationQuery_req_bits_datavalid; // @[MemBlock.scala 358:49]
  assign lsq_io_ldu_s2_storeLoadViolationQuery_1_req_bits_mask = LoadUnit_1_io_lsq_storeLoadViolationQuery_req_bits_mask
    ; // @[MemBlock.scala 358:49]
  assign lsq_io_ldu_s2_storeLoadViolationQuery_1_req_bits_paddr =
    LoadUnit_1_io_lsq_storeLoadViolationQuery_req_bits_paddr; // @[MemBlock.scala 358:49]
  assign lsq_io_ldu_s2_loadLoadViolationQuery_0_req_valid = LoadUnit_0_io_lsq_loadLoadViolationQuery_req_valid; // @[MemBlock.scala 357:48]
  assign lsq_io_ldu_s2_loadLoadViolationQuery_0_req_bits_uop_robIdx_flag =
    LoadUnit_0_io_lsq_loadLoadViolationQuery_req_bits_uop_robIdx_flag; // @[MemBlock.scala 357:48]
  assign lsq_io_ldu_s2_loadLoadViolationQuery_0_req_bits_uop_robIdx_value =
    LoadUnit_0_io_lsq_loadLoadViolationQuery_req_bits_uop_robIdx_value; // @[MemBlock.scala 357:48]
  assign lsq_io_ldu_s2_loadLoadViolationQuery_0_req_bits_uop_lqIdx_flag =
    LoadUnit_0_io_lsq_loadLoadViolationQuery_req_bits_uop_lqIdx_flag; // @[MemBlock.scala 357:48]
  assign lsq_io_ldu_s2_loadLoadViolationQuery_0_req_bits_uop_lqIdx_value =
    LoadUnit_0_io_lsq_loadLoadViolationQuery_req_bits_uop_lqIdx_value; // @[MemBlock.scala 357:48]
  assign lsq_io_ldu_s2_loadLoadViolationQuery_0_req_bits_index = LoadUnit_0_io_lsq_loadLoadViolationQuery_req_bits_index
    ; // @[MemBlock.scala 357:48]
  assign lsq_io_ldu_s2_loadLoadViolationQuery_0_req_bits_allocated =
    LoadUnit_0_io_lsq_loadLoadViolationQuery_req_bits_allocated; // @[MemBlock.scala 357:48]
  assign lsq_io_ldu_s2_loadLoadViolationQuery_0_req_bits_datavalid =
    LoadUnit_0_io_lsq_loadLoadViolationQuery_req_bits_datavalid; // @[MemBlock.scala 357:48]
  assign lsq_io_ldu_s2_loadLoadViolationQuery_0_req_bits_miss = LoadUnit_0_io_lsq_loadLoadViolationQuery_req_bits_miss; // @[MemBlock.scala 357:48]
  assign lsq_io_ldu_s2_loadLoadViolationQuery_0_req_bits_paddr = LoadUnit_0_io_lsq_loadLoadViolationQuery_req_bits_paddr
    ; // @[MemBlock.scala 357:48]
  assign lsq_io_ldu_s2_loadLoadViolationQuery_1_req_valid = LoadUnit_1_io_lsq_loadLoadViolationQuery_req_valid; // @[MemBlock.scala 357:48]
  assign lsq_io_ldu_s2_loadLoadViolationQuery_1_req_bits_uop_robIdx_flag =
    LoadUnit_1_io_lsq_loadLoadViolationQuery_req_bits_uop_robIdx_flag; // @[MemBlock.scala 357:48]
  assign lsq_io_ldu_s2_loadLoadViolationQuery_1_req_bits_uop_robIdx_value =
    LoadUnit_1_io_lsq_loadLoadViolationQuery_req_bits_uop_robIdx_value; // @[MemBlock.scala 357:48]
  assign lsq_io_ldu_s2_loadLoadViolationQuery_1_req_bits_uop_lqIdx_flag =
    LoadUnit_1_io_lsq_loadLoadViolationQuery_req_bits_uop_lqIdx_flag; // @[MemBlock.scala 357:48]
  assign lsq_io_ldu_s2_loadLoadViolationQuery_1_req_bits_uop_lqIdx_value =
    LoadUnit_1_io_lsq_loadLoadViolationQuery_req_bits_uop_lqIdx_value; // @[MemBlock.scala 357:48]
  assign lsq_io_ldu_s2_loadLoadViolationQuery_1_req_bits_index = LoadUnit_1_io_lsq_loadLoadViolationQuery_req_bits_index
    ; // @[MemBlock.scala 357:48]
  assign lsq_io_ldu_s2_loadLoadViolationQuery_1_req_bits_allocated =
    LoadUnit_1_io_lsq_loadLoadViolationQuery_req_bits_allocated; // @[MemBlock.scala 357:48]
  assign lsq_io_ldu_s2_loadLoadViolationQuery_1_req_bits_datavalid =
    LoadUnit_1_io_lsq_loadLoadViolationQuery_req_bits_datavalid; // @[MemBlock.scala 357:48]
  assign lsq_io_ldu_s2_loadLoadViolationQuery_1_req_bits_miss = LoadUnit_1_io_lsq_loadLoadViolationQuery_req_bits_miss; // @[MemBlock.scala 357:48]
  assign lsq_io_ldu_s2_loadLoadViolationQuery_1_req_bits_paddr = LoadUnit_1_io_lsq_loadLoadViolationQuery_req_bits_paddr
    ; // @[MemBlock.scala 357:48]
  assign lsq_io_ldu_s3_loadIn_0_valid = LoadUnit_0_io_lsq_loadIn_valid; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_0_bits_uop_cf_foldpc = LoadUnit_0_io_lsq_loadIn_bits_uop_cf_foldpc; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_0_bits_uop_cf_exceptionVec_4 = LoadUnit_0_io_lsq_loadIn_bits_uop_cf_exceptionVec_4; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_0_bits_uop_cf_exceptionVec_5 = LoadUnit_0_io_lsq_loadIn_bits_uop_cf_exceptionVec_5; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_0_bits_uop_cf_exceptionVec_13 = LoadUnit_0_io_lsq_loadIn_bits_uop_cf_exceptionVec_13; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_0_bits_uop_cf_trigger_backendEn_1 =
    LoadUnit_0_io_lsq_loadIn_bits_uop_cf_trigger_backendEn_1; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_0_bits_uop_cf_trigger_backendHit_0 =
    LoadUnit_0_io_lsq_loadIn_bits_uop_cf_trigger_backendHit_0; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_0_bits_uop_cf_trigger_backendHit_1 =
    LoadUnit_0_io_lsq_loadIn_bits_uop_cf_trigger_backendHit_1; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_0_bits_uop_cf_trigger_backendHit_4 =
    LoadUnit_0_io_lsq_loadIn_bits_uop_cf_trigger_backendHit_4; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_0_bits_uop_cf_waitForRobIdx_flag = LoadUnit_0_io_lsq_loadIn_bits_uop_cf_waitForRobIdx_flag
    ; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_0_bits_uop_cf_waitForRobIdx_value =
    LoadUnit_0_io_lsq_loadIn_bits_uop_cf_waitForRobIdx_value; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_0_bits_uop_cf_loadWaitBit = LoadUnit_0_io_lsq_loadIn_bits_uop_cf_loadWaitBit; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_0_bits_uop_cf_loadWaitStrict = LoadUnit_0_io_lsq_loadIn_bits_uop_cf_loadWaitStrict; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_0_bits_uop_cf_ftqPtr_flag = LoadUnit_0_io_lsq_loadIn_bits_uop_cf_ftqPtr_flag; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_0_bits_uop_cf_ftqPtr_value = LoadUnit_0_io_lsq_loadIn_bits_uop_cf_ftqPtr_value; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_0_bits_uop_cf_ftqOffset = LoadUnit_0_io_lsq_loadIn_bits_uop_cf_ftqOffset; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_0_bits_uop_ctrl_fuType = LoadUnit_0_io_lsq_loadIn_bits_uop_ctrl_fuType; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_0_bits_uop_ctrl_fuOpType = LoadUnit_0_io_lsq_loadIn_bits_uop_ctrl_fuOpType; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_0_bits_uop_ctrl_rfWen = LoadUnit_0_io_lsq_loadIn_bits_uop_ctrl_rfWen; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_0_bits_uop_ctrl_fpWen = LoadUnit_0_io_lsq_loadIn_bits_uop_ctrl_fpWen; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_0_bits_uop_ctrl_replayInst = LoadUnit_0_io_lsq_loadIn_bits_uop_ctrl_replayInst; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_0_bits_uop_pdest = LoadUnit_0_io_lsq_loadIn_bits_uop_pdest; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_0_bits_uop_robIdx_flag = LoadUnit_0_io_lsq_loadIn_bits_uop_robIdx_flag; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_0_bits_uop_robIdx_value = LoadUnit_0_io_lsq_loadIn_bits_uop_robIdx_value; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_0_bits_uop_lqIdx_flag = LoadUnit_0_io_lsq_loadIn_bits_uop_lqIdx_flag; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_0_bits_uop_lqIdx_value = LoadUnit_0_io_lsq_loadIn_bits_uop_lqIdx_value; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_0_bits_uop_sqIdx_flag = LoadUnit_0_io_lsq_loadIn_bits_uop_sqIdx_flag; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_0_bits_uop_sqIdx_value = LoadUnit_0_io_lsq_loadIn_bits_uop_sqIdx_value; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_0_bits_vaddr = LoadUnit_0_io_lsq_loadIn_bits_vaddr; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_0_bits_paddr = LoadUnit_0_io_lsq_loadIn_bits_paddr; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_0_bits_mask = LoadUnit_0_io_lsq_loadIn_bits_mask; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_0_bits_miss = LoadUnit_0_io_lsq_loadIn_bits_miss; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_0_bits_tlbMiss = LoadUnit_0_io_lsq_loadIn_bits_tlbMiss; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_0_bits_mmio = LoadUnit_0_io_lsq_loadIn_bits_mmio; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_0_bits_rarAllocated = LoadUnit_0_io_lsq_loadIn_bits_rarAllocated; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_0_bits_rarIndex = LoadUnit_0_io_lsq_loadIn_bits_rarIndex; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_0_bits_rawAllocated = LoadUnit_0_io_lsq_loadIn_bits_rawAllocated; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_0_bits_rawIndex = LoadUnit_0_io_lsq_loadIn_bits_rawIndex; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_0_bits_replayInfo_missMSHRId = LoadUnit_0_io_lsq_loadIn_bits_replayInfo_missMSHRId; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_0_bits_replayInfo_canForwardFullData =
    LoadUnit_0_io_lsq_loadIn_bits_replayInfo_canForwardFullData; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_0_bits_replayInfo_dataInvalidSqIdx_flag =
    LoadUnit_0_io_lsq_loadIn_bits_replayInfo_dataInvalidSqIdx_flag; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_0_bits_replayInfo_dataInvalidSqIdx_value =
    LoadUnit_0_io_lsq_loadIn_bits_replayInfo_dataInvalidSqIdx_value; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_0_bits_replayInfo_addrInvalidSqIdx_flag =
    LoadUnit_0_io_lsq_loadIn_bits_replayInfo_addrInvalidSqIdx_flag; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_0_bits_replayInfo_addrInvalidSqIdx_value =
    LoadUnit_0_io_lsq_loadIn_bits_replayInfo_addrInvalidSqIdx_value; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_0_bits_replayInfo_replayCarry_real_way_en =
    LoadUnit_0_io_lsq_loadIn_bits_replayInfo_replayCarry_real_way_en; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_0_bits_replayInfo_replayCarry_valid =
    LoadUnit_0_io_lsq_loadIn_bits_replayInfo_replayCarry_valid; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_0_bits_replayInfo_dataInLastBeat = LoadUnit_0_io_lsq_loadIn_bits_replayInfo_dataInLastBeat
    ; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_0_bits_replayInfo_cause_0 = LoadUnit_0_io_lsq_loadIn_bits_replayInfo_cause_0; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_0_bits_replayInfo_cause_1 = LoadUnit_0_io_lsq_loadIn_bits_replayInfo_cause_1; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_0_bits_replayInfo_cause_2 = LoadUnit_0_io_lsq_loadIn_bits_replayInfo_cause_2; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_0_bits_replayInfo_cause_3 = LoadUnit_0_io_lsq_loadIn_bits_replayInfo_cause_3; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_0_bits_replayInfo_cause_4 = LoadUnit_0_io_lsq_loadIn_bits_replayInfo_cause_4; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_0_bits_replayInfo_cause_5 = LoadUnit_0_io_lsq_loadIn_bits_replayInfo_cause_5; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_0_bits_replayInfo_cause_6 = LoadUnit_0_io_lsq_loadIn_bits_replayInfo_cause_6; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_0_bits_replayInfo_cause_7 = LoadUnit_0_io_lsq_loadIn_bits_replayInfo_cause_7; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_0_bits_lqDataWenDup_1 = LoadUnit_0_io_lsq_loadIn_bits_lqDataWenDup_1; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_0_bits_lqDataWenDup_2 = LoadUnit_0_io_lsq_loadIn_bits_lqDataWenDup_2; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_0_bits_lqDataWenDup_3 = LoadUnit_0_io_lsq_loadIn_bits_lqDataWenDup_3; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_0_bits_lqDataWenDup_5 = LoadUnit_0_io_lsq_loadIn_bits_lqDataWenDup_5; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_1_valid = LoadUnit_1_io_lsq_loadIn_valid; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_1_bits_uop_cf_foldpc = LoadUnit_1_io_lsq_loadIn_bits_uop_cf_foldpc; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_1_bits_uop_cf_exceptionVec_4 = LoadUnit_1_io_lsq_loadIn_bits_uop_cf_exceptionVec_4; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_1_bits_uop_cf_exceptionVec_5 = LoadUnit_1_io_lsq_loadIn_bits_uop_cf_exceptionVec_5; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_1_bits_uop_cf_exceptionVec_13 = LoadUnit_1_io_lsq_loadIn_bits_uop_cf_exceptionVec_13; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_1_bits_uop_cf_trigger_backendEn_1 =
    LoadUnit_1_io_lsq_loadIn_bits_uop_cf_trigger_backendEn_1; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_1_bits_uop_cf_trigger_backendHit_0 =
    LoadUnit_1_io_lsq_loadIn_bits_uop_cf_trigger_backendHit_0; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_1_bits_uop_cf_trigger_backendHit_1 =
    LoadUnit_1_io_lsq_loadIn_bits_uop_cf_trigger_backendHit_1; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_1_bits_uop_cf_trigger_backendHit_4 =
    LoadUnit_1_io_lsq_loadIn_bits_uop_cf_trigger_backendHit_4; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_1_bits_uop_cf_waitForRobIdx_flag = LoadUnit_1_io_lsq_loadIn_bits_uop_cf_waitForRobIdx_flag
    ; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_1_bits_uop_cf_waitForRobIdx_value =
    LoadUnit_1_io_lsq_loadIn_bits_uop_cf_waitForRobIdx_value; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_1_bits_uop_cf_loadWaitBit = LoadUnit_1_io_lsq_loadIn_bits_uop_cf_loadWaitBit; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_1_bits_uop_cf_loadWaitStrict = LoadUnit_1_io_lsq_loadIn_bits_uop_cf_loadWaitStrict; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_1_bits_uop_cf_ftqPtr_flag = LoadUnit_1_io_lsq_loadIn_bits_uop_cf_ftqPtr_flag; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_1_bits_uop_cf_ftqPtr_value = LoadUnit_1_io_lsq_loadIn_bits_uop_cf_ftqPtr_value; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_1_bits_uop_cf_ftqOffset = LoadUnit_1_io_lsq_loadIn_bits_uop_cf_ftqOffset; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_1_bits_uop_ctrl_fuType = LoadUnit_1_io_lsq_loadIn_bits_uop_ctrl_fuType; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_1_bits_uop_ctrl_fuOpType = LoadUnit_1_io_lsq_loadIn_bits_uop_ctrl_fuOpType; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_1_bits_uop_ctrl_rfWen = LoadUnit_1_io_lsq_loadIn_bits_uop_ctrl_rfWen; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_1_bits_uop_ctrl_fpWen = LoadUnit_1_io_lsq_loadIn_bits_uop_ctrl_fpWen; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_1_bits_uop_ctrl_replayInst = LoadUnit_1_io_lsq_loadIn_bits_uop_ctrl_replayInst; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_1_bits_uop_pdest = LoadUnit_1_io_lsq_loadIn_bits_uop_pdest; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_1_bits_uop_robIdx_flag = LoadUnit_1_io_lsq_loadIn_bits_uop_robIdx_flag; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_1_bits_uop_robIdx_value = LoadUnit_1_io_lsq_loadIn_bits_uop_robIdx_value; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_1_bits_uop_lqIdx_flag = LoadUnit_1_io_lsq_loadIn_bits_uop_lqIdx_flag; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_1_bits_uop_lqIdx_value = LoadUnit_1_io_lsq_loadIn_bits_uop_lqIdx_value; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_1_bits_uop_sqIdx_flag = LoadUnit_1_io_lsq_loadIn_bits_uop_sqIdx_flag; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_1_bits_uop_sqIdx_value = LoadUnit_1_io_lsq_loadIn_bits_uop_sqIdx_value; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_1_bits_vaddr = LoadUnit_1_io_lsq_loadIn_bits_vaddr; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_1_bits_paddr = LoadUnit_1_io_lsq_loadIn_bits_paddr; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_1_bits_mask = LoadUnit_1_io_lsq_loadIn_bits_mask; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_1_bits_miss = LoadUnit_1_io_lsq_loadIn_bits_miss; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_1_bits_tlbMiss = LoadUnit_1_io_lsq_loadIn_bits_tlbMiss; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_1_bits_mmio = LoadUnit_1_io_lsq_loadIn_bits_mmio; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_1_bits_rarAllocated = LoadUnit_1_io_lsq_loadIn_bits_rarAllocated; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_1_bits_rarIndex = LoadUnit_1_io_lsq_loadIn_bits_rarIndex; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_1_bits_rawAllocated = LoadUnit_1_io_lsq_loadIn_bits_rawAllocated; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_1_bits_rawIndex = LoadUnit_1_io_lsq_loadIn_bits_rawIndex; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_1_bits_replayInfo_missMSHRId = LoadUnit_1_io_lsq_loadIn_bits_replayInfo_missMSHRId; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_1_bits_replayInfo_canForwardFullData =
    LoadUnit_1_io_lsq_loadIn_bits_replayInfo_canForwardFullData; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_1_bits_replayInfo_dataInvalidSqIdx_flag =
    LoadUnit_1_io_lsq_loadIn_bits_replayInfo_dataInvalidSqIdx_flag; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_1_bits_replayInfo_dataInvalidSqIdx_value =
    LoadUnit_1_io_lsq_loadIn_bits_replayInfo_dataInvalidSqIdx_value; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_1_bits_replayInfo_addrInvalidSqIdx_flag =
    LoadUnit_1_io_lsq_loadIn_bits_replayInfo_addrInvalidSqIdx_flag; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_1_bits_replayInfo_addrInvalidSqIdx_value =
    LoadUnit_1_io_lsq_loadIn_bits_replayInfo_addrInvalidSqIdx_value; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_1_bits_replayInfo_replayCarry_real_way_en =
    LoadUnit_1_io_lsq_loadIn_bits_replayInfo_replayCarry_real_way_en; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_1_bits_replayInfo_replayCarry_valid =
    LoadUnit_1_io_lsq_loadIn_bits_replayInfo_replayCarry_valid; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_1_bits_replayInfo_dataInLastBeat = LoadUnit_1_io_lsq_loadIn_bits_replayInfo_dataInLastBeat
    ; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_1_bits_replayInfo_cause_0 = LoadUnit_1_io_lsq_loadIn_bits_replayInfo_cause_0; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_1_bits_replayInfo_cause_1 = LoadUnit_1_io_lsq_loadIn_bits_replayInfo_cause_1; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_1_bits_replayInfo_cause_2 = LoadUnit_1_io_lsq_loadIn_bits_replayInfo_cause_2; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_1_bits_replayInfo_cause_3 = LoadUnit_1_io_lsq_loadIn_bits_replayInfo_cause_3; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_1_bits_replayInfo_cause_4 = LoadUnit_1_io_lsq_loadIn_bits_replayInfo_cause_4; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_1_bits_replayInfo_cause_5 = LoadUnit_1_io_lsq_loadIn_bits_replayInfo_cause_5; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_1_bits_replayInfo_cause_6 = LoadUnit_1_io_lsq_loadIn_bits_replayInfo_cause_6; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_1_bits_replayInfo_cause_7 = LoadUnit_1_io_lsq_loadIn_bits_replayInfo_cause_7; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_1_bits_lqDataWenDup_1 = LoadUnit_1_io_lsq_loadIn_bits_lqDataWenDup_1; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_1_bits_lqDataWenDup_2 = LoadUnit_1_io_lsq_loadIn_bits_lqDataWenDup_2; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_1_bits_lqDataWenDup_3 = LoadUnit_1_io_lsq_loadIn_bits_lqDataWenDup_3; // @[MemBlock.scala 399:29]
  assign lsq_io_ldu_s3_loadIn_1_bits_lqDataWenDup_5 = LoadUnit_1_io_lsq_loadIn_bits_lqDataWenDup_5; // @[MemBlock.scala 399:29]
  assign lsq_io_sta_s0_storeMaskIn_0_valid = StoreUnit_0_io_storeMaskOut_valid; // @[MemBlock.scala 471:34]
  assign lsq_io_sta_s0_storeMaskIn_0_bits_sqIdx_value = StoreUnit_0_io_storeMaskOut_bits_sqIdx_value; // @[MemBlock.scala 471:34]
  assign lsq_io_sta_s0_storeMaskIn_0_bits_mask = StoreUnit_0_io_storeMaskOut_bits_mask; // @[MemBlock.scala 471:34]
  assign lsq_io_sta_s0_storeMaskIn_1_valid = StoreUnit_1_io_storeMaskOut_valid; // @[MemBlock.scala 471:34]
  assign lsq_io_sta_s0_storeMaskIn_1_bits_sqIdx_value = StoreUnit_1_io_storeMaskOut_bits_sqIdx_value; // @[MemBlock.scala 471:34]
  assign lsq_io_sta_s0_storeMaskIn_1_bits_mask = StoreUnit_1_io_storeMaskOut_bits_mask; // @[MemBlock.scala 471:34]
  assign lsq_io_sta_s1_storeAddrIn_0_valid = StoreUnit_0_io_lsq_valid; // @[MemBlock.scala 461:25]
  assign lsq_io_sta_s1_storeAddrIn_0_bits_uop_cf_ftqPtr_value = StoreUnit_0_io_lsq_bits_uop_cf_ftqPtr_value; // @[MemBlock.scala 461:25]
  assign lsq_io_sta_s1_storeAddrIn_0_bits_uop_cf_ftqOffset = StoreUnit_0_io_lsq_bits_uop_cf_ftqOffset; // @[MemBlock.scala 461:25]
  assign lsq_io_sta_s1_storeAddrIn_0_bits_uop_ctrl_fuOpType = StoreUnit_0_io_lsq_bits_uop_ctrl_fuOpType; // @[MemBlock.scala 461:25]
  assign lsq_io_sta_s1_storeAddrIn_0_bits_uop_robIdx_flag = StoreUnit_0_io_lsq_bits_uop_robIdx_flag; // @[MemBlock.scala 461:25]
  assign lsq_io_sta_s1_storeAddrIn_0_bits_uop_robIdx_value = StoreUnit_0_io_lsq_bits_uop_robIdx_value; // @[MemBlock.scala 461:25]
  assign lsq_io_sta_s1_storeAddrIn_0_bits_uop_sqIdx_flag = StoreUnit_0_io_lsq_bits_uop_sqIdx_flag; // @[MemBlock.scala 461:25]
  assign lsq_io_sta_s1_storeAddrIn_0_bits_uop_sqIdx_value = StoreUnit_0_io_lsq_bits_uop_sqIdx_value; // @[MemBlock.scala 461:25]
  assign lsq_io_sta_s1_storeAddrIn_0_bits_vaddr = StoreUnit_0_io_lsq_bits_vaddr; // @[MemBlock.scala 461:25]
  assign lsq_io_sta_s1_storeAddrIn_0_bits_paddr = StoreUnit_0_io_lsq_bits_paddr; // @[MemBlock.scala 461:25]
  assign lsq_io_sta_s1_storeAddrIn_0_bits_mask = StoreUnit_0_io_lsq_bits_mask; // @[MemBlock.scala 461:25]
  assign lsq_io_sta_s1_storeAddrIn_0_bits_wlineflag = StoreUnit_0_io_lsq_bits_wlineflag; // @[MemBlock.scala 461:25]
  assign lsq_io_sta_s1_storeAddrIn_0_bits_miss = StoreUnit_0_io_lsq_bits_miss; // @[MemBlock.scala 461:25]
  assign lsq_io_sta_s1_storeAddrIn_1_valid = StoreUnit_1_io_lsq_valid; // @[MemBlock.scala 461:25]
  assign lsq_io_sta_s1_storeAddrIn_1_bits_uop_cf_ftqPtr_value = StoreUnit_1_io_lsq_bits_uop_cf_ftqPtr_value; // @[MemBlock.scala 461:25]
  assign lsq_io_sta_s1_storeAddrIn_1_bits_uop_cf_ftqOffset = StoreUnit_1_io_lsq_bits_uop_cf_ftqOffset; // @[MemBlock.scala 461:25]
  assign lsq_io_sta_s1_storeAddrIn_1_bits_uop_ctrl_fuOpType = StoreUnit_1_io_lsq_bits_uop_ctrl_fuOpType; // @[MemBlock.scala 461:25]
  assign lsq_io_sta_s1_storeAddrIn_1_bits_uop_robIdx_flag = StoreUnit_1_io_lsq_bits_uop_robIdx_flag; // @[MemBlock.scala 461:25]
  assign lsq_io_sta_s1_storeAddrIn_1_bits_uop_robIdx_value = StoreUnit_1_io_lsq_bits_uop_robIdx_value; // @[MemBlock.scala 461:25]
  assign lsq_io_sta_s1_storeAddrIn_1_bits_uop_sqIdx_flag = StoreUnit_1_io_lsq_bits_uop_sqIdx_flag; // @[MemBlock.scala 461:25]
  assign lsq_io_sta_s1_storeAddrIn_1_bits_uop_sqIdx_value = StoreUnit_1_io_lsq_bits_uop_sqIdx_value; // @[MemBlock.scala 461:25]
  assign lsq_io_sta_s1_storeAddrIn_1_bits_vaddr = StoreUnit_1_io_lsq_bits_vaddr; // @[MemBlock.scala 461:25]
  assign lsq_io_sta_s1_storeAddrIn_1_bits_paddr = StoreUnit_1_io_lsq_bits_paddr; // @[MemBlock.scala 461:25]
  assign lsq_io_sta_s1_storeAddrIn_1_bits_mask = StoreUnit_1_io_lsq_bits_mask; // @[MemBlock.scala 461:25]
  assign lsq_io_sta_s1_storeAddrIn_1_bits_wlineflag = StoreUnit_1_io_lsq_bits_wlineflag; // @[MemBlock.scala 461:25]
  assign lsq_io_sta_s1_storeAddrIn_1_bits_miss = StoreUnit_1_io_lsq_bits_miss; // @[MemBlock.scala 461:25]
  assign lsq_io_sta_s2_storeAddrInRe_0_mmio = StoreUnit_0_io_lsq_replenish_mmio; // @[MemBlock.scala 462:26]
  assign lsq_io_sta_s2_storeAddrInRe_0_atomic = StoreUnit_0_io_lsq_replenish_atomic; // @[MemBlock.scala 462:26]
  assign lsq_io_sta_s2_storeAddrInRe_1_mmio = StoreUnit_1_io_lsq_replenish_mmio; // @[MemBlock.scala 462:26]
  assign lsq_io_sta_s2_storeAddrInRe_1_atomic = StoreUnit_1_io_lsq_replenish_atomic; // @[MemBlock.scala 462:26]
  assign lsq_io_std_s0_storeDataIn_0_valid = stdExeUnits_0_io_out_valid; // @[MemBlock.scala 474:34]
  assign lsq_io_std_s0_storeDataIn_0_bits_uop_ctrl_fuOpType = stdExeUnits_0_io_out_bits_uop_ctrl_fuOpType; // @[MemBlock.scala 474:34]
  assign lsq_io_std_s0_storeDataIn_0_bits_uop_sqIdx_flag = stdExeUnits_0_io_out_bits_uop_sqIdx_flag; // @[MemBlock.scala 474:34]
  assign lsq_io_std_s0_storeDataIn_0_bits_uop_sqIdx_value = stdExeUnits_0_io_out_bits_uop_sqIdx_value; // @[MemBlock.scala 474:34]
  assign lsq_io_std_s0_storeDataIn_0_bits_data = stdExeUnits_0_io_out_bits_data; // @[MemBlock.scala 474:34]
  assign lsq_io_std_s0_storeDataIn_1_valid = stdExeUnits_1_io_out_valid; // @[MemBlock.scala 474:34]
  assign lsq_io_std_s0_storeDataIn_1_bits_uop_ctrl_fuOpType = stdExeUnits_1_io_out_bits_uop_ctrl_fuOpType; // @[MemBlock.scala 474:34]
  assign lsq_io_std_s0_storeDataIn_1_bits_uop_sqIdx_flag = stdExeUnits_1_io_out_bits_uop_sqIdx_flag; // @[MemBlock.scala 474:34]
  assign lsq_io_std_s0_storeDataIn_1_bits_uop_sqIdx_value = stdExeUnits_1_io_out_bits_uop_sqIdx_value; // @[MemBlock.scala 474:34]
  assign lsq_io_std_s0_storeDataIn_1_bits_data = stdExeUnits_1_io_out_bits_data; // @[MemBlock.scala 474:34]
  assign lsq_io_loadOut_0_ready = LoadUnit_0_io_lsq_loadOut_ready; // @[MemBlock.scala 400:23]
  assign lsq_io_replay_0_ready = LoadUnit_0_io_replay_ready; // @[MemBlock.scala 396:28]
  assign lsq_io_replay_1_ready = LoadUnit_1_io_replay_ready; // @[MemBlock.scala 396:28]
  assign lsq_io_sbuffer_0_ready = sbuffer_io_in_0_ready; // @[MemBlock.scala 556:25]
  assign lsq_io_sbuffer_1_ready = sbuffer_io_in_1_ready; // @[MemBlock.scala 556:25]
  assign lsq_io_forward_0_vaddr = LoadUnit_0_io_lsq_forward_vaddr; // @[MemBlock.scala 350:33]
  assign lsq_io_forward_0_paddr = LoadUnit_0_io_lsq_forward_paddr; // @[MemBlock.scala 350:33]
  assign lsq_io_forward_0_uop_cf_waitForRobIdx_flag = LoadUnit_0_io_lsq_forward_uop_cf_waitForRobIdx_flag; // @[MemBlock.scala 350:33]
  assign lsq_io_forward_0_uop_cf_waitForRobIdx_value = LoadUnit_0_io_lsq_forward_uop_cf_waitForRobIdx_value; // @[MemBlock.scala 350:33]
  assign lsq_io_forward_0_uop_sqIdx_flag = LoadUnit_0_io_lsq_forward_uop_sqIdx_flag; // @[MemBlock.scala 350:33]
  assign lsq_io_forward_0_uop_sqIdx_value = LoadUnit_0_io_lsq_forward_uop_sqIdx_value; // @[MemBlock.scala 350:33]
  assign lsq_io_forward_0_valid = LoadUnit_0_io_lsq_forward_valid; // @[MemBlock.scala 350:33]
  assign lsq_io_forward_0_sqIdx_flag = LoadUnit_0_io_lsq_forward_sqIdx_flag; // @[MemBlock.scala 350:33]
  assign lsq_io_forward_0_sqIdxMask = LoadUnit_0_io_lsq_forward_sqIdxMask; // @[MemBlock.scala 350:33]
  assign lsq_io_forward_1_vaddr = LoadUnit_1_io_lsq_forward_vaddr; // @[MemBlock.scala 350:33]
  assign lsq_io_forward_1_paddr = LoadUnit_1_io_lsq_forward_paddr; // @[MemBlock.scala 350:33]
  assign lsq_io_forward_1_uop_cf_waitForRobIdx_flag = LoadUnit_1_io_lsq_forward_uop_cf_waitForRobIdx_flag; // @[MemBlock.scala 350:33]
  assign lsq_io_forward_1_uop_cf_waitForRobIdx_value = LoadUnit_1_io_lsq_forward_uop_cf_waitForRobIdx_value; // @[MemBlock.scala 350:33]
  assign lsq_io_forward_1_uop_sqIdx_flag = LoadUnit_1_io_lsq_forward_uop_sqIdx_flag; // @[MemBlock.scala 350:33]
  assign lsq_io_forward_1_uop_sqIdx_value = LoadUnit_1_io_lsq_forward_uop_sqIdx_value; // @[MemBlock.scala 350:33]
  assign lsq_io_forward_1_valid = LoadUnit_1_io_lsq_forward_valid; // @[MemBlock.scala 350:33]
  assign lsq_io_forward_1_sqIdx_flag = LoadUnit_1_io_lsq_forward_sqIdx_flag; // @[MemBlock.scala 350:33]
  assign lsq_io_forward_1_sqIdxMask = LoadUnit_1_io_lsq_forward_sqIdxMask; // @[MemBlock.scala 350:33]
  assign lsq_io_rob_scommit = io_lsqio_rob_scommit; // @[MemBlock.scala 539:25]
  assign lsq_io_rob_pendingld = io_lsqio_rob_pendingld; // @[MemBlock.scala 539:25]
  assign lsq_io_rob_pendingst = io_lsqio_rob_pendingst; // @[MemBlock.scala 539:25]
  assign lsq_io_rob_commit = io_lsqio_rob_commit; // @[MemBlock.scala 539:25]
  assign lsq_io_release_valid = dcache_io_lsu_release_valid; // @[MemBlock.scala 549:25]
  assign lsq_io_release_bits_paddr = dcache_io_lsu_release_bits_paddr; // @[MemBlock.scala 549:25]
  assign lsq_io_refill_valid = delayedDcacheRefill_valid; // @[MemBlock.scala 548:25]
  assign lsq_io_refill_bits_id = delayedDcacheRefill_bits_id; // @[MemBlock.scala 548:25]
  assign lsq_io_uncacheOutstanding = io_csrCtrl_uncache_write_outstanding_enable; // @[MemBlock.scala 536:29]
  assign lsq_io_uncache_req_ready = pipelineReg_io_in_ready; // @[MemCommon.scala 398:23]
  assign lsq_io_uncache_resp_valid = pipelineReg_1_io_out_valid; // @[MemCommon.scala 399:11]
  assign lsq_io_uncache_resp_bits_data = pipelineReg_1_io_out_bits_data; // @[MemCommon.scala 399:11]
  assign lsq_io_mmioStout_ready = lsq_io_mmioStout_valid & ~StoreUnit_0_io_stout_valid; // @[MemBlock.scala 514:32]
  assign lsq_io_exceptionAddr_isStore = io_lsqio_exceptionAddr_isStore; // @[MemBlock.scala 658:32]
  assign lsq_io_trigger_0_hitLoadAddrTriggerHitVec_0 = LoadUnit_0_io_lsq_trigger_hitLoadAddrTriggerHitVec_0; // @[MemBlock.scala 402:23]
  assign lsq_io_trigger_0_hitLoadAddrTriggerHitVec_1 = LoadUnit_0_io_lsq_trigger_hitLoadAddrTriggerHitVec_1; // @[MemBlock.scala 402:23]
  assign lsq_io_trigger_0_hitLoadAddrTriggerHitVec_2 = LoadUnit_0_io_lsq_trigger_hitLoadAddrTriggerHitVec_2; // @[MemBlock.scala 402:23]
  assign lsq_io_trigger_1_hitLoadAddrTriggerHitVec_0 = LoadUnit_1_io_lsq_trigger_hitLoadAddrTriggerHitVec_0; // @[MemBlock.scala 402:23]
  assign lsq_io_trigger_1_hitLoadAddrTriggerHitVec_1 = LoadUnit_1_io_lsq_trigger_hitLoadAddrTriggerHitVec_1; // @[MemBlock.scala 402:23]
  assign lsq_io_trigger_1_hitLoadAddrTriggerHitVec_2 = LoadUnit_1_io_lsq_trigger_hitLoadAddrTriggerHitVec_2; // @[MemBlock.scala 402:23]
  assign sbuffer_clock = clock;
  assign sbuffer_reset = reset;
  assign sbuffer_io_in_0_valid = lsq_io_sbuffer_0_valid; // @[MemBlock.scala 556:25]
  assign sbuffer_io_in_0_bits_addr = lsq_io_sbuffer_0_bits_addr; // @[MemBlock.scala 556:25]
  assign sbuffer_io_in_0_bits_data = lsq_io_sbuffer_0_bits_data; // @[MemBlock.scala 556:25]
  assign sbuffer_io_in_0_bits_mask = lsq_io_sbuffer_0_bits_mask; // @[MemBlock.scala 556:25]
  assign sbuffer_io_in_0_bits_vaddr = lsq_io_sbuffer_0_bits_vaddr; // @[MemBlock.scala 556:25]
  assign sbuffer_io_in_0_bits_wline = lsq_io_sbuffer_0_bits_wline; // @[MemBlock.scala 556:25]
  assign sbuffer_io_in_1_valid = lsq_io_sbuffer_1_valid; // @[MemBlock.scala 556:25]
  assign sbuffer_io_in_1_bits_addr = lsq_io_sbuffer_1_bits_addr; // @[MemBlock.scala 556:25]
  assign sbuffer_io_in_1_bits_data = lsq_io_sbuffer_1_bits_data; // @[MemBlock.scala 556:25]
  assign sbuffer_io_in_1_bits_mask = lsq_io_sbuffer_1_bits_mask; // @[MemBlock.scala 556:25]
  assign sbuffer_io_in_1_bits_vaddr = lsq_io_sbuffer_1_bits_vaddr; // @[MemBlock.scala 556:25]
  assign sbuffer_io_in_1_bits_wline = lsq_io_sbuffer_1_bits_wline; // @[MemBlock.scala 556:25]
  assign sbuffer_io_dcache_req_ready = dcache_io_lsu_store_req_ready; // @[MemBlock.scala 561:25]
  assign sbuffer_io_dcache_main_pipe_hit_resp_valid = dcache_io_lsu_store_main_pipe_hit_resp_valid; // @[MemBlock.scala 561:25]
  assign sbuffer_io_dcache_main_pipe_hit_resp_bits_id = dcache_io_lsu_store_main_pipe_hit_resp_bits_id; // @[MemBlock.scala 561:25]
  assign sbuffer_io_dcache_refill_hit_resp_valid = dcache_io_lsu_store_refill_hit_resp_valid; // @[MemBlock.scala 561:25]
  assign sbuffer_io_dcache_refill_hit_resp_bits_id = dcache_io_lsu_store_refill_hit_resp_bits_id; // @[MemBlock.scala 561:25]
  assign sbuffer_io_dcache_replay_resp_valid = dcache_io_lsu_store_replay_resp_valid; // @[MemBlock.scala 561:25]
  assign sbuffer_io_dcache_replay_resp_bits_id = dcache_io_lsu_store_replay_resp_bits_id; // @[MemBlock.scala 561:25]
  assign sbuffer_io_forward_0_vaddr = LoadUnit_0_io_sbuffer_vaddr; // @[MemBlock.scala 351:29]
  assign sbuffer_io_forward_0_paddr = LoadUnit_0_io_sbuffer_paddr; // @[MemBlock.scala 351:29]
  assign sbuffer_io_forward_0_valid = LoadUnit_0_io_sbuffer_valid; // @[MemBlock.scala 351:29]
  assign sbuffer_io_forward_1_vaddr = LoadUnit_1_io_sbuffer_vaddr; // @[MemBlock.scala 351:29]
  assign sbuffer_io_forward_1_paddr = LoadUnit_1_io_sbuffer_paddr; // @[MemBlock.scala 351:29]
  assign sbuffer_io_forward_1_valid = LoadUnit_1_io_sbuffer_valid; // @[MemBlock.scala 351:29]
  assign sbuffer_io_sqempty = lsq_io_sqEmpty; // @[MemBlock.scala 557:25]
  assign sbuffer_io_flush_valid = sbuffer_io_flush_valid_REG; // @[MemBlock.scala 572:26]
  assign sbuffer_io_csrCtrl_sbuffer_threshold = csrCtrl_delay_io_out_sbuffer_threshold; // @[MemBlock.scala 560:25]
  assign dtlb_ld_tlb_ld_clock = clock;
  assign dtlb_ld_tlb_ld_reset = reset;
  assign dtlb_ld_tlb_ld_io_sfence_valid = sfence_valid; // @[MemBlock.scala 245:24 260:21]
  assign dtlb_ld_tlb_ld_io_sfence_bits_rs1 = sfence_bits_rs1; // @[MemBlock.scala 245:24 260:21]
  assign dtlb_ld_tlb_ld_io_sfence_bits_rs2 = sfence_bits_rs2; // @[MemBlock.scala 245:24 260:21]
  assign dtlb_ld_tlb_ld_io_sfence_bits_addr = sfence_bits_addr; // @[MemBlock.scala 245:24 260:21]
  assign dtlb_ld_tlb_ld_io_sfence_bits_asid = sfence_bits_asid; // @[MemBlock.scala 245:24 260:21]
  assign dtlb_ld_tlb_ld_io_csr_satp_mode = tlbcsr_satp_mode; // @[MemBlock.scala 245:24 261:18]
  assign dtlb_ld_tlb_ld_io_csr_satp_asid = tlbcsr_satp_asid; // @[MemBlock.scala 245:24 261:18]
  assign dtlb_ld_tlb_ld_io_csr_satp_changed = tlbcsr_satp_changed; // @[MemBlock.scala 245:24 261:18]
  assign dtlb_ld_tlb_ld_io_csr_priv_mxr = tlbcsr_priv_mxr; // @[MemBlock.scala 245:24 261:18]
  assign dtlb_ld_tlb_ld_io_csr_priv_sum = tlbcsr_priv_sum; // @[MemBlock.scala 245:24 261:18]
  assign dtlb_ld_tlb_ld_io_csr_priv_dmode = tlbcsr_priv_dmode; // @[MemBlock.scala 245:24 261:18]
  assign dtlb_ld_tlb_ld_io_requestor_0_req_valid = state != 2'h0 ? atomicsUnit_io_dtlb_req_valid :
    LoadUnit_0_io_tlb_req_valid; // @[MemBlock.scala 363:25 639:29 643:25]
  assign dtlb_ld_tlb_ld_io_requestor_0_req_bits_vaddr = state != 2'h0 ? atomicsUnit_io_dtlb_req_bits_vaddr :
    LoadUnit_0_io_tlb_req_bits_vaddr; // @[MemBlock.scala 363:25 639:29 643:25]
  assign dtlb_ld_tlb_ld_io_requestor_0_req_bits_cmd = state != 2'h0 ? atomicsUnit_io_dtlb_req_bits_cmd :
    LoadUnit_0_io_tlb_req_bits_cmd; // @[MemBlock.scala 363:25 639:29 643:25]
  assign dtlb_ld_tlb_ld_io_requestor_0_req_bits_no_translate = state != 2'h0 ? 1'h0 :
    LoadUnit_0_io_tlb_req_bits_no_translate; // @[MemBlock.scala 363:25 639:29 643:25]
  assign dtlb_ld_tlb_ld_io_requestor_0_req_kill = state != 2'h0 ? 1'h0 : LoadUnit_0_io_tlb_req_kill; // @[MemBlock.scala 363:25 639:29 643:25]
  assign dtlb_ld_tlb_ld_io_requestor_1_req_valid = LoadUnit_1_io_tlb_req_valid; // @[MemBlock.scala 245:24 363:25]
  assign dtlb_ld_tlb_ld_io_requestor_1_req_bits_vaddr = LoadUnit_1_io_tlb_req_bits_vaddr; // @[MemBlock.scala 245:24 363:25]
  assign dtlb_ld_tlb_ld_io_requestor_1_req_bits_cmd = LoadUnit_1_io_tlb_req_bits_cmd; // @[MemBlock.scala 245:24 363:25]
  assign dtlb_ld_tlb_ld_io_requestor_1_req_bits_no_translate = LoadUnit_1_io_tlb_req_bits_no_translate; // @[MemBlock.scala 245:24 363:25]
  assign dtlb_ld_tlb_ld_io_requestor_1_req_kill = LoadUnit_1_io_tlb_req_kill; // @[MemBlock.scala 245:24 363:25]
  assign dtlb_ld_tlb_ld_io_ptw_resp_valid = ptw_resp_v & vector_hit; // @[MemBlock.scala 298:52]
  assign dtlb_ld_tlb_ld_io_ptw_resp_bits_entry_tag = ptw_resp_next_data_entry_tag; // @[MemBlock.scala 245:24 294:32]
  assign dtlb_ld_tlb_ld_io_ptw_resp_bits_entry_asid = ptw_resp_next_data_entry_asid; // @[MemBlock.scala 245:24 294:32]
  assign dtlb_ld_tlb_ld_io_ptw_resp_bits_entry_ppn = ptw_resp_next_data_entry_ppn; // @[MemBlock.scala 245:24 294:32]
  assign dtlb_ld_tlb_ld_io_ptw_resp_bits_entry_perm_d = ptw_resp_next_data_entry_perm_d; // @[MemBlock.scala 245:24 294:32]
  assign dtlb_ld_tlb_ld_io_ptw_resp_bits_entry_perm_a = ptw_resp_next_data_entry_perm_a; // @[MemBlock.scala 245:24 294:32]
  assign dtlb_ld_tlb_ld_io_ptw_resp_bits_entry_perm_g = ptw_resp_next_data_entry_perm_g; // @[MemBlock.scala 245:24 294:32]
  assign dtlb_ld_tlb_ld_io_ptw_resp_bits_entry_perm_u = ptw_resp_next_data_entry_perm_u; // @[MemBlock.scala 245:24 294:32]
  assign dtlb_ld_tlb_ld_io_ptw_resp_bits_entry_perm_x = ptw_resp_next_data_entry_perm_x; // @[MemBlock.scala 245:24 294:32]
  assign dtlb_ld_tlb_ld_io_ptw_resp_bits_entry_perm_w = ptw_resp_next_data_entry_perm_w; // @[MemBlock.scala 245:24 294:32]
  assign dtlb_ld_tlb_ld_io_ptw_resp_bits_entry_perm_r = ptw_resp_next_data_entry_perm_r; // @[MemBlock.scala 245:24 294:32]
  assign dtlb_ld_tlb_ld_io_ptw_resp_bits_entry_level = ptw_resp_next_data_entry_level; // @[MemBlock.scala 245:24 294:32]
  assign dtlb_ld_tlb_ld_io_ptw_resp_bits_pf = ptw_resp_next_data_pf; // @[MemBlock.scala 245:24 294:32]
  assign dtlb_ld_tlb_ld_io_ptw_resp_bits_af = ptw_resp_next_data_af; // @[MemBlock.scala 245:24 294:32]
  assign dtlb_ld_tlb_ld_io_ptw_replenish_c = pmp_check_ptw_io_resp_c; // @[MemBlock.scala 245:24 322:28]
  assign dtlb_ld_tlb_ld_io_ptw_replenish_atomic = pmp_check_ptw_io_resp_atomic; // @[MemBlock.scala 245:24 322:28]
  assign dtlb_ld_tlb_ld_io_ptw_replenish_x = pmp_check_ptw_io_resp_x; // @[MemBlock.scala 245:24 322:28]
  assign dtlb_ld_tlb_ld_io_ptw_replenish_w = pmp_check_ptw_io_resp_w; // @[MemBlock.scala 245:24 322:28]
  assign dtlb_ld_tlb_ld_io_ptw_replenish_r = pmp_check_ptw_io_resp_r; // @[MemBlock.scala 245:24 322:28]
  assign dtlb_st_tlb_st_clock = clock;
  assign dtlb_st_tlb_st_reset = reset;
  assign dtlb_st_tlb_st_io_sfence_valid = sfence_valid; // @[MemBlock.scala 249:24 260:21]
  assign dtlb_st_tlb_st_io_sfence_bits_rs1 = sfence_bits_rs1; // @[MemBlock.scala 249:24 260:21]
  assign dtlb_st_tlb_st_io_sfence_bits_rs2 = sfence_bits_rs2; // @[MemBlock.scala 249:24 260:21]
  assign dtlb_st_tlb_st_io_sfence_bits_addr = sfence_bits_addr; // @[MemBlock.scala 249:24 260:21]
  assign dtlb_st_tlb_st_io_sfence_bits_asid = sfence_bits_asid; // @[MemBlock.scala 249:24 260:21]
  assign dtlb_st_tlb_st_io_csr_satp_mode = tlbcsr_satp_mode; // @[MemBlock.scala 249:24 261:18]
  assign dtlb_st_tlb_st_io_csr_satp_asid = tlbcsr_satp_asid; // @[MemBlock.scala 249:24 261:18]
  assign dtlb_st_tlb_st_io_csr_satp_changed = tlbcsr_satp_changed; // @[MemBlock.scala 249:24 261:18]
  assign dtlb_st_tlb_st_io_csr_priv_sum = tlbcsr_priv_sum; // @[MemBlock.scala 249:24 261:18]
  assign dtlb_st_tlb_st_io_csr_priv_dmode = tlbcsr_priv_dmode; // @[MemBlock.scala 249:24 261:18]
  assign dtlb_st_tlb_st_io_requestor_0_req_valid = StoreUnit_0_io_tlb_req_valid; // @[MemBlock.scala 249:24 464:25]
  assign dtlb_st_tlb_st_io_requestor_0_req_bits_vaddr = StoreUnit_0_io_tlb_req_bits_vaddr; // @[MemBlock.scala 249:24 464:25]
  assign dtlb_st_tlb_st_io_requestor_1_req_valid = StoreUnit_1_io_tlb_req_valid; // @[MemBlock.scala 249:24 464:25]
  assign dtlb_st_tlb_st_io_requestor_1_req_bits_vaddr = StoreUnit_1_io_tlb_req_bits_vaddr; // @[MemBlock.scala 249:24 464:25]
  assign dtlb_st_tlb_st_io_ptw_resp_valid = ptw_resp_v & |vector_hit_hi; // @[MemBlock.scala 299:52]
  assign dtlb_st_tlb_st_io_ptw_resp_bits_entry_tag = ptw_resp_next_data_entry_tag; // @[MemBlock.scala 249:24 294:32]
  assign dtlb_st_tlb_st_io_ptw_resp_bits_entry_asid = ptw_resp_next_data_entry_asid; // @[MemBlock.scala 249:24 294:32]
  assign dtlb_st_tlb_st_io_ptw_resp_bits_entry_ppn = ptw_resp_next_data_entry_ppn; // @[MemBlock.scala 249:24 294:32]
  assign dtlb_st_tlb_st_io_ptw_resp_bits_entry_perm_d = ptw_resp_next_data_entry_perm_d; // @[MemBlock.scala 249:24 294:32]
  assign dtlb_st_tlb_st_io_ptw_resp_bits_entry_perm_a = ptw_resp_next_data_entry_perm_a; // @[MemBlock.scala 249:24 294:32]
  assign dtlb_st_tlb_st_io_ptw_resp_bits_entry_perm_g = ptw_resp_next_data_entry_perm_g; // @[MemBlock.scala 249:24 294:32]
  assign dtlb_st_tlb_st_io_ptw_resp_bits_entry_perm_u = ptw_resp_next_data_entry_perm_u; // @[MemBlock.scala 249:24 294:32]
  assign dtlb_st_tlb_st_io_ptw_resp_bits_entry_perm_x = ptw_resp_next_data_entry_perm_x; // @[MemBlock.scala 249:24 294:32]
  assign dtlb_st_tlb_st_io_ptw_resp_bits_entry_perm_w = ptw_resp_next_data_entry_perm_w; // @[MemBlock.scala 249:24 294:32]
  assign dtlb_st_tlb_st_io_ptw_resp_bits_entry_perm_r = ptw_resp_next_data_entry_perm_r; // @[MemBlock.scala 249:24 294:32]
  assign dtlb_st_tlb_st_io_ptw_resp_bits_entry_level = ptw_resp_next_data_entry_level; // @[MemBlock.scala 249:24 294:32]
  assign dtlb_st_tlb_st_io_ptw_resp_bits_pf = ptw_resp_next_data_pf; // @[MemBlock.scala 249:24 294:32]
  assign dtlb_st_tlb_st_io_ptw_resp_bits_af = ptw_resp_next_data_af; // @[MemBlock.scala 249:24 294:32]
  assign dtlb_st_tlb_st_io_ptw_replenish_c = pmp_check_ptw_io_resp_c; // @[MemBlock.scala 249:24 322:28]
  assign dtlb_st_tlb_st_io_ptw_replenish_atomic = pmp_check_ptw_io_resp_atomic; // @[MemBlock.scala 249:24 322:28]
  assign dtlb_st_tlb_st_io_ptw_replenish_x = pmp_check_ptw_io_resp_x; // @[MemBlock.scala 249:24 322:28]
  assign dtlb_st_tlb_st_io_ptw_replenish_w = pmp_check_ptw_io_resp_w; // @[MemBlock.scala 249:24 322:28]
  assign dtlb_st_tlb_st_io_ptw_replenish_r = pmp_check_ptw_io_resp_r; // @[MemBlock.scala 249:24 322:28]
  assign dtlb_prefetch_tlb_prefetch_clock = clock;
  assign dtlb_prefetch_tlb_prefetch_io_sfence_valid = sfence_valid; // @[MemBlock.scala 253:30 260:21]
  assign dtlb_prefetch_tlb_prefetch_io_sfence_bits_rs1 = sfence_bits_rs1; // @[MemBlock.scala 253:30 260:21]
  assign dtlb_prefetch_tlb_prefetch_io_sfence_bits_rs2 = sfence_bits_rs2; // @[MemBlock.scala 253:30 260:21]
  assign dtlb_prefetch_tlb_prefetch_io_sfence_bits_addr = sfence_bits_addr; // @[MemBlock.scala 253:30 260:21]
  assign dtlb_prefetch_tlb_prefetch_io_sfence_bits_asid = sfence_bits_asid; // @[MemBlock.scala 253:30 260:21]
  assign dtlb_prefetch_tlb_prefetch_io_csr_satp_mode = tlbcsr_satp_mode; // @[MemBlock.scala 253:30 261:18]
  assign dtlb_prefetch_tlb_prefetch_io_csr_satp_asid = tlbcsr_satp_asid; // @[MemBlock.scala 253:30 261:18]
  assign dtlb_prefetch_tlb_prefetch_io_csr_satp_changed = tlbcsr_satp_changed; // @[MemBlock.scala 253:30 261:18]
  assign dtlb_prefetch_tlb_prefetch_io_csr_priv_dmode = tlbcsr_priv_dmode; // @[MemBlock.scala 253:30 261:18]
  assign dtlb_prefetch_tlb_prefetch_io_ptw_resp_valid = ptw_resp_v & |ptw_resp_next_vector_4; // @[MemBlock.scala 300:58]
  assign dtlb_prefetch_tlb_prefetch_io_ptw_resp_bits_entry_tag = ptw_resp_next_data_entry_tag; // @[MemBlock.scala 253:30 294:32]
  assign dtlb_prefetch_tlb_prefetch_io_ptw_resp_bits_entry_asid = ptw_resp_next_data_entry_asid; // @[MemBlock.scala 253:30 294:32]
  assign dtlb_prefetch_tlb_prefetch_io_ptw_resp_bits_entry_ppn = ptw_resp_next_data_entry_ppn; // @[MemBlock.scala 253:30 294:32]
  assign dtlb_prefetch_tlb_prefetch_io_ptw_resp_bits_entry_level = ptw_resp_next_data_entry_level; // @[MemBlock.scala 253:30 294:32]
  assign pmp_clock = clock;
  assign pmp_reset = reset;
  assign pmp_io_distribute_csr_wvalid = csrCtrl_delay_io_out_distribute_csr_wvalid; // @[MemBlock.scala 312:25]
  assign pmp_io_distribute_csr_waddr = csrCtrl_delay_io_out_distribute_csr_waddr; // @[MemBlock.scala 312:25]
  assign pmp_io_distribute_csr_wdata = csrCtrl_delay_io_out_distribute_csr_wdata; // @[MemBlock.scala 312:25]
  assign PMPChecker_clock = clock;
  assign PMPChecker_io_check_env_mode = tlbcsr_priv_dmode; // @[MemBlock.scala 314:26 PMP.scala 465:15]
  assign PMPChecker_io_check_env_pmp_0_cfg_l = pmp_io_pmp_0_cfg_l; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_0_cfg_a = pmp_io_pmp_0_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_0_cfg_w = pmp_io_pmp_0_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_0_cfg_r = pmp_io_pmp_0_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_0_addr = pmp_io_pmp_0_addr; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_0_mask = pmp_io_pmp_0_mask; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_1_cfg_l = pmp_io_pmp_1_cfg_l; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_1_cfg_a = pmp_io_pmp_1_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_1_cfg_w = pmp_io_pmp_1_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_1_cfg_r = pmp_io_pmp_1_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_1_addr = pmp_io_pmp_1_addr; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_1_mask = pmp_io_pmp_1_mask; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_2_cfg_l = pmp_io_pmp_2_cfg_l; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_2_cfg_a = pmp_io_pmp_2_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_2_cfg_w = pmp_io_pmp_2_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_2_cfg_r = pmp_io_pmp_2_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_2_addr = pmp_io_pmp_2_addr; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_2_mask = pmp_io_pmp_2_mask; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_3_cfg_l = pmp_io_pmp_3_cfg_l; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_3_cfg_a = pmp_io_pmp_3_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_3_cfg_w = pmp_io_pmp_3_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_3_cfg_r = pmp_io_pmp_3_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_3_addr = pmp_io_pmp_3_addr; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_3_mask = pmp_io_pmp_3_mask; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_4_cfg_l = pmp_io_pmp_4_cfg_l; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_4_cfg_a = pmp_io_pmp_4_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_4_cfg_w = pmp_io_pmp_4_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_4_cfg_r = pmp_io_pmp_4_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_4_addr = pmp_io_pmp_4_addr; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_4_mask = pmp_io_pmp_4_mask; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_5_cfg_l = pmp_io_pmp_5_cfg_l; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_5_cfg_a = pmp_io_pmp_5_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_5_cfg_w = pmp_io_pmp_5_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_5_cfg_r = pmp_io_pmp_5_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_5_addr = pmp_io_pmp_5_addr; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_5_mask = pmp_io_pmp_5_mask; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_6_cfg_l = pmp_io_pmp_6_cfg_l; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_6_cfg_a = pmp_io_pmp_6_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_6_cfg_w = pmp_io_pmp_6_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_6_cfg_r = pmp_io_pmp_6_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_6_addr = pmp_io_pmp_6_addr; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_6_mask = pmp_io_pmp_6_mask; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_7_cfg_l = pmp_io_pmp_7_cfg_l; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_7_cfg_a = pmp_io_pmp_7_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_7_cfg_w = pmp_io_pmp_7_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_7_cfg_r = pmp_io_pmp_7_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_7_addr = pmp_io_pmp_7_addr; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_7_mask = pmp_io_pmp_7_mask; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_8_cfg_l = pmp_io_pmp_8_cfg_l; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_8_cfg_a = pmp_io_pmp_8_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_8_cfg_w = pmp_io_pmp_8_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_8_cfg_r = pmp_io_pmp_8_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_8_addr = pmp_io_pmp_8_addr; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_8_mask = pmp_io_pmp_8_mask; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_9_cfg_l = pmp_io_pmp_9_cfg_l; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_9_cfg_a = pmp_io_pmp_9_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_9_cfg_w = pmp_io_pmp_9_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_9_cfg_r = pmp_io_pmp_9_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_9_addr = pmp_io_pmp_9_addr; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_9_mask = pmp_io_pmp_9_mask; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_10_cfg_l = pmp_io_pmp_10_cfg_l; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_10_cfg_a = pmp_io_pmp_10_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_10_cfg_w = pmp_io_pmp_10_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_10_cfg_r = pmp_io_pmp_10_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_10_addr = pmp_io_pmp_10_addr; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_10_mask = pmp_io_pmp_10_mask; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_11_cfg_l = pmp_io_pmp_11_cfg_l; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_11_cfg_a = pmp_io_pmp_11_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_11_cfg_w = pmp_io_pmp_11_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_11_cfg_r = pmp_io_pmp_11_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_11_addr = pmp_io_pmp_11_addr; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_11_mask = pmp_io_pmp_11_mask; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_12_cfg_l = pmp_io_pmp_12_cfg_l; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_12_cfg_a = pmp_io_pmp_12_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_12_cfg_w = pmp_io_pmp_12_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_12_cfg_r = pmp_io_pmp_12_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_12_addr = pmp_io_pmp_12_addr; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_12_mask = pmp_io_pmp_12_mask; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_13_cfg_l = pmp_io_pmp_13_cfg_l; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_13_cfg_a = pmp_io_pmp_13_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_13_cfg_w = pmp_io_pmp_13_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_13_cfg_r = pmp_io_pmp_13_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_13_addr = pmp_io_pmp_13_addr; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_13_mask = pmp_io_pmp_13_mask; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_14_cfg_l = pmp_io_pmp_14_cfg_l; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_14_cfg_a = pmp_io_pmp_14_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_14_cfg_w = pmp_io_pmp_14_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_14_cfg_r = pmp_io_pmp_14_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_14_addr = pmp_io_pmp_14_addr; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_14_mask = pmp_io_pmp_14_mask; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_15_cfg_l = pmp_io_pmp_15_cfg_l; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_15_cfg_a = pmp_io_pmp_15_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_15_cfg_w = pmp_io_pmp_15_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_15_cfg_r = pmp_io_pmp_15_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_15_addr = pmp_io_pmp_15_addr; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pmp_15_mask = pmp_io_pmp_15_mask; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_io_check_env_pma_0_cfg_c = pmp_io_pma_0_cfg_c; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_0_cfg_atomic = pmp_io_pma_0_cfg_atomic; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_0_cfg_a = pmp_io_pma_0_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_0_cfg_w = pmp_io_pma_0_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_0_cfg_r = pmp_io_pma_0_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_0_addr = pmp_io_pma_0_addr; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_0_mask = pmp_io_pma_0_mask; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_1_cfg_c = pmp_io_pma_1_cfg_c; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_1_cfg_atomic = pmp_io_pma_1_cfg_atomic; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_1_cfg_a = pmp_io_pma_1_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_1_cfg_w = pmp_io_pma_1_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_1_cfg_r = pmp_io_pma_1_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_1_addr = pmp_io_pma_1_addr; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_1_mask = pmp_io_pma_1_mask; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_2_cfg_c = pmp_io_pma_2_cfg_c; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_2_cfg_atomic = pmp_io_pma_2_cfg_atomic; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_2_cfg_a = pmp_io_pma_2_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_2_cfg_w = pmp_io_pma_2_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_2_cfg_r = pmp_io_pma_2_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_2_addr = pmp_io_pma_2_addr; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_2_mask = pmp_io_pma_2_mask; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_3_cfg_c = pmp_io_pma_3_cfg_c; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_3_cfg_atomic = pmp_io_pma_3_cfg_atomic; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_3_cfg_a = pmp_io_pma_3_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_3_cfg_w = pmp_io_pma_3_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_3_cfg_r = pmp_io_pma_3_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_3_addr = pmp_io_pma_3_addr; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_3_mask = pmp_io_pma_3_mask; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_4_cfg_c = pmp_io_pma_4_cfg_c; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_4_cfg_atomic = pmp_io_pma_4_cfg_atomic; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_4_cfg_a = pmp_io_pma_4_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_4_cfg_w = pmp_io_pma_4_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_4_cfg_r = pmp_io_pma_4_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_4_addr = pmp_io_pma_4_addr; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_4_mask = pmp_io_pma_4_mask; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_5_cfg_c = pmp_io_pma_5_cfg_c; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_5_cfg_atomic = pmp_io_pma_5_cfg_atomic; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_5_cfg_a = pmp_io_pma_5_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_5_cfg_w = pmp_io_pma_5_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_5_cfg_r = pmp_io_pma_5_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_5_addr = pmp_io_pma_5_addr; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_5_mask = pmp_io_pma_5_mask; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_6_cfg_c = pmp_io_pma_6_cfg_c; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_6_cfg_atomic = pmp_io_pma_6_cfg_atomic; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_6_cfg_a = pmp_io_pma_6_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_6_cfg_w = pmp_io_pma_6_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_6_cfg_r = pmp_io_pma_6_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_6_addr = pmp_io_pma_6_addr; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_6_mask = pmp_io_pma_6_mask; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_7_cfg_c = pmp_io_pma_7_cfg_c; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_7_cfg_atomic = pmp_io_pma_7_cfg_atomic; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_7_cfg_a = pmp_io_pma_7_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_7_cfg_w = pmp_io_pma_7_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_7_cfg_r = pmp_io_pma_7_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_7_addr = pmp_io_pma_7_addr; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_7_mask = pmp_io_pma_7_mask; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_8_cfg_c = pmp_io_pma_8_cfg_c; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_8_cfg_atomic = pmp_io_pma_8_cfg_atomic; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_8_cfg_a = pmp_io_pma_8_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_8_cfg_w = pmp_io_pma_8_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_8_cfg_r = pmp_io_pma_8_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_8_addr = pmp_io_pma_8_addr; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_8_mask = pmp_io_pma_8_mask; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_9_cfg_c = pmp_io_pma_9_cfg_c; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_9_cfg_atomic = pmp_io_pma_9_cfg_atomic; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_9_cfg_a = pmp_io_pma_9_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_9_cfg_w = pmp_io_pma_9_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_9_cfg_r = pmp_io_pma_9_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_9_addr = pmp_io_pma_9_addr; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_9_mask = pmp_io_pma_9_mask; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_10_cfg_c = pmp_io_pma_10_cfg_c; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_10_cfg_atomic = pmp_io_pma_10_cfg_atomic; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_10_cfg_a = pmp_io_pma_10_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_10_cfg_w = pmp_io_pma_10_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_10_cfg_r = pmp_io_pma_10_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_10_addr = pmp_io_pma_10_addr; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_10_mask = pmp_io_pma_10_mask; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_11_cfg_c = pmp_io_pma_11_cfg_c; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_11_cfg_atomic = pmp_io_pma_11_cfg_atomic; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_11_cfg_a = pmp_io_pma_11_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_11_cfg_w = pmp_io_pma_11_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_11_cfg_r = pmp_io_pma_11_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_11_addr = pmp_io_pma_11_addr; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_11_mask = pmp_io_pma_11_mask; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_12_cfg_c = pmp_io_pma_12_cfg_c; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_12_cfg_atomic = pmp_io_pma_12_cfg_atomic; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_12_cfg_a = pmp_io_pma_12_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_12_cfg_w = pmp_io_pma_12_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_12_cfg_r = pmp_io_pma_12_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_12_addr = pmp_io_pma_12_addr; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_12_mask = pmp_io_pma_12_mask; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_13_cfg_c = pmp_io_pma_13_cfg_c; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_13_cfg_atomic = pmp_io_pma_13_cfg_atomic; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_13_cfg_a = pmp_io_pma_13_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_13_cfg_w = pmp_io_pma_13_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_13_cfg_r = pmp_io_pma_13_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_13_addr = pmp_io_pma_13_addr; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_13_mask = pmp_io_pma_13_mask; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_14_cfg_c = pmp_io_pma_14_cfg_c; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_14_cfg_atomic = pmp_io_pma_14_cfg_atomic; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_14_cfg_a = pmp_io_pma_14_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_14_cfg_w = pmp_io_pma_14_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_14_cfg_r = pmp_io_pma_14_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_14_addr = pmp_io_pma_14_addr; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_14_mask = pmp_io_pma_14_mask; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_15_cfg_c = pmp_io_pma_15_cfg_c; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_15_cfg_atomic = pmp_io_pma_15_cfg_atomic; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_15_cfg_a = pmp_io_pma_15_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_15_cfg_w = pmp_io_pma_15_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_15_cfg_r = pmp_io_pma_15_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_15_addr = pmp_io_pma_15_addr; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_check_env_pma_15_mask = pmp_io_pma_15_mask; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_io_req_valid = dtlb_ld_tlb_ld_io_pmp_0_valid; // @[MemBlock.scala 245:{24,24}]
  assign PMPChecker_io_req_bits_addr = dtlb_ld_tlb_ld_io_pmp_0_bits_addr; // @[MemBlock.scala 245:{24,24}]
  assign PMPChecker_io_req_bits_cmd = dtlb_ld_tlb_ld_io_pmp_0_bits_cmd; // @[MemBlock.scala 245:{24,24}]
  assign PMPChecker_1_clock = clock;
  assign PMPChecker_1_io_check_env_mode = tlbcsr_priv_dmode; // @[MemBlock.scala 314:26 PMP.scala 465:15]
  assign PMPChecker_1_io_check_env_pmp_0_cfg_l = pmp_io_pmp_0_cfg_l; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_0_cfg_a = pmp_io_pmp_0_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_0_cfg_w = pmp_io_pmp_0_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_0_cfg_r = pmp_io_pmp_0_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_0_addr = pmp_io_pmp_0_addr; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_0_mask = pmp_io_pmp_0_mask; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_1_cfg_l = pmp_io_pmp_1_cfg_l; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_1_cfg_a = pmp_io_pmp_1_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_1_cfg_w = pmp_io_pmp_1_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_1_cfg_r = pmp_io_pmp_1_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_1_addr = pmp_io_pmp_1_addr; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_1_mask = pmp_io_pmp_1_mask; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_2_cfg_l = pmp_io_pmp_2_cfg_l; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_2_cfg_a = pmp_io_pmp_2_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_2_cfg_w = pmp_io_pmp_2_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_2_cfg_r = pmp_io_pmp_2_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_2_addr = pmp_io_pmp_2_addr; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_2_mask = pmp_io_pmp_2_mask; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_3_cfg_l = pmp_io_pmp_3_cfg_l; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_3_cfg_a = pmp_io_pmp_3_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_3_cfg_w = pmp_io_pmp_3_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_3_cfg_r = pmp_io_pmp_3_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_3_addr = pmp_io_pmp_3_addr; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_3_mask = pmp_io_pmp_3_mask; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_4_cfg_l = pmp_io_pmp_4_cfg_l; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_4_cfg_a = pmp_io_pmp_4_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_4_cfg_w = pmp_io_pmp_4_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_4_cfg_r = pmp_io_pmp_4_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_4_addr = pmp_io_pmp_4_addr; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_4_mask = pmp_io_pmp_4_mask; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_5_cfg_l = pmp_io_pmp_5_cfg_l; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_5_cfg_a = pmp_io_pmp_5_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_5_cfg_w = pmp_io_pmp_5_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_5_cfg_r = pmp_io_pmp_5_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_5_addr = pmp_io_pmp_5_addr; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_5_mask = pmp_io_pmp_5_mask; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_6_cfg_l = pmp_io_pmp_6_cfg_l; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_6_cfg_a = pmp_io_pmp_6_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_6_cfg_w = pmp_io_pmp_6_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_6_cfg_r = pmp_io_pmp_6_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_6_addr = pmp_io_pmp_6_addr; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_6_mask = pmp_io_pmp_6_mask; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_7_cfg_l = pmp_io_pmp_7_cfg_l; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_7_cfg_a = pmp_io_pmp_7_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_7_cfg_w = pmp_io_pmp_7_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_7_cfg_r = pmp_io_pmp_7_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_7_addr = pmp_io_pmp_7_addr; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_7_mask = pmp_io_pmp_7_mask; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_8_cfg_l = pmp_io_pmp_8_cfg_l; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_8_cfg_a = pmp_io_pmp_8_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_8_cfg_w = pmp_io_pmp_8_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_8_cfg_r = pmp_io_pmp_8_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_8_addr = pmp_io_pmp_8_addr; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_8_mask = pmp_io_pmp_8_mask; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_9_cfg_l = pmp_io_pmp_9_cfg_l; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_9_cfg_a = pmp_io_pmp_9_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_9_cfg_w = pmp_io_pmp_9_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_9_cfg_r = pmp_io_pmp_9_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_9_addr = pmp_io_pmp_9_addr; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_9_mask = pmp_io_pmp_9_mask; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_10_cfg_l = pmp_io_pmp_10_cfg_l; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_10_cfg_a = pmp_io_pmp_10_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_10_cfg_w = pmp_io_pmp_10_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_10_cfg_r = pmp_io_pmp_10_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_10_addr = pmp_io_pmp_10_addr; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_10_mask = pmp_io_pmp_10_mask; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_11_cfg_l = pmp_io_pmp_11_cfg_l; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_11_cfg_a = pmp_io_pmp_11_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_11_cfg_w = pmp_io_pmp_11_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_11_cfg_r = pmp_io_pmp_11_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_11_addr = pmp_io_pmp_11_addr; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_11_mask = pmp_io_pmp_11_mask; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_12_cfg_l = pmp_io_pmp_12_cfg_l; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_12_cfg_a = pmp_io_pmp_12_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_12_cfg_w = pmp_io_pmp_12_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_12_cfg_r = pmp_io_pmp_12_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_12_addr = pmp_io_pmp_12_addr; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_12_mask = pmp_io_pmp_12_mask; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_13_cfg_l = pmp_io_pmp_13_cfg_l; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_13_cfg_a = pmp_io_pmp_13_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_13_cfg_w = pmp_io_pmp_13_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_13_cfg_r = pmp_io_pmp_13_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_13_addr = pmp_io_pmp_13_addr; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_13_mask = pmp_io_pmp_13_mask; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_14_cfg_l = pmp_io_pmp_14_cfg_l; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_14_cfg_a = pmp_io_pmp_14_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_14_cfg_w = pmp_io_pmp_14_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_14_cfg_r = pmp_io_pmp_14_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_14_addr = pmp_io_pmp_14_addr; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_14_mask = pmp_io_pmp_14_mask; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_15_cfg_l = pmp_io_pmp_15_cfg_l; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_15_cfg_a = pmp_io_pmp_15_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_15_cfg_w = pmp_io_pmp_15_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_15_cfg_r = pmp_io_pmp_15_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_15_addr = pmp_io_pmp_15_addr; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pmp_15_mask = pmp_io_pmp_15_mask; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_1_io_check_env_pma_0_cfg_c = pmp_io_pma_0_cfg_c; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_0_cfg_atomic = pmp_io_pma_0_cfg_atomic; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_0_cfg_a = pmp_io_pma_0_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_0_cfg_w = pmp_io_pma_0_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_0_cfg_r = pmp_io_pma_0_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_0_addr = pmp_io_pma_0_addr; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_0_mask = pmp_io_pma_0_mask; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_1_cfg_c = pmp_io_pma_1_cfg_c; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_1_cfg_atomic = pmp_io_pma_1_cfg_atomic; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_1_cfg_a = pmp_io_pma_1_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_1_cfg_w = pmp_io_pma_1_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_1_cfg_r = pmp_io_pma_1_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_1_addr = pmp_io_pma_1_addr; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_1_mask = pmp_io_pma_1_mask; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_2_cfg_c = pmp_io_pma_2_cfg_c; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_2_cfg_atomic = pmp_io_pma_2_cfg_atomic; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_2_cfg_a = pmp_io_pma_2_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_2_cfg_w = pmp_io_pma_2_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_2_cfg_r = pmp_io_pma_2_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_2_addr = pmp_io_pma_2_addr; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_2_mask = pmp_io_pma_2_mask; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_3_cfg_c = pmp_io_pma_3_cfg_c; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_3_cfg_atomic = pmp_io_pma_3_cfg_atomic; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_3_cfg_a = pmp_io_pma_3_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_3_cfg_w = pmp_io_pma_3_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_3_cfg_r = pmp_io_pma_3_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_3_addr = pmp_io_pma_3_addr; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_3_mask = pmp_io_pma_3_mask; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_4_cfg_c = pmp_io_pma_4_cfg_c; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_4_cfg_atomic = pmp_io_pma_4_cfg_atomic; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_4_cfg_a = pmp_io_pma_4_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_4_cfg_w = pmp_io_pma_4_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_4_cfg_r = pmp_io_pma_4_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_4_addr = pmp_io_pma_4_addr; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_4_mask = pmp_io_pma_4_mask; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_5_cfg_c = pmp_io_pma_5_cfg_c; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_5_cfg_atomic = pmp_io_pma_5_cfg_atomic; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_5_cfg_a = pmp_io_pma_5_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_5_cfg_w = pmp_io_pma_5_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_5_cfg_r = pmp_io_pma_5_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_5_addr = pmp_io_pma_5_addr; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_5_mask = pmp_io_pma_5_mask; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_6_cfg_c = pmp_io_pma_6_cfg_c; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_6_cfg_atomic = pmp_io_pma_6_cfg_atomic; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_6_cfg_a = pmp_io_pma_6_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_6_cfg_w = pmp_io_pma_6_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_6_cfg_r = pmp_io_pma_6_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_6_addr = pmp_io_pma_6_addr; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_6_mask = pmp_io_pma_6_mask; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_7_cfg_c = pmp_io_pma_7_cfg_c; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_7_cfg_atomic = pmp_io_pma_7_cfg_atomic; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_7_cfg_a = pmp_io_pma_7_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_7_cfg_w = pmp_io_pma_7_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_7_cfg_r = pmp_io_pma_7_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_7_addr = pmp_io_pma_7_addr; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_7_mask = pmp_io_pma_7_mask; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_8_cfg_c = pmp_io_pma_8_cfg_c; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_8_cfg_atomic = pmp_io_pma_8_cfg_atomic; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_8_cfg_a = pmp_io_pma_8_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_8_cfg_w = pmp_io_pma_8_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_8_cfg_r = pmp_io_pma_8_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_8_addr = pmp_io_pma_8_addr; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_8_mask = pmp_io_pma_8_mask; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_9_cfg_c = pmp_io_pma_9_cfg_c; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_9_cfg_atomic = pmp_io_pma_9_cfg_atomic; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_9_cfg_a = pmp_io_pma_9_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_9_cfg_w = pmp_io_pma_9_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_9_cfg_r = pmp_io_pma_9_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_9_addr = pmp_io_pma_9_addr; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_9_mask = pmp_io_pma_9_mask; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_10_cfg_c = pmp_io_pma_10_cfg_c; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_10_cfg_atomic = pmp_io_pma_10_cfg_atomic; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_10_cfg_a = pmp_io_pma_10_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_10_cfg_w = pmp_io_pma_10_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_10_cfg_r = pmp_io_pma_10_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_10_addr = pmp_io_pma_10_addr; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_10_mask = pmp_io_pma_10_mask; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_11_cfg_c = pmp_io_pma_11_cfg_c; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_11_cfg_atomic = pmp_io_pma_11_cfg_atomic; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_11_cfg_a = pmp_io_pma_11_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_11_cfg_w = pmp_io_pma_11_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_11_cfg_r = pmp_io_pma_11_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_11_addr = pmp_io_pma_11_addr; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_11_mask = pmp_io_pma_11_mask; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_12_cfg_c = pmp_io_pma_12_cfg_c; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_12_cfg_atomic = pmp_io_pma_12_cfg_atomic; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_12_cfg_a = pmp_io_pma_12_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_12_cfg_w = pmp_io_pma_12_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_12_cfg_r = pmp_io_pma_12_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_12_addr = pmp_io_pma_12_addr; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_12_mask = pmp_io_pma_12_mask; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_13_cfg_c = pmp_io_pma_13_cfg_c; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_13_cfg_atomic = pmp_io_pma_13_cfg_atomic; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_13_cfg_a = pmp_io_pma_13_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_13_cfg_w = pmp_io_pma_13_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_13_cfg_r = pmp_io_pma_13_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_13_addr = pmp_io_pma_13_addr; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_13_mask = pmp_io_pma_13_mask; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_14_cfg_c = pmp_io_pma_14_cfg_c; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_14_cfg_atomic = pmp_io_pma_14_cfg_atomic; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_14_cfg_a = pmp_io_pma_14_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_14_cfg_w = pmp_io_pma_14_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_14_cfg_r = pmp_io_pma_14_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_14_addr = pmp_io_pma_14_addr; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_14_mask = pmp_io_pma_14_mask; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_15_cfg_c = pmp_io_pma_15_cfg_c; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_15_cfg_atomic = pmp_io_pma_15_cfg_atomic; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_15_cfg_a = pmp_io_pma_15_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_15_cfg_w = pmp_io_pma_15_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_15_cfg_r = pmp_io_pma_15_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_15_addr = pmp_io_pma_15_addr; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_check_env_pma_15_mask = pmp_io_pma_15_mask; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_1_io_req_valid = dtlb_ld_tlb_ld_io_pmp_1_valid; // @[MemBlock.scala 245:{24,24}]
  assign PMPChecker_1_io_req_bits_addr = dtlb_ld_tlb_ld_io_pmp_1_bits_addr; // @[MemBlock.scala 245:{24,24}]
  assign PMPChecker_1_io_req_bits_cmd = dtlb_ld_tlb_ld_io_pmp_1_bits_cmd; // @[MemBlock.scala 245:{24,24}]
  assign PMPChecker_2_clock = clock;
  assign PMPChecker_2_io_check_env_mode = tlbcsr_priv_dmode; // @[MemBlock.scala 314:26 PMP.scala 465:15]
  assign PMPChecker_2_io_check_env_pmp_0_cfg_l = pmp_io_pmp_0_cfg_l; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_0_cfg_a = pmp_io_pmp_0_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_0_cfg_w = pmp_io_pmp_0_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_0_cfg_r = pmp_io_pmp_0_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_0_addr = pmp_io_pmp_0_addr; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_0_mask = pmp_io_pmp_0_mask; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_1_cfg_l = pmp_io_pmp_1_cfg_l; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_1_cfg_a = pmp_io_pmp_1_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_1_cfg_w = pmp_io_pmp_1_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_1_cfg_r = pmp_io_pmp_1_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_1_addr = pmp_io_pmp_1_addr; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_1_mask = pmp_io_pmp_1_mask; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_2_cfg_l = pmp_io_pmp_2_cfg_l; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_2_cfg_a = pmp_io_pmp_2_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_2_cfg_w = pmp_io_pmp_2_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_2_cfg_r = pmp_io_pmp_2_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_2_addr = pmp_io_pmp_2_addr; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_2_mask = pmp_io_pmp_2_mask; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_3_cfg_l = pmp_io_pmp_3_cfg_l; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_3_cfg_a = pmp_io_pmp_3_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_3_cfg_w = pmp_io_pmp_3_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_3_cfg_r = pmp_io_pmp_3_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_3_addr = pmp_io_pmp_3_addr; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_3_mask = pmp_io_pmp_3_mask; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_4_cfg_l = pmp_io_pmp_4_cfg_l; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_4_cfg_a = pmp_io_pmp_4_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_4_cfg_w = pmp_io_pmp_4_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_4_cfg_r = pmp_io_pmp_4_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_4_addr = pmp_io_pmp_4_addr; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_4_mask = pmp_io_pmp_4_mask; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_5_cfg_l = pmp_io_pmp_5_cfg_l; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_5_cfg_a = pmp_io_pmp_5_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_5_cfg_w = pmp_io_pmp_5_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_5_cfg_r = pmp_io_pmp_5_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_5_addr = pmp_io_pmp_5_addr; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_5_mask = pmp_io_pmp_5_mask; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_6_cfg_l = pmp_io_pmp_6_cfg_l; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_6_cfg_a = pmp_io_pmp_6_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_6_cfg_w = pmp_io_pmp_6_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_6_cfg_r = pmp_io_pmp_6_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_6_addr = pmp_io_pmp_6_addr; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_6_mask = pmp_io_pmp_6_mask; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_7_cfg_l = pmp_io_pmp_7_cfg_l; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_7_cfg_a = pmp_io_pmp_7_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_7_cfg_w = pmp_io_pmp_7_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_7_cfg_r = pmp_io_pmp_7_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_7_addr = pmp_io_pmp_7_addr; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_7_mask = pmp_io_pmp_7_mask; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_8_cfg_l = pmp_io_pmp_8_cfg_l; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_8_cfg_a = pmp_io_pmp_8_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_8_cfg_w = pmp_io_pmp_8_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_8_cfg_r = pmp_io_pmp_8_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_8_addr = pmp_io_pmp_8_addr; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_8_mask = pmp_io_pmp_8_mask; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_9_cfg_l = pmp_io_pmp_9_cfg_l; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_9_cfg_a = pmp_io_pmp_9_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_9_cfg_w = pmp_io_pmp_9_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_9_cfg_r = pmp_io_pmp_9_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_9_addr = pmp_io_pmp_9_addr; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_9_mask = pmp_io_pmp_9_mask; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_10_cfg_l = pmp_io_pmp_10_cfg_l; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_10_cfg_a = pmp_io_pmp_10_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_10_cfg_w = pmp_io_pmp_10_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_10_cfg_r = pmp_io_pmp_10_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_10_addr = pmp_io_pmp_10_addr; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_10_mask = pmp_io_pmp_10_mask; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_11_cfg_l = pmp_io_pmp_11_cfg_l; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_11_cfg_a = pmp_io_pmp_11_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_11_cfg_w = pmp_io_pmp_11_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_11_cfg_r = pmp_io_pmp_11_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_11_addr = pmp_io_pmp_11_addr; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_11_mask = pmp_io_pmp_11_mask; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_12_cfg_l = pmp_io_pmp_12_cfg_l; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_12_cfg_a = pmp_io_pmp_12_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_12_cfg_w = pmp_io_pmp_12_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_12_cfg_r = pmp_io_pmp_12_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_12_addr = pmp_io_pmp_12_addr; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_12_mask = pmp_io_pmp_12_mask; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_13_cfg_l = pmp_io_pmp_13_cfg_l; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_13_cfg_a = pmp_io_pmp_13_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_13_cfg_w = pmp_io_pmp_13_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_13_cfg_r = pmp_io_pmp_13_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_13_addr = pmp_io_pmp_13_addr; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_13_mask = pmp_io_pmp_13_mask; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_14_cfg_l = pmp_io_pmp_14_cfg_l; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_14_cfg_a = pmp_io_pmp_14_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_14_cfg_w = pmp_io_pmp_14_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_14_cfg_r = pmp_io_pmp_14_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_14_addr = pmp_io_pmp_14_addr; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_14_mask = pmp_io_pmp_14_mask; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_15_cfg_l = pmp_io_pmp_15_cfg_l; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_15_cfg_a = pmp_io_pmp_15_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_15_cfg_w = pmp_io_pmp_15_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_15_cfg_r = pmp_io_pmp_15_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_15_addr = pmp_io_pmp_15_addr; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pmp_15_mask = pmp_io_pmp_15_mask; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_2_io_check_env_pma_0_cfg_c = pmp_io_pma_0_cfg_c; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_0_cfg_atomic = pmp_io_pma_0_cfg_atomic; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_0_cfg_a = pmp_io_pma_0_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_0_cfg_w = pmp_io_pma_0_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_0_cfg_r = pmp_io_pma_0_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_0_addr = pmp_io_pma_0_addr; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_0_mask = pmp_io_pma_0_mask; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_1_cfg_c = pmp_io_pma_1_cfg_c; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_1_cfg_atomic = pmp_io_pma_1_cfg_atomic; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_1_cfg_a = pmp_io_pma_1_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_1_cfg_w = pmp_io_pma_1_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_1_cfg_r = pmp_io_pma_1_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_1_addr = pmp_io_pma_1_addr; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_1_mask = pmp_io_pma_1_mask; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_2_cfg_c = pmp_io_pma_2_cfg_c; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_2_cfg_atomic = pmp_io_pma_2_cfg_atomic; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_2_cfg_a = pmp_io_pma_2_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_2_cfg_w = pmp_io_pma_2_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_2_cfg_r = pmp_io_pma_2_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_2_addr = pmp_io_pma_2_addr; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_2_mask = pmp_io_pma_2_mask; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_3_cfg_c = pmp_io_pma_3_cfg_c; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_3_cfg_atomic = pmp_io_pma_3_cfg_atomic; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_3_cfg_a = pmp_io_pma_3_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_3_cfg_w = pmp_io_pma_3_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_3_cfg_r = pmp_io_pma_3_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_3_addr = pmp_io_pma_3_addr; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_3_mask = pmp_io_pma_3_mask; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_4_cfg_c = pmp_io_pma_4_cfg_c; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_4_cfg_atomic = pmp_io_pma_4_cfg_atomic; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_4_cfg_a = pmp_io_pma_4_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_4_cfg_w = pmp_io_pma_4_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_4_cfg_r = pmp_io_pma_4_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_4_addr = pmp_io_pma_4_addr; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_4_mask = pmp_io_pma_4_mask; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_5_cfg_c = pmp_io_pma_5_cfg_c; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_5_cfg_atomic = pmp_io_pma_5_cfg_atomic; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_5_cfg_a = pmp_io_pma_5_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_5_cfg_w = pmp_io_pma_5_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_5_cfg_r = pmp_io_pma_5_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_5_addr = pmp_io_pma_5_addr; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_5_mask = pmp_io_pma_5_mask; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_6_cfg_c = pmp_io_pma_6_cfg_c; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_6_cfg_atomic = pmp_io_pma_6_cfg_atomic; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_6_cfg_a = pmp_io_pma_6_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_6_cfg_w = pmp_io_pma_6_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_6_cfg_r = pmp_io_pma_6_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_6_addr = pmp_io_pma_6_addr; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_6_mask = pmp_io_pma_6_mask; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_7_cfg_c = pmp_io_pma_7_cfg_c; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_7_cfg_atomic = pmp_io_pma_7_cfg_atomic; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_7_cfg_a = pmp_io_pma_7_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_7_cfg_w = pmp_io_pma_7_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_7_cfg_r = pmp_io_pma_7_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_7_addr = pmp_io_pma_7_addr; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_7_mask = pmp_io_pma_7_mask; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_8_cfg_c = pmp_io_pma_8_cfg_c; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_8_cfg_atomic = pmp_io_pma_8_cfg_atomic; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_8_cfg_a = pmp_io_pma_8_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_8_cfg_w = pmp_io_pma_8_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_8_cfg_r = pmp_io_pma_8_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_8_addr = pmp_io_pma_8_addr; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_8_mask = pmp_io_pma_8_mask; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_9_cfg_c = pmp_io_pma_9_cfg_c; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_9_cfg_atomic = pmp_io_pma_9_cfg_atomic; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_9_cfg_a = pmp_io_pma_9_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_9_cfg_w = pmp_io_pma_9_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_9_cfg_r = pmp_io_pma_9_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_9_addr = pmp_io_pma_9_addr; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_9_mask = pmp_io_pma_9_mask; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_10_cfg_c = pmp_io_pma_10_cfg_c; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_10_cfg_atomic = pmp_io_pma_10_cfg_atomic; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_10_cfg_a = pmp_io_pma_10_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_10_cfg_w = pmp_io_pma_10_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_10_cfg_r = pmp_io_pma_10_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_10_addr = pmp_io_pma_10_addr; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_10_mask = pmp_io_pma_10_mask; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_11_cfg_c = pmp_io_pma_11_cfg_c; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_11_cfg_atomic = pmp_io_pma_11_cfg_atomic; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_11_cfg_a = pmp_io_pma_11_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_11_cfg_w = pmp_io_pma_11_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_11_cfg_r = pmp_io_pma_11_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_11_addr = pmp_io_pma_11_addr; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_11_mask = pmp_io_pma_11_mask; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_12_cfg_c = pmp_io_pma_12_cfg_c; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_12_cfg_atomic = pmp_io_pma_12_cfg_atomic; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_12_cfg_a = pmp_io_pma_12_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_12_cfg_w = pmp_io_pma_12_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_12_cfg_r = pmp_io_pma_12_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_12_addr = pmp_io_pma_12_addr; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_12_mask = pmp_io_pma_12_mask; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_13_cfg_c = pmp_io_pma_13_cfg_c; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_13_cfg_atomic = pmp_io_pma_13_cfg_atomic; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_13_cfg_a = pmp_io_pma_13_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_13_cfg_w = pmp_io_pma_13_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_13_cfg_r = pmp_io_pma_13_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_13_addr = pmp_io_pma_13_addr; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_13_mask = pmp_io_pma_13_mask; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_14_cfg_c = pmp_io_pma_14_cfg_c; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_14_cfg_atomic = pmp_io_pma_14_cfg_atomic; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_14_cfg_a = pmp_io_pma_14_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_14_cfg_w = pmp_io_pma_14_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_14_cfg_r = pmp_io_pma_14_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_14_addr = pmp_io_pma_14_addr; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_14_mask = pmp_io_pma_14_mask; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_15_cfg_c = pmp_io_pma_15_cfg_c; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_15_cfg_atomic = pmp_io_pma_15_cfg_atomic; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_15_cfg_a = pmp_io_pma_15_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_15_cfg_w = pmp_io_pma_15_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_15_cfg_r = pmp_io_pma_15_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_15_addr = pmp_io_pma_15_addr; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_check_env_pma_15_mask = pmp_io_pma_15_mask; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_2_io_req_valid = dtlb_st_tlb_st_io_pmp_0_valid; // @[MemBlock.scala 249:{24,24}]
  assign PMPChecker_2_io_req_bits_addr = dtlb_st_tlb_st_io_pmp_0_bits_addr; // @[MemBlock.scala 249:{24,24}]
  assign PMPChecker_2_io_req_bits_cmd = 3'h1; // @[MemBlock.scala 249:{24,24}]
  assign PMPChecker_3_clock = clock;
  assign PMPChecker_3_io_check_env_mode = tlbcsr_priv_dmode; // @[MemBlock.scala 314:26 PMP.scala 465:15]
  assign PMPChecker_3_io_check_env_pmp_0_cfg_l = pmp_io_pmp_0_cfg_l; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_0_cfg_a = pmp_io_pmp_0_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_0_cfg_w = pmp_io_pmp_0_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_0_cfg_r = pmp_io_pmp_0_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_0_addr = pmp_io_pmp_0_addr; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_0_mask = pmp_io_pmp_0_mask; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_1_cfg_l = pmp_io_pmp_1_cfg_l; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_1_cfg_a = pmp_io_pmp_1_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_1_cfg_w = pmp_io_pmp_1_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_1_cfg_r = pmp_io_pmp_1_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_1_addr = pmp_io_pmp_1_addr; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_1_mask = pmp_io_pmp_1_mask; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_2_cfg_l = pmp_io_pmp_2_cfg_l; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_2_cfg_a = pmp_io_pmp_2_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_2_cfg_w = pmp_io_pmp_2_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_2_cfg_r = pmp_io_pmp_2_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_2_addr = pmp_io_pmp_2_addr; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_2_mask = pmp_io_pmp_2_mask; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_3_cfg_l = pmp_io_pmp_3_cfg_l; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_3_cfg_a = pmp_io_pmp_3_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_3_cfg_w = pmp_io_pmp_3_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_3_cfg_r = pmp_io_pmp_3_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_3_addr = pmp_io_pmp_3_addr; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_3_mask = pmp_io_pmp_3_mask; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_4_cfg_l = pmp_io_pmp_4_cfg_l; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_4_cfg_a = pmp_io_pmp_4_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_4_cfg_w = pmp_io_pmp_4_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_4_cfg_r = pmp_io_pmp_4_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_4_addr = pmp_io_pmp_4_addr; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_4_mask = pmp_io_pmp_4_mask; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_5_cfg_l = pmp_io_pmp_5_cfg_l; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_5_cfg_a = pmp_io_pmp_5_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_5_cfg_w = pmp_io_pmp_5_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_5_cfg_r = pmp_io_pmp_5_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_5_addr = pmp_io_pmp_5_addr; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_5_mask = pmp_io_pmp_5_mask; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_6_cfg_l = pmp_io_pmp_6_cfg_l; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_6_cfg_a = pmp_io_pmp_6_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_6_cfg_w = pmp_io_pmp_6_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_6_cfg_r = pmp_io_pmp_6_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_6_addr = pmp_io_pmp_6_addr; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_6_mask = pmp_io_pmp_6_mask; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_7_cfg_l = pmp_io_pmp_7_cfg_l; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_7_cfg_a = pmp_io_pmp_7_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_7_cfg_w = pmp_io_pmp_7_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_7_cfg_r = pmp_io_pmp_7_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_7_addr = pmp_io_pmp_7_addr; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_7_mask = pmp_io_pmp_7_mask; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_8_cfg_l = pmp_io_pmp_8_cfg_l; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_8_cfg_a = pmp_io_pmp_8_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_8_cfg_w = pmp_io_pmp_8_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_8_cfg_r = pmp_io_pmp_8_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_8_addr = pmp_io_pmp_8_addr; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_8_mask = pmp_io_pmp_8_mask; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_9_cfg_l = pmp_io_pmp_9_cfg_l; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_9_cfg_a = pmp_io_pmp_9_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_9_cfg_w = pmp_io_pmp_9_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_9_cfg_r = pmp_io_pmp_9_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_9_addr = pmp_io_pmp_9_addr; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_9_mask = pmp_io_pmp_9_mask; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_10_cfg_l = pmp_io_pmp_10_cfg_l; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_10_cfg_a = pmp_io_pmp_10_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_10_cfg_w = pmp_io_pmp_10_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_10_cfg_r = pmp_io_pmp_10_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_10_addr = pmp_io_pmp_10_addr; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_10_mask = pmp_io_pmp_10_mask; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_11_cfg_l = pmp_io_pmp_11_cfg_l; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_11_cfg_a = pmp_io_pmp_11_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_11_cfg_w = pmp_io_pmp_11_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_11_cfg_r = pmp_io_pmp_11_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_11_addr = pmp_io_pmp_11_addr; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_11_mask = pmp_io_pmp_11_mask; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_12_cfg_l = pmp_io_pmp_12_cfg_l; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_12_cfg_a = pmp_io_pmp_12_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_12_cfg_w = pmp_io_pmp_12_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_12_cfg_r = pmp_io_pmp_12_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_12_addr = pmp_io_pmp_12_addr; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_12_mask = pmp_io_pmp_12_mask; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_13_cfg_l = pmp_io_pmp_13_cfg_l; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_13_cfg_a = pmp_io_pmp_13_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_13_cfg_w = pmp_io_pmp_13_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_13_cfg_r = pmp_io_pmp_13_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_13_addr = pmp_io_pmp_13_addr; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_13_mask = pmp_io_pmp_13_mask; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_14_cfg_l = pmp_io_pmp_14_cfg_l; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_14_cfg_a = pmp_io_pmp_14_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_14_cfg_w = pmp_io_pmp_14_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_14_cfg_r = pmp_io_pmp_14_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_14_addr = pmp_io_pmp_14_addr; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_14_mask = pmp_io_pmp_14_mask; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_15_cfg_l = pmp_io_pmp_15_cfg_l; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_15_cfg_a = pmp_io_pmp_15_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_15_cfg_w = pmp_io_pmp_15_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_15_cfg_r = pmp_io_pmp_15_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_15_addr = pmp_io_pmp_15_addr; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pmp_15_mask = pmp_io_pmp_15_mask; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_3_io_check_env_pma_0_cfg_c = pmp_io_pma_0_cfg_c; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_0_cfg_atomic = pmp_io_pma_0_cfg_atomic; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_0_cfg_a = pmp_io_pma_0_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_0_cfg_w = pmp_io_pma_0_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_0_cfg_r = pmp_io_pma_0_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_0_addr = pmp_io_pma_0_addr; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_0_mask = pmp_io_pma_0_mask; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_1_cfg_c = pmp_io_pma_1_cfg_c; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_1_cfg_atomic = pmp_io_pma_1_cfg_atomic; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_1_cfg_a = pmp_io_pma_1_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_1_cfg_w = pmp_io_pma_1_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_1_cfg_r = pmp_io_pma_1_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_1_addr = pmp_io_pma_1_addr; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_1_mask = pmp_io_pma_1_mask; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_2_cfg_c = pmp_io_pma_2_cfg_c; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_2_cfg_atomic = pmp_io_pma_2_cfg_atomic; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_2_cfg_a = pmp_io_pma_2_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_2_cfg_w = pmp_io_pma_2_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_2_cfg_r = pmp_io_pma_2_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_2_addr = pmp_io_pma_2_addr; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_2_mask = pmp_io_pma_2_mask; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_3_cfg_c = pmp_io_pma_3_cfg_c; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_3_cfg_atomic = pmp_io_pma_3_cfg_atomic; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_3_cfg_a = pmp_io_pma_3_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_3_cfg_w = pmp_io_pma_3_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_3_cfg_r = pmp_io_pma_3_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_3_addr = pmp_io_pma_3_addr; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_3_mask = pmp_io_pma_3_mask; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_4_cfg_c = pmp_io_pma_4_cfg_c; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_4_cfg_atomic = pmp_io_pma_4_cfg_atomic; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_4_cfg_a = pmp_io_pma_4_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_4_cfg_w = pmp_io_pma_4_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_4_cfg_r = pmp_io_pma_4_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_4_addr = pmp_io_pma_4_addr; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_4_mask = pmp_io_pma_4_mask; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_5_cfg_c = pmp_io_pma_5_cfg_c; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_5_cfg_atomic = pmp_io_pma_5_cfg_atomic; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_5_cfg_a = pmp_io_pma_5_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_5_cfg_w = pmp_io_pma_5_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_5_cfg_r = pmp_io_pma_5_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_5_addr = pmp_io_pma_5_addr; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_5_mask = pmp_io_pma_5_mask; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_6_cfg_c = pmp_io_pma_6_cfg_c; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_6_cfg_atomic = pmp_io_pma_6_cfg_atomic; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_6_cfg_a = pmp_io_pma_6_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_6_cfg_w = pmp_io_pma_6_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_6_cfg_r = pmp_io_pma_6_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_6_addr = pmp_io_pma_6_addr; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_6_mask = pmp_io_pma_6_mask; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_7_cfg_c = pmp_io_pma_7_cfg_c; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_7_cfg_atomic = pmp_io_pma_7_cfg_atomic; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_7_cfg_a = pmp_io_pma_7_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_7_cfg_w = pmp_io_pma_7_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_7_cfg_r = pmp_io_pma_7_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_7_addr = pmp_io_pma_7_addr; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_7_mask = pmp_io_pma_7_mask; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_8_cfg_c = pmp_io_pma_8_cfg_c; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_8_cfg_atomic = pmp_io_pma_8_cfg_atomic; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_8_cfg_a = pmp_io_pma_8_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_8_cfg_w = pmp_io_pma_8_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_8_cfg_r = pmp_io_pma_8_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_8_addr = pmp_io_pma_8_addr; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_8_mask = pmp_io_pma_8_mask; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_9_cfg_c = pmp_io_pma_9_cfg_c; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_9_cfg_atomic = pmp_io_pma_9_cfg_atomic; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_9_cfg_a = pmp_io_pma_9_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_9_cfg_w = pmp_io_pma_9_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_9_cfg_r = pmp_io_pma_9_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_9_addr = pmp_io_pma_9_addr; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_9_mask = pmp_io_pma_9_mask; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_10_cfg_c = pmp_io_pma_10_cfg_c; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_10_cfg_atomic = pmp_io_pma_10_cfg_atomic; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_10_cfg_a = pmp_io_pma_10_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_10_cfg_w = pmp_io_pma_10_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_10_cfg_r = pmp_io_pma_10_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_10_addr = pmp_io_pma_10_addr; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_10_mask = pmp_io_pma_10_mask; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_11_cfg_c = pmp_io_pma_11_cfg_c; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_11_cfg_atomic = pmp_io_pma_11_cfg_atomic; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_11_cfg_a = pmp_io_pma_11_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_11_cfg_w = pmp_io_pma_11_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_11_cfg_r = pmp_io_pma_11_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_11_addr = pmp_io_pma_11_addr; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_11_mask = pmp_io_pma_11_mask; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_12_cfg_c = pmp_io_pma_12_cfg_c; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_12_cfg_atomic = pmp_io_pma_12_cfg_atomic; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_12_cfg_a = pmp_io_pma_12_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_12_cfg_w = pmp_io_pma_12_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_12_cfg_r = pmp_io_pma_12_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_12_addr = pmp_io_pma_12_addr; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_12_mask = pmp_io_pma_12_mask; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_13_cfg_c = pmp_io_pma_13_cfg_c; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_13_cfg_atomic = pmp_io_pma_13_cfg_atomic; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_13_cfg_a = pmp_io_pma_13_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_13_cfg_w = pmp_io_pma_13_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_13_cfg_r = pmp_io_pma_13_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_13_addr = pmp_io_pma_13_addr; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_13_mask = pmp_io_pma_13_mask; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_14_cfg_c = pmp_io_pma_14_cfg_c; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_14_cfg_atomic = pmp_io_pma_14_cfg_atomic; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_14_cfg_a = pmp_io_pma_14_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_14_cfg_w = pmp_io_pma_14_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_14_cfg_r = pmp_io_pma_14_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_14_addr = pmp_io_pma_14_addr; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_14_mask = pmp_io_pma_14_mask; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_15_cfg_c = pmp_io_pma_15_cfg_c; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_15_cfg_atomic = pmp_io_pma_15_cfg_atomic; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_15_cfg_a = pmp_io_pma_15_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_15_cfg_w = pmp_io_pma_15_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_15_cfg_r = pmp_io_pma_15_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_15_addr = pmp_io_pma_15_addr; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_check_env_pma_15_mask = pmp_io_pma_15_mask; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_3_io_req_valid = dtlb_st_tlb_st_io_pmp_1_valid; // @[MemBlock.scala 249:{24,24}]
  assign PMPChecker_3_io_req_bits_addr = dtlb_st_tlb_st_io_pmp_1_bits_addr; // @[MemBlock.scala 249:{24,24}]
  assign PMPChecker_3_io_req_bits_cmd = 3'h1; // @[MemBlock.scala 249:{24,24}]
  assign PMPChecker_4_clock = clock;
  assign PMPChecker_4_io_check_env_mode = tlbcsr_priv_dmode; // @[MemBlock.scala 314:26 PMP.scala 465:15]
  assign PMPChecker_4_io_check_env_pmp_0_cfg_l = pmp_io_pmp_0_cfg_l; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_0_cfg_a = pmp_io_pmp_0_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_0_cfg_w = pmp_io_pmp_0_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_0_cfg_r = pmp_io_pmp_0_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_0_addr = pmp_io_pmp_0_addr; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_0_mask = pmp_io_pmp_0_mask; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_1_cfg_l = pmp_io_pmp_1_cfg_l; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_1_cfg_a = pmp_io_pmp_1_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_1_cfg_w = pmp_io_pmp_1_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_1_cfg_r = pmp_io_pmp_1_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_1_addr = pmp_io_pmp_1_addr; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_1_mask = pmp_io_pmp_1_mask; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_2_cfg_l = pmp_io_pmp_2_cfg_l; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_2_cfg_a = pmp_io_pmp_2_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_2_cfg_w = pmp_io_pmp_2_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_2_cfg_r = pmp_io_pmp_2_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_2_addr = pmp_io_pmp_2_addr; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_2_mask = pmp_io_pmp_2_mask; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_3_cfg_l = pmp_io_pmp_3_cfg_l; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_3_cfg_a = pmp_io_pmp_3_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_3_cfg_w = pmp_io_pmp_3_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_3_cfg_r = pmp_io_pmp_3_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_3_addr = pmp_io_pmp_3_addr; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_3_mask = pmp_io_pmp_3_mask; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_4_cfg_l = pmp_io_pmp_4_cfg_l; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_4_cfg_a = pmp_io_pmp_4_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_4_cfg_w = pmp_io_pmp_4_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_4_cfg_r = pmp_io_pmp_4_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_4_addr = pmp_io_pmp_4_addr; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_4_mask = pmp_io_pmp_4_mask; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_5_cfg_l = pmp_io_pmp_5_cfg_l; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_5_cfg_a = pmp_io_pmp_5_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_5_cfg_w = pmp_io_pmp_5_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_5_cfg_r = pmp_io_pmp_5_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_5_addr = pmp_io_pmp_5_addr; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_5_mask = pmp_io_pmp_5_mask; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_6_cfg_l = pmp_io_pmp_6_cfg_l; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_6_cfg_a = pmp_io_pmp_6_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_6_cfg_w = pmp_io_pmp_6_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_6_cfg_r = pmp_io_pmp_6_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_6_addr = pmp_io_pmp_6_addr; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_6_mask = pmp_io_pmp_6_mask; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_7_cfg_l = pmp_io_pmp_7_cfg_l; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_7_cfg_a = pmp_io_pmp_7_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_7_cfg_w = pmp_io_pmp_7_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_7_cfg_r = pmp_io_pmp_7_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_7_addr = pmp_io_pmp_7_addr; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_7_mask = pmp_io_pmp_7_mask; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_8_cfg_l = pmp_io_pmp_8_cfg_l; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_8_cfg_a = pmp_io_pmp_8_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_8_cfg_w = pmp_io_pmp_8_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_8_cfg_r = pmp_io_pmp_8_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_8_addr = pmp_io_pmp_8_addr; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_8_mask = pmp_io_pmp_8_mask; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_9_cfg_l = pmp_io_pmp_9_cfg_l; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_9_cfg_a = pmp_io_pmp_9_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_9_cfg_w = pmp_io_pmp_9_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_9_cfg_r = pmp_io_pmp_9_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_9_addr = pmp_io_pmp_9_addr; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_9_mask = pmp_io_pmp_9_mask; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_10_cfg_l = pmp_io_pmp_10_cfg_l; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_10_cfg_a = pmp_io_pmp_10_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_10_cfg_w = pmp_io_pmp_10_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_10_cfg_r = pmp_io_pmp_10_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_10_addr = pmp_io_pmp_10_addr; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_10_mask = pmp_io_pmp_10_mask; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_11_cfg_l = pmp_io_pmp_11_cfg_l; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_11_cfg_a = pmp_io_pmp_11_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_11_cfg_w = pmp_io_pmp_11_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_11_cfg_r = pmp_io_pmp_11_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_11_addr = pmp_io_pmp_11_addr; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_11_mask = pmp_io_pmp_11_mask; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_12_cfg_l = pmp_io_pmp_12_cfg_l; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_12_cfg_a = pmp_io_pmp_12_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_12_cfg_w = pmp_io_pmp_12_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_12_cfg_r = pmp_io_pmp_12_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_12_addr = pmp_io_pmp_12_addr; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_12_mask = pmp_io_pmp_12_mask; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_13_cfg_l = pmp_io_pmp_13_cfg_l; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_13_cfg_a = pmp_io_pmp_13_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_13_cfg_w = pmp_io_pmp_13_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_13_cfg_r = pmp_io_pmp_13_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_13_addr = pmp_io_pmp_13_addr; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_13_mask = pmp_io_pmp_13_mask; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_14_cfg_l = pmp_io_pmp_14_cfg_l; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_14_cfg_a = pmp_io_pmp_14_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_14_cfg_w = pmp_io_pmp_14_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_14_cfg_r = pmp_io_pmp_14_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_14_addr = pmp_io_pmp_14_addr; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_14_mask = pmp_io_pmp_14_mask; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_15_cfg_l = pmp_io_pmp_15_cfg_l; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_15_cfg_a = pmp_io_pmp_15_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_15_cfg_w = pmp_io_pmp_15_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_15_cfg_r = pmp_io_pmp_15_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_15_addr = pmp_io_pmp_15_addr; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pmp_15_mask = pmp_io_pmp_15_mask; // @[MemBlock.scala 314:26 PMP.scala 466:14]
  assign PMPChecker_4_io_check_env_pma_0_cfg_c = pmp_io_pma_0_cfg_c; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_0_cfg_atomic = pmp_io_pma_0_cfg_atomic; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_0_cfg_a = pmp_io_pma_0_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_0_cfg_w = pmp_io_pma_0_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_0_cfg_r = pmp_io_pma_0_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_0_addr = pmp_io_pma_0_addr; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_0_mask = pmp_io_pma_0_mask; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_1_cfg_c = pmp_io_pma_1_cfg_c; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_1_cfg_atomic = pmp_io_pma_1_cfg_atomic; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_1_cfg_a = pmp_io_pma_1_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_1_cfg_w = pmp_io_pma_1_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_1_cfg_r = pmp_io_pma_1_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_1_addr = pmp_io_pma_1_addr; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_1_mask = pmp_io_pma_1_mask; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_2_cfg_c = pmp_io_pma_2_cfg_c; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_2_cfg_atomic = pmp_io_pma_2_cfg_atomic; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_2_cfg_a = pmp_io_pma_2_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_2_cfg_w = pmp_io_pma_2_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_2_cfg_r = pmp_io_pma_2_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_2_addr = pmp_io_pma_2_addr; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_2_mask = pmp_io_pma_2_mask; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_3_cfg_c = pmp_io_pma_3_cfg_c; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_3_cfg_atomic = pmp_io_pma_3_cfg_atomic; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_3_cfg_a = pmp_io_pma_3_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_3_cfg_w = pmp_io_pma_3_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_3_cfg_r = pmp_io_pma_3_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_3_addr = pmp_io_pma_3_addr; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_3_mask = pmp_io_pma_3_mask; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_4_cfg_c = pmp_io_pma_4_cfg_c; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_4_cfg_atomic = pmp_io_pma_4_cfg_atomic; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_4_cfg_a = pmp_io_pma_4_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_4_cfg_w = pmp_io_pma_4_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_4_cfg_r = pmp_io_pma_4_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_4_addr = pmp_io_pma_4_addr; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_4_mask = pmp_io_pma_4_mask; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_5_cfg_c = pmp_io_pma_5_cfg_c; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_5_cfg_atomic = pmp_io_pma_5_cfg_atomic; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_5_cfg_a = pmp_io_pma_5_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_5_cfg_w = pmp_io_pma_5_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_5_cfg_r = pmp_io_pma_5_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_5_addr = pmp_io_pma_5_addr; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_5_mask = pmp_io_pma_5_mask; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_6_cfg_c = pmp_io_pma_6_cfg_c; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_6_cfg_atomic = pmp_io_pma_6_cfg_atomic; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_6_cfg_a = pmp_io_pma_6_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_6_cfg_w = pmp_io_pma_6_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_6_cfg_r = pmp_io_pma_6_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_6_addr = pmp_io_pma_6_addr; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_6_mask = pmp_io_pma_6_mask; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_7_cfg_c = pmp_io_pma_7_cfg_c; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_7_cfg_atomic = pmp_io_pma_7_cfg_atomic; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_7_cfg_a = pmp_io_pma_7_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_7_cfg_w = pmp_io_pma_7_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_7_cfg_r = pmp_io_pma_7_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_7_addr = pmp_io_pma_7_addr; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_7_mask = pmp_io_pma_7_mask; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_8_cfg_c = pmp_io_pma_8_cfg_c; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_8_cfg_atomic = pmp_io_pma_8_cfg_atomic; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_8_cfg_a = pmp_io_pma_8_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_8_cfg_w = pmp_io_pma_8_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_8_cfg_r = pmp_io_pma_8_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_8_addr = pmp_io_pma_8_addr; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_8_mask = pmp_io_pma_8_mask; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_9_cfg_c = pmp_io_pma_9_cfg_c; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_9_cfg_atomic = pmp_io_pma_9_cfg_atomic; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_9_cfg_a = pmp_io_pma_9_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_9_cfg_w = pmp_io_pma_9_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_9_cfg_r = pmp_io_pma_9_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_9_addr = pmp_io_pma_9_addr; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_9_mask = pmp_io_pma_9_mask; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_10_cfg_c = pmp_io_pma_10_cfg_c; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_10_cfg_atomic = pmp_io_pma_10_cfg_atomic; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_10_cfg_a = pmp_io_pma_10_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_10_cfg_w = pmp_io_pma_10_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_10_cfg_r = pmp_io_pma_10_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_10_addr = pmp_io_pma_10_addr; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_10_mask = pmp_io_pma_10_mask; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_11_cfg_c = pmp_io_pma_11_cfg_c; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_11_cfg_atomic = pmp_io_pma_11_cfg_atomic; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_11_cfg_a = pmp_io_pma_11_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_11_cfg_w = pmp_io_pma_11_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_11_cfg_r = pmp_io_pma_11_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_11_addr = pmp_io_pma_11_addr; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_11_mask = pmp_io_pma_11_mask; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_12_cfg_c = pmp_io_pma_12_cfg_c; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_12_cfg_atomic = pmp_io_pma_12_cfg_atomic; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_12_cfg_a = pmp_io_pma_12_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_12_cfg_w = pmp_io_pma_12_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_12_cfg_r = pmp_io_pma_12_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_12_addr = pmp_io_pma_12_addr; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_12_mask = pmp_io_pma_12_mask; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_13_cfg_c = pmp_io_pma_13_cfg_c; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_13_cfg_atomic = pmp_io_pma_13_cfg_atomic; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_13_cfg_a = pmp_io_pma_13_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_13_cfg_w = pmp_io_pma_13_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_13_cfg_r = pmp_io_pma_13_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_13_addr = pmp_io_pma_13_addr; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_13_mask = pmp_io_pma_13_mask; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_14_cfg_c = pmp_io_pma_14_cfg_c; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_14_cfg_atomic = pmp_io_pma_14_cfg_atomic; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_14_cfg_a = pmp_io_pma_14_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_14_cfg_w = pmp_io_pma_14_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_14_cfg_r = pmp_io_pma_14_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_14_addr = pmp_io_pma_14_addr; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_14_mask = pmp_io_pma_14_mask; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_15_cfg_c = pmp_io_pma_15_cfg_c; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_15_cfg_atomic = pmp_io_pma_15_cfg_atomic; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_15_cfg_a = pmp_io_pma_15_cfg_a; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_15_cfg_w = pmp_io_pma_15_cfg_w; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_15_cfg_r = pmp_io_pma_15_cfg_r; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_15_addr = pmp_io_pma_15_addr; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_check_env_pma_15_mask = pmp_io_pma_15_mask; // @[MemBlock.scala 314:26 PMP.scala 467:14]
  assign PMPChecker_4_io_req_valid = dtlb_prefetch_tlb_prefetch_io_pmp_0_valid; // @[MemBlock.scala 253:{30,30}]
  assign PMPChecker_4_io_req_bits_addr = dtlb_prefetch_tlb_prefetch_io_pmp_0_bits_addr; // @[MemBlock.scala 253:{30,30}]
  assign PMPChecker_4_io_req_bits_cmd = 3'h0; // @[MemBlock.scala 253:{30,30}]
  assign pmp_check_ptw_clock = clock;
  assign pmp_check_ptw_reset = reset;
  assign pmp_check_ptw_io_check_env_mode = tlbcsr_priv_dmode; // @[PMP.scala 465:15]
  assign pmp_check_ptw_io_check_env_pmp_0_cfg_l = pmp_io_pmp_0_cfg_l; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_0_cfg_a = pmp_io_pmp_0_cfg_a; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_0_cfg_x = pmp_io_pmp_0_cfg_x; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_0_cfg_w = pmp_io_pmp_0_cfg_w; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_0_cfg_r = pmp_io_pmp_0_cfg_r; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_0_addr = pmp_io_pmp_0_addr; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_0_mask = pmp_io_pmp_0_mask; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_1_cfg_l = pmp_io_pmp_1_cfg_l; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_1_cfg_a = pmp_io_pmp_1_cfg_a; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_1_cfg_x = pmp_io_pmp_1_cfg_x; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_1_cfg_w = pmp_io_pmp_1_cfg_w; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_1_cfg_r = pmp_io_pmp_1_cfg_r; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_1_addr = pmp_io_pmp_1_addr; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_1_mask = pmp_io_pmp_1_mask; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_2_cfg_l = pmp_io_pmp_2_cfg_l; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_2_cfg_a = pmp_io_pmp_2_cfg_a; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_2_cfg_x = pmp_io_pmp_2_cfg_x; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_2_cfg_w = pmp_io_pmp_2_cfg_w; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_2_cfg_r = pmp_io_pmp_2_cfg_r; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_2_addr = pmp_io_pmp_2_addr; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_2_mask = pmp_io_pmp_2_mask; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_3_cfg_l = pmp_io_pmp_3_cfg_l; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_3_cfg_a = pmp_io_pmp_3_cfg_a; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_3_cfg_x = pmp_io_pmp_3_cfg_x; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_3_cfg_w = pmp_io_pmp_3_cfg_w; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_3_cfg_r = pmp_io_pmp_3_cfg_r; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_3_addr = pmp_io_pmp_3_addr; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_3_mask = pmp_io_pmp_3_mask; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_4_cfg_l = pmp_io_pmp_4_cfg_l; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_4_cfg_a = pmp_io_pmp_4_cfg_a; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_4_cfg_x = pmp_io_pmp_4_cfg_x; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_4_cfg_w = pmp_io_pmp_4_cfg_w; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_4_cfg_r = pmp_io_pmp_4_cfg_r; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_4_addr = pmp_io_pmp_4_addr; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_4_mask = pmp_io_pmp_4_mask; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_5_cfg_l = pmp_io_pmp_5_cfg_l; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_5_cfg_a = pmp_io_pmp_5_cfg_a; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_5_cfg_x = pmp_io_pmp_5_cfg_x; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_5_cfg_w = pmp_io_pmp_5_cfg_w; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_5_cfg_r = pmp_io_pmp_5_cfg_r; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_5_addr = pmp_io_pmp_5_addr; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_5_mask = pmp_io_pmp_5_mask; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_6_cfg_l = pmp_io_pmp_6_cfg_l; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_6_cfg_a = pmp_io_pmp_6_cfg_a; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_6_cfg_x = pmp_io_pmp_6_cfg_x; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_6_cfg_w = pmp_io_pmp_6_cfg_w; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_6_cfg_r = pmp_io_pmp_6_cfg_r; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_6_addr = pmp_io_pmp_6_addr; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_6_mask = pmp_io_pmp_6_mask; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_7_cfg_l = pmp_io_pmp_7_cfg_l; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_7_cfg_a = pmp_io_pmp_7_cfg_a; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_7_cfg_x = pmp_io_pmp_7_cfg_x; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_7_cfg_w = pmp_io_pmp_7_cfg_w; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_7_cfg_r = pmp_io_pmp_7_cfg_r; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_7_addr = pmp_io_pmp_7_addr; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_7_mask = pmp_io_pmp_7_mask; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_8_cfg_l = pmp_io_pmp_8_cfg_l; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_8_cfg_a = pmp_io_pmp_8_cfg_a; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_8_cfg_x = pmp_io_pmp_8_cfg_x; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_8_cfg_w = pmp_io_pmp_8_cfg_w; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_8_cfg_r = pmp_io_pmp_8_cfg_r; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_8_addr = pmp_io_pmp_8_addr; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_8_mask = pmp_io_pmp_8_mask; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_9_cfg_l = pmp_io_pmp_9_cfg_l; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_9_cfg_a = pmp_io_pmp_9_cfg_a; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_9_cfg_x = pmp_io_pmp_9_cfg_x; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_9_cfg_w = pmp_io_pmp_9_cfg_w; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_9_cfg_r = pmp_io_pmp_9_cfg_r; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_9_addr = pmp_io_pmp_9_addr; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_9_mask = pmp_io_pmp_9_mask; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_10_cfg_l = pmp_io_pmp_10_cfg_l; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_10_cfg_a = pmp_io_pmp_10_cfg_a; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_10_cfg_x = pmp_io_pmp_10_cfg_x; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_10_cfg_w = pmp_io_pmp_10_cfg_w; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_10_cfg_r = pmp_io_pmp_10_cfg_r; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_10_addr = pmp_io_pmp_10_addr; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_10_mask = pmp_io_pmp_10_mask; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_11_cfg_l = pmp_io_pmp_11_cfg_l; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_11_cfg_a = pmp_io_pmp_11_cfg_a; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_11_cfg_x = pmp_io_pmp_11_cfg_x; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_11_cfg_w = pmp_io_pmp_11_cfg_w; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_11_cfg_r = pmp_io_pmp_11_cfg_r; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_11_addr = pmp_io_pmp_11_addr; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_11_mask = pmp_io_pmp_11_mask; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_12_cfg_l = pmp_io_pmp_12_cfg_l; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_12_cfg_a = pmp_io_pmp_12_cfg_a; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_12_cfg_x = pmp_io_pmp_12_cfg_x; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_12_cfg_w = pmp_io_pmp_12_cfg_w; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_12_cfg_r = pmp_io_pmp_12_cfg_r; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_12_addr = pmp_io_pmp_12_addr; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_12_mask = pmp_io_pmp_12_mask; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_13_cfg_l = pmp_io_pmp_13_cfg_l; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_13_cfg_a = pmp_io_pmp_13_cfg_a; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_13_cfg_x = pmp_io_pmp_13_cfg_x; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_13_cfg_w = pmp_io_pmp_13_cfg_w; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_13_cfg_r = pmp_io_pmp_13_cfg_r; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_13_addr = pmp_io_pmp_13_addr; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_13_mask = pmp_io_pmp_13_mask; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_14_cfg_l = pmp_io_pmp_14_cfg_l; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_14_cfg_a = pmp_io_pmp_14_cfg_a; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_14_cfg_x = pmp_io_pmp_14_cfg_x; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_14_cfg_w = pmp_io_pmp_14_cfg_w; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_14_cfg_r = pmp_io_pmp_14_cfg_r; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_14_addr = pmp_io_pmp_14_addr; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_14_mask = pmp_io_pmp_14_mask; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_15_cfg_l = pmp_io_pmp_15_cfg_l; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_15_cfg_a = pmp_io_pmp_15_cfg_a; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_15_cfg_x = pmp_io_pmp_15_cfg_x; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_15_cfg_w = pmp_io_pmp_15_cfg_w; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_15_cfg_r = pmp_io_pmp_15_cfg_r; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_15_addr = pmp_io_pmp_15_addr; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pmp_15_mask = pmp_io_pmp_15_mask; // @[PMP.scala 466:14]
  assign pmp_check_ptw_io_check_env_pma_0_cfg_c = pmp_io_pma_0_cfg_c; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_0_cfg_atomic = pmp_io_pma_0_cfg_atomic; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_0_cfg_a = pmp_io_pma_0_cfg_a; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_0_cfg_x = pmp_io_pma_0_cfg_x; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_0_cfg_w = pmp_io_pma_0_cfg_w; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_0_cfg_r = pmp_io_pma_0_cfg_r; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_0_addr = pmp_io_pma_0_addr; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_0_mask = pmp_io_pma_0_mask; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_1_cfg_c = pmp_io_pma_1_cfg_c; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_1_cfg_atomic = pmp_io_pma_1_cfg_atomic; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_1_cfg_a = pmp_io_pma_1_cfg_a; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_1_cfg_x = pmp_io_pma_1_cfg_x; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_1_cfg_w = pmp_io_pma_1_cfg_w; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_1_cfg_r = pmp_io_pma_1_cfg_r; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_1_addr = pmp_io_pma_1_addr; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_1_mask = pmp_io_pma_1_mask; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_2_cfg_c = pmp_io_pma_2_cfg_c; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_2_cfg_atomic = pmp_io_pma_2_cfg_atomic; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_2_cfg_a = pmp_io_pma_2_cfg_a; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_2_cfg_x = pmp_io_pma_2_cfg_x; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_2_cfg_w = pmp_io_pma_2_cfg_w; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_2_cfg_r = pmp_io_pma_2_cfg_r; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_2_addr = pmp_io_pma_2_addr; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_2_mask = pmp_io_pma_2_mask; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_3_cfg_c = pmp_io_pma_3_cfg_c; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_3_cfg_atomic = pmp_io_pma_3_cfg_atomic; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_3_cfg_a = pmp_io_pma_3_cfg_a; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_3_cfg_x = pmp_io_pma_3_cfg_x; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_3_cfg_w = pmp_io_pma_3_cfg_w; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_3_cfg_r = pmp_io_pma_3_cfg_r; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_3_addr = pmp_io_pma_3_addr; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_3_mask = pmp_io_pma_3_mask; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_4_cfg_c = pmp_io_pma_4_cfg_c; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_4_cfg_atomic = pmp_io_pma_4_cfg_atomic; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_4_cfg_a = pmp_io_pma_4_cfg_a; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_4_cfg_x = pmp_io_pma_4_cfg_x; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_4_cfg_w = pmp_io_pma_4_cfg_w; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_4_cfg_r = pmp_io_pma_4_cfg_r; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_4_addr = pmp_io_pma_4_addr; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_4_mask = pmp_io_pma_4_mask; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_5_cfg_c = pmp_io_pma_5_cfg_c; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_5_cfg_atomic = pmp_io_pma_5_cfg_atomic; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_5_cfg_a = pmp_io_pma_5_cfg_a; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_5_cfg_x = pmp_io_pma_5_cfg_x; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_5_cfg_w = pmp_io_pma_5_cfg_w; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_5_cfg_r = pmp_io_pma_5_cfg_r; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_5_addr = pmp_io_pma_5_addr; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_5_mask = pmp_io_pma_5_mask; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_6_cfg_c = pmp_io_pma_6_cfg_c; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_6_cfg_atomic = pmp_io_pma_6_cfg_atomic; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_6_cfg_a = pmp_io_pma_6_cfg_a; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_6_cfg_x = pmp_io_pma_6_cfg_x; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_6_cfg_w = pmp_io_pma_6_cfg_w; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_6_cfg_r = pmp_io_pma_6_cfg_r; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_6_addr = pmp_io_pma_6_addr; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_6_mask = pmp_io_pma_6_mask; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_7_cfg_c = pmp_io_pma_7_cfg_c; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_7_cfg_atomic = pmp_io_pma_7_cfg_atomic; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_7_cfg_a = pmp_io_pma_7_cfg_a; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_7_cfg_x = pmp_io_pma_7_cfg_x; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_7_cfg_w = pmp_io_pma_7_cfg_w; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_7_cfg_r = pmp_io_pma_7_cfg_r; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_7_addr = pmp_io_pma_7_addr; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_7_mask = pmp_io_pma_7_mask; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_8_cfg_c = pmp_io_pma_8_cfg_c; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_8_cfg_atomic = pmp_io_pma_8_cfg_atomic; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_8_cfg_a = pmp_io_pma_8_cfg_a; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_8_cfg_x = pmp_io_pma_8_cfg_x; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_8_cfg_w = pmp_io_pma_8_cfg_w; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_8_cfg_r = pmp_io_pma_8_cfg_r; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_8_addr = pmp_io_pma_8_addr; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_8_mask = pmp_io_pma_8_mask; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_9_cfg_c = pmp_io_pma_9_cfg_c; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_9_cfg_atomic = pmp_io_pma_9_cfg_atomic; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_9_cfg_a = pmp_io_pma_9_cfg_a; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_9_cfg_x = pmp_io_pma_9_cfg_x; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_9_cfg_w = pmp_io_pma_9_cfg_w; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_9_cfg_r = pmp_io_pma_9_cfg_r; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_9_addr = pmp_io_pma_9_addr; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_9_mask = pmp_io_pma_9_mask; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_10_cfg_c = pmp_io_pma_10_cfg_c; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_10_cfg_atomic = pmp_io_pma_10_cfg_atomic; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_10_cfg_a = pmp_io_pma_10_cfg_a; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_10_cfg_x = pmp_io_pma_10_cfg_x; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_10_cfg_w = pmp_io_pma_10_cfg_w; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_10_cfg_r = pmp_io_pma_10_cfg_r; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_10_addr = pmp_io_pma_10_addr; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_10_mask = pmp_io_pma_10_mask; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_11_cfg_c = pmp_io_pma_11_cfg_c; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_11_cfg_atomic = pmp_io_pma_11_cfg_atomic; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_11_cfg_a = pmp_io_pma_11_cfg_a; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_11_cfg_x = pmp_io_pma_11_cfg_x; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_11_cfg_w = pmp_io_pma_11_cfg_w; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_11_cfg_r = pmp_io_pma_11_cfg_r; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_11_addr = pmp_io_pma_11_addr; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_11_mask = pmp_io_pma_11_mask; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_12_cfg_c = pmp_io_pma_12_cfg_c; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_12_cfg_atomic = pmp_io_pma_12_cfg_atomic; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_12_cfg_a = pmp_io_pma_12_cfg_a; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_12_cfg_x = pmp_io_pma_12_cfg_x; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_12_cfg_w = pmp_io_pma_12_cfg_w; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_12_cfg_r = pmp_io_pma_12_cfg_r; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_12_addr = pmp_io_pma_12_addr; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_12_mask = pmp_io_pma_12_mask; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_13_cfg_c = pmp_io_pma_13_cfg_c; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_13_cfg_atomic = pmp_io_pma_13_cfg_atomic; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_13_cfg_a = pmp_io_pma_13_cfg_a; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_13_cfg_x = pmp_io_pma_13_cfg_x; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_13_cfg_w = pmp_io_pma_13_cfg_w; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_13_cfg_r = pmp_io_pma_13_cfg_r; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_13_addr = pmp_io_pma_13_addr; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_13_mask = pmp_io_pma_13_mask; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_14_cfg_c = pmp_io_pma_14_cfg_c; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_14_cfg_atomic = pmp_io_pma_14_cfg_atomic; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_14_cfg_a = pmp_io_pma_14_cfg_a; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_14_cfg_x = pmp_io_pma_14_cfg_x; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_14_cfg_w = pmp_io_pma_14_cfg_w; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_14_cfg_r = pmp_io_pma_14_cfg_r; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_14_addr = pmp_io_pma_14_addr; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_14_mask = pmp_io_pma_14_mask; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_15_cfg_c = pmp_io_pma_15_cfg_c; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_15_cfg_atomic = pmp_io_pma_15_cfg_atomic; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_15_cfg_a = pmp_io_pma_15_cfg_a; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_15_cfg_x = pmp_io_pma_15_cfg_x; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_15_cfg_w = pmp_io_pma_15_cfg_w; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_15_cfg_r = pmp_io_pma_15_cfg_r; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_15_addr = pmp_io_pma_15_addr; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_check_env_pma_15_mask = pmp_io_pma_15_mask; // @[PMP.scala 467:14]
  assign pmp_check_ptw_io_req_valid = io_ptw_resp_valid; // @[PMP.scala 506:20]
  assign pmp_check_ptw_io_req_bits_addr = {io_ptw_resp_bits_data_entry_ppn,12'h0}; // @[Cat.scala 31:58]
  assign pipelineReg_clock = clock;
  assign pipelineReg_reset = reset;
  assign pipelineReg_io_in_valid = lsq_io_uncache_req_valid; // @[MemCommon.scala 398:23]
  assign pipelineReg_io_in_bits_cmd = lsq_io_uncache_req_bits_cmd; // @[MemCommon.scala 398:23]
  assign pipelineReg_io_in_bits_addr = lsq_io_uncache_req_bits_addr; // @[MemCommon.scala 398:23]
  assign pipelineReg_io_in_bits_data = lsq_io_uncache_req_bits_data; // @[MemCommon.scala 398:23]
  assign pipelineReg_io_in_bits_mask = lsq_io_uncache_req_bits_mask; // @[MemCommon.scala 398:23]
  assign pipelineReg_io_in_bits_atomic = lsq_io_uncache_req_bits_atomic; // @[MemCommon.scala 398:23]
  assign pipelineReg_io_out_ready = uncache_io_lsq_req_ready; // @[MemCommon.scala 399:11]
  assign pipelineReg_1_clock = clock;
  assign pipelineReg_1_reset = reset;
  assign pipelineReg_1_io_in_valid = uncache_io_lsq_resp_valid; // @[MemCommon.scala 398:23]
  assign pipelineReg_1_io_in_bits_data = uncache_io_lsq_resp_bits_data; // @[MemCommon.scala 398:23]
  assign delay_clock = clock;
  assign delay_io_in = redirect_next_valid_REG; // @[BitUtils.scala 26:20 28:18]
  assign pfevent_clock = clock;
  assign pfevent_reset = reset;
  assign pfevent_io_distribute_csr_wvalid = csrCtrl_delay_io_out_distribute_csr_wvalid; // @[MemBlock.scala 688:29]
  assign pfevent_io_distribute_csr_waddr = csrCtrl_delay_io_out_distribute_csr_waddr; // @[MemBlock.scala 688:29]
  assign pfevent_io_distribute_csr_wdata = csrCtrl_delay_io_out_distribute_csr_wdata; // @[MemBlock.scala 688:29]
  assign hpm_clock = clock;
  assign hpm_io_hpm_event_0 = pfevent_io_hpmevent_16; // @[PerfCounterUtils.scala 256:22]
  assign hpm_io_hpm_event_1 = pfevent_io_hpmevent_17; // @[PerfCounterUtils.scala 256:22]
  assign hpm_io_hpm_event_2 = pfevent_io_hpmevent_18; // @[PerfCounterUtils.scala 256:22]
  assign hpm_io_hpm_event_3 = pfevent_io_hpmevent_19; // @[PerfCounterUtils.scala 256:22]
  assign hpm_io_hpm_event_4 = pfevent_io_hpmevent_20; // @[PerfCounterUtils.scala 256:22]
  assign hpm_io_hpm_event_5 = pfevent_io_hpmevent_21; // @[PerfCounterUtils.scala 256:22]
  assign hpm_io_hpm_event_6 = pfevent_io_hpmevent_22; // @[PerfCounterUtils.scala 256:22]
  assign hpm_io_hpm_event_7 = pfevent_io_hpmevent_23; // @[PerfCounterUtils.scala 256:22]
  assign hpm_io_events_sets_0_value = {{4'd0}, ldDeqCount}; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_1_value = {{3'd0}, stDeqCount}; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_2_value = LoadUnit_0_io_perf_0_value; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_3_value = LoadUnit_0_io_perf_1_value; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_4_value = LoadUnit_0_io_perf_2_value; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_5_value = LoadUnit_0_io_perf_3_value; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_6_value = LoadUnit_0_io_perf_4_value; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_7_value = LoadUnit_0_io_perf_5_value; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_8_value = LoadUnit_0_io_perf_6_value; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_9_value = LoadUnit_1_io_perf_0_value; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_10_value = LoadUnit_1_io_perf_1_value; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_11_value = LoadUnit_1_io_perf_2_value; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_12_value = LoadUnit_1_io_perf_3_value; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_13_value = LoadUnit_1_io_perf_4_value; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_14_value = LoadUnit_1_io_perf_5_value; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_15_value = LoadUnit_1_io_perf_6_value; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_16_value = sbuffer_io_perf_0_value; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_17_value = sbuffer_io_perf_1_value; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_18_value = sbuffer_io_perf_2_value; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_19_value = sbuffer_io_perf_3_value; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_20_value = sbuffer_io_perf_4_value; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_21_value = sbuffer_io_perf_5_value; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_22_value = sbuffer_io_perf_6_value; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_23_value = sbuffer_io_perf_7_value; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_24_value = sbuffer_io_perf_8_value; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_25_value = sbuffer_io_perf_9_value; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_26_value = sbuffer_io_perf_10_value; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_27_value = sbuffer_io_perf_11_value; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_28_value = sbuffer_io_perf_12_value; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_29_value = sbuffer_io_perf_13_value; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_30_value = sbuffer_io_perf_14_value; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_31_value = sbuffer_io_perf_15_value; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_32_value = sbuffer_io_perf_16_value; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_33_value = lsq_io_perf_0_value; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_34_value = lsq_io_perf_1_value; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_35_value = lsq_io_perf_2_value; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_36_value = lsq_io_perf_3_value; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_37_value = lsq_io_perf_4_value; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_38_value = lsq_io_perf_5_value; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_39_value = lsq_io_perf_6_value; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_40_value = lsq_io_perf_7_value; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_41_value = lsq_io_perf_8_value; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_42_value = lsq_io_perf_9_value; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_43_value = lsq_io_perf_10_value; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_44_value = lsq_io_perf_11_value; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_45_value = lsq_io_perf_12_value; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_46_value = lsq_io_perf_13_value; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_47_value = lsq_io_perf_14_value; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_48_value = lsq_io_perf_15_value; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_49_value = lsq_io_perf_16_value; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_50_value = lsq_io_perf_17_value; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_51_value = lsq_io_perf_18_value; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_52_value = lsq_io_perf_19_value; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_53_value = lsq_io_perf_20_value; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_54_value = lsq_io_perf_21_value; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_55_value = lsq_io_perf_22_value; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_56_value = lsq_io_perf_23_value; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_57_value = lsq_io_perf_24_value; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_58_value = lsq_io_perf_25_value; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_59_value = lsq_io_perf_26_value; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_60_value = lsq_io_perf_27_value; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_61_value = lsq_io_perf_28_value; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_62_value = lsq_io_perf_29_value; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_63_value = dcache_io_perf_0_value; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_64_value = dcache_io_perf_1_value; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_65_value = dcache_io_perf_2_value; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_66_value = dcache_io_perf_3_value; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_67_value = dcache_io_perf_4_value; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_68_value = dcache_io_perf_5_value; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_69_value = dcache_io_perf_6_value; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_70_value = dcache_io_perf_7_value; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_71_value = dcache_io_perf_8_value; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_72_value = dcache_io_perf_9_value; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_73_value = dcache_io_perf_10_value; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_74_value = dcache_io_perf_11_value; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_75_value = dcache_io_perf_12_value; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_76_value = dcache_io_perf_13_value; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_77_value = dcache_io_perf_14_value; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_78_value = dcache_io_perf_15_value; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_79_value = dcache_io_perf_16_value; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_80_value = dcache_io_perf_17_value; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_81_value = dcache_io_perf_18_value; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_82_value = dcache_io_perf_19_value; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_83_value = dcache_io_perf_20_value; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_84_value = dcache_io_perf_21_value; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_85_value = dcache_io_perf_22_value; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_86_value = dcache_io_perf_23_value; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_87_value = dcache_io_perf_24_value; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_88_value = dcache_io_perf_25_value; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_89_value = dcache_io_perf_26_value; // @[MemBlock.scala 696:50]
  assign hpm_io_events_sets_90_value = io_perfEventsPTW_0_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_91_value = io_perfEventsPTW_1_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_92_value = io_perfEventsPTW_2_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_93_value = io_perfEventsPTW_3_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_94_value = io_perfEventsPTW_4_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_95_value = io_perfEventsPTW_5_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_96_value = io_perfEventsPTW_6_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_97_value = io_perfEventsPTW_7_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_98_value = io_perfEventsPTW_8_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_99_value = io_perfEventsPTW_9_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_100_value = io_perfEventsPTW_10_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_101_value = io_perfEventsPTW_11_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_102_value = io_perfEventsPTW_12_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_103_value = io_perfEventsPTW_13_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_104_value = io_perfEventsPTW_14_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_105_value = io_perfEventsPTW_15_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_106_value = io_perfEventsPTW_16_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_107_value = io_perfEventsPTW_17_value; // @[PerfCounterUtils.scala 257:24]
  assign hpm_io_events_sets_108_value = io_perfEventsPTW_18_value; // @[PerfCounterUtils.scala 257:24]
  always @(posedge clock) begin
    if (io_redirect_valid) begin // @[Reg.scala 17:18]
      redirect_next_bits_rrobIdx_flag <= io_redirect_bits_robIdx_flag; // @[Reg.scala 17:22]
    end
    if (io_redirect_valid) begin // @[Reg.scala 17:18]
      redirect_next_bits_rrobIdx_value <= io_redirect_bits_robIdx_value; // @[Reg.scala 17:22]
    end
    if (io_redirect_valid) begin // @[Reg.scala 17:18]
      redirect_next_bits_rlevel <= io_redirect_bits_level; // @[Reg.scala 17:22]
    end
    delayedDcacheRefill_valid <= dcache_io_lsu_lsq_valid; // @[MemBlock.scala 127:36]
    delayedDcacheRefill_bits_id <= dcache_io_lsu_lsq_bits_id; // @[MemBlock.scala 127:36]
    io_csrUpdate_REG_wvalid <= dcache_io_csr_update_wvalid; // @[MemBlock.scala 132:26]
    io_csrUpdate_REG_waddr <= dcache_io_csr_update_waddr; // @[MemBlock.scala 132:26]
    io_csrUpdate_REG_wdata <= dcache_io_csr_update_wdata; // @[MemBlock.scala 132:26]
    io_error_REG_paddr <= dcache_io_error_paddr; // @[MemBlock.scala 133:30]
    io_error_REG_report_to_beu <= dcache_io_error_report_to_beu; // @[MemBlock.scala 133:30]
    io_error_REG_1_paddr <= io_error_REG_paddr; // @[MemBlock.scala 133:22]
    io_error_REG_1_report_to_beu <= io_error_REG_report_to_beu; // @[MemBlock.scala 133:22]
    sfence_REG_valid <= io_sfence_valid; // @[MemBlock.scala 243:31]
    sfence_REG_bits_rs1 <= io_sfence_bits_rs1; // @[MemBlock.scala 243:31]
    sfence_REG_bits_rs2 <= io_sfence_bits_rs2; // @[MemBlock.scala 243:31]
    sfence_REG_bits_addr <= io_sfence_bits_addr; // @[MemBlock.scala 243:31]
    sfence_REG_bits_asid <= io_sfence_bits_asid; // @[MemBlock.scala 243:31]
    sfence_valid <= sfence_REG_valid; // @[MemBlock.scala 243:23]
    sfence_bits_rs1 <= sfence_REG_bits_rs1; // @[MemBlock.scala 243:23]
    sfence_bits_rs2 <= sfence_REG_bits_rs2; // @[MemBlock.scala 243:23]
    sfence_bits_addr <= sfence_REG_bits_addr; // @[MemBlock.scala 243:23]
    sfence_bits_asid <= sfence_REG_bits_asid; // @[MemBlock.scala 243:23]
    tlbcsr_REG_satp_mode <= io_tlbCsr_satp_mode; // @[MemBlock.scala 244:31]
    tlbcsr_REG_satp_asid <= io_tlbCsr_satp_asid; // @[MemBlock.scala 244:31]
    tlbcsr_REG_satp_changed <= io_tlbCsr_satp_changed; // @[MemBlock.scala 244:31]
    tlbcsr_REG_priv_mxr <= io_tlbCsr_priv_mxr; // @[MemBlock.scala 244:31]
    tlbcsr_REG_priv_sum <= io_tlbCsr_priv_sum; // @[MemBlock.scala 244:31]
    tlbcsr_REG_priv_dmode <= io_tlbCsr_priv_dmode; // @[MemBlock.scala 244:31]
    tlbcsr_satp_mode <= tlbcsr_REG_satp_mode; // @[MemBlock.scala 244:23]
    tlbcsr_satp_asid <= tlbcsr_REG_satp_asid; // @[MemBlock.scala 244:23]
    tlbcsr_satp_changed <= tlbcsr_REG_satp_changed; // @[MemBlock.scala 244:23]
    tlbcsr_priv_mxr <= tlbcsr_REG_priv_mxr; // @[MemBlock.scala 244:23]
    tlbcsr_priv_sum <= tlbcsr_REG_priv_sum; // @[MemBlock.scala 244:23]
    tlbcsr_priv_dmode <= tlbcsr_REG_priv_dmode; // @[MemBlock.scala 244:23]
    if (io_ptw_resp_valid) begin // @[Reg.scala 17:18]
      ptw_resp_next_data_entry_tag <= io_ptw_resp_bits_data_entry_tag; // @[Reg.scala 17:22]
    end
    if (io_ptw_resp_valid) begin // @[Reg.scala 17:18]
      ptw_resp_next_data_entry_asid <= io_ptw_resp_bits_data_entry_asid; // @[Reg.scala 17:22]
    end
    if (io_ptw_resp_valid) begin // @[Reg.scala 17:18]
      ptw_resp_next_data_entry_ppn <= io_ptw_resp_bits_data_entry_ppn; // @[Reg.scala 17:22]
    end
    if (io_ptw_resp_valid) begin // @[Reg.scala 17:18]
      ptw_resp_next_data_entry_perm_d <= io_ptw_resp_bits_data_entry_perm_d; // @[Reg.scala 17:22]
    end
    if (io_ptw_resp_valid) begin // @[Reg.scala 17:18]
      ptw_resp_next_data_entry_perm_a <= io_ptw_resp_bits_data_entry_perm_a; // @[Reg.scala 17:22]
    end
    if (io_ptw_resp_valid) begin // @[Reg.scala 17:18]
      ptw_resp_next_data_entry_perm_g <= io_ptw_resp_bits_data_entry_perm_g; // @[Reg.scala 17:22]
    end
    if (io_ptw_resp_valid) begin // @[Reg.scala 17:18]
      ptw_resp_next_data_entry_perm_u <= io_ptw_resp_bits_data_entry_perm_u; // @[Reg.scala 17:22]
    end
    if (io_ptw_resp_valid) begin // @[Reg.scala 17:18]
      ptw_resp_next_data_entry_perm_x <= io_ptw_resp_bits_data_entry_perm_x; // @[Reg.scala 17:22]
    end
    if (io_ptw_resp_valid) begin // @[Reg.scala 17:18]
      ptw_resp_next_data_entry_perm_w <= io_ptw_resp_bits_data_entry_perm_w; // @[Reg.scala 17:22]
    end
    if (io_ptw_resp_valid) begin // @[Reg.scala 17:18]
      ptw_resp_next_data_entry_perm_r <= io_ptw_resp_bits_data_entry_perm_r; // @[Reg.scala 17:22]
    end
    if (io_ptw_resp_valid) begin // @[Reg.scala 17:18]
      ptw_resp_next_data_entry_level <= io_ptw_resp_bits_data_entry_level; // @[Reg.scala 17:22]
    end
    if (io_ptw_resp_valid) begin // @[Reg.scala 17:18]
      ptw_resp_next_data_pf <= io_ptw_resp_bits_data_pf; // @[Reg.scala 17:22]
    end
    if (io_ptw_resp_valid) begin // @[Reg.scala 17:18]
      ptw_resp_next_data_af <= io_ptw_resp_bits_data_af; // @[Reg.scala 17:22]
    end
    if (io_ptw_resp_valid) begin // @[Reg.scala 17:18]
      ptw_resp_next_vector_0 <= io_ptw_resp_bits_vector_0; // @[Reg.scala 17:22]
    end
    if (io_ptw_resp_valid) begin // @[Reg.scala 17:18]
      ptw_resp_next_vector_1 <= io_ptw_resp_bits_vector_1; // @[Reg.scala 17:22]
    end
    if (io_ptw_resp_valid) begin // @[Reg.scala 17:18]
      ptw_resp_next_vector_2 <= io_ptw_resp_bits_vector_2; // @[Reg.scala 17:22]
    end
    if (io_ptw_resp_valid) begin // @[Reg.scala 17:18]
      ptw_resp_next_vector_3 <= io_ptw_resp_bits_vector_3; // @[Reg.scala 17:22]
    end
    if (io_ptw_resp_valid) begin // @[Reg.scala 17:18]
      ptw_resp_next_vector_4 <= io_ptw_resp_bits_vector_4; // @[Reg.scala 17:22]
    end
    io_fenceToSbuffer_sbIsEmpty_REG <= sbuffer_io_flush_empty & uncache_io_flush_empty; // @[MemBlock.scala 566:42]
    sbuffer_io_flush_valid_REG <= io_fenceToSbuffer_flushSb | atomicsUnit_io_flush_sbuffer_valid; // @[MemBlock.scala 572:48]
    if (atomicsUnit_io_exceptionAddr_valid) begin // @[Reg.scala 17:18]
      atomicsExceptionAddress <= atomicsUnit_io_exceptionAddr_bits; // @[Reg.scala 17:22]
    end
    if (atomicsException) begin // @[MemBlock.scala 668:46]
      io_lsqio_exceptionAddr_vaddr_REG <= atomicsExceptionAddress;
    end else begin
      io_lsqio_exceptionAddr_vaddr_REG <= lsq_io_exceptionAddr_vaddr;
    end
    io_perf_0_value_REG <= hpm_io_perf_0_value; // @[PerfCounterUtils.scala 188:35]
    io_perf_0_value_REG_1 <= io_perf_0_value_REG; // @[PerfCounterUtils.scala 188:27]
    io_perf_1_value_REG <= hpm_io_perf_1_value; // @[PerfCounterUtils.scala 188:35]
    io_perf_1_value_REG_1 <= io_perf_1_value_REG; // @[PerfCounterUtils.scala 188:27]
    io_perf_2_value_REG <= hpm_io_perf_2_value; // @[PerfCounterUtils.scala 188:35]
    io_perf_2_value_REG_1 <= io_perf_2_value_REG; // @[PerfCounterUtils.scala 188:27]
    io_perf_3_value_REG <= hpm_io_perf_3_value; // @[PerfCounterUtils.scala 188:35]
    io_perf_3_value_REG_1 <= io_perf_3_value_REG; // @[PerfCounterUtils.scala 188:27]
    io_perf_4_value_REG <= hpm_io_perf_4_value; // @[PerfCounterUtils.scala 188:35]
    io_perf_4_value_REG_1 <= io_perf_4_value_REG; // @[PerfCounterUtils.scala 188:27]
    io_perf_5_value_REG <= hpm_io_perf_5_value; // @[PerfCounterUtils.scala 188:35]
    io_perf_5_value_REG_1 <= io_perf_5_value_REG; // @[PerfCounterUtils.scala 188:27]
    io_perf_6_value_REG <= hpm_io_perf_6_value; // @[PerfCounterUtils.scala 188:35]
    io_perf_6_value_REG_1 <= io_perf_6_value_REG; // @[PerfCounterUtils.scala 188:27]
    io_perf_7_value_REG <= hpm_io_perf_7_value; // @[PerfCounterUtils.scala 188:35]
    io_perf_7_value_REG_1 <= io_perf_7_value_REG; // @[PerfCounterUtils.scala 188:27]
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BitUtils.scala 28:28]
      redirect_next_valid_REG <= 1'h0; // @[BitUtils.scala 28:28]
    end else begin
      redirect_next_valid_REG <= io_redirect_valid; // @[BitUtils.scala 28:28]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[MemBlock.scala 281:46]
      ptw_resp_v <= 1'h0;
    end else begin
      ptw_resp_v <= io_ptw_resp_valid & ~(sfence_valid & tlbcsr_satp_changed);
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[MemBlock.scala 328:37]
      tdata_0_matchType <= 2'h0; // @[MemBlock.scala 324:22 329:{44,44}]
    end else if (csrCtrl_delay_io_out_mem_trigger_t_valid) begin // @[MemBlock.scala 324:22]
      if (3'h0 == csrCtrl_delay_io_out_mem_trigger_t_bits_addr) begin
        tdata_0_matchType <= _tdata_csrCtrl_delay_io_out_mem_trigger_t_bits_addr_matchType;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[MemBlock.scala 328:37]
      tdata_0_select <= 1'h0; // @[MemBlock.scala 324:22 329:{44,44}]
    end else if (csrCtrl_delay_io_out_mem_trigger_t_valid) begin // @[MemBlock.scala 324:22]
      if (3'h0 == csrCtrl_delay_io_out_mem_trigger_t_bits_addr) begin
        tdata_0_select <= csrCtrl_delay_io_out_mem_trigger_t_bits_tdata_select;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[MemBlock.scala 328:37]
      tdata_0_chain <= 1'h0; // @[MemBlock.scala 324:22 329:{44,44}]
    end else if (csrCtrl_delay_io_out_mem_trigger_t_valid) begin // @[MemBlock.scala 324:22]
      if (3'h0 == csrCtrl_delay_io_out_mem_trigger_t_bits_addr) begin
        tdata_0_chain <= csrCtrl_delay_io_out_mem_trigger_t_bits_tdata_chain;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[MemBlock.scala 328:37]
      tdata_0_tdata2 <= 64'h0; // @[MemBlock.scala 324:22 329:{44,44}]
    end else if (csrCtrl_delay_io_out_mem_trigger_t_valid) begin // @[MemBlock.scala 324:22]
      if (3'h0 == csrCtrl_delay_io_out_mem_trigger_t_bits_addr) begin
        tdata_0_tdata2 <= _tdata_csrCtrl_delay_io_out_mem_trigger_t_bits_addr_tdata2;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[MemBlock.scala 328:37]
      tdata_1_matchType <= 2'h0; // @[MemBlock.scala 324:22 329:{44,44}]
    end else if (csrCtrl_delay_io_out_mem_trigger_t_valid) begin // @[MemBlock.scala 324:22]
      if (3'h1 == csrCtrl_delay_io_out_mem_trigger_t_bits_addr) begin
        tdata_1_matchType <= _tdata_csrCtrl_delay_io_out_mem_trigger_t_bits_addr_matchType;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[MemBlock.scala 328:37]
      tdata_1_select <= 1'h0; // @[MemBlock.scala 324:22 329:{44,44}]
    end else if (csrCtrl_delay_io_out_mem_trigger_t_valid) begin // @[MemBlock.scala 324:22]
      if (3'h1 == csrCtrl_delay_io_out_mem_trigger_t_bits_addr) begin
        tdata_1_select <= csrCtrl_delay_io_out_mem_trigger_t_bits_tdata_select;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[MemBlock.scala 328:37]
      tdata_1_tdata2 <= 64'h0; // @[MemBlock.scala 324:22 329:{44,44}]
    end else if (csrCtrl_delay_io_out_mem_trigger_t_valid) begin // @[MemBlock.scala 324:22]
      if (3'h1 == csrCtrl_delay_io_out_mem_trigger_t_bits_addr) begin
        tdata_1_tdata2 <= _tdata_csrCtrl_delay_io_out_mem_trigger_t_bits_addr_tdata2;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[MemBlock.scala 328:37]
      tdata_2_matchType <= 2'h0; // @[MemBlock.scala 324:22 329:{44,44}]
    end else if (csrCtrl_delay_io_out_mem_trigger_t_valid) begin // @[MemBlock.scala 324:22]
      if (3'h2 == csrCtrl_delay_io_out_mem_trigger_t_bits_addr) begin
        tdata_2_matchType <= _tdata_csrCtrl_delay_io_out_mem_trigger_t_bits_addr_matchType;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[MemBlock.scala 328:37]
      tdata_2_select <= 1'h0; // @[MemBlock.scala 324:22 329:{44,44}]
    end else if (csrCtrl_delay_io_out_mem_trigger_t_valid) begin // @[MemBlock.scala 324:22]
      if (3'h2 == csrCtrl_delay_io_out_mem_trigger_t_bits_addr) begin
        tdata_2_select <= csrCtrl_delay_io_out_mem_trigger_t_bits_tdata_select;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[MemBlock.scala 328:37]
      tdata_2_chain <= 1'h0; // @[MemBlock.scala 324:22 329:{44,44}]
    end else if (csrCtrl_delay_io_out_mem_trigger_t_valid) begin // @[MemBlock.scala 324:22]
      if (3'h2 == csrCtrl_delay_io_out_mem_trigger_t_bits_addr) begin
        tdata_2_chain <= csrCtrl_delay_io_out_mem_trigger_t_bits_tdata_chain;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[MemBlock.scala 328:37]
      tdata_2_tdata2 <= 64'h0; // @[MemBlock.scala 324:22 329:{44,44}]
    end else if (csrCtrl_delay_io_out_mem_trigger_t_valid) begin // @[MemBlock.scala 324:22]
      if (3'h2 == csrCtrl_delay_io_out_mem_trigger_t_bits_addr) begin
        tdata_2_tdata2 <= _tdata_csrCtrl_delay_io_out_mem_trigger_t_bits_addr_tdata2;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[MemBlock.scala 328:37]
      tdata_3_matchType <= 2'h0; // @[MemBlock.scala 324:22 329:{44,44}]
    end else if (csrCtrl_delay_io_out_mem_trigger_t_valid) begin // @[MemBlock.scala 324:22]
      if (3'h3 == csrCtrl_delay_io_out_mem_trigger_t_bits_addr) begin
        tdata_3_matchType <= _tdata_csrCtrl_delay_io_out_mem_trigger_t_bits_addr_matchType;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[MemBlock.scala 328:37]
      tdata_3_select <= 1'h0; // @[MemBlock.scala 324:22 329:{44,44}]
    end else if (csrCtrl_delay_io_out_mem_trigger_t_valid) begin // @[MemBlock.scala 324:22]
      if (3'h3 == csrCtrl_delay_io_out_mem_trigger_t_bits_addr) begin
        tdata_3_select <= csrCtrl_delay_io_out_mem_trigger_t_bits_tdata_select;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[MemBlock.scala 328:37]
      tdata_3_tdata2 <= 64'h0; // @[MemBlock.scala 324:22 329:{44,44}]
    end else if (csrCtrl_delay_io_out_mem_trigger_t_valid) begin // @[MemBlock.scala 324:22]
      if (3'h3 == csrCtrl_delay_io_out_mem_trigger_t_bits_addr) begin
        tdata_3_tdata2 <= _tdata_csrCtrl_delay_io_out_mem_trigger_t_bits_addr_tdata2;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[MemBlock.scala 328:37]
      tdata_4_matchType <= 2'h0; // @[MemBlock.scala 324:22 329:{44,44}]
    end else if (csrCtrl_delay_io_out_mem_trigger_t_valid) begin // @[MemBlock.scala 324:22]
      if (3'h4 == csrCtrl_delay_io_out_mem_trigger_t_bits_addr) begin
        tdata_4_matchType <= _tdata_csrCtrl_delay_io_out_mem_trigger_t_bits_addr_matchType;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[MemBlock.scala 328:37]
      tdata_4_select <= 1'h0; // @[MemBlock.scala 324:22 329:{44,44}]
    end else if (csrCtrl_delay_io_out_mem_trigger_t_valid) begin // @[MemBlock.scala 324:22]
      if (3'h4 == csrCtrl_delay_io_out_mem_trigger_t_bits_addr) begin
        tdata_4_select <= csrCtrl_delay_io_out_mem_trigger_t_bits_tdata_select;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[MemBlock.scala 328:37]
      tdata_4_tdata2 <= 64'h0; // @[MemBlock.scala 324:22 329:{44,44}]
    end else if (csrCtrl_delay_io_out_mem_trigger_t_valid) begin // @[MemBlock.scala 324:22]
      if (3'h4 == csrCtrl_delay_io_out_mem_trigger_t_bits_addr) begin
        tdata_4_tdata2 <= _tdata_csrCtrl_delay_io_out_mem_trigger_t_bits_addr_tdata2;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[MemBlock.scala 328:37]
      tdata_5_matchType <= 2'h0; // @[MemBlock.scala 324:22 329:{44,44}]
    end else if (csrCtrl_delay_io_out_mem_trigger_t_valid) begin // @[MemBlock.scala 324:22]
      if (3'h5 == csrCtrl_delay_io_out_mem_trigger_t_bits_addr) begin
        tdata_5_matchType <= _tdata_csrCtrl_delay_io_out_mem_trigger_t_bits_addr_matchType;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[MemBlock.scala 328:37]
      tdata_5_select <= 1'h0; // @[MemBlock.scala 324:22 329:{44,44}]
    end else if (csrCtrl_delay_io_out_mem_trigger_t_valid) begin // @[MemBlock.scala 324:22]
      if (3'h5 == csrCtrl_delay_io_out_mem_trigger_t_bits_addr) begin
        tdata_5_select <= csrCtrl_delay_io_out_mem_trigger_t_bits_tdata_select;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[MemBlock.scala 328:37]
      tdata_5_tdata2 <= 64'h0; // @[MemBlock.scala 324:22 329:{44,44}]
    end else if (csrCtrl_delay_io_out_mem_trigger_t_valid) begin // @[MemBlock.scala 324:22]
      if (3'h5 == csrCtrl_delay_io_out_mem_trigger_t_bits_addr) begin
        tdata_5_tdata2 <= _tdata_csrCtrl_delay_io_out_mem_trigger_t_bits_addr_tdata2;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[MemBlock.scala 327:{21,21}]
      tEnable_0 <= 1'h0;
    end else begin
      tEnable_0 <= csrCtrl_delay_io_out_trigger_enable_2;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[MemBlock.scala 327:{21,21}]
      tEnable_1 <= 1'h0;
    end else begin
      tEnable_1 <= csrCtrl_delay_io_out_trigger_enable_3;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[MemBlock.scala 327:{21,21}]
      tEnable_2 <= 1'h0;
    end else begin
      tEnable_2 <= csrCtrl_delay_io_out_trigger_enable_4;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[MemBlock.scala 327:{21,21}]
      tEnable_3 <= 1'h0;
    end else begin
      tEnable_3 <= csrCtrl_delay_io_out_trigger_enable_5;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[MemBlock.scala 327:{21,21}]
      tEnable_4 <= 1'h0;
    end else begin
      tEnable_4 <= csrCtrl_delay_io_out_trigger_enable_7;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[MemBlock.scala 327:{21,21}]
      tEnable_5 <= 1'h0;
    end else begin
      tEnable_5 <= csrCtrl_delay_io_out_trigger_enable_9;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[MemBlock.scala 610:35]
      state <= 2'h0; // @[MemBlock.scala 612:11]
    end else if (atomicsUnit_io_out_valid) begin // @[MemBlock.scala 602:63]
      state <= 2'h0; // @[MemBlock.scala 606:11]
    end else if (st_atomics_1) begin // @[MemBlock.scala 602:63]
      state <= 2'h2; // @[MemBlock.scala 606:11]
    end else if (st_atomics_0) begin // @[MemBlock.scala 590:22]
      state <= 2'h1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[MemBlock.scala 662:57]
      atomicsException <= 1'h0; // @[MemBlock.scala 663:22]
    end else if (delay_io_out & atomicsException) begin
      atomicsException <= 1'h0;
    end else begin
      atomicsException <= _GEN_670;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  redirect_next_valid_REG = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  redirect_next_bits_rrobIdx_flag = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  redirect_next_bits_rrobIdx_value = _RAND_2[4:0];
  _RAND_3 = {1{`RANDOM}};
  redirect_next_bits_rlevel = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  delayedDcacheRefill_valid = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  delayedDcacheRefill_bits_id = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  io_csrUpdate_REG_wvalid = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  io_csrUpdate_REG_waddr = _RAND_7[11:0];
  _RAND_8 = {2{`RANDOM}};
  io_csrUpdate_REG_wdata = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  io_error_REG_paddr = _RAND_9[35:0];
  _RAND_10 = {1{`RANDOM}};
  io_error_REG_report_to_beu = _RAND_10[0:0];
  _RAND_11 = {2{`RANDOM}};
  io_error_REG_1_paddr = _RAND_11[35:0];
  _RAND_12 = {1{`RANDOM}};
  io_error_REG_1_report_to_beu = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  sfence_REG_valid = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  sfence_REG_bits_rs1 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  sfence_REG_bits_rs2 = _RAND_15[0:0];
  _RAND_16 = {2{`RANDOM}};
  sfence_REG_bits_addr = _RAND_16[38:0];
  _RAND_17 = {1{`RANDOM}};
  sfence_REG_bits_asid = _RAND_17[15:0];
  _RAND_18 = {1{`RANDOM}};
  sfence_valid = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  sfence_bits_rs1 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  sfence_bits_rs2 = _RAND_20[0:0];
  _RAND_21 = {2{`RANDOM}};
  sfence_bits_addr = _RAND_21[38:0];
  _RAND_22 = {1{`RANDOM}};
  sfence_bits_asid = _RAND_22[15:0];
  _RAND_23 = {1{`RANDOM}};
  tlbcsr_REG_satp_mode = _RAND_23[3:0];
  _RAND_24 = {1{`RANDOM}};
  tlbcsr_REG_satp_asid = _RAND_24[15:0];
  _RAND_25 = {1{`RANDOM}};
  tlbcsr_REG_satp_changed = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  tlbcsr_REG_priv_mxr = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  tlbcsr_REG_priv_sum = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  tlbcsr_REG_priv_dmode = _RAND_28[1:0];
  _RAND_29 = {1{`RANDOM}};
  tlbcsr_satp_mode = _RAND_29[3:0];
  _RAND_30 = {1{`RANDOM}};
  tlbcsr_satp_asid = _RAND_30[15:0];
  _RAND_31 = {1{`RANDOM}};
  tlbcsr_satp_changed = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  tlbcsr_priv_mxr = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  tlbcsr_priv_sum = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  tlbcsr_priv_dmode = _RAND_34[1:0];
  _RAND_35 = {1{`RANDOM}};
  ptw_resp_next_data_entry_tag = _RAND_35[26:0];
  _RAND_36 = {1{`RANDOM}};
  ptw_resp_next_data_entry_asid = _RAND_36[15:0];
  _RAND_37 = {1{`RANDOM}};
  ptw_resp_next_data_entry_ppn = _RAND_37[23:0];
  _RAND_38 = {1{`RANDOM}};
  ptw_resp_next_data_entry_perm_d = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  ptw_resp_next_data_entry_perm_a = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  ptw_resp_next_data_entry_perm_g = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  ptw_resp_next_data_entry_perm_u = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  ptw_resp_next_data_entry_perm_x = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  ptw_resp_next_data_entry_perm_w = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  ptw_resp_next_data_entry_perm_r = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  ptw_resp_next_data_entry_level = _RAND_45[1:0];
  _RAND_46 = {1{`RANDOM}};
  ptw_resp_next_data_pf = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  ptw_resp_next_data_af = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  ptw_resp_next_vector_0 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  ptw_resp_next_vector_1 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  ptw_resp_next_vector_2 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  ptw_resp_next_vector_3 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  ptw_resp_next_vector_4 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  ptw_resp_v = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  tdata_0_matchType = _RAND_54[1:0];
  _RAND_55 = {1{`RANDOM}};
  tdata_0_select = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  tdata_0_chain = _RAND_56[0:0];
  _RAND_57 = {2{`RANDOM}};
  tdata_0_tdata2 = _RAND_57[63:0];
  _RAND_58 = {1{`RANDOM}};
  tdata_1_matchType = _RAND_58[1:0];
  _RAND_59 = {1{`RANDOM}};
  tdata_1_select = _RAND_59[0:0];
  _RAND_60 = {2{`RANDOM}};
  tdata_1_tdata2 = _RAND_60[63:0];
  _RAND_61 = {1{`RANDOM}};
  tdata_2_matchType = _RAND_61[1:0];
  _RAND_62 = {1{`RANDOM}};
  tdata_2_select = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  tdata_2_chain = _RAND_63[0:0];
  _RAND_64 = {2{`RANDOM}};
  tdata_2_tdata2 = _RAND_64[63:0];
  _RAND_65 = {1{`RANDOM}};
  tdata_3_matchType = _RAND_65[1:0];
  _RAND_66 = {1{`RANDOM}};
  tdata_3_select = _RAND_66[0:0];
  _RAND_67 = {2{`RANDOM}};
  tdata_3_tdata2 = _RAND_67[63:0];
  _RAND_68 = {1{`RANDOM}};
  tdata_4_matchType = _RAND_68[1:0];
  _RAND_69 = {1{`RANDOM}};
  tdata_4_select = _RAND_69[0:0];
  _RAND_70 = {2{`RANDOM}};
  tdata_4_tdata2 = _RAND_70[63:0];
  _RAND_71 = {1{`RANDOM}};
  tdata_5_matchType = _RAND_71[1:0];
  _RAND_72 = {1{`RANDOM}};
  tdata_5_select = _RAND_72[0:0];
  _RAND_73 = {2{`RANDOM}};
  tdata_5_tdata2 = _RAND_73[63:0];
  _RAND_74 = {1{`RANDOM}};
  tEnable_0 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  tEnable_1 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  tEnable_2 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  tEnable_3 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  tEnable_4 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  tEnable_5 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  io_fenceToSbuffer_sbIsEmpty_REG = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  sbuffer_io_flush_valid_REG = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  state = _RAND_82[1:0];
  _RAND_83 = {1{`RANDOM}};
  atomicsException = _RAND_83[0:0];
  _RAND_84 = {2{`RANDOM}};
  atomicsExceptionAddress = _RAND_84[38:0];
  _RAND_85 = {2{`RANDOM}};
  io_lsqio_exceptionAddr_vaddr_REG = _RAND_85[38:0];
  _RAND_86 = {1{`RANDOM}};
  io_perf_0_value_REG = _RAND_86[5:0];
  _RAND_87 = {1{`RANDOM}};
  io_perf_0_value_REG_1 = _RAND_87[5:0];
  _RAND_88 = {1{`RANDOM}};
  io_perf_1_value_REG = _RAND_88[5:0];
  _RAND_89 = {1{`RANDOM}};
  io_perf_1_value_REG_1 = _RAND_89[5:0];
  _RAND_90 = {1{`RANDOM}};
  io_perf_2_value_REG = _RAND_90[5:0];
  _RAND_91 = {1{`RANDOM}};
  io_perf_2_value_REG_1 = _RAND_91[5:0];
  _RAND_92 = {1{`RANDOM}};
  io_perf_3_value_REG = _RAND_92[5:0];
  _RAND_93 = {1{`RANDOM}};
  io_perf_3_value_REG_1 = _RAND_93[5:0];
  _RAND_94 = {1{`RANDOM}};
  io_perf_4_value_REG = _RAND_94[5:0];
  _RAND_95 = {1{`RANDOM}};
  io_perf_4_value_REG_1 = _RAND_95[5:0];
  _RAND_96 = {1{`RANDOM}};
  io_perf_5_value_REG = _RAND_96[5:0];
  _RAND_97 = {1{`RANDOM}};
  io_perf_5_value_REG_1 = _RAND_97[5:0];
  _RAND_98 = {1{`RANDOM}};
  io_perf_6_value_REG = _RAND_98[5:0];
  _RAND_99 = {1{`RANDOM}};
  io_perf_6_value_REG_1 = _RAND_99[5:0];
  _RAND_100 = {1{`RANDOM}};
  io_perf_7_value_REG = _RAND_100[5:0];
  _RAND_101 = {1{`RANDOM}};
  io_perf_7_value_REG_1 = _RAND_101[5:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    redirect_next_valid_REG = 1'h0;
  end
  if (reset) begin
    ptw_resp_v = 1'h0;
  end
  if (reset) begin
    tdata_0_matchType = 2'h0;
  end
  if (reset) begin
    tdata_0_select = 1'h0;
  end
  if (reset) begin
    tdata_0_chain = 1'h0;
  end
  if (reset) begin
    tdata_0_tdata2 = 64'h0;
  end
  if (reset) begin
    tdata_1_matchType = 2'h0;
  end
  if (reset) begin
    tdata_1_select = 1'h0;
  end
  if (reset) begin
    tdata_1_tdata2 = 64'h0;
  end
  if (reset) begin
    tdata_2_matchType = 2'h0;
  end
  if (reset) begin
    tdata_2_select = 1'h0;
  end
  if (reset) begin
    tdata_2_chain = 1'h0;
  end
  if (reset) begin
    tdata_2_tdata2 = 64'h0;
  end
  if (reset) begin
    tdata_3_matchType = 2'h0;
  end
  if (reset) begin
    tdata_3_select = 1'h0;
  end
  if (reset) begin
    tdata_3_tdata2 = 64'h0;
  end
  if (reset) begin
    tdata_4_matchType = 2'h0;
  end
  if (reset) begin
    tdata_4_select = 1'h0;
  end
  if (reset) begin
    tdata_4_tdata2 = 64'h0;
  end
  if (reset) begin
    tdata_5_matchType = 2'h0;
  end
  if (reset) begin
    tdata_5_select = 1'h0;
  end
  if (reset) begin
    tdata_5_tdata2 = 64'h0;
  end
  if (reset) begin
    tEnable_0 = 1'h0;
  end
  if (reset) begin
    tEnable_1 = 1'h0;
  end
  if (reset) begin
    tEnable_2 = 1'h0;
  end
  if (reset) begin
    tEnable_3 = 1'h0;
  end
  if (reset) begin
    tEnable_4 = 1'h0;
  end
  if (reset) begin
    tEnable_5 = 1'h0;
  end
  if (reset) begin
    state = 2'h0;
  end
  if (reset) begin
    atomicsException = 1'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule

