module bosc_mbist_controller_L1L2_dfx_top(
  input          io_mbist_ijtag_tck,
  input          io_mbist_ijtag_reset,
  input          io_mbist_ijtag_ce,
  input          io_mbist_ijtag_se,
  input          io_mbist_ijtag_ue,
  input          io_mbist_ijtag_sel,
  input          io_mbist_ijtag_si,
  output         io_mbist_ijtag_so,
  output         io_mbist_ijtag_diag_done,
  output [10:0]  io_hd2prf_out_trim_fuse,
  output [1:0]   io_hd2prf_out_sleep_fuse,
  output [19:0]  io_hsuspsr_out_trim_fuse,
  output [1:0]   io_hsuspsr_out_sleep_fuse,
  output [19:0]  io_uhdusplr_out_trim_fuse,
  output [1:0]   io_uhdusplr_out_sleep_fuse,
  output [19:0]  io_hduspsr_out_trim_fuse,
  output [1:0]   io_hduspsr_out_sleep_fuse,
  input  [10:0]  io_hd2prf_in_trim_fuse,
  input  [1:0]   io_hd2prf_in_sleep_fuse,
  input  [19:0]  io_hsuspsr_in_trim_fuse,
  input  [1:0]   io_hsuspsr_in_sleep_fuse,
  input  [19:0]  io_uhdusplr_in_trim_fuse,
  input  [1:0]   io_uhdusplr_in_sleep_fuse,
  input  [19:0]  io_hduspsr_in_trim_fuse,
  input  [1:0]   io_hduspsr_in_sleep_fuse,
  input          io_xsx_fscan_in_bypsel,
  input          io_xsx_fscan_in_wdis_b,
  input          io_xsx_fscan_in_rdis_b,
  input          io_xsx_fscan_in_init_en,
  input          io_xsx_fscan_in_init_val,
  input          io_xsl2_fscan_in_bypsel,
  input          io_xsl2_fscan_in_wdis_b,
  input          io_xsl2_fscan_in_rdis_b,
  input          io_xsl2_fscan_in_init_en,
  input          io_xsl2_fscan_in_init_val,
  input          io_fscan_clkungate,
  input          io_clock,
  output [4:0]   io_L1_SRAM_array,
  output         io_L1_SRAM_all,
  output         io_L1_SRAM_req,
  input          io_L1_SRAM_ack,
  output         io_L1_SRAM_writeen,
  output [15:0]  io_L1_SRAM_be,
  output [9:0]   io_L1_SRAM_addr,
  output [159:0] io_L1_SRAM_indata,
  output         io_L1_SRAM_readen,
  input  [159:0] io_L1_SRAM_outdata,
  output [7:0]   io_L1_RF_array,
  output         io_L1_RF_all,
  output         io_L1_RF_req,
  input          io_L1_RF_ack,
  output         io_L1_RF_writeen,
  output [7:0]   io_L1_RF_be,
  output [11:0]  io_L1_RF_addr,
  output [255:0] io_L1_RF_indata,
  output         io_L1_RF_readen,
  output [11:0]  io_L1_RF_addr_rd,
  input  [255:0] io_L1_RF_outdata,
  output [6:0]   io_L2_SRAM_array,
  output         io_L2_SRAM_all,
  output         io_L2_SRAM_req,
  input          io_L2_SRAM_ack,
  output         io_L2_SRAM_writeen,
  output [7:0]   io_L2_SRAM_be,
  output [10:0]  io_L2_SRAM_addr,
  output [175:0] io_L2_SRAM_indata,
  output         io_L2_SRAM_readen,
  input  [175:0] io_L2_SRAM_outdata,
  output [3:0]   io_L2_RF_array,
  output         io_L2_RF_all,
  output         io_L2_RF_req,
  input          io_L2_RF_ack,
  output         io_L2_RF_writeen,
  output [9:0]   io_L2_RF_be,
  output [8:0]   io_L2_RF_addr,
  output [229:0] io_L2_RF_indata,
  output         io_L2_RF_readen,
  output [8:0]   io_L2_RF_addr_rd,
  input  [229:0] io_L2_RF_outdata,
  output         io_fscan_ram_L1_bypsel,
  output         io_fscan_ram_L1_wdis_b,
  output         io_fscan_ram_L1_rdis_b,
  output         io_fscan_ram_L1_init_en,
  output         io_fscan_ram_L1_init_val,
  output         io_fscan_ram_L1_clkungate,
  output         io_fscan_ram_L2_bypsel,
  output         io_fscan_ram_L2_wdis_b,
  output         io_fscan_ram_L2_rdis_b,
  output         io_fscan_ram_L2_init_en,
  output         io_fscan_ram_L2_init_val,
  output         io_fscan_ram_L2_clkungate
);
  mbist_controller_L1L2_dfx_wrap mbistControllerCoreWithL2 ( // @[XSTile.scala 291:45]
    .i_L1L2_mbist_ijtag_tck(io_mbist_ijtag_tck),
    .i_L1L2_mbist_ijtag_reset(io_mbist_ijtag_reset),
    .i_L1L2_mbist_ijtag_ce(io_mbist_ijtag_ce),
    .i_L1L2_mbist_ijtag_se(io_mbist_ijtag_se),
    .i_L1L2_mbist_ijtag_ue(io_mbist_ijtag_ue),
    .i_L1L2_mbist_ijtag_sel(io_mbist_ijtag_sel),
    .i_L1L2_mbist_ijtag_si(io_mbist_ijtag_si),
    .o_L1L2_mbist_ijtag_so(io_mbist_ijtag_so),
    .o_L1L2_aary_mbist_diag_done(io_mbist_ijtag_diag_done),
    .o_L1L2_hd2prf_trim_fuse_out(io_hd2prf_out_trim_fuse),
    .o_L1L2_hd2prf_sleep_fuse_out(io_hd2prf_out_sleep_fuse),
    .o_L1L2_hsuspsr_trim_fuse_out(io_hsuspsr_out_trim_fuse),
    .o_L1L2_hsuspsr_sleep_fuse_out(io_hsuspsr_out_sleep_fuse),
    .o_L1L2_hduspsr_trim_fuse_out(io_hduspsr_out_trim_fuse),
    .o_L1L2_hduspsr_sleep_fuse_out(io_hduspsr_out_sleep_fuse),
    .i_L1L2_hd2prf_trim_fuse_in(io_hd2prf_in_trim_fuse),
    .i_L1L2_hd2prf_sleep_fuse_in(io_hd2prf_in_sleep_fuse),
    .i_L1L2_hsuspsr_trim_fuse_in(io_hsuspsr_in_trim_fuse),
    .i_L1L2_hsuspsr_sleep_fuse_in(io_hsuspsr_in_sleep_fuse),
    .i_L1L2_hduspsr_trim_fuse_in(io_hduspsr_in_trim_fuse),
    .i_L1L2_hduspsr_sleep_fuse_in(io_hduspsr_in_sleep_fuse),
    .i_xsx_fscan_ram_bypsel(io_xsx_fscan_in_bypsel),
    .i_xsx_fscan_ram_wdis_b(io_xsx_fscan_in_wdis_b),
    .i_xsx_fscan_ram_rdis_b(io_xsx_fscan_in_rdis_b),
    .i_xsx_fscan_ram_init_en(io_xsx_fscan_in_init_en),
    .i_xsx_fscan_ram_init_val(io_xsx_fscan_in_init_val),
    .i_xsl2_fscan_ram_bypsel(io_xsl2_fscan_in_bypsel),
    .i_xsl2_fscan_ram_wdis_b(io_xsl2_fscan_in_wdis_b),
    .i_xsl2_fscan_ram_rdis_b(io_xsl2_fscan_in_rdis_b),
    .i_xsl2_fscan_ram_init_en(io_xsl2_fscan_in_init_en),
    .i_xsl2_fscan_ram_init_val(io_xsl2_fscan_in_init_val),
    .i_fscan_clkungate(io_fscan_clkungate),
    .core_with_l2_clock(io_clock),
    .o_L1_sram_mbist_array(io_L1_SRAM_array),
    .o_L1_sram_mbist_all(io_L1_SRAM_all),
    .o_L1_sram_mbist_req(io_L1_SRAM_req),
    .i_L1_sram_mbist_ack(io_L1_SRAM_ack),
    .o_L1_sram_mbist_writeen(io_L1_SRAM_writeen),
    .o_L1_sram_mbist_be(io_L1_SRAM_be),
    .o_L1_sram_mbist_addr(io_L1_SRAM_addr),
    .o_L1_sram_mbist_indata(io_L1_SRAM_indata),
    .o_L1_sram_mbist_readen(io_L1_SRAM_readen),
    .i_L1_sram_mbist_outdata(io_L1_SRAM_outdata),
    .o_L1_rf_mbist_array(io_L1_RF_array),
    .o_L1_rf_mbist_all(io_L1_RF_all),
    .o_L1_rf_mbist_req(io_L1_RF_req),
    .i_L1_rf_mbist_ack(io_L1_RF_ack),
    .o_L1_rf_mbist_writeen(io_L1_RF_writeen),
    .o_L1_rf_mbist_be(io_L1_RF_be),
    .o_L1_rf_mbist_addr(io_L1_RF_addr),
    .o_L1_rf_mbist_indata(io_L1_RF_indata),
    .o_L1_rf_mbist_readen(io_L1_RF_readen),
    .o_L1_rf_mbist_addr_rd(io_L1_RF_addr_rd),
    .i_L1_rf_mbist_outdata(io_L1_RF_outdata),
    .o_L2_sram_mbist_array(io_L2_SRAM_array),
    .o_L2_sram_mbist_all(io_L2_SRAM_all),
    .o_L2_sram_mbist_req(io_L2_SRAM_req),
    .i_L2_sram_mbist_ack(io_L2_SRAM_ack),
    .o_L2_sram_mbist_writeen(io_L2_SRAM_writeen),
    .o_L2_sram_mbist_be(io_L2_SRAM_be),
    .o_L2_sram_mbist_addr(io_L2_SRAM_addr),
    .o_L2_sram_mbist_indata(io_L2_SRAM_indata),
    .o_L2_sram_mbist_readen(io_L2_SRAM_readen),
    .i_L2_sram_mbist_outdata(io_L2_SRAM_outdata),
    .o_L2_rf_mbist_array(io_L2_RF_array),
    .o_L2_rf_mbist_all(io_L2_RF_all),
    .o_L2_rf_mbist_req(io_L2_RF_req),
    .i_L2_rf_mbist_ack(io_L2_RF_ack),
    .o_L2_rf_mbist_writeen(io_L2_RF_writeen),
    .o_L2_rf_mbist_be(io_L2_RF_be),
    .o_L2_rf_mbist_addr(io_L2_RF_addr),
    .o_L2_rf_mbist_indata(io_L2_RF_indata),
    .o_L2_rf_mbist_readen(io_L2_RF_readen),
    .o_L2_rf_mbist_addr_rd(io_L2_RF_addr_rd),
    .i_L2_rf_mbist_outdata(io_L2_RF_outdata),
    .o_L1_fscan_ram_bypsel(io_fscan_ram_L1_bypsel),
    .o_L1_fscan_ram_wdis_b(io_fscan_ram_L1_wdis_b),
    .o_L1_fscan_ram_rdis_b(io_fscan_ram_L1_rdis_b),
    .o_L1_fscan_ram_init_en(io_fscan_ram_L1_init_en),
    .o_L1_fscan_ram_init_val(io_fscan_ram_L1_init_val),
    .o_L1_fscan_clkungate(io_fscan_ram_L1_clkungate),
    .o_L2_fscan_ram_bypsel(io_fscan_ram_L2_bypsel),
    .o_L2_fscan_ram_wdis_b(io_fscan_ram_L2_wdis_b),
    .o_L2_fscan_ram_rdis_b(io_fscan_ram_L2_rdis_b),
    .o_L2_fscan_ram_init_en(io_fscan_ram_L2_init_en),
    .o_L2_fscan_ram_init_val(io_fscan_ram_L2_init_val),
    .o_L2_fscan_clkungate(io_fscan_ram_L2_clkungate)
  );
  assign io_uhdusplr_out_trim_fuse = 20'h0;
  assign io_uhdusplr_out_sleep_fuse = 2'h0;
endmodule

