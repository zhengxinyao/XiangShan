module LZA_4(
  input  [106:0] io_a,
  input  [106:0] io_b,
  output [106:0] io_f
);
  wire  k_0 = ~io_a[0] & ~io_b[0]; // @[LZA.scala 19:21]
  wire  p_1 = io_a[1] ^ io_b[1]; // @[LZA.scala 18:18]
  wire  k_1 = ~io_a[1] & ~io_b[1]; // @[LZA.scala 19:21]
  wire  f_1 = p_1 ^ ~k_0; // @[LZA.scala 23:20]
  wire  p_2 = io_a[2] ^ io_b[2]; // @[LZA.scala 18:18]
  wire  k_2 = ~io_a[2] & ~io_b[2]; // @[LZA.scala 19:21]
  wire  f_2 = p_2 ^ ~k_1; // @[LZA.scala 23:20]
  wire  p_3 = io_a[3] ^ io_b[3]; // @[LZA.scala 18:18]
  wire  k_3 = ~io_a[3] & ~io_b[3]; // @[LZA.scala 19:21]
  wire  f_3 = p_3 ^ ~k_2; // @[LZA.scala 23:20]
  wire  p_4 = io_a[4] ^ io_b[4]; // @[LZA.scala 18:18]
  wire  k_4 = ~io_a[4] & ~io_b[4]; // @[LZA.scala 19:21]
  wire  f_4 = p_4 ^ ~k_3; // @[LZA.scala 23:20]
  wire  p_5 = io_a[5] ^ io_b[5]; // @[LZA.scala 18:18]
  wire  k_5 = ~io_a[5] & ~io_b[5]; // @[LZA.scala 19:21]
  wire  f_5 = p_5 ^ ~k_4; // @[LZA.scala 23:20]
  wire  p_6 = io_a[6] ^ io_b[6]; // @[LZA.scala 18:18]
  wire  k_6 = ~io_a[6] & ~io_b[6]; // @[LZA.scala 19:21]
  wire  f_6 = p_6 ^ ~k_5; // @[LZA.scala 23:20]
  wire  p_7 = io_a[7] ^ io_b[7]; // @[LZA.scala 18:18]
  wire  k_7 = ~io_a[7] & ~io_b[7]; // @[LZA.scala 19:21]
  wire  f_7 = p_7 ^ ~k_6; // @[LZA.scala 23:20]
  wire  p_8 = io_a[8] ^ io_b[8]; // @[LZA.scala 18:18]
  wire  k_8 = ~io_a[8] & ~io_b[8]; // @[LZA.scala 19:21]
  wire  f_8 = p_8 ^ ~k_7; // @[LZA.scala 23:20]
  wire  p_9 = io_a[9] ^ io_b[9]; // @[LZA.scala 18:18]
  wire  k_9 = ~io_a[9] & ~io_b[9]; // @[LZA.scala 19:21]
  wire  f_9 = p_9 ^ ~k_8; // @[LZA.scala 23:20]
  wire  p_10 = io_a[10] ^ io_b[10]; // @[LZA.scala 18:18]
  wire  k_10 = ~io_a[10] & ~io_b[10]; // @[LZA.scala 19:21]
  wire  f_10 = p_10 ^ ~k_9; // @[LZA.scala 23:20]
  wire  p_11 = io_a[11] ^ io_b[11]; // @[LZA.scala 18:18]
  wire  k_11 = ~io_a[11] & ~io_b[11]; // @[LZA.scala 19:21]
  wire  f_11 = p_11 ^ ~k_10; // @[LZA.scala 23:20]
  wire  p_12 = io_a[12] ^ io_b[12]; // @[LZA.scala 18:18]
  wire  k_12 = ~io_a[12] & ~io_b[12]; // @[LZA.scala 19:21]
  wire  f_12 = p_12 ^ ~k_11; // @[LZA.scala 23:20]
  wire  p_13 = io_a[13] ^ io_b[13]; // @[LZA.scala 18:18]
  wire  k_13 = ~io_a[13] & ~io_b[13]; // @[LZA.scala 19:21]
  wire  f_13 = p_13 ^ ~k_12; // @[LZA.scala 23:20]
  wire  p_14 = io_a[14] ^ io_b[14]; // @[LZA.scala 18:18]
  wire  k_14 = ~io_a[14] & ~io_b[14]; // @[LZA.scala 19:21]
  wire  f_14 = p_14 ^ ~k_13; // @[LZA.scala 23:20]
  wire  p_15 = io_a[15] ^ io_b[15]; // @[LZA.scala 18:18]
  wire  k_15 = ~io_a[15] & ~io_b[15]; // @[LZA.scala 19:21]
  wire  f_15 = p_15 ^ ~k_14; // @[LZA.scala 23:20]
  wire  p_16 = io_a[16] ^ io_b[16]; // @[LZA.scala 18:18]
  wire  k_16 = ~io_a[16] & ~io_b[16]; // @[LZA.scala 19:21]
  wire  f_16 = p_16 ^ ~k_15; // @[LZA.scala 23:20]
  wire  p_17 = io_a[17] ^ io_b[17]; // @[LZA.scala 18:18]
  wire  k_17 = ~io_a[17] & ~io_b[17]; // @[LZA.scala 19:21]
  wire  f_17 = p_17 ^ ~k_16; // @[LZA.scala 23:20]
  wire  p_18 = io_a[18] ^ io_b[18]; // @[LZA.scala 18:18]
  wire  k_18 = ~io_a[18] & ~io_b[18]; // @[LZA.scala 19:21]
  wire  f_18 = p_18 ^ ~k_17; // @[LZA.scala 23:20]
  wire  p_19 = io_a[19] ^ io_b[19]; // @[LZA.scala 18:18]
  wire  k_19 = ~io_a[19] & ~io_b[19]; // @[LZA.scala 19:21]
  wire  f_19 = p_19 ^ ~k_18; // @[LZA.scala 23:20]
  wire  p_20 = io_a[20] ^ io_b[20]; // @[LZA.scala 18:18]
  wire  k_20 = ~io_a[20] & ~io_b[20]; // @[LZA.scala 19:21]
  wire  f_20 = p_20 ^ ~k_19; // @[LZA.scala 23:20]
  wire  p_21 = io_a[21] ^ io_b[21]; // @[LZA.scala 18:18]
  wire  k_21 = ~io_a[21] & ~io_b[21]; // @[LZA.scala 19:21]
  wire  f_21 = p_21 ^ ~k_20; // @[LZA.scala 23:20]
  wire  p_22 = io_a[22] ^ io_b[22]; // @[LZA.scala 18:18]
  wire  k_22 = ~io_a[22] & ~io_b[22]; // @[LZA.scala 19:21]
  wire  f_22 = p_22 ^ ~k_21; // @[LZA.scala 23:20]
  wire  p_23 = io_a[23] ^ io_b[23]; // @[LZA.scala 18:18]
  wire  k_23 = ~io_a[23] & ~io_b[23]; // @[LZA.scala 19:21]
  wire  f_23 = p_23 ^ ~k_22; // @[LZA.scala 23:20]
  wire  p_24 = io_a[24] ^ io_b[24]; // @[LZA.scala 18:18]
  wire  k_24 = ~io_a[24] & ~io_b[24]; // @[LZA.scala 19:21]
  wire  f_24 = p_24 ^ ~k_23; // @[LZA.scala 23:20]
  wire  p_25 = io_a[25] ^ io_b[25]; // @[LZA.scala 18:18]
  wire  k_25 = ~io_a[25] & ~io_b[25]; // @[LZA.scala 19:21]
  wire  f_25 = p_25 ^ ~k_24; // @[LZA.scala 23:20]
  wire  p_26 = io_a[26] ^ io_b[26]; // @[LZA.scala 18:18]
  wire  k_26 = ~io_a[26] & ~io_b[26]; // @[LZA.scala 19:21]
  wire  f_26 = p_26 ^ ~k_25; // @[LZA.scala 23:20]
  wire  p_27 = io_a[27] ^ io_b[27]; // @[LZA.scala 18:18]
  wire  k_27 = ~io_a[27] & ~io_b[27]; // @[LZA.scala 19:21]
  wire  f_27 = p_27 ^ ~k_26; // @[LZA.scala 23:20]
  wire  p_28 = io_a[28] ^ io_b[28]; // @[LZA.scala 18:18]
  wire  k_28 = ~io_a[28] & ~io_b[28]; // @[LZA.scala 19:21]
  wire  f_28 = p_28 ^ ~k_27; // @[LZA.scala 23:20]
  wire  p_29 = io_a[29] ^ io_b[29]; // @[LZA.scala 18:18]
  wire  k_29 = ~io_a[29] & ~io_b[29]; // @[LZA.scala 19:21]
  wire  f_29 = p_29 ^ ~k_28; // @[LZA.scala 23:20]
  wire  p_30 = io_a[30] ^ io_b[30]; // @[LZA.scala 18:18]
  wire  k_30 = ~io_a[30] & ~io_b[30]; // @[LZA.scala 19:21]
  wire  f_30 = p_30 ^ ~k_29; // @[LZA.scala 23:20]
  wire  p_31 = io_a[31] ^ io_b[31]; // @[LZA.scala 18:18]
  wire  k_31 = ~io_a[31] & ~io_b[31]; // @[LZA.scala 19:21]
  wire  f_31 = p_31 ^ ~k_30; // @[LZA.scala 23:20]
  wire  p_32 = io_a[32] ^ io_b[32]; // @[LZA.scala 18:18]
  wire  k_32 = ~io_a[32] & ~io_b[32]; // @[LZA.scala 19:21]
  wire  f_32 = p_32 ^ ~k_31; // @[LZA.scala 23:20]
  wire  p_33 = io_a[33] ^ io_b[33]; // @[LZA.scala 18:18]
  wire  k_33 = ~io_a[33] & ~io_b[33]; // @[LZA.scala 19:21]
  wire  f_33 = p_33 ^ ~k_32; // @[LZA.scala 23:20]
  wire  p_34 = io_a[34] ^ io_b[34]; // @[LZA.scala 18:18]
  wire  k_34 = ~io_a[34] & ~io_b[34]; // @[LZA.scala 19:21]
  wire  f_34 = p_34 ^ ~k_33; // @[LZA.scala 23:20]
  wire  p_35 = io_a[35] ^ io_b[35]; // @[LZA.scala 18:18]
  wire  k_35 = ~io_a[35] & ~io_b[35]; // @[LZA.scala 19:21]
  wire  f_35 = p_35 ^ ~k_34; // @[LZA.scala 23:20]
  wire  p_36 = io_a[36] ^ io_b[36]; // @[LZA.scala 18:18]
  wire  k_36 = ~io_a[36] & ~io_b[36]; // @[LZA.scala 19:21]
  wire  f_36 = p_36 ^ ~k_35; // @[LZA.scala 23:20]
  wire  p_37 = io_a[37] ^ io_b[37]; // @[LZA.scala 18:18]
  wire  k_37 = ~io_a[37] & ~io_b[37]; // @[LZA.scala 19:21]
  wire  f_37 = p_37 ^ ~k_36; // @[LZA.scala 23:20]
  wire  p_38 = io_a[38] ^ io_b[38]; // @[LZA.scala 18:18]
  wire  k_38 = ~io_a[38] & ~io_b[38]; // @[LZA.scala 19:21]
  wire  f_38 = p_38 ^ ~k_37; // @[LZA.scala 23:20]
  wire  p_39 = io_a[39] ^ io_b[39]; // @[LZA.scala 18:18]
  wire  k_39 = ~io_a[39] & ~io_b[39]; // @[LZA.scala 19:21]
  wire  f_39 = p_39 ^ ~k_38; // @[LZA.scala 23:20]
  wire  p_40 = io_a[40] ^ io_b[40]; // @[LZA.scala 18:18]
  wire  k_40 = ~io_a[40] & ~io_b[40]; // @[LZA.scala 19:21]
  wire  f_40 = p_40 ^ ~k_39; // @[LZA.scala 23:20]
  wire  p_41 = io_a[41] ^ io_b[41]; // @[LZA.scala 18:18]
  wire  k_41 = ~io_a[41] & ~io_b[41]; // @[LZA.scala 19:21]
  wire  f_41 = p_41 ^ ~k_40; // @[LZA.scala 23:20]
  wire  p_42 = io_a[42] ^ io_b[42]; // @[LZA.scala 18:18]
  wire  k_42 = ~io_a[42] & ~io_b[42]; // @[LZA.scala 19:21]
  wire  f_42 = p_42 ^ ~k_41; // @[LZA.scala 23:20]
  wire  p_43 = io_a[43] ^ io_b[43]; // @[LZA.scala 18:18]
  wire  k_43 = ~io_a[43] & ~io_b[43]; // @[LZA.scala 19:21]
  wire  f_43 = p_43 ^ ~k_42; // @[LZA.scala 23:20]
  wire  p_44 = io_a[44] ^ io_b[44]; // @[LZA.scala 18:18]
  wire  k_44 = ~io_a[44] & ~io_b[44]; // @[LZA.scala 19:21]
  wire  f_44 = p_44 ^ ~k_43; // @[LZA.scala 23:20]
  wire  p_45 = io_a[45] ^ io_b[45]; // @[LZA.scala 18:18]
  wire  k_45 = ~io_a[45] & ~io_b[45]; // @[LZA.scala 19:21]
  wire  f_45 = p_45 ^ ~k_44; // @[LZA.scala 23:20]
  wire  p_46 = io_a[46] ^ io_b[46]; // @[LZA.scala 18:18]
  wire  k_46 = ~io_a[46] & ~io_b[46]; // @[LZA.scala 19:21]
  wire  f_46 = p_46 ^ ~k_45; // @[LZA.scala 23:20]
  wire  p_47 = io_a[47] ^ io_b[47]; // @[LZA.scala 18:18]
  wire  k_47 = ~io_a[47] & ~io_b[47]; // @[LZA.scala 19:21]
  wire  f_47 = p_47 ^ ~k_46; // @[LZA.scala 23:20]
  wire  p_48 = io_a[48] ^ io_b[48]; // @[LZA.scala 18:18]
  wire  k_48 = ~io_a[48] & ~io_b[48]; // @[LZA.scala 19:21]
  wire  f_48 = p_48 ^ ~k_47; // @[LZA.scala 23:20]
  wire  p_49 = io_a[49] ^ io_b[49]; // @[LZA.scala 18:18]
  wire  k_49 = ~io_a[49] & ~io_b[49]; // @[LZA.scala 19:21]
  wire  f_49 = p_49 ^ ~k_48; // @[LZA.scala 23:20]
  wire  p_50 = io_a[50] ^ io_b[50]; // @[LZA.scala 18:18]
  wire  k_50 = ~io_a[50] & ~io_b[50]; // @[LZA.scala 19:21]
  wire  f_50 = p_50 ^ ~k_49; // @[LZA.scala 23:20]
  wire  p_51 = io_a[51] ^ io_b[51]; // @[LZA.scala 18:18]
  wire  k_51 = ~io_a[51] & ~io_b[51]; // @[LZA.scala 19:21]
  wire  f_51 = p_51 ^ ~k_50; // @[LZA.scala 23:20]
  wire  p_52 = io_a[52] ^ io_b[52]; // @[LZA.scala 18:18]
  wire  k_52 = ~io_a[52] & ~io_b[52]; // @[LZA.scala 19:21]
  wire  f_52 = p_52 ^ ~k_51; // @[LZA.scala 23:20]
  wire  p_53 = io_a[53] ^ io_b[53]; // @[LZA.scala 18:18]
  wire  k_53 = ~io_a[53] & ~io_b[53]; // @[LZA.scala 19:21]
  wire  f_53 = p_53 ^ ~k_52; // @[LZA.scala 23:20]
  wire  p_54 = io_a[54] ^ io_b[54]; // @[LZA.scala 18:18]
  wire  k_54 = ~io_a[54] & ~io_b[54]; // @[LZA.scala 19:21]
  wire  f_54 = p_54 ^ ~k_53; // @[LZA.scala 23:20]
  wire  p_55 = io_a[55] ^ io_b[55]; // @[LZA.scala 18:18]
  wire  k_55 = ~io_a[55] & ~io_b[55]; // @[LZA.scala 19:21]
  wire  f_55 = p_55 ^ ~k_54; // @[LZA.scala 23:20]
  wire  p_56 = io_a[56] ^ io_b[56]; // @[LZA.scala 18:18]
  wire  k_56 = ~io_a[56] & ~io_b[56]; // @[LZA.scala 19:21]
  wire  f_56 = p_56 ^ ~k_55; // @[LZA.scala 23:20]
  wire  p_57 = io_a[57] ^ io_b[57]; // @[LZA.scala 18:18]
  wire  k_57 = ~io_a[57] & ~io_b[57]; // @[LZA.scala 19:21]
  wire  f_57 = p_57 ^ ~k_56; // @[LZA.scala 23:20]
  wire  p_58 = io_a[58] ^ io_b[58]; // @[LZA.scala 18:18]
  wire  k_58 = ~io_a[58] & ~io_b[58]; // @[LZA.scala 19:21]
  wire  f_58 = p_58 ^ ~k_57; // @[LZA.scala 23:20]
  wire  p_59 = io_a[59] ^ io_b[59]; // @[LZA.scala 18:18]
  wire  k_59 = ~io_a[59] & ~io_b[59]; // @[LZA.scala 19:21]
  wire  f_59 = p_59 ^ ~k_58; // @[LZA.scala 23:20]
  wire  p_60 = io_a[60] ^ io_b[60]; // @[LZA.scala 18:18]
  wire  k_60 = ~io_a[60] & ~io_b[60]; // @[LZA.scala 19:21]
  wire  f_60 = p_60 ^ ~k_59; // @[LZA.scala 23:20]
  wire  p_61 = io_a[61] ^ io_b[61]; // @[LZA.scala 18:18]
  wire  k_61 = ~io_a[61] & ~io_b[61]; // @[LZA.scala 19:21]
  wire  f_61 = p_61 ^ ~k_60; // @[LZA.scala 23:20]
  wire  p_62 = io_a[62] ^ io_b[62]; // @[LZA.scala 18:18]
  wire  k_62 = ~io_a[62] & ~io_b[62]; // @[LZA.scala 19:21]
  wire  f_62 = p_62 ^ ~k_61; // @[LZA.scala 23:20]
  wire  p_63 = io_a[63] ^ io_b[63]; // @[LZA.scala 18:18]
  wire  k_63 = ~io_a[63] & ~io_b[63]; // @[LZA.scala 19:21]
  wire  f_63 = p_63 ^ ~k_62; // @[LZA.scala 23:20]
  wire  p_64 = io_a[64] ^ io_b[64]; // @[LZA.scala 18:18]
  wire  k_64 = ~io_a[64] & ~io_b[64]; // @[LZA.scala 19:21]
  wire  f_64 = p_64 ^ ~k_63; // @[LZA.scala 23:20]
  wire  p_65 = io_a[65] ^ io_b[65]; // @[LZA.scala 18:18]
  wire  k_65 = ~io_a[65] & ~io_b[65]; // @[LZA.scala 19:21]
  wire  f_65 = p_65 ^ ~k_64; // @[LZA.scala 23:20]
  wire  p_66 = io_a[66] ^ io_b[66]; // @[LZA.scala 18:18]
  wire  k_66 = ~io_a[66] & ~io_b[66]; // @[LZA.scala 19:21]
  wire  f_66 = p_66 ^ ~k_65; // @[LZA.scala 23:20]
  wire  p_67 = io_a[67] ^ io_b[67]; // @[LZA.scala 18:18]
  wire  k_67 = ~io_a[67] & ~io_b[67]; // @[LZA.scala 19:21]
  wire  f_67 = p_67 ^ ~k_66; // @[LZA.scala 23:20]
  wire  p_68 = io_a[68] ^ io_b[68]; // @[LZA.scala 18:18]
  wire  k_68 = ~io_a[68] & ~io_b[68]; // @[LZA.scala 19:21]
  wire  f_68 = p_68 ^ ~k_67; // @[LZA.scala 23:20]
  wire  p_69 = io_a[69] ^ io_b[69]; // @[LZA.scala 18:18]
  wire  k_69 = ~io_a[69] & ~io_b[69]; // @[LZA.scala 19:21]
  wire  f_69 = p_69 ^ ~k_68; // @[LZA.scala 23:20]
  wire  p_70 = io_a[70] ^ io_b[70]; // @[LZA.scala 18:18]
  wire  k_70 = ~io_a[70] & ~io_b[70]; // @[LZA.scala 19:21]
  wire  f_70 = p_70 ^ ~k_69; // @[LZA.scala 23:20]
  wire  p_71 = io_a[71] ^ io_b[71]; // @[LZA.scala 18:18]
  wire  k_71 = ~io_a[71] & ~io_b[71]; // @[LZA.scala 19:21]
  wire  f_71 = p_71 ^ ~k_70; // @[LZA.scala 23:20]
  wire  p_72 = io_a[72] ^ io_b[72]; // @[LZA.scala 18:18]
  wire  k_72 = ~io_a[72] & ~io_b[72]; // @[LZA.scala 19:21]
  wire  f_72 = p_72 ^ ~k_71; // @[LZA.scala 23:20]
  wire  p_73 = io_a[73] ^ io_b[73]; // @[LZA.scala 18:18]
  wire  k_73 = ~io_a[73] & ~io_b[73]; // @[LZA.scala 19:21]
  wire  f_73 = p_73 ^ ~k_72; // @[LZA.scala 23:20]
  wire  p_74 = io_a[74] ^ io_b[74]; // @[LZA.scala 18:18]
  wire  k_74 = ~io_a[74] & ~io_b[74]; // @[LZA.scala 19:21]
  wire  f_74 = p_74 ^ ~k_73; // @[LZA.scala 23:20]
  wire  p_75 = io_a[75] ^ io_b[75]; // @[LZA.scala 18:18]
  wire  k_75 = ~io_a[75] & ~io_b[75]; // @[LZA.scala 19:21]
  wire  f_75 = p_75 ^ ~k_74; // @[LZA.scala 23:20]
  wire  p_76 = io_a[76] ^ io_b[76]; // @[LZA.scala 18:18]
  wire  k_76 = ~io_a[76] & ~io_b[76]; // @[LZA.scala 19:21]
  wire  f_76 = p_76 ^ ~k_75; // @[LZA.scala 23:20]
  wire  p_77 = io_a[77] ^ io_b[77]; // @[LZA.scala 18:18]
  wire  k_77 = ~io_a[77] & ~io_b[77]; // @[LZA.scala 19:21]
  wire  f_77 = p_77 ^ ~k_76; // @[LZA.scala 23:20]
  wire  p_78 = io_a[78] ^ io_b[78]; // @[LZA.scala 18:18]
  wire  k_78 = ~io_a[78] & ~io_b[78]; // @[LZA.scala 19:21]
  wire  f_78 = p_78 ^ ~k_77; // @[LZA.scala 23:20]
  wire  p_79 = io_a[79] ^ io_b[79]; // @[LZA.scala 18:18]
  wire  k_79 = ~io_a[79] & ~io_b[79]; // @[LZA.scala 19:21]
  wire  f_79 = p_79 ^ ~k_78; // @[LZA.scala 23:20]
  wire  p_80 = io_a[80] ^ io_b[80]; // @[LZA.scala 18:18]
  wire  k_80 = ~io_a[80] & ~io_b[80]; // @[LZA.scala 19:21]
  wire  f_80 = p_80 ^ ~k_79; // @[LZA.scala 23:20]
  wire  p_81 = io_a[81] ^ io_b[81]; // @[LZA.scala 18:18]
  wire  k_81 = ~io_a[81] & ~io_b[81]; // @[LZA.scala 19:21]
  wire  f_81 = p_81 ^ ~k_80; // @[LZA.scala 23:20]
  wire  p_82 = io_a[82] ^ io_b[82]; // @[LZA.scala 18:18]
  wire  k_82 = ~io_a[82] & ~io_b[82]; // @[LZA.scala 19:21]
  wire  f_82 = p_82 ^ ~k_81; // @[LZA.scala 23:20]
  wire  p_83 = io_a[83] ^ io_b[83]; // @[LZA.scala 18:18]
  wire  k_83 = ~io_a[83] & ~io_b[83]; // @[LZA.scala 19:21]
  wire  f_83 = p_83 ^ ~k_82; // @[LZA.scala 23:20]
  wire  p_84 = io_a[84] ^ io_b[84]; // @[LZA.scala 18:18]
  wire  k_84 = ~io_a[84] & ~io_b[84]; // @[LZA.scala 19:21]
  wire  f_84 = p_84 ^ ~k_83; // @[LZA.scala 23:20]
  wire  p_85 = io_a[85] ^ io_b[85]; // @[LZA.scala 18:18]
  wire  k_85 = ~io_a[85] & ~io_b[85]; // @[LZA.scala 19:21]
  wire  f_85 = p_85 ^ ~k_84; // @[LZA.scala 23:20]
  wire  p_86 = io_a[86] ^ io_b[86]; // @[LZA.scala 18:18]
  wire  k_86 = ~io_a[86] & ~io_b[86]; // @[LZA.scala 19:21]
  wire  f_86 = p_86 ^ ~k_85; // @[LZA.scala 23:20]
  wire  p_87 = io_a[87] ^ io_b[87]; // @[LZA.scala 18:18]
  wire  k_87 = ~io_a[87] & ~io_b[87]; // @[LZA.scala 19:21]
  wire  f_87 = p_87 ^ ~k_86; // @[LZA.scala 23:20]
  wire  p_88 = io_a[88] ^ io_b[88]; // @[LZA.scala 18:18]
  wire  k_88 = ~io_a[88] & ~io_b[88]; // @[LZA.scala 19:21]
  wire  f_88 = p_88 ^ ~k_87; // @[LZA.scala 23:20]
  wire  p_89 = io_a[89] ^ io_b[89]; // @[LZA.scala 18:18]
  wire  k_89 = ~io_a[89] & ~io_b[89]; // @[LZA.scala 19:21]
  wire  f_89 = p_89 ^ ~k_88; // @[LZA.scala 23:20]
  wire  p_90 = io_a[90] ^ io_b[90]; // @[LZA.scala 18:18]
  wire  k_90 = ~io_a[90] & ~io_b[90]; // @[LZA.scala 19:21]
  wire  f_90 = p_90 ^ ~k_89; // @[LZA.scala 23:20]
  wire  p_91 = io_a[91] ^ io_b[91]; // @[LZA.scala 18:18]
  wire  k_91 = ~io_a[91] & ~io_b[91]; // @[LZA.scala 19:21]
  wire  f_91 = p_91 ^ ~k_90; // @[LZA.scala 23:20]
  wire  p_92 = io_a[92] ^ io_b[92]; // @[LZA.scala 18:18]
  wire  k_92 = ~io_a[92] & ~io_b[92]; // @[LZA.scala 19:21]
  wire  f_92 = p_92 ^ ~k_91; // @[LZA.scala 23:20]
  wire  p_93 = io_a[93] ^ io_b[93]; // @[LZA.scala 18:18]
  wire  k_93 = ~io_a[93] & ~io_b[93]; // @[LZA.scala 19:21]
  wire  f_93 = p_93 ^ ~k_92; // @[LZA.scala 23:20]
  wire  p_94 = io_a[94] ^ io_b[94]; // @[LZA.scala 18:18]
  wire  k_94 = ~io_a[94] & ~io_b[94]; // @[LZA.scala 19:21]
  wire  f_94 = p_94 ^ ~k_93; // @[LZA.scala 23:20]
  wire  p_95 = io_a[95] ^ io_b[95]; // @[LZA.scala 18:18]
  wire  k_95 = ~io_a[95] & ~io_b[95]; // @[LZA.scala 19:21]
  wire  f_95 = p_95 ^ ~k_94; // @[LZA.scala 23:20]
  wire  p_96 = io_a[96] ^ io_b[96]; // @[LZA.scala 18:18]
  wire  k_96 = ~io_a[96] & ~io_b[96]; // @[LZA.scala 19:21]
  wire  f_96 = p_96 ^ ~k_95; // @[LZA.scala 23:20]
  wire  p_97 = io_a[97] ^ io_b[97]; // @[LZA.scala 18:18]
  wire  k_97 = ~io_a[97] & ~io_b[97]; // @[LZA.scala 19:21]
  wire  f_97 = p_97 ^ ~k_96; // @[LZA.scala 23:20]
  wire  p_98 = io_a[98] ^ io_b[98]; // @[LZA.scala 18:18]
  wire  k_98 = ~io_a[98] & ~io_b[98]; // @[LZA.scala 19:21]
  wire  f_98 = p_98 ^ ~k_97; // @[LZA.scala 23:20]
  wire  p_99 = io_a[99] ^ io_b[99]; // @[LZA.scala 18:18]
  wire  k_99 = ~io_a[99] & ~io_b[99]; // @[LZA.scala 19:21]
  wire  f_99 = p_99 ^ ~k_98; // @[LZA.scala 23:20]
  wire  p_100 = io_a[100] ^ io_b[100]; // @[LZA.scala 18:18]
  wire  k_100 = ~io_a[100] & ~io_b[100]; // @[LZA.scala 19:21]
  wire  f_100 = p_100 ^ ~k_99; // @[LZA.scala 23:20]
  wire  p_101 = io_a[101] ^ io_b[101]; // @[LZA.scala 18:18]
  wire  k_101 = ~io_a[101] & ~io_b[101]; // @[LZA.scala 19:21]
  wire  f_101 = p_101 ^ ~k_100; // @[LZA.scala 23:20]
  wire  p_102 = io_a[102] ^ io_b[102]; // @[LZA.scala 18:18]
  wire  k_102 = ~io_a[102] & ~io_b[102]; // @[LZA.scala 19:21]
  wire  f_102 = p_102 ^ ~k_101; // @[LZA.scala 23:20]
  wire  p_103 = io_a[103] ^ io_b[103]; // @[LZA.scala 18:18]
  wire  k_103 = ~io_a[103] & ~io_b[103]; // @[LZA.scala 19:21]
  wire  f_103 = p_103 ^ ~k_102; // @[LZA.scala 23:20]
  wire  p_104 = io_a[104] ^ io_b[104]; // @[LZA.scala 18:18]
  wire  k_104 = ~io_a[104] & ~io_b[104]; // @[LZA.scala 19:21]
  wire  f_104 = p_104 ^ ~k_103; // @[LZA.scala 23:20]
  wire  p_105 = io_a[105] ^ io_b[105]; // @[LZA.scala 18:18]
  wire  k_105 = ~io_a[105] & ~io_b[105]; // @[LZA.scala 19:21]
  wire  f_105 = p_105 ^ ~k_104; // @[LZA.scala 23:20]
  wire  p_106 = io_a[106] ^ io_b[106]; // @[LZA.scala 18:18]
  wire  f_106 = p_106 ^ ~k_105; // @[LZA.scala 23:20]
  wire [5:0] io_f_lo_lo_lo_lo = {f_5,f_4,f_3,f_2,f_1,1'h0}; // @[Cat.scala 31:58]
  wire [12:0] io_f_lo_lo_lo = {f_12,f_11,f_10,f_9,f_8,f_7,f_6,io_f_lo_lo_lo_lo}; // @[Cat.scala 31:58]
  wire [5:0] io_f_lo_lo_hi_lo = {f_18,f_17,f_16,f_15,f_14,f_13}; // @[Cat.scala 31:58]
  wire [25:0] io_f_lo_lo = {f_25,f_24,f_23,f_22,f_21,f_20,f_19,io_f_lo_lo_hi_lo,io_f_lo_lo_lo}; // @[Cat.scala 31:58]
  wire [5:0] io_f_lo_hi_lo_lo = {f_31,f_30,f_29,f_28,f_27,f_26}; // @[Cat.scala 31:58]
  wire [12:0] io_f_lo_hi_lo = {f_38,f_37,f_36,f_35,f_34,f_33,f_32,io_f_lo_hi_lo_lo}; // @[Cat.scala 31:58]
  wire [6:0] io_f_lo_hi_hi_lo = {f_45,f_44,f_43,f_42,f_41,f_40,f_39}; // @[Cat.scala 31:58]
  wire [52:0] io_f_lo = {f_52,f_51,f_50,f_49,f_48,f_47,f_46,io_f_lo_hi_hi_lo,io_f_lo_hi_lo,io_f_lo_lo}; // @[Cat.scala 31:58]
  wire [5:0] io_f_hi_lo_lo_lo = {f_58,f_57,f_56,f_55,f_54,f_53}; // @[Cat.scala 31:58]
  wire [12:0] io_f_hi_lo_lo = {f_65,f_64,f_63,f_62,f_61,f_60,f_59,io_f_hi_lo_lo_lo}; // @[Cat.scala 31:58]
  wire [6:0] io_f_hi_lo_hi_lo = {f_72,f_71,f_70,f_69,f_68,f_67,f_66}; // @[Cat.scala 31:58]
  wire [26:0] io_f_hi_lo = {f_79,f_78,f_77,f_76,f_75,f_74,f_73,io_f_hi_lo_hi_lo,io_f_hi_lo_lo}; // @[Cat.scala 31:58]
  wire [5:0] io_f_hi_hi_lo_lo = {f_85,f_84,f_83,f_82,f_81,f_80}; // @[Cat.scala 31:58]
  wire [12:0] io_f_hi_hi_lo = {f_92,f_91,f_90,f_89,f_88,f_87,f_86,io_f_hi_hi_lo_lo}; // @[Cat.scala 31:58]
  wire [6:0] io_f_hi_hi_hi_lo = {f_99,f_98,f_97,f_96,f_95,f_94,f_93}; // @[Cat.scala 31:58]
  wire [53:0] io_f_hi = {f_106,f_105,f_104,f_103,f_102,f_101,f_100,io_f_hi_hi_hi_lo,io_f_hi_hi_lo,io_f_hi_lo}; // @[Cat.scala 31:58]
  assign io_f = {io_f_hi,io_f_lo}; // @[Cat.scala 31:58]
endmodule

