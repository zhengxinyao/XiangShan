module LazyModule(
  output  auto_source_out_0,
  output  auto_source_out_1,
  output  auto_source_out_2,
  output  auto_source_out_3,
  output  auto_source_out_4,
  output  auto_source_out_5,
  output  auto_source_out_6,
  output  auto_source_out_7,
  output  auto_source_out_8,
  output  auto_source_out_9,
  output  auto_source_out_10,
  output  auto_source_out_11,
  output  auto_source_out_12,
  output  auto_source_out_13,
  output  auto_source_out_14,
  output  auto_source_out_15,
  output  auto_source_out_16,
  output  auto_source_out_17,
  output  auto_source_out_18,
  output  auto_source_out_19,
  output  auto_source_out_20,
  output  auto_source_out_21,
  output  auto_source_out_22,
  output  auto_source_out_23,
  output  auto_source_out_24,
  output  auto_source_out_25,
  output  auto_source_out_26,
  output  auto_source_out_27,
  output  auto_source_out_28,
  output  auto_source_out_29,
  output  auto_source_out_30,
  output  auto_source_out_31,
  output  auto_source_out_32,
  output  auto_source_out_33,
  output  auto_source_out_34,
  output  auto_source_out_35,
  output  auto_source_out_36,
  output  auto_source_out_37,
  output  auto_source_out_38,
  output  auto_source_out_39,
  output  auto_source_out_40,
  output  auto_source_out_41,
  output  auto_source_out_42,
  output  auto_source_out_43,
  output  auto_source_out_44,
  output  auto_source_out_45,
  output  auto_source_out_46,
  output  auto_source_out_47,
  output  auto_source_out_48,
  output  auto_source_out_49,
  output  auto_source_out_50,
  output  auto_source_out_51,
  output  auto_source_out_52,
  output  auto_source_out_53,
  output  auto_source_out_54,
  output  auto_source_out_55,
  output  auto_source_out_56,
  output  auto_source_out_57,
  output  auto_source_out_58,
  output  auto_source_out_59,
  output  auto_source_out_60,
  output  auto_source_out_61,
  output  auto_source_out_62,
  output  auto_source_out_63,
  input   in_0,
  input   in_1,
  input   in_2,
  input   in_3,
  input   in_4,
  input   in_5,
  input   in_6,
  input   in_7,
  input   in_8,
  input   in_9,
  input   in_10,
  input   in_11,
  input   in_12,
  input   in_13,
  input   in_14,
  input   in_15,
  input   in_16,
  input   in_17,
  input   in_18,
  input   in_19,
  input   in_20,
  input   in_21,
  input   in_22,
  input   in_23,
  input   in_24,
  input   in_25,
  input   in_26,
  input   in_27,
  input   in_28,
  input   in_29,
  input   in_30,
  input   in_31,
  input   in_32,
  input   in_33,
  input   in_34,
  input   in_35,
  input   in_36,
  input   in_37,
  input   in_38,
  input   in_39,
  input   in_40,
  input   in_41,
  input   in_42,
  input   in_43,
  input   in_44,
  input   in_45,
  input   in_46,
  input   in_47,
  input   in_48,
  input   in_49,
  input   in_50,
  input   in_51,
  input   in_52,
  input   in_53,
  input   in_54,
  input   in_55,
  input   in_56,
  input   in_57,
  input   in_58,
  input   in_59,
  input   in_60,
  input   in_61,
  input   in_62,
  input   in_63
);
  assign auto_source_out_0 = in_0; // @[Nodes.scala 1207:84 SoC.scala 263:64]
  assign auto_source_out_1 = in_1; // @[Nodes.scala 1207:84 SoC.scala 263:64]
  assign auto_source_out_2 = in_2; // @[Nodes.scala 1207:84 SoC.scala 263:64]
  assign auto_source_out_3 = in_3; // @[Nodes.scala 1207:84 SoC.scala 263:64]
  assign auto_source_out_4 = in_4; // @[Nodes.scala 1207:84 SoC.scala 263:64]
  assign auto_source_out_5 = in_5; // @[Nodes.scala 1207:84 SoC.scala 263:64]
  assign auto_source_out_6 = in_6; // @[Nodes.scala 1207:84 SoC.scala 263:64]
  assign auto_source_out_7 = in_7; // @[Nodes.scala 1207:84 SoC.scala 263:64]
  assign auto_source_out_8 = in_8; // @[Nodes.scala 1207:84 SoC.scala 263:64]
  assign auto_source_out_9 = in_9; // @[Nodes.scala 1207:84 SoC.scala 263:64]
  assign auto_source_out_10 = in_10; // @[Nodes.scala 1207:84 SoC.scala 263:64]
  assign auto_source_out_11 = in_11; // @[Nodes.scala 1207:84 SoC.scala 263:64]
  assign auto_source_out_12 = in_12; // @[Nodes.scala 1207:84 SoC.scala 263:64]
  assign auto_source_out_13 = in_13; // @[Nodes.scala 1207:84 SoC.scala 263:64]
  assign auto_source_out_14 = in_14; // @[Nodes.scala 1207:84 SoC.scala 263:64]
  assign auto_source_out_15 = in_15; // @[Nodes.scala 1207:84 SoC.scala 263:64]
  assign auto_source_out_16 = in_16; // @[Nodes.scala 1207:84 SoC.scala 263:64]
  assign auto_source_out_17 = in_17; // @[Nodes.scala 1207:84 SoC.scala 263:64]
  assign auto_source_out_18 = in_18; // @[Nodes.scala 1207:84 SoC.scala 263:64]
  assign auto_source_out_19 = in_19; // @[Nodes.scala 1207:84 SoC.scala 263:64]
  assign auto_source_out_20 = in_20; // @[Nodes.scala 1207:84 SoC.scala 263:64]
  assign auto_source_out_21 = in_21; // @[Nodes.scala 1207:84 SoC.scala 263:64]
  assign auto_source_out_22 = in_22; // @[Nodes.scala 1207:84 SoC.scala 263:64]
  assign auto_source_out_23 = in_23; // @[Nodes.scala 1207:84 SoC.scala 263:64]
  assign auto_source_out_24 = in_24; // @[Nodes.scala 1207:84 SoC.scala 263:64]
  assign auto_source_out_25 = in_25; // @[Nodes.scala 1207:84 SoC.scala 263:64]
  assign auto_source_out_26 = in_26; // @[Nodes.scala 1207:84 SoC.scala 263:64]
  assign auto_source_out_27 = in_27; // @[Nodes.scala 1207:84 SoC.scala 263:64]
  assign auto_source_out_28 = in_28; // @[Nodes.scala 1207:84 SoC.scala 263:64]
  assign auto_source_out_29 = in_29; // @[Nodes.scala 1207:84 SoC.scala 263:64]
  assign auto_source_out_30 = in_30; // @[Nodes.scala 1207:84 SoC.scala 263:64]
  assign auto_source_out_31 = in_31; // @[Nodes.scala 1207:84 SoC.scala 263:64]
  assign auto_source_out_32 = in_32; // @[Nodes.scala 1207:84 SoC.scala 263:64]
  assign auto_source_out_33 = in_33; // @[Nodes.scala 1207:84 SoC.scala 263:64]
  assign auto_source_out_34 = in_34; // @[Nodes.scala 1207:84 SoC.scala 263:64]
  assign auto_source_out_35 = in_35; // @[Nodes.scala 1207:84 SoC.scala 263:64]
  assign auto_source_out_36 = in_36; // @[Nodes.scala 1207:84 SoC.scala 263:64]
  assign auto_source_out_37 = in_37; // @[Nodes.scala 1207:84 SoC.scala 263:64]
  assign auto_source_out_38 = in_38; // @[Nodes.scala 1207:84 SoC.scala 263:64]
  assign auto_source_out_39 = in_39; // @[Nodes.scala 1207:84 SoC.scala 263:64]
  assign auto_source_out_40 = in_40; // @[Nodes.scala 1207:84 SoC.scala 263:64]
  assign auto_source_out_41 = in_41; // @[Nodes.scala 1207:84 SoC.scala 263:64]
  assign auto_source_out_42 = in_42; // @[Nodes.scala 1207:84 SoC.scala 263:64]
  assign auto_source_out_43 = in_43; // @[Nodes.scala 1207:84 SoC.scala 263:64]
  assign auto_source_out_44 = in_44; // @[Nodes.scala 1207:84 SoC.scala 263:64]
  assign auto_source_out_45 = in_45; // @[Nodes.scala 1207:84 SoC.scala 263:64]
  assign auto_source_out_46 = in_46; // @[Nodes.scala 1207:84 SoC.scala 263:64]
  assign auto_source_out_47 = in_47; // @[Nodes.scala 1207:84 SoC.scala 263:64]
  assign auto_source_out_48 = in_48; // @[Nodes.scala 1207:84 SoC.scala 263:64]
  assign auto_source_out_49 = in_49; // @[Nodes.scala 1207:84 SoC.scala 263:64]
  assign auto_source_out_50 = in_50; // @[Nodes.scala 1207:84 SoC.scala 263:64]
  assign auto_source_out_51 = in_51; // @[Nodes.scala 1207:84 SoC.scala 263:64]
  assign auto_source_out_52 = in_52; // @[Nodes.scala 1207:84 SoC.scala 263:64]
  assign auto_source_out_53 = in_53; // @[Nodes.scala 1207:84 SoC.scala 263:64]
  assign auto_source_out_54 = in_54; // @[Nodes.scala 1207:84 SoC.scala 263:64]
  assign auto_source_out_55 = in_55; // @[Nodes.scala 1207:84 SoC.scala 263:64]
  assign auto_source_out_56 = in_56; // @[Nodes.scala 1207:84 SoC.scala 263:64]
  assign auto_source_out_57 = in_57; // @[Nodes.scala 1207:84 SoC.scala 263:64]
  assign auto_source_out_58 = in_58; // @[Nodes.scala 1207:84 SoC.scala 263:64]
  assign auto_source_out_59 = in_59; // @[Nodes.scala 1207:84 SoC.scala 263:64]
  assign auto_source_out_60 = in_60; // @[Nodes.scala 1207:84 SoC.scala 263:64]
  assign auto_source_out_61 = in_61; // @[Nodes.scala 1207:84 SoC.scala 263:64]
  assign auto_source_out_62 = in_62; // @[Nodes.scala 1207:84 SoC.scala 263:64]
  assign auto_source_out_63 = in_63; // @[Nodes.scala 1207:84 SoC.scala 263:64]
endmodule

