module Multiplier(
  input          clock,
  input  [53:0]  io_a,
  input  [53:0]  io_b,
  input          io_regEnables_0,
  output [107:0] io_result
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
`endif // RANDOMIZE_REG_INIT
  wire  c22_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_1_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_1_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_1_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_1_io_out_1; // @[Multiplier.scala 73:25]
  wire  c32_io_in_0; // @[Multiplier.scala 78:25]
  wire  c32_io_in_1; // @[Multiplier.scala 78:25]
  wire  c32_io_in_2; // @[Multiplier.scala 78:25]
  wire  c32_io_out_0; // @[Multiplier.scala 78:25]
  wire  c32_io_out_1; // @[Multiplier.scala 78:25]
  wire  c32_1_io_in_0; // @[Multiplier.scala 78:25]
  wire  c32_1_io_in_1; // @[Multiplier.scala 78:25]
  wire  c32_1_io_in_2; // @[Multiplier.scala 78:25]
  wire  c32_1_io_out_0; // @[Multiplier.scala 78:25]
  wire  c32_1_io_out_1; // @[Multiplier.scala 78:25]
  wire  c53_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_1_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_1_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_1_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_1_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_1_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_1_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_1_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_1_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_2_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_2_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_2_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_2_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_2_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_2_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_2_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_2_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_3_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_3_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_3_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_3_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_3_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_3_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_3_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_3_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_4_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_4_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_4_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_4_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_4_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_4_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_4_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_4_io_out_2; // @[Multiplier.scala 83:25]
  wire  c22_2_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_2_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_2_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_2_io_out_1; // @[Multiplier.scala 73:25]
  wire  c53_5_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_5_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_5_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_5_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_5_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_5_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_5_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_5_io_out_2; // @[Multiplier.scala 83:25]
  wire  c22_3_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_3_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_3_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_3_io_out_1; // @[Multiplier.scala 73:25]
  wire  c53_6_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_6_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_6_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_6_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_6_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_6_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_6_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_6_io_out_2; // @[Multiplier.scala 83:25]
  wire  c32_2_io_in_0; // @[Multiplier.scala 78:25]
  wire  c32_2_io_in_1; // @[Multiplier.scala 78:25]
  wire  c32_2_io_in_2; // @[Multiplier.scala 78:25]
  wire  c32_2_io_out_0; // @[Multiplier.scala 78:25]
  wire  c32_2_io_out_1; // @[Multiplier.scala 78:25]
  wire  c53_7_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_7_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_7_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_7_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_7_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_7_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_7_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_7_io_out_2; // @[Multiplier.scala 83:25]
  wire  c32_3_io_in_0; // @[Multiplier.scala 78:25]
  wire  c32_3_io_in_1; // @[Multiplier.scala 78:25]
  wire  c32_3_io_in_2; // @[Multiplier.scala 78:25]
  wire  c32_3_io_out_0; // @[Multiplier.scala 78:25]
  wire  c32_3_io_out_1; // @[Multiplier.scala 78:25]
  wire  c53_8_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_8_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_8_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_8_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_8_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_8_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_8_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_8_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_9_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_9_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_9_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_9_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_9_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_9_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_9_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_9_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_10_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_10_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_10_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_10_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_10_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_10_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_10_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_10_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_11_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_11_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_11_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_11_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_11_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_11_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_11_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_11_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_12_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_12_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_12_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_12_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_12_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_12_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_12_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_12_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_13_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_13_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_13_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_13_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_13_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_13_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_13_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_13_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_14_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_14_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_14_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_14_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_14_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_14_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_14_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_14_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_15_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_15_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_15_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_15_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_15_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_15_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_15_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_15_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_16_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_16_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_16_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_16_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_16_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_16_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_16_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_16_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_17_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_17_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_17_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_17_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_17_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_17_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_17_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_17_io_out_2; // @[Multiplier.scala 83:25]
  wire  c22_4_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_4_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_4_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_4_io_out_1; // @[Multiplier.scala 73:25]
  wire  c53_18_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_18_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_18_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_18_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_18_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_18_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_18_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_18_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_19_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_19_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_19_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_19_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_19_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_19_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_19_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_19_io_out_2; // @[Multiplier.scala 83:25]
  wire  c22_5_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_5_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_5_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_5_io_out_1; // @[Multiplier.scala 73:25]
  wire  c53_20_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_20_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_20_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_20_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_20_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_20_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_20_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_20_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_21_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_21_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_21_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_21_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_21_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_21_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_21_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_21_io_out_2; // @[Multiplier.scala 83:25]
  wire  c32_4_io_in_0; // @[Multiplier.scala 78:25]
  wire  c32_4_io_in_1; // @[Multiplier.scala 78:25]
  wire  c32_4_io_in_2; // @[Multiplier.scala 78:25]
  wire  c32_4_io_out_0; // @[Multiplier.scala 78:25]
  wire  c32_4_io_out_1; // @[Multiplier.scala 78:25]
  wire  c53_22_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_22_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_22_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_22_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_22_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_22_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_22_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_22_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_23_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_23_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_23_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_23_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_23_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_23_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_23_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_23_io_out_2; // @[Multiplier.scala 83:25]
  wire  c32_5_io_in_0; // @[Multiplier.scala 78:25]
  wire  c32_5_io_in_1; // @[Multiplier.scala 78:25]
  wire  c32_5_io_in_2; // @[Multiplier.scala 78:25]
  wire  c32_5_io_out_0; // @[Multiplier.scala 78:25]
  wire  c32_5_io_out_1; // @[Multiplier.scala 78:25]
  wire  c53_24_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_24_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_24_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_24_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_24_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_24_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_24_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_24_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_25_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_25_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_25_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_25_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_25_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_25_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_25_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_25_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_26_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_26_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_26_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_26_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_26_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_26_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_26_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_26_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_27_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_27_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_27_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_27_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_27_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_27_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_27_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_27_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_28_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_28_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_28_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_28_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_28_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_28_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_28_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_28_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_29_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_29_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_29_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_29_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_29_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_29_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_29_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_29_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_30_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_30_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_30_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_30_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_30_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_30_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_30_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_30_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_31_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_31_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_31_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_31_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_31_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_31_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_31_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_31_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_32_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_32_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_32_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_32_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_32_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_32_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_32_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_32_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_33_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_33_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_33_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_33_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_33_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_33_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_33_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_33_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_34_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_34_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_34_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_34_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_34_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_34_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_34_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_34_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_35_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_35_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_35_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_35_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_35_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_35_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_35_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_35_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_36_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_36_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_36_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_36_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_36_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_36_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_36_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_36_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_37_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_37_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_37_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_37_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_37_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_37_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_37_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_37_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_38_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_38_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_38_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_38_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_38_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_38_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_38_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_38_io_out_2; // @[Multiplier.scala 83:25]
  wire  c22_6_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_6_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_6_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_6_io_out_1; // @[Multiplier.scala 73:25]
  wire  c53_39_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_39_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_39_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_39_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_39_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_39_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_39_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_39_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_40_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_40_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_40_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_40_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_40_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_40_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_40_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_40_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_41_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_41_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_41_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_41_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_41_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_41_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_41_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_41_io_out_2; // @[Multiplier.scala 83:25]
  wire  c22_7_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_7_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_7_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_7_io_out_1; // @[Multiplier.scala 73:25]
  wire  c53_42_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_42_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_42_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_42_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_42_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_42_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_42_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_42_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_43_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_43_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_43_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_43_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_43_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_43_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_43_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_43_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_44_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_44_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_44_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_44_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_44_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_44_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_44_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_44_io_out_2; // @[Multiplier.scala 83:25]
  wire  c32_6_io_in_0; // @[Multiplier.scala 78:25]
  wire  c32_6_io_in_1; // @[Multiplier.scala 78:25]
  wire  c32_6_io_in_2; // @[Multiplier.scala 78:25]
  wire  c32_6_io_out_0; // @[Multiplier.scala 78:25]
  wire  c32_6_io_out_1; // @[Multiplier.scala 78:25]
  wire  c53_45_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_45_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_45_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_45_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_45_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_45_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_45_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_45_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_46_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_46_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_46_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_46_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_46_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_46_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_46_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_46_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_47_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_47_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_47_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_47_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_47_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_47_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_47_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_47_io_out_2; // @[Multiplier.scala 83:25]
  wire  c32_7_io_in_0; // @[Multiplier.scala 78:25]
  wire  c32_7_io_in_1; // @[Multiplier.scala 78:25]
  wire  c32_7_io_in_2; // @[Multiplier.scala 78:25]
  wire  c32_7_io_out_0; // @[Multiplier.scala 78:25]
  wire  c32_7_io_out_1; // @[Multiplier.scala 78:25]
  wire  c53_48_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_48_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_48_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_48_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_48_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_48_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_48_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_48_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_49_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_49_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_49_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_49_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_49_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_49_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_49_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_49_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_50_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_50_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_50_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_50_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_50_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_50_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_50_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_50_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_51_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_51_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_51_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_51_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_51_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_51_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_51_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_51_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_52_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_52_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_52_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_52_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_52_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_52_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_52_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_52_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_53_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_53_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_53_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_53_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_53_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_53_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_53_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_53_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_54_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_54_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_54_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_54_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_54_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_54_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_54_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_54_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_55_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_55_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_55_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_55_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_55_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_55_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_55_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_55_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_56_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_56_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_56_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_56_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_56_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_56_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_56_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_56_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_57_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_57_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_57_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_57_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_57_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_57_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_57_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_57_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_58_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_58_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_58_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_58_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_58_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_58_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_58_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_58_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_59_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_59_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_59_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_59_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_59_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_59_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_59_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_59_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_60_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_60_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_60_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_60_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_60_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_60_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_60_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_60_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_61_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_61_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_61_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_61_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_61_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_61_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_61_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_61_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_62_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_62_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_62_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_62_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_62_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_62_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_62_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_62_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_63_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_63_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_63_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_63_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_63_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_63_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_63_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_63_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_64_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_64_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_64_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_64_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_64_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_64_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_64_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_64_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_65_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_65_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_65_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_65_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_65_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_65_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_65_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_65_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_66_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_66_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_66_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_66_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_66_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_66_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_66_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_66_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_67_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_67_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_67_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_67_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_67_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_67_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_67_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_67_io_out_2; // @[Multiplier.scala 83:25]
  wire  c22_8_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_8_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_8_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_8_io_out_1; // @[Multiplier.scala 73:25]
  wire  c53_68_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_68_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_68_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_68_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_68_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_68_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_68_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_68_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_69_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_69_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_69_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_69_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_69_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_69_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_69_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_69_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_70_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_70_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_70_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_70_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_70_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_70_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_70_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_70_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_71_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_71_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_71_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_71_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_71_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_71_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_71_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_71_io_out_2; // @[Multiplier.scala 83:25]
  wire  c22_9_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_9_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_9_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_9_io_out_1; // @[Multiplier.scala 73:25]
  wire  c53_72_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_72_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_72_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_72_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_72_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_72_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_72_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_72_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_73_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_73_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_73_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_73_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_73_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_73_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_73_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_73_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_74_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_74_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_74_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_74_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_74_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_74_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_74_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_74_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_75_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_75_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_75_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_75_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_75_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_75_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_75_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_75_io_out_2; // @[Multiplier.scala 83:25]
  wire  c32_8_io_in_0; // @[Multiplier.scala 78:25]
  wire  c32_8_io_in_1; // @[Multiplier.scala 78:25]
  wire  c32_8_io_in_2; // @[Multiplier.scala 78:25]
  wire  c32_8_io_out_0; // @[Multiplier.scala 78:25]
  wire  c32_8_io_out_1; // @[Multiplier.scala 78:25]
  wire  c53_76_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_76_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_76_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_76_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_76_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_76_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_76_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_76_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_77_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_77_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_77_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_77_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_77_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_77_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_77_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_77_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_78_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_78_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_78_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_78_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_78_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_78_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_78_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_78_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_79_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_79_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_79_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_79_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_79_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_79_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_79_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_79_io_out_2; // @[Multiplier.scala 83:25]
  wire  c32_9_io_in_0; // @[Multiplier.scala 78:25]
  wire  c32_9_io_in_1; // @[Multiplier.scala 78:25]
  wire  c32_9_io_in_2; // @[Multiplier.scala 78:25]
  wire  c32_9_io_out_0; // @[Multiplier.scala 78:25]
  wire  c32_9_io_out_1; // @[Multiplier.scala 78:25]
  wire  c53_80_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_80_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_80_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_80_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_80_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_80_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_80_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_80_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_81_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_81_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_81_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_81_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_81_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_81_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_81_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_81_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_82_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_82_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_82_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_82_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_82_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_82_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_82_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_82_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_83_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_83_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_83_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_83_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_83_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_83_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_83_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_83_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_84_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_84_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_84_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_84_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_84_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_84_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_84_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_84_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_85_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_85_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_85_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_85_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_85_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_85_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_85_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_85_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_86_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_86_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_86_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_86_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_86_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_86_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_86_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_86_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_87_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_87_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_87_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_87_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_87_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_87_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_87_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_87_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_88_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_88_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_88_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_88_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_88_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_88_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_88_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_88_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_89_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_89_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_89_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_89_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_89_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_89_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_89_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_89_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_90_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_90_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_90_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_90_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_90_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_90_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_90_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_90_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_91_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_91_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_91_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_91_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_91_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_91_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_91_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_91_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_92_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_92_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_92_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_92_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_92_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_92_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_92_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_92_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_93_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_93_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_93_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_93_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_93_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_93_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_93_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_93_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_94_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_94_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_94_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_94_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_94_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_94_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_94_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_94_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_95_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_95_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_95_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_95_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_95_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_95_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_95_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_95_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_96_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_96_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_96_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_96_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_96_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_96_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_96_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_96_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_97_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_97_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_97_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_97_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_97_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_97_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_97_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_97_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_98_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_98_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_98_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_98_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_98_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_98_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_98_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_98_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_99_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_99_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_99_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_99_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_99_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_99_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_99_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_99_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_100_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_100_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_100_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_100_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_100_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_100_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_100_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_100_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_101_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_101_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_101_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_101_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_101_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_101_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_101_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_101_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_102_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_102_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_102_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_102_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_102_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_102_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_102_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_102_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_103_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_103_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_103_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_103_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_103_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_103_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_103_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_103_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_104_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_104_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_104_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_104_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_104_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_104_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_104_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_104_io_out_2; // @[Multiplier.scala 83:25]
  wire  c22_10_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_10_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_10_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_10_io_out_1; // @[Multiplier.scala 73:25]
  wire  c53_105_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_105_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_105_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_105_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_105_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_105_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_105_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_105_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_106_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_106_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_106_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_106_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_106_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_106_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_106_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_106_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_107_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_107_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_107_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_107_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_107_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_107_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_107_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_107_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_108_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_108_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_108_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_108_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_108_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_108_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_108_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_108_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_109_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_109_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_109_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_109_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_109_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_109_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_109_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_109_io_out_2; // @[Multiplier.scala 83:25]
  wire  c22_11_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_11_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_11_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_11_io_out_1; // @[Multiplier.scala 73:25]
  wire  c53_110_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_110_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_110_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_110_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_110_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_110_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_110_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_110_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_111_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_111_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_111_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_111_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_111_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_111_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_111_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_111_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_112_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_112_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_112_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_112_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_112_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_112_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_112_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_112_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_113_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_113_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_113_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_113_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_113_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_113_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_113_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_113_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_114_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_114_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_114_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_114_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_114_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_114_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_114_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_114_io_out_2; // @[Multiplier.scala 83:25]
  wire  c32_10_io_in_0; // @[Multiplier.scala 78:25]
  wire  c32_10_io_in_1; // @[Multiplier.scala 78:25]
  wire  c32_10_io_in_2; // @[Multiplier.scala 78:25]
  wire  c32_10_io_out_0; // @[Multiplier.scala 78:25]
  wire  c32_10_io_out_1; // @[Multiplier.scala 78:25]
  wire  c53_115_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_115_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_115_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_115_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_115_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_115_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_115_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_115_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_116_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_116_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_116_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_116_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_116_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_116_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_116_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_116_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_117_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_117_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_117_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_117_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_117_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_117_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_117_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_117_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_118_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_118_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_118_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_118_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_118_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_118_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_118_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_118_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_119_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_119_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_119_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_119_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_119_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_119_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_119_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_119_io_out_2; // @[Multiplier.scala 83:25]
  wire  c32_11_io_in_0; // @[Multiplier.scala 78:25]
  wire  c32_11_io_in_1; // @[Multiplier.scala 78:25]
  wire  c32_11_io_in_2; // @[Multiplier.scala 78:25]
  wire  c32_11_io_out_0; // @[Multiplier.scala 78:25]
  wire  c32_11_io_out_1; // @[Multiplier.scala 78:25]
  wire  c53_120_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_120_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_120_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_120_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_120_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_120_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_120_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_120_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_121_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_121_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_121_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_121_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_121_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_121_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_121_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_121_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_122_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_122_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_122_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_122_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_122_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_122_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_122_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_122_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_123_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_123_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_123_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_123_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_123_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_123_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_123_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_123_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_124_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_124_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_124_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_124_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_124_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_124_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_124_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_124_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_125_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_125_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_125_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_125_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_125_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_125_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_125_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_125_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_126_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_126_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_126_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_126_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_126_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_126_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_126_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_126_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_127_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_127_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_127_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_127_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_127_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_127_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_127_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_127_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_128_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_128_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_128_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_128_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_128_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_128_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_128_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_128_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_129_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_129_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_129_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_129_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_129_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_129_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_129_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_129_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_130_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_130_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_130_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_130_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_130_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_130_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_130_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_130_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_131_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_131_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_131_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_131_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_131_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_131_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_131_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_131_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_132_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_132_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_132_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_132_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_132_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_132_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_132_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_132_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_133_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_133_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_133_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_133_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_133_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_133_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_133_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_133_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_134_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_134_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_134_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_134_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_134_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_134_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_134_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_134_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_135_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_135_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_135_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_135_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_135_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_135_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_135_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_135_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_136_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_136_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_136_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_136_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_136_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_136_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_136_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_136_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_137_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_137_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_137_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_137_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_137_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_137_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_137_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_137_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_138_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_138_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_138_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_138_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_138_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_138_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_138_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_138_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_139_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_139_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_139_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_139_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_139_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_139_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_139_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_139_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_140_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_140_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_140_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_140_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_140_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_140_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_140_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_140_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_141_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_141_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_141_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_141_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_141_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_141_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_141_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_141_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_142_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_142_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_142_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_142_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_142_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_142_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_142_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_142_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_143_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_143_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_143_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_143_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_143_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_143_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_143_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_143_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_144_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_144_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_144_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_144_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_144_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_144_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_144_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_144_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_145_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_145_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_145_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_145_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_145_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_145_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_145_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_145_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_146_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_146_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_146_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_146_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_146_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_146_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_146_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_146_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_147_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_147_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_147_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_147_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_147_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_147_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_147_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_147_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_148_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_148_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_148_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_148_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_148_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_148_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_148_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_148_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_149_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_149_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_149_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_149_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_149_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_149_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_149_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_149_io_out_2; // @[Multiplier.scala 83:25]
  wire  c22_12_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_12_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_12_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_12_io_out_1; // @[Multiplier.scala 73:25]
  wire  c53_150_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_150_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_150_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_150_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_150_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_150_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_150_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_150_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_151_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_151_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_151_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_151_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_151_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_151_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_151_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_151_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_152_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_152_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_152_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_152_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_152_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_152_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_152_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_152_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_153_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_153_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_153_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_153_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_153_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_153_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_153_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_153_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_154_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_154_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_154_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_154_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_154_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_154_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_154_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_154_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_155_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_155_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_155_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_155_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_155_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_155_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_155_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_155_io_out_2; // @[Multiplier.scala 83:25]
  wire  c22_13_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_13_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_13_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_13_io_out_1; // @[Multiplier.scala 73:25]
  wire  c53_156_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_156_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_156_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_156_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_156_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_156_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_156_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_156_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_157_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_157_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_157_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_157_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_157_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_157_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_157_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_157_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_158_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_158_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_158_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_158_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_158_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_158_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_158_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_158_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_159_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_159_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_159_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_159_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_159_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_159_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_159_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_159_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_160_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_160_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_160_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_160_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_160_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_160_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_160_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_160_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_161_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_161_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_161_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_161_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_161_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_161_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_161_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_161_io_out_2; // @[Multiplier.scala 83:25]
  wire  c32_12_io_in_0; // @[Multiplier.scala 78:25]
  wire  c32_12_io_in_1; // @[Multiplier.scala 78:25]
  wire  c32_12_io_in_2; // @[Multiplier.scala 78:25]
  wire  c32_12_io_out_0; // @[Multiplier.scala 78:25]
  wire  c32_12_io_out_1; // @[Multiplier.scala 78:25]
  wire  c53_162_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_162_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_162_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_162_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_162_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_162_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_162_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_162_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_163_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_163_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_163_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_163_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_163_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_163_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_163_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_163_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_164_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_164_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_164_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_164_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_164_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_164_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_164_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_164_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_165_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_165_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_165_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_165_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_165_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_165_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_165_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_165_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_166_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_166_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_166_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_166_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_166_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_166_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_166_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_166_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_167_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_167_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_167_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_167_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_167_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_167_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_167_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_167_io_out_2; // @[Multiplier.scala 83:25]
  wire  c32_13_io_in_0; // @[Multiplier.scala 78:25]
  wire  c32_13_io_in_1; // @[Multiplier.scala 78:25]
  wire  c32_13_io_in_2; // @[Multiplier.scala 78:25]
  wire  c32_13_io_out_0; // @[Multiplier.scala 78:25]
  wire  c32_13_io_out_1; // @[Multiplier.scala 78:25]
  wire  c53_168_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_168_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_168_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_168_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_168_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_168_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_168_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_168_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_169_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_169_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_169_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_169_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_169_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_169_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_169_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_169_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_170_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_170_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_170_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_170_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_170_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_170_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_170_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_170_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_171_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_171_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_171_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_171_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_171_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_171_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_171_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_171_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_172_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_172_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_172_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_172_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_172_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_172_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_172_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_172_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_173_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_173_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_173_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_173_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_173_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_173_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_173_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_173_io_out_2; // @[Multiplier.scala 83:25]
  wire  c32_14_io_in_0; // @[Multiplier.scala 78:25]
  wire  c32_14_io_in_1; // @[Multiplier.scala 78:25]
  wire  c32_14_io_in_2; // @[Multiplier.scala 78:25]
  wire  c32_14_io_out_0; // @[Multiplier.scala 78:25]
  wire  c32_14_io_out_1; // @[Multiplier.scala 78:25]
  wire  c53_174_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_174_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_174_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_174_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_174_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_174_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_174_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_174_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_175_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_175_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_175_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_175_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_175_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_175_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_175_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_175_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_176_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_176_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_176_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_176_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_176_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_176_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_176_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_176_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_177_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_177_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_177_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_177_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_177_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_177_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_177_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_177_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_178_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_178_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_178_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_178_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_178_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_178_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_178_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_178_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_179_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_179_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_179_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_179_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_179_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_179_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_179_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_179_io_out_2; // @[Multiplier.scala 83:25]
  wire  c32_15_io_in_0; // @[Multiplier.scala 78:25]
  wire  c32_15_io_in_1; // @[Multiplier.scala 78:25]
  wire  c32_15_io_in_2; // @[Multiplier.scala 78:25]
  wire  c32_15_io_out_0; // @[Multiplier.scala 78:25]
  wire  c32_15_io_out_1; // @[Multiplier.scala 78:25]
  wire  c53_180_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_180_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_180_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_180_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_180_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_180_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_180_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_180_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_181_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_181_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_181_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_181_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_181_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_181_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_181_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_181_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_182_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_182_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_182_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_182_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_182_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_182_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_182_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_182_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_183_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_183_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_183_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_183_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_183_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_183_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_183_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_183_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_184_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_184_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_184_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_184_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_184_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_184_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_184_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_184_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_185_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_185_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_185_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_185_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_185_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_185_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_185_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_185_io_out_2; // @[Multiplier.scala 83:25]
  wire  c32_16_io_in_0; // @[Multiplier.scala 78:25]
  wire  c32_16_io_in_1; // @[Multiplier.scala 78:25]
  wire  c32_16_io_in_2; // @[Multiplier.scala 78:25]
  wire  c32_16_io_out_0; // @[Multiplier.scala 78:25]
  wire  c32_16_io_out_1; // @[Multiplier.scala 78:25]
  wire  c53_186_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_186_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_186_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_186_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_186_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_186_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_186_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_186_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_187_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_187_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_187_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_187_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_187_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_187_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_187_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_187_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_188_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_188_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_188_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_188_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_188_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_188_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_188_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_188_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_189_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_189_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_189_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_189_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_189_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_189_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_189_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_189_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_190_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_190_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_190_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_190_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_190_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_190_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_190_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_190_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_191_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_191_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_191_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_191_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_191_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_191_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_191_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_191_io_out_2; // @[Multiplier.scala 83:25]
  wire  c32_17_io_in_0; // @[Multiplier.scala 78:25]
  wire  c32_17_io_in_1; // @[Multiplier.scala 78:25]
  wire  c32_17_io_in_2; // @[Multiplier.scala 78:25]
  wire  c32_17_io_out_0; // @[Multiplier.scala 78:25]
  wire  c32_17_io_out_1; // @[Multiplier.scala 78:25]
  wire  c53_192_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_192_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_192_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_192_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_192_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_192_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_192_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_192_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_193_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_193_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_193_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_193_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_193_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_193_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_193_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_193_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_194_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_194_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_194_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_194_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_194_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_194_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_194_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_194_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_195_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_195_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_195_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_195_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_195_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_195_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_195_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_195_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_196_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_196_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_196_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_196_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_196_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_196_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_196_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_196_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_197_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_197_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_197_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_197_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_197_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_197_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_197_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_197_io_out_2; // @[Multiplier.scala 83:25]
  wire  c32_18_io_in_0; // @[Multiplier.scala 78:25]
  wire  c32_18_io_in_1; // @[Multiplier.scala 78:25]
  wire  c32_18_io_in_2; // @[Multiplier.scala 78:25]
  wire  c32_18_io_out_0; // @[Multiplier.scala 78:25]
  wire  c32_18_io_out_1; // @[Multiplier.scala 78:25]
  wire  c53_198_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_198_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_198_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_198_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_198_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_198_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_198_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_198_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_199_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_199_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_199_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_199_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_199_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_199_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_199_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_199_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_200_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_200_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_200_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_200_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_200_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_200_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_200_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_200_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_201_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_201_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_201_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_201_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_201_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_201_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_201_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_201_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_202_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_202_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_202_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_202_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_202_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_202_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_202_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_202_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_203_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_203_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_203_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_203_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_203_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_203_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_203_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_203_io_out_2; // @[Multiplier.scala 83:25]
  wire  c32_19_io_in_0; // @[Multiplier.scala 78:25]
  wire  c32_19_io_in_1; // @[Multiplier.scala 78:25]
  wire  c32_19_io_in_2; // @[Multiplier.scala 78:25]
  wire  c32_19_io_out_0; // @[Multiplier.scala 78:25]
  wire  c32_19_io_out_1; // @[Multiplier.scala 78:25]
  wire  c53_204_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_204_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_204_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_204_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_204_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_204_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_204_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_204_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_205_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_205_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_205_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_205_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_205_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_205_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_205_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_205_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_206_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_206_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_206_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_206_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_206_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_206_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_206_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_206_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_207_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_207_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_207_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_207_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_207_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_207_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_207_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_207_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_208_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_208_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_208_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_208_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_208_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_208_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_208_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_208_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_209_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_209_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_209_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_209_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_209_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_209_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_209_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_209_io_out_2; // @[Multiplier.scala 83:25]
  wire  c22_14_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_14_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_14_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_14_io_out_1; // @[Multiplier.scala 73:25]
  wire  c53_210_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_210_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_210_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_210_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_210_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_210_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_210_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_210_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_211_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_211_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_211_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_211_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_211_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_211_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_211_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_211_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_212_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_212_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_212_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_212_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_212_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_212_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_212_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_212_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_213_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_213_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_213_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_213_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_213_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_213_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_213_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_213_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_214_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_214_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_214_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_214_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_214_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_214_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_214_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_214_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_215_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_215_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_215_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_215_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_215_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_215_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_215_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_215_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_216_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_216_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_216_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_216_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_216_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_216_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_216_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_216_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_217_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_217_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_217_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_217_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_217_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_217_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_217_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_217_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_218_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_218_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_218_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_218_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_218_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_218_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_218_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_218_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_219_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_219_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_219_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_219_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_219_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_219_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_219_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_219_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_220_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_220_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_220_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_220_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_220_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_220_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_220_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_220_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_221_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_221_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_221_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_221_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_221_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_221_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_221_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_221_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_222_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_222_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_222_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_222_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_222_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_222_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_222_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_222_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_223_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_223_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_223_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_223_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_223_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_223_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_223_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_223_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_224_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_224_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_224_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_224_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_224_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_224_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_224_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_224_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_225_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_225_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_225_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_225_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_225_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_225_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_225_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_225_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_226_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_226_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_226_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_226_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_226_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_226_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_226_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_226_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_227_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_227_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_227_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_227_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_227_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_227_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_227_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_227_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_228_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_228_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_228_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_228_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_228_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_228_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_228_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_228_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_229_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_229_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_229_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_229_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_229_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_229_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_229_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_229_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_230_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_230_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_230_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_230_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_230_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_230_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_230_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_230_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_231_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_231_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_231_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_231_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_231_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_231_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_231_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_231_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_232_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_232_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_232_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_232_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_232_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_232_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_232_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_232_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_233_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_233_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_233_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_233_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_233_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_233_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_233_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_233_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_234_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_234_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_234_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_234_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_234_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_234_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_234_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_234_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_235_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_235_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_235_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_235_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_235_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_235_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_235_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_235_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_236_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_236_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_236_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_236_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_236_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_236_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_236_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_236_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_237_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_237_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_237_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_237_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_237_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_237_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_237_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_237_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_238_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_238_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_238_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_238_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_238_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_238_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_238_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_238_io_out_2; // @[Multiplier.scala 83:25]
  wire  c32_20_io_in_0; // @[Multiplier.scala 78:25]
  wire  c32_20_io_in_1; // @[Multiplier.scala 78:25]
  wire  c32_20_io_in_2; // @[Multiplier.scala 78:25]
  wire  c32_20_io_out_0; // @[Multiplier.scala 78:25]
  wire  c32_20_io_out_1; // @[Multiplier.scala 78:25]
  wire  c53_239_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_239_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_239_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_239_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_239_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_239_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_239_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_239_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_240_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_240_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_240_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_240_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_240_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_240_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_240_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_240_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_241_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_241_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_241_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_241_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_241_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_241_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_241_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_241_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_242_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_242_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_242_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_242_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_242_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_242_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_242_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_242_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_243_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_243_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_243_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_243_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_243_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_243_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_243_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_243_io_out_2; // @[Multiplier.scala 83:25]
  wire  c32_21_io_in_0; // @[Multiplier.scala 78:25]
  wire  c32_21_io_in_1; // @[Multiplier.scala 78:25]
  wire  c32_21_io_in_2; // @[Multiplier.scala 78:25]
  wire  c32_21_io_out_0; // @[Multiplier.scala 78:25]
  wire  c32_21_io_out_1; // @[Multiplier.scala 78:25]
  wire  c53_244_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_244_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_244_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_244_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_244_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_244_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_244_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_244_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_245_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_245_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_245_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_245_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_245_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_245_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_245_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_245_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_246_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_246_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_246_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_246_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_246_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_246_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_246_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_246_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_247_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_247_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_247_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_247_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_247_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_247_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_247_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_247_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_248_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_248_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_248_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_248_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_248_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_248_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_248_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_248_io_out_2; // @[Multiplier.scala 83:25]
  wire  c22_15_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_15_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_15_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_15_io_out_1; // @[Multiplier.scala 73:25]
  wire  c53_249_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_249_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_249_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_249_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_249_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_249_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_249_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_249_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_250_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_250_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_250_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_250_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_250_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_250_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_250_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_250_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_251_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_251_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_251_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_251_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_251_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_251_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_251_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_251_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_252_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_252_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_252_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_252_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_252_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_252_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_252_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_252_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_253_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_253_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_253_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_253_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_253_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_253_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_253_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_253_io_out_2; // @[Multiplier.scala 83:25]
  wire  c22_16_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_16_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_16_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_16_io_out_1; // @[Multiplier.scala 73:25]
  wire  c53_254_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_254_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_254_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_254_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_254_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_254_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_254_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_254_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_255_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_255_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_255_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_255_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_255_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_255_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_255_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_255_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_256_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_256_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_256_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_256_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_256_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_256_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_256_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_256_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_257_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_257_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_257_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_257_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_257_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_257_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_257_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_257_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_258_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_258_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_258_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_258_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_258_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_258_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_258_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_258_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_259_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_259_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_259_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_259_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_259_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_259_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_259_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_259_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_260_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_260_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_260_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_260_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_260_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_260_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_260_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_260_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_261_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_261_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_261_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_261_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_261_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_261_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_261_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_261_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_262_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_262_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_262_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_262_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_262_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_262_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_262_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_262_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_263_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_263_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_263_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_263_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_263_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_263_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_263_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_263_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_264_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_264_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_264_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_264_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_264_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_264_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_264_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_264_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_265_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_265_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_265_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_265_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_265_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_265_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_265_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_265_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_266_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_266_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_266_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_266_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_266_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_266_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_266_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_266_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_267_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_267_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_267_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_267_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_267_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_267_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_267_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_267_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_268_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_268_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_268_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_268_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_268_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_268_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_268_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_268_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_269_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_269_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_269_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_269_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_269_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_269_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_269_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_269_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_270_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_270_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_270_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_270_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_270_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_270_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_270_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_270_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_271_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_271_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_271_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_271_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_271_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_271_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_271_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_271_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_272_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_272_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_272_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_272_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_272_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_272_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_272_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_272_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_273_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_273_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_273_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_273_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_273_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_273_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_273_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_273_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_274_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_274_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_274_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_274_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_274_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_274_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_274_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_274_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_275_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_275_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_275_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_275_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_275_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_275_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_275_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_275_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_276_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_276_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_276_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_276_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_276_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_276_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_276_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_276_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_277_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_277_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_277_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_277_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_277_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_277_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_277_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_277_io_out_2; // @[Multiplier.scala 83:25]
  wire  c32_22_io_in_0; // @[Multiplier.scala 78:25]
  wire  c32_22_io_in_1; // @[Multiplier.scala 78:25]
  wire  c32_22_io_in_2; // @[Multiplier.scala 78:25]
  wire  c32_22_io_out_0; // @[Multiplier.scala 78:25]
  wire  c32_22_io_out_1; // @[Multiplier.scala 78:25]
  wire  c53_278_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_278_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_278_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_278_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_278_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_278_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_278_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_278_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_279_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_279_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_279_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_279_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_279_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_279_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_279_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_279_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_280_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_280_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_280_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_280_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_280_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_280_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_280_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_280_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_281_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_281_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_281_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_281_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_281_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_281_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_281_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_281_io_out_2; // @[Multiplier.scala 83:25]
  wire  c32_23_io_in_0; // @[Multiplier.scala 78:25]
  wire  c32_23_io_in_1; // @[Multiplier.scala 78:25]
  wire  c32_23_io_in_2; // @[Multiplier.scala 78:25]
  wire  c32_23_io_out_0; // @[Multiplier.scala 78:25]
  wire  c32_23_io_out_1; // @[Multiplier.scala 78:25]
  wire  c53_282_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_282_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_282_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_282_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_282_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_282_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_282_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_282_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_283_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_283_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_283_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_283_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_283_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_283_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_283_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_283_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_284_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_284_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_284_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_284_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_284_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_284_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_284_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_284_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_285_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_285_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_285_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_285_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_285_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_285_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_285_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_285_io_out_2; // @[Multiplier.scala 83:25]
  wire  c22_17_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_17_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_17_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_17_io_out_1; // @[Multiplier.scala 73:25]
  wire  c53_286_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_286_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_286_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_286_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_286_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_286_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_286_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_286_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_287_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_287_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_287_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_287_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_287_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_287_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_287_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_287_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_288_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_288_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_288_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_288_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_288_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_288_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_288_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_288_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_289_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_289_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_289_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_289_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_289_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_289_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_289_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_289_io_out_2; // @[Multiplier.scala 83:25]
  wire  c22_18_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_18_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_18_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_18_io_out_1; // @[Multiplier.scala 73:25]
  wire  c53_290_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_290_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_290_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_290_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_290_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_290_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_290_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_290_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_291_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_291_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_291_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_291_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_291_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_291_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_291_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_291_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_292_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_292_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_292_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_292_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_292_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_292_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_292_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_292_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_293_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_293_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_293_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_293_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_293_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_293_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_293_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_293_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_294_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_294_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_294_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_294_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_294_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_294_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_294_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_294_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_295_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_295_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_295_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_295_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_295_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_295_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_295_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_295_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_296_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_296_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_296_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_296_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_296_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_296_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_296_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_296_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_297_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_297_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_297_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_297_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_297_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_297_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_297_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_297_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_298_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_298_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_298_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_298_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_298_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_298_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_298_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_298_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_299_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_299_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_299_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_299_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_299_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_299_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_299_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_299_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_300_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_300_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_300_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_300_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_300_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_300_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_300_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_300_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_301_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_301_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_301_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_301_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_301_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_301_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_301_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_301_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_302_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_302_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_302_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_302_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_302_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_302_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_302_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_302_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_303_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_303_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_303_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_303_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_303_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_303_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_303_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_303_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_304_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_304_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_304_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_304_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_304_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_304_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_304_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_304_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_305_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_305_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_305_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_305_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_305_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_305_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_305_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_305_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_306_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_306_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_306_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_306_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_306_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_306_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_306_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_306_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_307_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_307_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_307_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_307_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_307_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_307_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_307_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_307_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_308_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_308_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_308_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_308_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_308_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_308_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_308_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_308_io_out_2; // @[Multiplier.scala 83:25]
  wire  c32_24_io_in_0; // @[Multiplier.scala 78:25]
  wire  c32_24_io_in_1; // @[Multiplier.scala 78:25]
  wire  c32_24_io_in_2; // @[Multiplier.scala 78:25]
  wire  c32_24_io_out_0; // @[Multiplier.scala 78:25]
  wire  c32_24_io_out_1; // @[Multiplier.scala 78:25]
  wire  c53_309_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_309_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_309_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_309_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_309_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_309_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_309_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_309_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_310_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_310_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_310_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_310_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_310_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_310_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_310_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_310_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_311_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_311_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_311_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_311_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_311_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_311_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_311_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_311_io_out_2; // @[Multiplier.scala 83:25]
  wire  c32_25_io_in_0; // @[Multiplier.scala 78:25]
  wire  c32_25_io_in_1; // @[Multiplier.scala 78:25]
  wire  c32_25_io_in_2; // @[Multiplier.scala 78:25]
  wire  c32_25_io_out_0; // @[Multiplier.scala 78:25]
  wire  c32_25_io_out_1; // @[Multiplier.scala 78:25]
  wire  c53_312_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_312_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_312_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_312_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_312_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_312_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_312_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_312_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_313_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_313_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_313_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_313_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_313_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_313_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_313_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_313_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_314_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_314_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_314_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_314_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_314_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_314_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_314_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_314_io_out_2; // @[Multiplier.scala 83:25]
  wire  c22_19_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_19_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_19_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_19_io_out_1; // @[Multiplier.scala 73:25]
  wire  c53_315_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_315_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_315_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_315_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_315_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_315_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_315_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_315_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_316_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_316_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_316_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_316_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_316_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_316_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_316_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_316_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_317_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_317_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_317_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_317_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_317_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_317_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_317_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_317_io_out_2; // @[Multiplier.scala 83:25]
  wire  c22_20_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_20_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_20_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_20_io_out_1; // @[Multiplier.scala 73:25]
  wire  c53_318_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_318_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_318_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_318_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_318_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_318_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_318_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_318_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_319_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_319_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_319_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_319_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_319_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_319_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_319_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_319_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_320_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_320_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_320_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_320_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_320_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_320_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_320_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_320_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_321_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_321_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_321_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_321_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_321_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_321_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_321_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_321_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_322_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_322_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_322_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_322_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_322_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_322_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_322_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_322_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_323_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_323_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_323_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_323_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_323_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_323_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_323_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_323_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_324_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_324_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_324_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_324_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_324_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_324_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_324_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_324_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_325_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_325_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_325_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_325_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_325_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_325_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_325_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_325_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_326_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_326_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_326_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_326_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_326_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_326_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_326_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_326_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_327_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_327_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_327_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_327_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_327_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_327_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_327_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_327_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_328_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_328_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_328_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_328_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_328_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_328_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_328_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_328_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_329_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_329_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_329_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_329_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_329_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_329_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_329_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_329_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_330_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_330_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_330_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_330_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_330_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_330_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_330_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_330_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_331_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_331_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_331_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_331_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_331_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_331_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_331_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_331_io_out_2; // @[Multiplier.scala 83:25]
  wire  c32_26_io_in_0; // @[Multiplier.scala 78:25]
  wire  c32_26_io_in_1; // @[Multiplier.scala 78:25]
  wire  c32_26_io_in_2; // @[Multiplier.scala 78:25]
  wire  c32_26_io_out_0; // @[Multiplier.scala 78:25]
  wire  c32_26_io_out_1; // @[Multiplier.scala 78:25]
  wire  c53_332_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_332_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_332_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_332_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_332_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_332_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_332_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_332_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_333_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_333_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_333_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_333_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_333_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_333_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_333_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_333_io_out_2; // @[Multiplier.scala 83:25]
  wire  c32_27_io_in_0; // @[Multiplier.scala 78:25]
  wire  c32_27_io_in_1; // @[Multiplier.scala 78:25]
  wire  c32_27_io_in_2; // @[Multiplier.scala 78:25]
  wire  c32_27_io_out_0; // @[Multiplier.scala 78:25]
  wire  c32_27_io_out_1; // @[Multiplier.scala 78:25]
  wire  c53_334_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_334_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_334_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_334_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_334_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_334_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_334_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_334_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_335_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_335_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_335_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_335_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_335_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_335_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_335_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_335_io_out_2; // @[Multiplier.scala 83:25]
  wire  c22_21_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_21_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_21_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_21_io_out_1; // @[Multiplier.scala 73:25]
  wire  c53_336_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_336_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_336_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_336_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_336_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_336_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_336_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_336_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_337_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_337_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_337_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_337_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_337_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_337_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_337_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_337_io_out_2; // @[Multiplier.scala 83:25]
  wire  c22_22_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_22_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_22_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_22_io_out_1; // @[Multiplier.scala 73:25]
  wire  c53_338_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_338_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_338_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_338_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_338_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_338_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_338_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_338_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_339_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_339_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_339_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_339_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_339_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_339_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_339_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_339_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_340_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_340_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_340_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_340_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_340_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_340_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_340_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_340_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_341_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_341_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_341_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_341_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_341_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_341_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_341_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_341_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_342_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_342_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_342_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_342_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_342_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_342_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_342_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_342_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_343_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_343_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_343_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_343_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_343_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_343_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_343_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_343_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_344_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_344_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_344_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_344_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_344_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_344_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_344_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_344_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_345_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_345_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_345_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_345_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_345_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_345_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_345_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_345_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_346_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_346_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_346_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_346_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_346_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_346_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_346_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_346_io_out_2; // @[Multiplier.scala 83:25]
  wire  c32_28_io_in_0; // @[Multiplier.scala 78:25]
  wire  c32_28_io_in_1; // @[Multiplier.scala 78:25]
  wire  c32_28_io_in_2; // @[Multiplier.scala 78:25]
  wire  c32_28_io_out_0; // @[Multiplier.scala 78:25]
  wire  c32_28_io_out_1; // @[Multiplier.scala 78:25]
  wire  c53_347_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_347_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_347_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_347_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_347_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_347_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_347_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_347_io_out_2; // @[Multiplier.scala 83:25]
  wire  c32_29_io_in_0; // @[Multiplier.scala 78:25]
  wire  c32_29_io_in_1; // @[Multiplier.scala 78:25]
  wire  c32_29_io_in_2; // @[Multiplier.scala 78:25]
  wire  c32_29_io_out_0; // @[Multiplier.scala 78:25]
  wire  c32_29_io_out_1; // @[Multiplier.scala 78:25]
  wire  c53_348_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_348_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_348_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_348_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_348_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_348_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_348_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_348_io_out_2; // @[Multiplier.scala 83:25]
  wire  c22_23_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_23_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_23_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_23_io_out_1; // @[Multiplier.scala 73:25]
  wire  c53_349_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_349_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_349_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_349_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_349_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_349_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_349_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_349_io_out_2; // @[Multiplier.scala 83:25]
  wire  c22_24_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_24_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_24_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_24_io_out_1; // @[Multiplier.scala 73:25]
  wire  c53_350_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_350_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_350_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_350_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_350_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_350_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_350_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_350_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_351_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_351_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_351_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_351_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_351_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_351_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_351_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_351_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_352_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_352_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_352_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_352_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_352_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_352_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_352_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_352_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_353_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_353_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_353_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_353_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_353_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_353_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_353_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_353_io_out_2; // @[Multiplier.scala 83:25]
  wire  c32_30_io_in_0; // @[Multiplier.scala 78:25]
  wire  c32_30_io_in_1; // @[Multiplier.scala 78:25]
  wire  c32_30_io_in_2; // @[Multiplier.scala 78:25]
  wire  c32_30_io_out_0; // @[Multiplier.scala 78:25]
  wire  c32_30_io_out_1; // @[Multiplier.scala 78:25]
  wire  c32_31_io_in_0; // @[Multiplier.scala 78:25]
  wire  c32_31_io_in_1; // @[Multiplier.scala 78:25]
  wire  c32_31_io_in_2; // @[Multiplier.scala 78:25]
  wire  c32_31_io_out_0; // @[Multiplier.scala 78:25]
  wire  c32_31_io_out_1; // @[Multiplier.scala 78:25]
  wire  c22_25_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_25_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_25_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_25_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_26_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_26_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_26_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_26_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_27_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_27_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_27_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_27_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_28_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_28_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_28_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_28_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_29_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_29_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_29_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_29_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_30_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_30_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_30_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_30_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_31_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_31_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_31_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_31_io_out_1; // @[Multiplier.scala 73:25]
  wire  c32_32_io_in_0; // @[Multiplier.scala 78:25]
  wire  c32_32_io_in_1; // @[Multiplier.scala 78:25]
  wire  c32_32_io_in_2; // @[Multiplier.scala 78:25]
  wire  c32_32_io_out_0; // @[Multiplier.scala 78:25]
  wire  c32_32_io_out_1; // @[Multiplier.scala 78:25]
  wire  c32_33_io_in_0; // @[Multiplier.scala 78:25]
  wire  c32_33_io_in_1; // @[Multiplier.scala 78:25]
  wire  c32_33_io_in_2; // @[Multiplier.scala 78:25]
  wire  c32_33_io_out_0; // @[Multiplier.scala 78:25]
  wire  c32_33_io_out_1; // @[Multiplier.scala 78:25]
  wire  c32_34_io_in_0; // @[Multiplier.scala 78:25]
  wire  c32_34_io_in_1; // @[Multiplier.scala 78:25]
  wire  c32_34_io_in_2; // @[Multiplier.scala 78:25]
  wire  c32_34_io_out_0; // @[Multiplier.scala 78:25]
  wire  c32_34_io_out_1; // @[Multiplier.scala 78:25]
  wire  c53_354_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_354_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_354_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_354_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_354_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_354_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_354_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_354_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_355_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_355_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_355_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_355_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_355_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_355_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_355_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_355_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_356_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_356_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_356_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_356_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_356_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_356_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_356_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_356_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_357_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_357_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_357_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_357_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_357_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_357_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_357_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_357_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_358_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_358_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_358_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_358_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_358_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_358_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_358_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_358_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_359_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_359_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_359_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_359_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_359_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_359_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_359_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_359_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_360_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_360_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_360_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_360_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_360_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_360_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_360_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_360_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_361_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_361_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_361_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_361_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_361_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_361_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_361_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_361_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_362_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_362_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_362_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_362_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_362_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_362_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_362_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_362_io_out_2; // @[Multiplier.scala 83:25]
  wire  c22_32_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_32_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_32_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_32_io_out_1; // @[Multiplier.scala 73:25]
  wire  c53_363_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_363_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_363_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_363_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_363_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_363_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_363_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_363_io_out_2; // @[Multiplier.scala 83:25]
  wire  c22_33_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_33_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_33_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_33_io_out_1; // @[Multiplier.scala 73:25]
  wire  c53_364_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_364_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_364_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_364_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_364_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_364_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_364_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_364_io_out_2; // @[Multiplier.scala 83:25]
  wire  c22_34_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_34_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_34_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_34_io_out_1; // @[Multiplier.scala 73:25]
  wire  c53_365_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_365_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_365_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_365_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_365_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_365_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_365_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_365_io_out_2; // @[Multiplier.scala 83:25]
  wire  c22_35_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_35_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_35_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_35_io_out_1; // @[Multiplier.scala 73:25]
  wire  c53_366_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_366_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_366_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_366_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_366_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_366_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_366_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_366_io_out_2; // @[Multiplier.scala 83:25]
  wire  c22_36_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_36_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_36_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_36_io_out_1; // @[Multiplier.scala 73:25]
  wire  c53_367_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_367_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_367_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_367_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_367_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_367_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_367_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_367_io_out_2; // @[Multiplier.scala 83:25]
  wire  c32_35_io_in_0; // @[Multiplier.scala 78:25]
  wire  c32_35_io_in_1; // @[Multiplier.scala 78:25]
  wire  c32_35_io_in_2; // @[Multiplier.scala 78:25]
  wire  c32_35_io_out_0; // @[Multiplier.scala 78:25]
  wire  c32_35_io_out_1; // @[Multiplier.scala 78:25]
  wire  c53_368_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_368_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_368_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_368_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_368_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_368_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_368_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_368_io_out_2; // @[Multiplier.scala 83:25]
  wire  c32_36_io_in_0; // @[Multiplier.scala 78:25]
  wire  c32_36_io_in_1; // @[Multiplier.scala 78:25]
  wire  c32_36_io_in_2; // @[Multiplier.scala 78:25]
  wire  c32_36_io_out_0; // @[Multiplier.scala 78:25]
  wire  c32_36_io_out_1; // @[Multiplier.scala 78:25]
  wire  c53_369_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_369_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_369_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_369_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_369_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_369_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_369_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_369_io_out_2; // @[Multiplier.scala 83:25]
  wire  c32_37_io_in_0; // @[Multiplier.scala 78:25]
  wire  c32_37_io_in_1; // @[Multiplier.scala 78:25]
  wire  c32_37_io_in_2; // @[Multiplier.scala 78:25]
  wire  c32_37_io_out_0; // @[Multiplier.scala 78:25]
  wire  c32_37_io_out_1; // @[Multiplier.scala 78:25]
  wire  c53_370_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_370_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_370_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_370_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_370_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_370_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_370_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_370_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_371_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_371_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_371_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_371_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_371_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_371_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_371_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_371_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_372_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_372_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_372_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_372_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_372_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_372_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_372_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_372_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_373_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_373_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_373_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_373_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_373_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_373_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_373_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_373_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_374_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_374_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_374_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_374_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_374_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_374_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_374_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_374_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_375_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_375_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_375_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_375_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_375_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_375_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_375_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_375_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_376_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_376_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_376_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_376_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_376_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_376_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_376_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_376_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_377_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_377_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_377_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_377_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_377_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_377_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_377_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_377_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_378_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_378_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_378_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_378_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_378_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_378_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_378_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_378_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_379_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_379_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_379_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_379_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_379_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_379_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_379_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_379_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_380_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_380_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_380_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_380_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_380_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_380_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_380_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_380_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_381_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_381_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_381_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_381_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_381_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_381_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_381_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_381_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_382_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_382_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_382_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_382_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_382_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_382_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_382_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_382_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_383_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_383_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_383_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_383_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_383_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_383_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_383_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_383_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_384_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_384_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_384_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_384_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_384_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_384_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_384_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_384_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_385_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_385_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_385_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_385_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_385_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_385_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_385_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_385_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_386_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_386_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_386_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_386_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_386_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_386_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_386_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_386_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_387_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_387_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_387_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_387_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_387_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_387_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_387_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_387_io_out_2; // @[Multiplier.scala 83:25]
  wire  c22_37_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_37_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_37_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_37_io_out_1; // @[Multiplier.scala 73:25]
  wire  c53_388_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_388_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_388_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_388_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_388_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_388_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_388_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_388_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_389_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_389_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_389_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_389_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_389_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_389_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_389_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_389_io_out_2; // @[Multiplier.scala 83:25]
  wire  c22_38_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_38_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_38_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_38_io_out_1; // @[Multiplier.scala 73:25]
  wire  c53_390_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_390_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_390_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_390_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_390_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_390_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_390_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_390_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_391_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_391_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_391_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_391_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_391_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_391_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_391_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_391_io_out_2; // @[Multiplier.scala 83:25]
  wire  c22_39_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_39_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_39_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_39_io_out_1; // @[Multiplier.scala 73:25]
  wire  c53_392_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_392_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_392_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_392_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_392_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_392_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_392_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_392_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_393_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_393_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_393_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_393_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_393_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_393_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_393_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_393_io_out_2; // @[Multiplier.scala 83:25]
  wire  c22_40_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_40_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_40_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_40_io_out_1; // @[Multiplier.scala 73:25]
  wire  c53_394_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_394_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_394_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_394_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_394_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_394_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_394_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_394_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_395_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_395_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_395_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_395_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_395_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_395_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_395_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_395_io_out_2; // @[Multiplier.scala 83:25]
  wire  c22_41_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_41_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_41_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_41_io_out_1; // @[Multiplier.scala 73:25]
  wire  c53_396_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_396_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_396_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_396_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_396_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_396_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_396_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_396_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_397_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_397_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_397_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_397_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_397_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_397_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_397_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_397_io_out_2; // @[Multiplier.scala 83:25]
  wire  c32_38_io_in_0; // @[Multiplier.scala 78:25]
  wire  c32_38_io_in_1; // @[Multiplier.scala 78:25]
  wire  c32_38_io_in_2; // @[Multiplier.scala 78:25]
  wire  c32_38_io_out_0; // @[Multiplier.scala 78:25]
  wire  c32_38_io_out_1; // @[Multiplier.scala 78:25]
  wire  c53_398_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_398_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_398_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_398_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_398_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_398_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_398_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_398_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_399_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_399_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_399_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_399_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_399_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_399_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_399_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_399_io_out_2; // @[Multiplier.scala 83:25]
  wire  c32_39_io_in_0; // @[Multiplier.scala 78:25]
  wire  c32_39_io_in_1; // @[Multiplier.scala 78:25]
  wire  c32_39_io_in_2; // @[Multiplier.scala 78:25]
  wire  c32_39_io_out_0; // @[Multiplier.scala 78:25]
  wire  c32_39_io_out_1; // @[Multiplier.scala 78:25]
  wire  c53_400_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_400_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_400_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_400_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_400_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_400_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_400_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_400_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_401_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_401_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_401_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_401_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_401_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_401_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_401_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_401_io_out_2; // @[Multiplier.scala 83:25]
  wire  c32_40_io_in_0; // @[Multiplier.scala 78:25]
  wire  c32_40_io_in_1; // @[Multiplier.scala 78:25]
  wire  c32_40_io_in_2; // @[Multiplier.scala 78:25]
  wire  c32_40_io_out_0; // @[Multiplier.scala 78:25]
  wire  c32_40_io_out_1; // @[Multiplier.scala 78:25]
  wire  c53_402_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_402_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_402_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_402_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_402_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_402_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_402_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_402_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_403_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_403_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_403_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_403_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_403_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_403_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_403_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_403_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_404_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_404_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_404_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_404_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_404_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_404_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_404_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_404_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_405_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_405_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_405_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_405_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_405_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_405_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_405_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_405_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_406_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_406_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_406_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_406_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_406_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_406_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_406_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_406_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_407_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_407_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_407_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_407_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_407_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_407_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_407_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_407_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_408_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_408_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_408_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_408_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_408_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_408_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_408_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_408_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_409_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_409_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_409_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_409_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_409_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_409_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_409_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_409_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_410_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_410_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_410_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_410_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_410_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_410_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_410_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_410_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_411_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_411_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_411_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_411_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_411_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_411_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_411_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_411_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_412_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_412_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_412_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_412_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_412_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_412_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_412_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_412_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_413_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_413_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_413_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_413_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_413_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_413_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_413_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_413_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_414_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_414_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_414_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_414_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_414_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_414_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_414_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_414_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_415_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_415_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_415_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_415_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_415_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_415_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_415_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_415_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_416_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_416_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_416_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_416_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_416_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_416_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_416_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_416_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_417_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_417_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_417_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_417_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_417_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_417_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_417_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_417_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_418_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_418_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_418_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_418_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_418_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_418_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_418_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_418_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_419_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_419_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_419_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_419_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_419_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_419_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_419_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_419_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_420_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_420_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_420_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_420_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_420_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_420_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_420_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_420_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_421_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_421_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_421_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_421_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_421_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_421_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_421_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_421_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_422_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_422_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_422_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_422_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_422_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_422_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_422_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_422_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_423_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_423_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_423_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_423_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_423_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_423_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_423_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_423_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_424_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_424_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_424_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_424_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_424_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_424_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_424_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_424_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_425_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_425_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_425_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_425_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_425_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_425_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_425_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_425_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_426_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_426_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_426_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_426_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_426_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_426_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_426_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_426_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_427_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_427_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_427_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_427_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_427_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_427_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_427_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_427_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_428_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_428_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_428_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_428_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_428_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_428_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_428_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_428_io_out_2; // @[Multiplier.scala 83:25]
  wire  c22_42_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_42_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_42_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_42_io_out_1; // @[Multiplier.scala 73:25]
  wire  c53_429_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_429_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_429_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_429_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_429_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_429_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_429_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_429_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_430_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_430_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_430_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_430_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_430_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_430_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_430_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_430_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_431_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_431_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_431_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_431_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_431_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_431_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_431_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_431_io_out_2; // @[Multiplier.scala 83:25]
  wire  c22_43_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_43_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_43_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_43_io_out_1; // @[Multiplier.scala 73:25]
  wire  c53_432_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_432_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_432_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_432_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_432_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_432_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_432_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_432_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_433_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_433_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_433_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_433_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_433_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_433_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_433_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_433_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_434_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_434_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_434_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_434_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_434_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_434_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_434_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_434_io_out_2; // @[Multiplier.scala 83:25]
  wire  c22_44_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_44_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_44_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_44_io_out_1; // @[Multiplier.scala 73:25]
  wire  c53_435_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_435_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_435_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_435_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_435_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_435_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_435_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_435_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_436_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_436_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_436_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_436_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_436_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_436_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_436_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_436_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_437_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_437_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_437_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_437_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_437_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_437_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_437_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_437_io_out_2; // @[Multiplier.scala 83:25]
  wire  c22_45_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_45_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_45_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_45_io_out_1; // @[Multiplier.scala 73:25]
  wire  c53_438_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_438_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_438_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_438_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_438_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_438_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_438_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_438_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_439_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_439_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_439_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_439_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_439_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_439_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_439_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_439_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_440_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_440_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_440_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_440_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_440_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_440_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_440_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_440_io_out_2; // @[Multiplier.scala 83:25]
  wire  c22_46_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_46_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_46_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_46_io_out_1; // @[Multiplier.scala 73:25]
  wire  c53_441_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_441_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_441_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_441_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_441_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_441_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_441_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_441_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_442_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_442_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_442_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_442_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_442_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_442_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_442_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_442_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_443_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_443_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_443_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_443_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_443_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_443_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_443_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_443_io_out_2; // @[Multiplier.scala 83:25]
  wire  c22_47_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_47_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_47_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_47_io_out_1; // @[Multiplier.scala 73:25]
  wire  c53_444_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_444_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_444_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_444_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_444_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_444_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_444_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_444_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_445_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_445_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_445_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_445_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_445_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_445_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_445_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_445_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_446_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_446_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_446_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_446_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_446_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_446_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_446_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_446_io_out_2; // @[Multiplier.scala 83:25]
  wire  c22_48_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_48_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_48_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_48_io_out_1; // @[Multiplier.scala 73:25]
  wire  c53_447_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_447_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_447_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_447_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_447_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_447_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_447_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_447_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_448_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_448_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_448_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_448_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_448_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_448_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_448_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_448_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_449_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_449_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_449_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_449_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_449_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_449_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_449_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_449_io_out_2; // @[Multiplier.scala 83:25]
  wire  c22_49_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_49_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_49_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_49_io_out_1; // @[Multiplier.scala 73:25]
  wire  c53_450_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_450_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_450_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_450_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_450_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_450_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_450_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_450_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_451_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_451_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_451_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_451_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_451_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_451_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_451_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_451_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_452_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_452_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_452_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_452_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_452_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_452_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_452_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_452_io_out_2; // @[Multiplier.scala 83:25]
  wire  c22_50_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_50_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_50_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_50_io_out_1; // @[Multiplier.scala 73:25]
  wire  c53_453_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_453_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_453_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_453_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_453_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_453_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_453_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_453_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_454_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_454_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_454_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_454_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_454_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_454_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_454_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_454_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_455_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_455_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_455_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_455_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_455_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_455_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_455_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_455_io_out_2; // @[Multiplier.scala 83:25]
  wire  c22_51_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_51_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_51_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_51_io_out_1; // @[Multiplier.scala 73:25]
  wire  c53_456_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_456_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_456_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_456_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_456_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_456_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_456_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_456_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_457_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_457_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_457_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_457_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_457_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_457_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_457_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_457_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_458_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_458_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_458_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_458_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_458_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_458_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_458_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_458_io_out_2; // @[Multiplier.scala 83:25]
  wire  c22_52_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_52_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_52_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_52_io_out_1; // @[Multiplier.scala 73:25]
  wire  c53_459_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_459_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_459_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_459_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_459_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_459_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_459_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_459_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_460_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_460_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_460_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_460_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_460_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_460_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_460_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_460_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_461_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_461_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_461_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_461_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_461_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_461_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_461_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_461_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_462_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_462_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_462_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_462_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_462_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_462_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_462_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_462_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_463_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_463_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_463_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_463_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_463_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_463_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_463_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_463_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_464_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_464_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_464_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_464_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_464_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_464_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_464_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_464_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_465_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_465_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_465_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_465_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_465_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_465_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_465_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_465_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_466_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_466_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_466_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_466_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_466_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_466_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_466_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_466_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_467_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_467_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_467_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_467_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_467_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_467_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_467_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_467_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_468_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_468_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_468_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_468_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_468_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_468_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_468_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_468_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_469_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_469_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_469_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_469_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_469_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_469_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_469_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_469_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_470_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_470_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_470_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_470_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_470_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_470_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_470_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_470_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_471_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_471_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_471_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_471_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_471_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_471_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_471_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_471_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_472_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_472_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_472_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_472_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_472_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_472_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_472_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_472_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_473_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_473_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_473_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_473_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_473_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_473_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_473_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_473_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_474_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_474_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_474_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_474_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_474_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_474_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_474_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_474_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_475_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_475_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_475_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_475_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_475_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_475_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_475_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_475_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_476_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_476_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_476_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_476_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_476_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_476_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_476_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_476_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_477_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_477_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_477_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_477_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_477_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_477_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_477_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_477_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_478_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_478_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_478_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_478_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_478_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_478_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_478_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_478_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_479_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_479_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_479_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_479_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_479_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_479_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_479_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_479_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_480_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_480_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_480_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_480_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_480_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_480_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_480_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_480_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_481_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_481_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_481_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_481_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_481_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_481_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_481_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_481_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_482_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_482_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_482_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_482_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_482_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_482_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_482_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_482_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_483_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_483_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_483_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_483_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_483_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_483_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_483_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_483_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_484_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_484_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_484_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_484_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_484_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_484_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_484_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_484_io_out_2; // @[Multiplier.scala 83:25]
  wire  c32_41_io_in_0; // @[Multiplier.scala 78:25]
  wire  c32_41_io_in_1; // @[Multiplier.scala 78:25]
  wire  c32_41_io_in_2; // @[Multiplier.scala 78:25]
  wire  c32_41_io_out_0; // @[Multiplier.scala 78:25]
  wire  c32_41_io_out_1; // @[Multiplier.scala 78:25]
  wire  c53_485_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_485_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_485_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_485_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_485_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_485_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_485_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_485_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_486_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_486_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_486_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_486_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_486_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_486_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_486_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_486_io_out_2; // @[Multiplier.scala 83:25]
  wire  c22_53_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_53_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_53_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_53_io_out_1; // @[Multiplier.scala 73:25]
  wire  c53_487_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_487_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_487_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_487_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_487_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_487_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_487_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_487_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_488_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_488_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_488_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_488_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_488_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_488_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_488_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_488_io_out_2; // @[Multiplier.scala 83:25]
  wire  c22_54_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_54_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_54_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_54_io_out_1; // @[Multiplier.scala 73:25]
  wire  c53_489_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_489_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_489_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_489_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_489_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_489_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_489_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_489_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_490_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_490_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_490_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_490_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_490_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_490_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_490_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_490_io_out_2; // @[Multiplier.scala 83:25]
  wire  c32_42_io_in_0; // @[Multiplier.scala 78:25]
  wire  c32_42_io_in_1; // @[Multiplier.scala 78:25]
  wire  c32_42_io_in_2; // @[Multiplier.scala 78:25]
  wire  c32_42_io_out_0; // @[Multiplier.scala 78:25]
  wire  c32_42_io_out_1; // @[Multiplier.scala 78:25]
  wire  c53_491_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_491_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_491_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_491_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_491_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_491_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_491_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_491_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_492_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_492_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_492_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_492_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_492_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_492_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_492_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_492_io_out_2; // @[Multiplier.scala 83:25]
  wire  c22_55_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_55_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_55_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_55_io_out_1; // @[Multiplier.scala 73:25]
  wire  c53_493_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_493_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_493_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_493_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_493_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_493_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_493_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_493_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_494_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_494_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_494_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_494_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_494_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_494_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_494_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_494_io_out_2; // @[Multiplier.scala 83:25]
  wire  c22_56_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_56_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_56_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_56_io_out_1; // @[Multiplier.scala 73:25]
  wire  c53_495_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_495_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_495_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_495_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_495_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_495_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_495_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_495_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_496_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_496_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_496_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_496_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_496_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_496_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_496_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_496_io_out_2; // @[Multiplier.scala 83:25]
  wire  c22_57_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_57_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_57_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_57_io_out_1; // @[Multiplier.scala 73:25]
  wire  c53_497_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_497_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_497_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_497_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_497_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_497_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_497_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_497_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_498_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_498_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_498_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_498_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_498_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_498_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_498_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_498_io_out_2; // @[Multiplier.scala 83:25]
  wire  c22_58_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_58_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_58_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_58_io_out_1; // @[Multiplier.scala 73:25]
  wire  c53_499_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_499_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_499_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_499_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_499_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_499_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_499_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_499_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_500_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_500_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_500_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_500_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_500_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_500_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_500_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_500_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_501_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_501_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_501_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_501_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_501_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_501_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_501_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_501_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_502_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_502_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_502_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_502_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_502_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_502_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_502_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_502_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_503_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_503_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_503_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_503_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_503_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_503_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_503_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_503_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_504_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_504_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_504_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_504_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_504_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_504_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_504_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_504_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_505_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_505_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_505_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_505_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_505_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_505_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_505_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_505_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_506_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_506_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_506_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_506_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_506_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_506_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_506_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_506_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_507_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_507_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_507_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_507_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_507_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_507_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_507_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_507_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_508_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_508_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_508_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_508_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_508_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_508_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_508_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_508_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_509_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_509_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_509_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_509_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_509_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_509_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_509_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_509_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_510_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_510_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_510_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_510_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_510_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_510_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_510_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_510_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_511_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_511_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_511_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_511_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_511_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_511_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_511_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_511_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_512_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_512_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_512_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_512_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_512_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_512_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_512_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_512_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_513_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_513_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_513_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_513_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_513_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_513_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_513_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_513_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_514_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_514_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_514_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_514_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_514_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_514_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_514_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_514_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_515_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_515_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_515_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_515_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_515_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_515_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_515_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_515_io_out_2; // @[Multiplier.scala 83:25]
  wire  c32_43_io_in_0; // @[Multiplier.scala 78:25]
  wire  c32_43_io_in_1; // @[Multiplier.scala 78:25]
  wire  c32_43_io_in_2; // @[Multiplier.scala 78:25]
  wire  c32_43_io_out_0; // @[Multiplier.scala 78:25]
  wire  c32_43_io_out_1; // @[Multiplier.scala 78:25]
  wire  c53_516_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_516_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_516_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_516_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_516_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_516_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_516_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_516_io_out_2; // @[Multiplier.scala 83:25]
  wire  c22_59_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_59_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_59_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_59_io_out_1; // @[Multiplier.scala 73:25]
  wire  c53_517_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_517_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_517_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_517_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_517_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_517_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_517_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_517_io_out_2; // @[Multiplier.scala 83:25]
  wire  c22_60_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_60_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_60_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_60_io_out_1; // @[Multiplier.scala 73:25]
  wire  c53_518_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_518_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_518_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_518_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_518_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_518_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_518_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_518_io_out_2; // @[Multiplier.scala 83:25]
  wire  c32_44_io_in_0; // @[Multiplier.scala 78:25]
  wire  c32_44_io_in_1; // @[Multiplier.scala 78:25]
  wire  c32_44_io_in_2; // @[Multiplier.scala 78:25]
  wire  c32_44_io_out_0; // @[Multiplier.scala 78:25]
  wire  c32_44_io_out_1; // @[Multiplier.scala 78:25]
  wire  c53_519_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_519_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_519_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_519_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_519_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_519_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_519_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_519_io_out_2; // @[Multiplier.scala 83:25]
  wire  c22_61_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_61_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_61_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_61_io_out_1; // @[Multiplier.scala 73:25]
  wire  c53_520_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_520_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_520_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_520_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_520_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_520_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_520_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_520_io_out_2; // @[Multiplier.scala 83:25]
  wire  c22_62_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_62_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_62_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_62_io_out_1; // @[Multiplier.scala 73:25]
  wire  c53_521_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_521_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_521_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_521_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_521_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_521_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_521_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_521_io_out_2; // @[Multiplier.scala 83:25]
  wire  c22_63_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_63_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_63_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_63_io_out_1; // @[Multiplier.scala 73:25]
  wire  c53_522_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_522_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_522_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_522_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_522_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_522_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_522_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_522_io_out_2; // @[Multiplier.scala 83:25]
  wire  c22_64_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_64_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_64_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_64_io_out_1; // @[Multiplier.scala 73:25]
  wire  c53_523_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_523_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_523_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_523_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_523_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_523_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_523_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_523_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_524_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_524_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_524_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_524_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_524_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_524_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_524_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_524_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_525_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_525_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_525_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_525_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_525_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_525_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_525_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_525_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_526_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_526_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_526_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_526_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_526_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_526_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_526_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_526_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_527_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_527_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_527_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_527_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_527_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_527_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_527_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_527_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_528_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_528_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_528_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_528_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_528_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_528_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_528_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_528_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_529_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_529_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_529_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_529_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_529_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_529_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_529_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_529_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_530_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_530_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_530_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_530_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_530_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_530_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_530_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_530_io_out_2; // @[Multiplier.scala 83:25]
  wire  c32_45_io_in_0; // @[Multiplier.scala 78:25]
  wire  c32_45_io_in_1; // @[Multiplier.scala 78:25]
  wire  c32_45_io_in_2; // @[Multiplier.scala 78:25]
  wire  c32_45_io_out_0; // @[Multiplier.scala 78:25]
  wire  c32_45_io_out_1; // @[Multiplier.scala 78:25]
  wire  c22_65_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_65_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_65_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_65_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_66_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_66_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_66_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_66_io_out_1; // @[Multiplier.scala 73:25]
  wire  c32_46_io_in_0; // @[Multiplier.scala 78:25]
  wire  c32_46_io_in_1; // @[Multiplier.scala 78:25]
  wire  c32_46_io_in_2; // @[Multiplier.scala 78:25]
  wire  c32_46_io_out_0; // @[Multiplier.scala 78:25]
  wire  c32_46_io_out_1; // @[Multiplier.scala 78:25]
  wire  c22_67_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_67_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_67_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_67_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_68_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_68_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_68_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_68_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_69_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_69_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_69_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_69_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_70_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_70_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_70_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_70_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_71_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_71_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_71_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_71_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_72_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_72_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_72_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_72_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_73_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_73_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_73_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_73_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_74_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_74_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_74_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_74_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_75_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_75_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_75_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_75_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_76_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_76_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_76_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_76_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_77_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_77_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_77_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_77_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_78_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_78_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_78_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_78_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_79_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_79_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_79_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_79_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_80_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_80_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_80_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_80_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_81_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_81_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_81_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_81_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_82_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_82_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_82_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_82_io_out_1; // @[Multiplier.scala 73:25]
  wire  c32_47_io_in_0; // @[Multiplier.scala 78:25]
  wire  c32_47_io_in_1; // @[Multiplier.scala 78:25]
  wire  c32_47_io_in_2; // @[Multiplier.scala 78:25]
  wire  c32_47_io_out_0; // @[Multiplier.scala 78:25]
  wire  c32_47_io_out_1; // @[Multiplier.scala 78:25]
  wire  c32_48_io_in_0; // @[Multiplier.scala 78:25]
  wire  c32_48_io_in_1; // @[Multiplier.scala 78:25]
  wire  c32_48_io_in_2; // @[Multiplier.scala 78:25]
  wire  c32_48_io_out_0; // @[Multiplier.scala 78:25]
  wire  c32_48_io_out_1; // @[Multiplier.scala 78:25]
  wire  c32_49_io_in_0; // @[Multiplier.scala 78:25]
  wire  c32_49_io_in_1; // @[Multiplier.scala 78:25]
  wire  c32_49_io_in_2; // @[Multiplier.scala 78:25]
  wire  c32_49_io_out_0; // @[Multiplier.scala 78:25]
  wire  c32_49_io_out_1; // @[Multiplier.scala 78:25]
  wire  c32_50_io_in_0; // @[Multiplier.scala 78:25]
  wire  c32_50_io_in_1; // @[Multiplier.scala 78:25]
  wire  c32_50_io_in_2; // @[Multiplier.scala 78:25]
  wire  c32_50_io_out_0; // @[Multiplier.scala 78:25]
  wire  c32_50_io_out_1; // @[Multiplier.scala 78:25]
  wire  c53_531_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_531_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_531_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_531_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_531_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_531_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_531_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_531_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_532_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_532_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_532_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_532_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_532_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_532_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_532_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_532_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_533_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_533_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_533_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_533_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_533_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_533_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_533_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_533_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_534_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_534_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_534_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_534_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_534_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_534_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_534_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_534_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_535_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_535_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_535_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_535_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_535_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_535_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_535_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_535_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_536_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_536_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_536_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_536_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_536_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_536_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_536_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_536_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_537_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_537_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_537_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_537_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_537_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_537_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_537_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_537_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_538_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_538_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_538_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_538_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_538_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_538_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_538_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_538_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_539_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_539_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_539_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_539_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_539_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_539_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_539_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_539_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_540_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_540_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_540_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_540_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_540_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_540_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_540_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_540_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_541_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_541_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_541_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_541_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_541_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_541_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_541_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_541_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_542_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_542_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_542_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_542_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_542_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_542_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_542_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_542_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_543_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_543_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_543_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_543_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_543_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_543_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_543_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_543_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_544_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_544_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_544_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_544_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_544_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_544_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_544_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_544_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_545_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_545_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_545_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_545_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_545_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_545_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_545_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_545_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_546_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_546_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_546_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_546_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_546_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_546_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_546_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_546_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_547_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_547_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_547_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_547_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_547_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_547_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_547_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_547_io_out_2; // @[Multiplier.scala 83:25]
  wire  c22_83_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_83_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_83_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_83_io_out_1; // @[Multiplier.scala 73:25]
  wire  c53_548_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_548_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_548_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_548_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_548_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_548_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_548_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_548_io_out_2; // @[Multiplier.scala 83:25]
  wire  c22_84_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_84_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_84_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_84_io_out_1; // @[Multiplier.scala 73:25]
  wire  c53_549_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_549_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_549_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_549_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_549_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_549_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_549_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_549_io_out_2; // @[Multiplier.scala 83:25]
  wire  c22_85_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_85_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_85_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_85_io_out_1; // @[Multiplier.scala 73:25]
  wire  c53_550_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_550_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_550_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_550_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_550_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_550_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_550_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_550_io_out_2; // @[Multiplier.scala 83:25]
  wire  c22_86_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_86_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_86_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_86_io_out_1; // @[Multiplier.scala 73:25]
  wire  c53_551_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_551_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_551_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_551_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_551_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_551_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_551_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_551_io_out_2; // @[Multiplier.scala 83:25]
  wire  c22_87_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_87_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_87_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_87_io_out_1; // @[Multiplier.scala 73:25]
  wire  c53_552_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_552_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_552_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_552_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_552_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_552_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_552_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_552_io_out_2; // @[Multiplier.scala 83:25]
  wire  c22_88_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_88_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_88_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_88_io_out_1; // @[Multiplier.scala 73:25]
  wire  c53_553_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_553_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_553_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_553_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_553_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_553_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_553_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_553_io_out_2; // @[Multiplier.scala 83:25]
  wire  c22_89_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_89_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_89_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_89_io_out_1; // @[Multiplier.scala 73:25]
  wire  c53_554_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_554_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_554_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_554_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_554_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_554_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_554_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_554_io_out_2; // @[Multiplier.scala 83:25]
  wire  c22_90_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_90_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_90_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_90_io_out_1; // @[Multiplier.scala 73:25]
  wire  c53_555_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_555_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_555_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_555_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_555_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_555_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_555_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_555_io_out_2; // @[Multiplier.scala 83:25]
  wire  c22_91_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_91_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_91_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_91_io_out_1; // @[Multiplier.scala 73:25]
  wire  c53_556_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_556_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_556_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_556_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_556_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_556_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_556_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_556_io_out_2; // @[Multiplier.scala 83:25]
  wire  c22_92_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_92_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_92_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_92_io_out_1; // @[Multiplier.scala 73:25]
  wire  c53_557_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_557_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_557_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_557_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_557_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_557_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_557_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_557_io_out_2; // @[Multiplier.scala 83:25]
  wire  c22_93_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_93_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_93_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_93_io_out_1; // @[Multiplier.scala 73:25]
  wire  c53_558_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_558_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_558_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_558_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_558_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_558_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_558_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_558_io_out_2; // @[Multiplier.scala 83:25]
  wire  c22_94_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_94_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_94_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_94_io_out_1; // @[Multiplier.scala 73:25]
  wire  c53_559_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_559_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_559_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_559_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_559_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_559_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_559_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_559_io_out_2; // @[Multiplier.scala 83:25]
  wire  c32_51_io_in_0; // @[Multiplier.scala 78:25]
  wire  c32_51_io_in_1; // @[Multiplier.scala 78:25]
  wire  c32_51_io_in_2; // @[Multiplier.scala 78:25]
  wire  c32_51_io_out_0; // @[Multiplier.scala 78:25]
  wire  c32_51_io_out_1; // @[Multiplier.scala 78:25]
  wire  c53_560_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_560_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_560_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_560_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_560_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_560_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_560_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_560_io_out_2; // @[Multiplier.scala 83:25]
  wire  c32_52_io_in_0; // @[Multiplier.scala 78:25]
  wire  c32_52_io_in_1; // @[Multiplier.scala 78:25]
  wire  c32_52_io_in_2; // @[Multiplier.scala 78:25]
  wire  c32_52_io_out_0; // @[Multiplier.scala 78:25]
  wire  c32_52_io_out_1; // @[Multiplier.scala 78:25]
  wire  c53_561_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_561_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_561_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_561_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_561_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_561_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_561_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_561_io_out_2; // @[Multiplier.scala 83:25]
  wire  c32_53_io_in_0; // @[Multiplier.scala 78:25]
  wire  c32_53_io_in_1; // @[Multiplier.scala 78:25]
  wire  c32_53_io_in_2; // @[Multiplier.scala 78:25]
  wire  c32_53_io_out_0; // @[Multiplier.scala 78:25]
  wire  c32_53_io_out_1; // @[Multiplier.scala 78:25]
  wire  c53_562_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_562_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_562_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_562_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_562_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_562_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_562_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_562_io_out_2; // @[Multiplier.scala 83:25]
  wire  c32_54_io_in_0; // @[Multiplier.scala 78:25]
  wire  c32_54_io_in_1; // @[Multiplier.scala 78:25]
  wire  c32_54_io_in_2; // @[Multiplier.scala 78:25]
  wire  c32_54_io_out_0; // @[Multiplier.scala 78:25]
  wire  c32_54_io_out_1; // @[Multiplier.scala 78:25]
  wire  c53_563_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_563_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_563_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_563_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_563_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_563_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_563_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_563_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_564_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_564_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_564_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_564_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_564_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_564_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_564_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_564_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_565_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_565_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_565_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_565_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_565_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_565_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_565_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_565_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_566_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_566_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_566_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_566_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_566_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_566_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_566_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_566_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_567_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_567_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_567_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_567_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_567_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_567_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_567_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_567_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_568_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_568_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_568_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_568_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_568_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_568_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_568_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_568_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_569_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_569_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_569_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_569_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_569_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_569_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_569_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_569_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_570_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_570_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_570_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_570_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_570_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_570_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_570_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_570_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_571_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_571_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_571_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_571_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_571_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_571_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_571_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_571_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_572_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_572_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_572_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_572_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_572_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_572_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_572_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_572_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_573_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_573_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_573_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_573_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_573_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_573_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_573_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_573_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_574_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_574_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_574_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_574_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_574_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_574_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_574_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_574_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_575_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_575_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_575_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_575_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_575_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_575_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_575_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_575_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_576_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_576_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_576_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_576_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_576_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_576_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_576_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_576_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_577_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_577_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_577_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_577_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_577_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_577_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_577_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_577_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_578_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_578_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_578_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_578_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_578_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_578_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_578_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_578_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_579_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_579_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_579_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_579_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_579_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_579_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_579_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_579_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_580_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_580_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_580_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_580_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_580_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_580_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_580_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_580_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_581_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_581_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_581_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_581_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_581_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_581_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_581_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_581_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_582_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_582_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_582_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_582_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_582_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_582_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_582_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_582_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_583_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_583_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_583_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_583_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_583_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_583_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_583_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_583_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_584_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_584_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_584_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_584_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_584_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_584_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_584_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_584_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_585_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_585_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_585_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_585_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_585_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_585_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_585_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_585_io_out_2; // @[Multiplier.scala 83:25]
  wire  c22_95_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_95_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_95_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_95_io_out_1; // @[Multiplier.scala 73:25]
  wire  c53_586_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_586_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_586_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_586_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_586_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_586_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_586_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_586_io_out_2; // @[Multiplier.scala 83:25]
  wire  c22_96_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_96_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_96_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_96_io_out_1; // @[Multiplier.scala 73:25]
  wire  c53_587_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_587_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_587_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_587_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_587_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_587_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_587_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_587_io_out_2; // @[Multiplier.scala 83:25]
  wire  c32_55_io_in_0; // @[Multiplier.scala 78:25]
  wire  c32_55_io_in_1; // @[Multiplier.scala 78:25]
  wire  c32_55_io_in_2; // @[Multiplier.scala 78:25]
  wire  c32_55_io_out_0; // @[Multiplier.scala 78:25]
  wire  c32_55_io_out_1; // @[Multiplier.scala 78:25]
  wire  c53_588_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_588_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_588_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_588_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_588_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_588_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_588_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_588_io_out_2; // @[Multiplier.scala 83:25]
  wire  c22_97_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_97_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_97_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_97_io_out_1; // @[Multiplier.scala 73:25]
  wire  c53_589_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_589_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_589_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_589_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_589_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_589_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_589_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_589_io_out_2; // @[Multiplier.scala 83:25]
  wire  c22_98_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_98_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_98_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_98_io_out_1; // @[Multiplier.scala 73:25]
  wire  c53_590_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_590_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_590_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_590_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_590_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_590_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_590_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_590_io_out_2; // @[Multiplier.scala 83:25]
  wire  c22_99_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_99_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_99_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_99_io_out_1; // @[Multiplier.scala 73:25]
  wire  c53_591_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_591_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_591_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_591_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_591_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_591_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_591_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_591_io_out_2; // @[Multiplier.scala 83:25]
  wire  c22_100_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_100_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_100_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_100_io_out_1; // @[Multiplier.scala 73:25]
  wire  c53_592_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_592_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_592_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_592_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_592_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_592_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_592_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_592_io_out_2; // @[Multiplier.scala 83:25]
  wire  c32_56_io_in_0; // @[Multiplier.scala 78:25]
  wire  c32_56_io_in_1; // @[Multiplier.scala 78:25]
  wire  c32_56_io_in_2; // @[Multiplier.scala 78:25]
  wire  c32_56_io_out_0; // @[Multiplier.scala 78:25]
  wire  c32_56_io_out_1; // @[Multiplier.scala 78:25]
  wire  c53_593_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_593_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_593_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_593_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_593_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_593_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_593_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_593_io_out_2; // @[Multiplier.scala 83:25]
  wire  c22_101_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_101_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_101_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_101_io_out_1; // @[Multiplier.scala 73:25]
  wire  c53_594_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_594_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_594_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_594_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_594_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_594_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_594_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_594_io_out_2; // @[Multiplier.scala 83:25]
  wire  c22_102_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_102_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_102_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_102_io_out_1; // @[Multiplier.scala 73:25]
  wire  c53_595_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_595_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_595_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_595_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_595_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_595_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_595_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_595_io_out_2; // @[Multiplier.scala 83:25]
  wire  c22_103_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_103_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_103_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_103_io_out_1; // @[Multiplier.scala 73:25]
  wire  c53_596_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_596_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_596_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_596_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_596_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_596_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_596_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_596_io_out_2; // @[Multiplier.scala 83:25]
  wire  c22_104_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_104_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_104_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_104_io_out_1; // @[Multiplier.scala 73:25]
  wire  c53_597_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_597_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_597_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_597_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_597_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_597_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_597_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_597_io_out_2; // @[Multiplier.scala 83:25]
  wire  c22_105_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_105_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_105_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_105_io_out_1; // @[Multiplier.scala 73:25]
  wire  c53_598_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_598_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_598_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_598_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_598_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_598_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_598_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_598_io_out_2; // @[Multiplier.scala 83:25]
  wire  c22_106_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_106_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_106_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_106_io_out_1; // @[Multiplier.scala 73:25]
  wire  c53_599_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_599_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_599_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_599_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_599_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_599_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_599_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_599_io_out_2; // @[Multiplier.scala 83:25]
  wire  c22_107_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_107_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_107_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_107_io_out_1; // @[Multiplier.scala 73:25]
  wire  c53_600_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_600_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_600_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_600_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_600_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_600_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_600_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_600_io_out_2; // @[Multiplier.scala 83:25]
  wire  c22_108_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_108_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_108_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_108_io_out_1; // @[Multiplier.scala 73:25]
  wire  c53_601_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_601_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_601_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_601_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_601_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_601_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_601_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_601_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_602_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_602_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_602_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_602_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_602_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_602_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_602_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_602_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_603_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_603_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_603_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_603_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_603_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_603_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_603_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_603_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_604_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_604_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_604_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_604_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_604_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_604_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_604_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_604_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_605_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_605_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_605_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_605_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_605_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_605_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_605_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_605_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_606_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_606_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_606_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_606_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_606_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_606_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_606_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_606_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_607_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_607_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_607_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_607_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_607_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_607_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_607_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_607_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_608_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_608_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_608_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_608_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_608_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_608_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_608_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_608_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_609_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_609_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_609_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_609_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_609_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_609_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_609_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_609_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_610_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_610_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_610_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_610_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_610_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_610_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_610_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_610_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_611_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_611_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_611_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_611_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_611_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_611_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_611_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_611_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_612_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_612_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_612_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_612_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_612_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_612_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_612_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_612_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_613_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_613_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_613_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_613_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_613_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_613_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_613_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_613_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_614_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_614_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_614_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_614_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_614_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_614_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_614_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_614_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_615_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_615_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_615_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_615_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_615_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_615_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_615_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_615_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_616_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_616_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_616_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_616_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_616_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_616_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_616_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_616_io_out_2; // @[Multiplier.scala 83:25]
  wire  c22_109_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_109_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_109_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_109_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_110_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_110_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_110_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_110_io_out_1; // @[Multiplier.scala 73:25]
  wire  c32_57_io_in_0; // @[Multiplier.scala 78:25]
  wire  c32_57_io_in_1; // @[Multiplier.scala 78:25]
  wire  c32_57_io_in_2; // @[Multiplier.scala 78:25]
  wire  c32_57_io_out_0; // @[Multiplier.scala 78:25]
  wire  c32_57_io_out_1; // @[Multiplier.scala 78:25]
  wire  c22_111_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_111_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_111_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_111_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_112_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_112_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_112_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_112_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_113_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_113_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_113_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_113_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_114_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_114_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_114_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_114_io_out_1; // @[Multiplier.scala 73:25]
  wire  c32_58_io_in_0; // @[Multiplier.scala 78:25]
  wire  c32_58_io_in_1; // @[Multiplier.scala 78:25]
  wire  c32_58_io_in_2; // @[Multiplier.scala 78:25]
  wire  c32_58_io_out_0; // @[Multiplier.scala 78:25]
  wire  c32_58_io_out_1; // @[Multiplier.scala 78:25]
  wire  c22_115_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_115_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_115_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_115_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_116_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_116_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_116_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_116_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_117_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_117_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_117_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_117_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_118_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_118_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_118_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_118_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_119_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_119_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_119_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_119_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_120_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_120_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_120_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_120_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_121_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_121_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_121_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_121_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_122_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_122_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_122_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_122_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_123_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_123_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_123_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_123_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_124_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_124_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_124_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_124_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_125_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_125_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_125_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_125_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_126_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_126_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_126_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_126_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_127_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_127_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_127_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_127_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_128_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_128_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_128_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_128_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_129_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_129_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_129_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_129_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_130_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_130_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_130_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_130_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_131_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_131_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_131_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_131_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_132_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_132_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_132_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_132_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_133_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_133_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_133_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_133_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_134_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_134_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_134_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_134_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_135_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_135_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_135_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_135_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_136_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_136_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_136_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_136_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_137_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_137_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_137_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_137_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_138_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_138_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_138_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_138_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_139_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_139_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_139_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_139_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_140_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_140_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_140_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_140_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_141_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_141_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_141_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_141_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_142_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_142_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_142_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_142_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_143_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_143_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_143_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_143_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_144_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_144_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_144_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_144_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_145_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_145_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_145_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_145_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_146_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_146_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_146_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_146_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_147_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_147_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_147_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_147_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_148_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_148_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_148_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_148_io_out_1; // @[Multiplier.scala 73:25]
  wire  c32_59_io_in_0; // @[Multiplier.scala 78:25]
  wire  c32_59_io_in_1; // @[Multiplier.scala 78:25]
  wire  c32_59_io_in_2; // @[Multiplier.scala 78:25]
  wire  c32_59_io_out_0; // @[Multiplier.scala 78:25]
  wire  c32_59_io_out_1; // @[Multiplier.scala 78:25]
  wire  c32_60_io_in_0; // @[Multiplier.scala 78:25]
  wire  c32_60_io_in_1; // @[Multiplier.scala 78:25]
  wire  c32_60_io_in_2; // @[Multiplier.scala 78:25]
  wire  c32_60_io_out_0; // @[Multiplier.scala 78:25]
  wire  c32_60_io_out_1; // @[Multiplier.scala 78:25]
  wire  c32_61_io_in_0; // @[Multiplier.scala 78:25]
  wire  c32_61_io_in_1; // @[Multiplier.scala 78:25]
  wire  c32_61_io_in_2; // @[Multiplier.scala 78:25]
  wire  c32_61_io_out_0; // @[Multiplier.scala 78:25]
  wire  c32_61_io_out_1; // @[Multiplier.scala 78:25]
  wire  c32_62_io_in_0; // @[Multiplier.scala 78:25]
  wire  c32_62_io_in_1; // @[Multiplier.scala 78:25]
  wire  c32_62_io_in_2; // @[Multiplier.scala 78:25]
  wire  c32_62_io_out_0; // @[Multiplier.scala 78:25]
  wire  c32_62_io_out_1; // @[Multiplier.scala 78:25]
  wire  c32_63_io_in_0; // @[Multiplier.scala 78:25]
  wire  c32_63_io_in_1; // @[Multiplier.scala 78:25]
  wire  c32_63_io_in_2; // @[Multiplier.scala 78:25]
  wire  c32_63_io_out_0; // @[Multiplier.scala 78:25]
  wire  c32_63_io_out_1; // @[Multiplier.scala 78:25]
  wire  c53_617_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_617_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_617_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_617_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_617_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_617_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_617_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_617_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_618_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_618_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_618_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_618_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_618_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_618_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_618_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_618_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_619_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_619_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_619_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_619_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_619_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_619_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_619_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_619_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_620_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_620_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_620_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_620_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_620_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_620_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_620_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_620_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_621_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_621_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_621_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_621_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_621_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_621_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_621_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_621_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_622_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_622_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_622_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_622_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_622_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_622_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_622_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_622_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_623_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_623_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_623_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_623_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_623_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_623_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_623_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_623_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_624_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_624_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_624_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_624_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_624_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_624_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_624_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_624_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_625_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_625_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_625_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_625_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_625_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_625_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_625_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_625_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_626_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_626_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_626_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_626_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_626_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_626_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_626_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_626_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_627_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_627_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_627_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_627_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_627_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_627_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_627_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_627_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_628_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_628_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_628_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_628_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_628_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_628_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_628_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_628_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_629_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_629_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_629_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_629_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_629_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_629_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_629_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_629_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_630_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_630_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_630_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_630_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_630_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_630_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_630_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_630_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_631_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_631_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_631_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_631_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_631_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_631_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_631_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_631_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_632_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_632_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_632_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_632_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_632_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_632_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_632_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_632_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_633_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_633_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_633_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_633_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_633_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_633_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_633_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_633_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_634_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_634_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_634_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_634_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_634_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_634_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_634_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_634_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_635_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_635_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_635_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_635_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_635_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_635_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_635_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_635_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_636_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_636_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_636_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_636_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_636_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_636_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_636_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_636_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_637_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_637_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_637_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_637_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_637_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_637_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_637_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_637_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_638_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_638_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_638_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_638_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_638_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_638_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_638_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_638_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_639_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_639_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_639_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_639_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_639_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_639_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_639_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_639_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_640_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_640_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_640_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_640_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_640_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_640_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_640_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_640_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_641_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_641_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_641_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_641_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_641_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_641_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_641_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_641_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_642_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_642_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_642_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_642_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_642_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_642_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_642_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_642_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_643_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_643_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_643_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_643_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_643_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_643_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_643_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_643_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_644_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_644_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_644_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_644_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_644_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_644_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_644_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_644_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_645_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_645_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_645_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_645_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_645_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_645_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_645_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_645_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_646_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_646_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_646_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_646_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_646_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_646_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_646_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_646_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_647_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_647_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_647_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_647_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_647_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_647_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_647_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_647_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_648_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_648_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_648_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_648_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_648_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_648_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_648_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_648_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_649_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_649_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_649_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_649_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_649_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_649_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_649_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_649_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_650_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_650_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_650_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_650_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_650_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_650_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_650_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_650_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_651_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_651_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_651_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_651_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_651_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_651_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_651_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_651_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_652_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_652_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_652_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_652_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_652_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_652_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_652_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_652_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_653_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_653_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_653_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_653_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_653_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_653_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_653_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_653_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_654_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_654_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_654_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_654_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_654_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_654_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_654_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_654_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_655_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_655_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_655_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_655_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_655_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_655_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_655_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_655_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_656_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_656_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_656_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_656_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_656_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_656_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_656_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_656_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_657_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_657_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_657_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_657_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_657_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_657_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_657_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_657_io_out_2; // @[Multiplier.scala 83:25]
  wire  c53_658_io_in_0; // @[Multiplier.scala 83:25]
  wire  c53_658_io_in_1; // @[Multiplier.scala 83:25]
  wire  c53_658_io_in_2; // @[Multiplier.scala 83:25]
  wire  c53_658_io_in_3; // @[Multiplier.scala 83:25]
  wire  c53_658_io_in_4; // @[Multiplier.scala 83:25]
  wire  c53_658_io_out_0; // @[Multiplier.scala 83:25]
  wire  c53_658_io_out_1; // @[Multiplier.scala 83:25]
  wire  c53_658_io_out_2; // @[Multiplier.scala 83:25]
  wire  c32_64_io_in_0; // @[Multiplier.scala 78:25]
  wire  c32_64_io_in_1; // @[Multiplier.scala 78:25]
  wire  c32_64_io_in_2; // @[Multiplier.scala 78:25]
  wire  c32_64_io_out_0; // @[Multiplier.scala 78:25]
  wire  c32_64_io_out_1; // @[Multiplier.scala 78:25]
  wire  c22_149_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_149_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_149_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_149_io_out_1; // @[Multiplier.scala 73:25]
  wire  c32_65_io_in_0; // @[Multiplier.scala 78:25]
  wire  c32_65_io_in_1; // @[Multiplier.scala 78:25]
  wire  c32_65_io_in_2; // @[Multiplier.scala 78:25]
  wire  c32_65_io_out_0; // @[Multiplier.scala 78:25]
  wire  c32_65_io_out_1; // @[Multiplier.scala 78:25]
  wire  c22_150_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_150_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_150_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_150_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_151_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_151_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_151_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_151_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_152_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_152_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_152_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_152_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_153_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_153_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_153_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_153_io_out_1; // @[Multiplier.scala 73:25]
  wire  c32_66_io_in_0; // @[Multiplier.scala 78:25]
  wire  c32_66_io_in_1; // @[Multiplier.scala 78:25]
  wire  c32_66_io_in_2; // @[Multiplier.scala 78:25]
  wire  c32_66_io_out_0; // @[Multiplier.scala 78:25]
  wire  c32_66_io_out_1; // @[Multiplier.scala 78:25]
  wire  c22_154_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_154_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_154_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_154_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_155_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_155_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_155_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_155_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_156_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_156_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_156_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_156_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_157_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_157_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_157_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_157_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_158_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_158_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_158_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_158_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_159_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_159_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_159_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_159_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_160_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_160_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_160_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_160_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_161_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_161_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_161_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_161_io_out_1; // @[Multiplier.scala 73:25]
  wire  c32_67_io_in_0; // @[Multiplier.scala 78:25]
  wire  c32_67_io_in_1; // @[Multiplier.scala 78:25]
  wire  c32_67_io_in_2; // @[Multiplier.scala 78:25]
  wire  c32_67_io_out_0; // @[Multiplier.scala 78:25]
  wire  c32_67_io_out_1; // @[Multiplier.scala 78:25]
  wire  c22_162_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_162_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_162_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_162_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_163_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_163_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_163_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_163_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_164_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_164_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_164_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_164_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_165_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_165_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_165_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_165_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_166_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_166_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_166_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_166_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_167_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_167_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_167_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_167_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_168_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_168_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_168_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_168_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_169_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_169_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_169_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_169_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_170_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_170_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_170_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_170_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_171_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_171_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_171_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_171_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_172_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_172_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_172_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_172_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_173_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_173_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_173_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_173_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_174_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_174_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_174_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_174_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_175_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_175_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_175_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_175_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_176_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_176_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_176_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_176_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_177_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_177_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_177_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_177_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_178_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_178_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_178_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_178_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_179_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_179_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_179_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_179_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_180_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_180_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_180_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_180_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_181_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_181_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_181_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_181_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_182_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_182_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_182_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_182_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_183_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_183_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_183_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_183_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_184_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_184_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_184_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_184_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_185_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_185_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_185_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_185_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_186_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_186_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_186_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_186_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_187_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_187_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_187_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_187_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_188_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_188_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_188_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_188_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_189_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_189_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_189_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_189_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_190_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_190_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_190_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_190_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_191_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_191_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_191_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_191_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_192_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_192_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_192_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_192_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_193_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_193_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_193_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_193_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_194_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_194_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_194_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_194_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_195_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_195_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_195_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_195_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_196_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_196_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_196_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_196_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_197_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_197_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_197_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_197_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_198_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_198_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_198_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_198_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_199_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_199_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_199_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_199_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_200_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_200_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_200_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_200_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_201_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_201_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_201_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_201_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_202_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_202_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_202_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_202_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_203_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_203_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_203_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_203_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_204_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_204_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_204_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_204_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_205_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_205_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_205_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_205_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_206_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_206_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_206_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_206_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_207_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_207_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_207_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_207_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_208_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_208_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_208_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_208_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_209_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_209_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_209_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_209_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_210_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_210_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_210_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_210_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_211_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_211_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_211_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_211_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_212_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_212_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_212_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_212_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_213_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_213_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_213_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_213_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_214_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_214_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_214_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_214_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_215_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_215_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_215_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_215_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_216_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_216_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_216_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_216_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_217_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_217_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_217_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_217_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_218_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_218_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_218_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_218_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_219_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_219_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_219_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_219_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_220_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_220_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_220_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_220_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_221_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_221_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_221_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_221_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_222_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_222_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_222_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_222_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_223_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_223_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_223_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_223_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_224_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_224_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_224_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_224_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_225_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_225_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_225_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_225_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_226_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_226_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_226_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_226_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_227_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_227_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_227_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_227_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_228_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_228_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_228_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_228_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_229_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_229_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_229_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_229_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_230_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_230_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_230_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_230_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_231_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_231_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_231_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_231_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_232_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_232_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_232_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_232_io_out_1; // @[Multiplier.scala 73:25]
  wire  c32_68_io_in_0; // @[Multiplier.scala 78:25]
  wire  c32_68_io_in_1; // @[Multiplier.scala 78:25]
  wire  c32_68_io_in_2; // @[Multiplier.scala 78:25]
  wire  c32_68_io_out_0; // @[Multiplier.scala 78:25]
  wire  c32_68_io_out_1; // @[Multiplier.scala 78:25]
  wire  c22_233_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_233_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_233_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_233_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_234_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_234_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_234_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_234_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_235_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_235_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_235_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_235_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_236_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_236_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_236_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_236_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_237_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_237_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_237_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_237_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_238_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_238_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_238_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_238_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_239_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_239_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_239_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_239_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_240_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_240_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_240_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_240_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_241_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_241_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_241_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_241_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_242_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_242_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_242_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_242_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_243_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_243_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_243_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_243_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_244_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_244_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_244_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_244_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_245_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_245_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_245_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_245_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_246_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_246_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_246_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_246_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_247_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_247_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_247_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_247_io_out_1; // @[Multiplier.scala 73:25]
  wire  c32_69_io_in_0; // @[Multiplier.scala 78:25]
  wire  c32_69_io_in_1; // @[Multiplier.scala 78:25]
  wire  c32_69_io_in_2; // @[Multiplier.scala 78:25]
  wire  c32_69_io_out_0; // @[Multiplier.scala 78:25]
  wire  c32_69_io_out_1; // @[Multiplier.scala 78:25]
  wire  c22_248_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_248_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_248_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_248_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_249_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_249_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_249_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_249_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_250_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_250_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_250_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_250_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_251_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_251_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_251_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_251_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_252_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_252_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_252_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_252_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_253_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_253_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_253_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_253_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_254_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_254_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_254_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_254_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_255_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_255_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_255_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_255_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_256_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_256_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_256_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_256_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_257_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_257_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_257_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_257_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_258_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_258_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_258_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_258_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_259_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_259_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_259_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_259_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_260_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_260_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_260_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_260_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_261_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_261_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_261_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_261_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_262_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_262_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_262_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_262_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_263_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_263_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_263_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_263_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_264_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_264_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_264_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_264_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_265_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_265_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_265_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_265_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_266_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_266_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_266_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_266_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_267_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_267_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_267_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_267_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_268_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_268_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_268_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_268_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_269_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_269_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_269_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_269_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_270_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_270_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_270_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_270_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_271_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_271_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_271_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_271_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_272_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_272_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_272_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_272_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_273_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_273_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_273_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_273_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_274_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_274_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_274_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_274_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_275_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_275_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_275_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_275_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_276_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_276_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_276_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_276_io_out_1; // @[Multiplier.scala 73:25]
  wire  c22_277_io_in_0; // @[Multiplier.scala 73:25]
  wire  c22_277_io_in_1; // @[Multiplier.scala 73:25]
  wire  c22_277_io_out_0; // @[Multiplier.scala 73:25]
  wire  c22_277_io_out_1; // @[Multiplier.scala 73:25]
  wire  b_sext_signBit = io_b[53]; // @[Multiplier.scala 9:20]
  wire [54:0] b_sext = {b_sext_signBit,io_b}; // @[Cat.scala 31:58]
  wire [55:0] _bx2_T = {b_sext, 1'h0}; // @[Multiplier.scala 26:17]
  wire [54:0] neg_b = ~b_sext; // @[Multiplier.scala 27:13]
  wire [55:0] _neg_bx2_T = {neg_b, 1'h0}; // @[Multiplier.scala 28:20]
  wire [2:0] x = {io_a[1:0],1'h0}; // @[Cat.scala 31:58]
  wire [54:0] _pp_temp_T_1 = 3'h1 == x ? b_sext : 55'h0; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_3 = 3'h2 == x ? b_sext : _pp_temp_T_1; // @[Mux.scala 81:58]
  wire [54:0] bx2 = _bx2_T[54:0]; // @[Multiplier.scala 24:41 26:7]
  wire [54:0] _pp_temp_T_5 = 3'h3 == x ? bx2 : _pp_temp_T_3; // @[Mux.scala 81:58]
  wire [54:0] neg_bx2 = _neg_bx2_T[54:0]; // @[Multiplier.scala 24:41 28:11]
  wire [54:0] _pp_temp_T_7 = 3'h4 == x ? neg_bx2 : _pp_temp_T_5; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_9 = 3'h5 == x ? neg_b : _pp_temp_T_7; // @[Mux.scala 81:58]
  wire [54:0] pp_temp = 3'h6 == x ? neg_b : _pp_temp_T_9; // @[Mux.scala 81:58]
  wire  s = pp_temp[54]; // @[Multiplier.scala 43:20]
  wire  _T = ~s; // @[Multiplier.scala 52:14]
  wire [57:0] pp = {_T,s,s,pp_temp}; // @[Cat.scala 31:58]
  wire [2:0] x_1 = io_a[3:1]; // @[Multiplier.scala 34:90]
  wire [54:0] _pp_temp_T_12 = 3'h1 == x_1 ? b_sext : 55'h0; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_14 = 3'h2 == x_1 ? b_sext : _pp_temp_T_12; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_16 = 3'h3 == x_1 ? bx2 : _pp_temp_T_14; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_18 = 3'h4 == x_1 ? neg_bx2 : _pp_temp_T_16; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_20 = 3'h5 == x_1 ? neg_b : _pp_temp_T_18; // @[Mux.scala 81:58]
  wire [54:0] pp_temp_1 = 3'h6 == x_1 ? neg_b : _pp_temp_T_20; // @[Mux.scala 81:58]
  wire  s_1 = pp_temp_1[54]; // @[Multiplier.scala 43:20]
  wire [1:0] _t_T_6 = 3'h4 == x ? 2'h2 : 2'h0; // @[Mux.scala 81:58]
  wire [1:0] _t_T_8 = 3'h5 == x ? 2'h1 : _t_T_6; // @[Mux.scala 81:58]
  wire [1:0] t_1 = 3'h6 == x ? 2'h1 : _t_T_8; // @[Mux.scala 81:58]
  wire  _T_59 = ~s_1; // @[Multiplier.scala 56:24]
  wire [58:0] pp_1 = {1'h1,_T_59,pp_temp_1,t_1}; // @[Cat.scala 31:58]
  wire [2:0] x_2 = io_a[5:3]; // @[Multiplier.scala 34:90]
  wire [54:0] _pp_temp_T_23 = 3'h1 == x_2 ? b_sext : 55'h0; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_25 = 3'h2 == x_2 ? b_sext : _pp_temp_T_23; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_27 = 3'h3 == x_2 ? bx2 : _pp_temp_T_25; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_29 = 3'h4 == x_2 ? neg_bx2 : _pp_temp_T_27; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_31 = 3'h5 == x_2 ? neg_b : _pp_temp_T_29; // @[Mux.scala 81:58]
  wire [54:0] pp_temp_2 = 3'h6 == x_2 ? neg_b : _pp_temp_T_31; // @[Mux.scala 81:58]
  wire  s_2 = pp_temp_2[54]; // @[Multiplier.scala 43:20]
  wire [1:0] _t_T_11 = 3'h4 == x_1 ? 2'h2 : 2'h0; // @[Mux.scala 81:58]
  wire [1:0] _t_T_13 = 3'h5 == x_1 ? 2'h1 : _t_T_11; // @[Mux.scala 81:58]
  wire [1:0] t_2 = 3'h6 == x_1 ? 2'h1 : _t_T_13; // @[Mux.scala 81:58]
  wire  _T_119 = ~s_2; // @[Multiplier.scala 56:24]
  wire [58:0] pp_2 = {1'h1,_T_119,pp_temp_2,t_2}; // @[Cat.scala 31:58]
  wire [2:0] x_3 = io_a[7:5]; // @[Multiplier.scala 34:90]
  wire [54:0] _pp_temp_T_34 = 3'h1 == x_3 ? b_sext : 55'h0; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_36 = 3'h2 == x_3 ? b_sext : _pp_temp_T_34; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_38 = 3'h3 == x_3 ? bx2 : _pp_temp_T_36; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_40 = 3'h4 == x_3 ? neg_bx2 : _pp_temp_T_38; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_42 = 3'h5 == x_3 ? neg_b : _pp_temp_T_40; // @[Mux.scala 81:58]
  wire [54:0] pp_temp_3 = 3'h6 == x_3 ? neg_b : _pp_temp_T_42; // @[Mux.scala 81:58]
  wire  s_3 = pp_temp_3[54]; // @[Multiplier.scala 43:20]
  wire [1:0] _t_T_16 = 3'h4 == x_2 ? 2'h2 : 2'h0; // @[Mux.scala 81:58]
  wire [1:0] _t_T_18 = 3'h5 == x_2 ? 2'h1 : _t_T_16; // @[Mux.scala 81:58]
  wire [1:0] t_3 = 3'h6 == x_2 ? 2'h1 : _t_T_18; // @[Mux.scala 81:58]
  wire  _T_179 = ~s_3; // @[Multiplier.scala 56:24]
  wire [58:0] pp_3 = {1'h1,_T_179,pp_temp_3,t_3}; // @[Cat.scala 31:58]
  wire [2:0] x_4 = io_a[9:7]; // @[Multiplier.scala 34:90]
  wire [54:0] _pp_temp_T_45 = 3'h1 == x_4 ? b_sext : 55'h0; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_47 = 3'h2 == x_4 ? b_sext : _pp_temp_T_45; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_49 = 3'h3 == x_4 ? bx2 : _pp_temp_T_47; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_51 = 3'h4 == x_4 ? neg_bx2 : _pp_temp_T_49; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_53 = 3'h5 == x_4 ? neg_b : _pp_temp_T_51; // @[Mux.scala 81:58]
  wire [54:0] pp_temp_4 = 3'h6 == x_4 ? neg_b : _pp_temp_T_53; // @[Mux.scala 81:58]
  wire  s_4 = pp_temp_4[54]; // @[Multiplier.scala 43:20]
  wire [1:0] _t_T_21 = 3'h4 == x_3 ? 2'h2 : 2'h0; // @[Mux.scala 81:58]
  wire [1:0] _t_T_23 = 3'h5 == x_3 ? 2'h1 : _t_T_21; // @[Mux.scala 81:58]
  wire [1:0] t_4 = 3'h6 == x_3 ? 2'h1 : _t_T_23; // @[Mux.scala 81:58]
  wire  _T_239 = ~s_4; // @[Multiplier.scala 56:24]
  wire [58:0] pp_4 = {1'h1,_T_239,pp_temp_4,t_4}; // @[Cat.scala 31:58]
  wire [2:0] x_5 = io_a[11:9]; // @[Multiplier.scala 34:90]
  wire [54:0] _pp_temp_T_56 = 3'h1 == x_5 ? b_sext : 55'h0; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_58 = 3'h2 == x_5 ? b_sext : _pp_temp_T_56; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_60 = 3'h3 == x_5 ? bx2 : _pp_temp_T_58; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_62 = 3'h4 == x_5 ? neg_bx2 : _pp_temp_T_60; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_64 = 3'h5 == x_5 ? neg_b : _pp_temp_T_62; // @[Mux.scala 81:58]
  wire [54:0] pp_temp_5 = 3'h6 == x_5 ? neg_b : _pp_temp_T_64; // @[Mux.scala 81:58]
  wire  s_5 = pp_temp_5[54]; // @[Multiplier.scala 43:20]
  wire [1:0] _t_T_26 = 3'h4 == x_4 ? 2'h2 : 2'h0; // @[Mux.scala 81:58]
  wire [1:0] _t_T_28 = 3'h5 == x_4 ? 2'h1 : _t_T_26; // @[Mux.scala 81:58]
  wire [1:0] t_5 = 3'h6 == x_4 ? 2'h1 : _t_T_28; // @[Mux.scala 81:58]
  wire  _T_299 = ~s_5; // @[Multiplier.scala 56:24]
  wire [58:0] pp_5 = {1'h1,_T_299,pp_temp_5,t_5}; // @[Cat.scala 31:58]
  wire [2:0] x_6 = io_a[13:11]; // @[Multiplier.scala 34:90]
  wire [54:0] _pp_temp_T_67 = 3'h1 == x_6 ? b_sext : 55'h0; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_69 = 3'h2 == x_6 ? b_sext : _pp_temp_T_67; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_71 = 3'h3 == x_6 ? bx2 : _pp_temp_T_69; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_73 = 3'h4 == x_6 ? neg_bx2 : _pp_temp_T_71; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_75 = 3'h5 == x_6 ? neg_b : _pp_temp_T_73; // @[Mux.scala 81:58]
  wire [54:0] pp_temp_6 = 3'h6 == x_6 ? neg_b : _pp_temp_T_75; // @[Mux.scala 81:58]
  wire  s_6 = pp_temp_6[54]; // @[Multiplier.scala 43:20]
  wire [1:0] _t_T_31 = 3'h4 == x_5 ? 2'h2 : 2'h0; // @[Mux.scala 81:58]
  wire [1:0] _t_T_33 = 3'h5 == x_5 ? 2'h1 : _t_T_31; // @[Mux.scala 81:58]
  wire [1:0] t_6 = 3'h6 == x_5 ? 2'h1 : _t_T_33; // @[Mux.scala 81:58]
  wire  _T_359 = ~s_6; // @[Multiplier.scala 56:24]
  wire [58:0] pp_6 = {1'h1,_T_359,pp_temp_6,t_6}; // @[Cat.scala 31:58]
  wire [2:0] x_7 = io_a[15:13]; // @[Multiplier.scala 34:90]
  wire [54:0] _pp_temp_T_78 = 3'h1 == x_7 ? b_sext : 55'h0; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_80 = 3'h2 == x_7 ? b_sext : _pp_temp_T_78; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_82 = 3'h3 == x_7 ? bx2 : _pp_temp_T_80; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_84 = 3'h4 == x_7 ? neg_bx2 : _pp_temp_T_82; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_86 = 3'h5 == x_7 ? neg_b : _pp_temp_T_84; // @[Mux.scala 81:58]
  wire [54:0] pp_temp_7 = 3'h6 == x_7 ? neg_b : _pp_temp_T_86; // @[Mux.scala 81:58]
  wire  s_7 = pp_temp_7[54]; // @[Multiplier.scala 43:20]
  wire [1:0] _t_T_36 = 3'h4 == x_6 ? 2'h2 : 2'h0; // @[Mux.scala 81:58]
  wire [1:0] _t_T_38 = 3'h5 == x_6 ? 2'h1 : _t_T_36; // @[Mux.scala 81:58]
  wire [1:0] t_7 = 3'h6 == x_6 ? 2'h1 : _t_T_38; // @[Mux.scala 81:58]
  wire  _T_419 = ~s_7; // @[Multiplier.scala 56:24]
  wire [58:0] pp_7 = {1'h1,_T_419,pp_temp_7,t_7}; // @[Cat.scala 31:58]
  wire [2:0] x_8 = io_a[17:15]; // @[Multiplier.scala 34:90]
  wire [54:0] _pp_temp_T_89 = 3'h1 == x_8 ? b_sext : 55'h0; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_91 = 3'h2 == x_8 ? b_sext : _pp_temp_T_89; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_93 = 3'h3 == x_8 ? bx2 : _pp_temp_T_91; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_95 = 3'h4 == x_8 ? neg_bx2 : _pp_temp_T_93; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_97 = 3'h5 == x_8 ? neg_b : _pp_temp_T_95; // @[Mux.scala 81:58]
  wire [54:0] pp_temp_8 = 3'h6 == x_8 ? neg_b : _pp_temp_T_97; // @[Mux.scala 81:58]
  wire  s_8 = pp_temp_8[54]; // @[Multiplier.scala 43:20]
  wire [1:0] _t_T_41 = 3'h4 == x_7 ? 2'h2 : 2'h0; // @[Mux.scala 81:58]
  wire [1:0] _t_T_43 = 3'h5 == x_7 ? 2'h1 : _t_T_41; // @[Mux.scala 81:58]
  wire [1:0] t_8 = 3'h6 == x_7 ? 2'h1 : _t_T_43; // @[Mux.scala 81:58]
  wire  _T_479 = ~s_8; // @[Multiplier.scala 56:24]
  wire [58:0] pp_8 = {1'h1,_T_479,pp_temp_8,t_8}; // @[Cat.scala 31:58]
  wire [2:0] x_9 = io_a[19:17]; // @[Multiplier.scala 34:90]
  wire [54:0] _pp_temp_T_100 = 3'h1 == x_9 ? b_sext : 55'h0; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_102 = 3'h2 == x_9 ? b_sext : _pp_temp_T_100; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_104 = 3'h3 == x_9 ? bx2 : _pp_temp_T_102; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_106 = 3'h4 == x_9 ? neg_bx2 : _pp_temp_T_104; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_108 = 3'h5 == x_9 ? neg_b : _pp_temp_T_106; // @[Mux.scala 81:58]
  wire [54:0] pp_temp_9 = 3'h6 == x_9 ? neg_b : _pp_temp_T_108; // @[Mux.scala 81:58]
  wire  s_9 = pp_temp_9[54]; // @[Multiplier.scala 43:20]
  wire [1:0] _t_T_46 = 3'h4 == x_8 ? 2'h2 : 2'h0; // @[Mux.scala 81:58]
  wire [1:0] _t_T_48 = 3'h5 == x_8 ? 2'h1 : _t_T_46; // @[Mux.scala 81:58]
  wire [1:0] t_9 = 3'h6 == x_8 ? 2'h1 : _t_T_48; // @[Mux.scala 81:58]
  wire  _T_539 = ~s_9; // @[Multiplier.scala 56:24]
  wire [58:0] pp_9 = {1'h1,_T_539,pp_temp_9,t_9}; // @[Cat.scala 31:58]
  wire [2:0] x_10 = io_a[21:19]; // @[Multiplier.scala 34:90]
  wire [54:0] _pp_temp_T_111 = 3'h1 == x_10 ? b_sext : 55'h0; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_113 = 3'h2 == x_10 ? b_sext : _pp_temp_T_111; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_115 = 3'h3 == x_10 ? bx2 : _pp_temp_T_113; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_117 = 3'h4 == x_10 ? neg_bx2 : _pp_temp_T_115; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_119 = 3'h5 == x_10 ? neg_b : _pp_temp_T_117; // @[Mux.scala 81:58]
  wire [54:0] pp_temp_10 = 3'h6 == x_10 ? neg_b : _pp_temp_T_119; // @[Mux.scala 81:58]
  wire  s_10 = pp_temp_10[54]; // @[Multiplier.scala 43:20]
  wire [1:0] _t_T_51 = 3'h4 == x_9 ? 2'h2 : 2'h0; // @[Mux.scala 81:58]
  wire [1:0] _t_T_53 = 3'h5 == x_9 ? 2'h1 : _t_T_51; // @[Mux.scala 81:58]
  wire [1:0] t_10 = 3'h6 == x_9 ? 2'h1 : _t_T_53; // @[Mux.scala 81:58]
  wire  _T_599 = ~s_10; // @[Multiplier.scala 56:24]
  wire [58:0] pp_10 = {1'h1,_T_599,pp_temp_10,t_10}; // @[Cat.scala 31:58]
  wire [2:0] x_11 = io_a[23:21]; // @[Multiplier.scala 34:90]
  wire [54:0] _pp_temp_T_122 = 3'h1 == x_11 ? b_sext : 55'h0; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_124 = 3'h2 == x_11 ? b_sext : _pp_temp_T_122; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_126 = 3'h3 == x_11 ? bx2 : _pp_temp_T_124; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_128 = 3'h4 == x_11 ? neg_bx2 : _pp_temp_T_126; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_130 = 3'h5 == x_11 ? neg_b : _pp_temp_T_128; // @[Mux.scala 81:58]
  wire [54:0] pp_temp_11 = 3'h6 == x_11 ? neg_b : _pp_temp_T_130; // @[Mux.scala 81:58]
  wire  s_11 = pp_temp_11[54]; // @[Multiplier.scala 43:20]
  wire [1:0] _t_T_56 = 3'h4 == x_10 ? 2'h2 : 2'h0; // @[Mux.scala 81:58]
  wire [1:0] _t_T_58 = 3'h5 == x_10 ? 2'h1 : _t_T_56; // @[Mux.scala 81:58]
  wire [1:0] t_11 = 3'h6 == x_10 ? 2'h1 : _t_T_58; // @[Mux.scala 81:58]
  wire  _T_659 = ~s_11; // @[Multiplier.scala 56:24]
  wire [58:0] pp_11 = {1'h1,_T_659,pp_temp_11,t_11}; // @[Cat.scala 31:58]
  wire [2:0] x_12 = io_a[25:23]; // @[Multiplier.scala 34:90]
  wire [54:0] _pp_temp_T_133 = 3'h1 == x_12 ? b_sext : 55'h0; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_135 = 3'h2 == x_12 ? b_sext : _pp_temp_T_133; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_137 = 3'h3 == x_12 ? bx2 : _pp_temp_T_135; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_139 = 3'h4 == x_12 ? neg_bx2 : _pp_temp_T_137; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_141 = 3'h5 == x_12 ? neg_b : _pp_temp_T_139; // @[Mux.scala 81:58]
  wire [54:0] pp_temp_12 = 3'h6 == x_12 ? neg_b : _pp_temp_T_141; // @[Mux.scala 81:58]
  wire  s_12 = pp_temp_12[54]; // @[Multiplier.scala 43:20]
  wire [1:0] _t_T_61 = 3'h4 == x_11 ? 2'h2 : 2'h0; // @[Mux.scala 81:58]
  wire [1:0] _t_T_63 = 3'h5 == x_11 ? 2'h1 : _t_T_61; // @[Mux.scala 81:58]
  wire [1:0] t_12 = 3'h6 == x_11 ? 2'h1 : _t_T_63; // @[Mux.scala 81:58]
  wire  _T_719 = ~s_12; // @[Multiplier.scala 56:24]
  wire [58:0] pp_12 = {1'h1,_T_719,pp_temp_12,t_12}; // @[Cat.scala 31:58]
  wire [2:0] x_13 = io_a[27:25]; // @[Multiplier.scala 34:90]
  wire [54:0] _pp_temp_T_144 = 3'h1 == x_13 ? b_sext : 55'h0; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_146 = 3'h2 == x_13 ? b_sext : _pp_temp_T_144; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_148 = 3'h3 == x_13 ? bx2 : _pp_temp_T_146; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_150 = 3'h4 == x_13 ? neg_bx2 : _pp_temp_T_148; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_152 = 3'h5 == x_13 ? neg_b : _pp_temp_T_150; // @[Mux.scala 81:58]
  wire [54:0] pp_temp_13 = 3'h6 == x_13 ? neg_b : _pp_temp_T_152; // @[Mux.scala 81:58]
  wire  s_13 = pp_temp_13[54]; // @[Multiplier.scala 43:20]
  wire [1:0] _t_T_66 = 3'h4 == x_12 ? 2'h2 : 2'h0; // @[Mux.scala 81:58]
  wire [1:0] _t_T_68 = 3'h5 == x_12 ? 2'h1 : _t_T_66; // @[Mux.scala 81:58]
  wire [1:0] t_13 = 3'h6 == x_12 ? 2'h1 : _t_T_68; // @[Mux.scala 81:58]
  wire  _T_779 = ~s_13; // @[Multiplier.scala 56:24]
  wire [58:0] pp_13 = {1'h1,_T_779,pp_temp_13,t_13}; // @[Cat.scala 31:58]
  wire [2:0] x_14 = io_a[29:27]; // @[Multiplier.scala 34:90]
  wire [54:0] _pp_temp_T_155 = 3'h1 == x_14 ? b_sext : 55'h0; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_157 = 3'h2 == x_14 ? b_sext : _pp_temp_T_155; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_159 = 3'h3 == x_14 ? bx2 : _pp_temp_T_157; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_161 = 3'h4 == x_14 ? neg_bx2 : _pp_temp_T_159; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_163 = 3'h5 == x_14 ? neg_b : _pp_temp_T_161; // @[Mux.scala 81:58]
  wire [54:0] pp_temp_14 = 3'h6 == x_14 ? neg_b : _pp_temp_T_163; // @[Mux.scala 81:58]
  wire  s_14 = pp_temp_14[54]; // @[Multiplier.scala 43:20]
  wire [1:0] _t_T_71 = 3'h4 == x_13 ? 2'h2 : 2'h0; // @[Mux.scala 81:58]
  wire [1:0] _t_T_73 = 3'h5 == x_13 ? 2'h1 : _t_T_71; // @[Mux.scala 81:58]
  wire [1:0] t_14 = 3'h6 == x_13 ? 2'h1 : _t_T_73; // @[Mux.scala 81:58]
  wire  _T_839 = ~s_14; // @[Multiplier.scala 56:24]
  wire [58:0] pp_14 = {1'h1,_T_839,pp_temp_14,t_14}; // @[Cat.scala 31:58]
  wire [2:0] x_15 = io_a[31:29]; // @[Multiplier.scala 34:90]
  wire [54:0] _pp_temp_T_166 = 3'h1 == x_15 ? b_sext : 55'h0; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_168 = 3'h2 == x_15 ? b_sext : _pp_temp_T_166; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_170 = 3'h3 == x_15 ? bx2 : _pp_temp_T_168; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_172 = 3'h4 == x_15 ? neg_bx2 : _pp_temp_T_170; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_174 = 3'h5 == x_15 ? neg_b : _pp_temp_T_172; // @[Mux.scala 81:58]
  wire [54:0] pp_temp_15 = 3'h6 == x_15 ? neg_b : _pp_temp_T_174; // @[Mux.scala 81:58]
  wire  s_15 = pp_temp_15[54]; // @[Multiplier.scala 43:20]
  wire [1:0] _t_T_76 = 3'h4 == x_14 ? 2'h2 : 2'h0; // @[Mux.scala 81:58]
  wire [1:0] _t_T_78 = 3'h5 == x_14 ? 2'h1 : _t_T_76; // @[Mux.scala 81:58]
  wire [1:0] t_15 = 3'h6 == x_14 ? 2'h1 : _t_T_78; // @[Mux.scala 81:58]
  wire  _T_899 = ~s_15; // @[Multiplier.scala 56:24]
  wire [58:0] pp_15 = {1'h1,_T_899,pp_temp_15,t_15}; // @[Cat.scala 31:58]
  wire [2:0] x_16 = io_a[33:31]; // @[Multiplier.scala 34:90]
  wire [54:0] _pp_temp_T_177 = 3'h1 == x_16 ? b_sext : 55'h0; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_179 = 3'h2 == x_16 ? b_sext : _pp_temp_T_177; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_181 = 3'h3 == x_16 ? bx2 : _pp_temp_T_179; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_183 = 3'h4 == x_16 ? neg_bx2 : _pp_temp_T_181; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_185 = 3'h5 == x_16 ? neg_b : _pp_temp_T_183; // @[Mux.scala 81:58]
  wire [54:0] pp_temp_16 = 3'h6 == x_16 ? neg_b : _pp_temp_T_185; // @[Mux.scala 81:58]
  wire  s_16 = pp_temp_16[54]; // @[Multiplier.scala 43:20]
  wire [1:0] _t_T_81 = 3'h4 == x_15 ? 2'h2 : 2'h0; // @[Mux.scala 81:58]
  wire [1:0] _t_T_83 = 3'h5 == x_15 ? 2'h1 : _t_T_81; // @[Mux.scala 81:58]
  wire [1:0] t_16 = 3'h6 == x_15 ? 2'h1 : _t_T_83; // @[Mux.scala 81:58]
  wire  _T_959 = ~s_16; // @[Multiplier.scala 56:24]
  wire [58:0] pp_16 = {1'h1,_T_959,pp_temp_16,t_16}; // @[Cat.scala 31:58]
  wire [2:0] x_17 = io_a[35:33]; // @[Multiplier.scala 34:90]
  wire [54:0] _pp_temp_T_188 = 3'h1 == x_17 ? b_sext : 55'h0; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_190 = 3'h2 == x_17 ? b_sext : _pp_temp_T_188; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_192 = 3'h3 == x_17 ? bx2 : _pp_temp_T_190; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_194 = 3'h4 == x_17 ? neg_bx2 : _pp_temp_T_192; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_196 = 3'h5 == x_17 ? neg_b : _pp_temp_T_194; // @[Mux.scala 81:58]
  wire [54:0] pp_temp_17 = 3'h6 == x_17 ? neg_b : _pp_temp_T_196; // @[Mux.scala 81:58]
  wire  s_17 = pp_temp_17[54]; // @[Multiplier.scala 43:20]
  wire [1:0] _t_T_86 = 3'h4 == x_16 ? 2'h2 : 2'h0; // @[Mux.scala 81:58]
  wire [1:0] _t_T_88 = 3'h5 == x_16 ? 2'h1 : _t_T_86; // @[Mux.scala 81:58]
  wire [1:0] t_17 = 3'h6 == x_16 ? 2'h1 : _t_T_88; // @[Mux.scala 81:58]
  wire  _T_1019 = ~s_17; // @[Multiplier.scala 56:24]
  wire [58:0] pp_17 = {1'h1,_T_1019,pp_temp_17,t_17}; // @[Cat.scala 31:58]
  wire [2:0] x_18 = io_a[37:35]; // @[Multiplier.scala 34:90]
  wire [54:0] _pp_temp_T_199 = 3'h1 == x_18 ? b_sext : 55'h0; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_201 = 3'h2 == x_18 ? b_sext : _pp_temp_T_199; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_203 = 3'h3 == x_18 ? bx2 : _pp_temp_T_201; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_205 = 3'h4 == x_18 ? neg_bx2 : _pp_temp_T_203; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_207 = 3'h5 == x_18 ? neg_b : _pp_temp_T_205; // @[Mux.scala 81:58]
  wire [54:0] pp_temp_18 = 3'h6 == x_18 ? neg_b : _pp_temp_T_207; // @[Mux.scala 81:58]
  wire  s_18 = pp_temp_18[54]; // @[Multiplier.scala 43:20]
  wire [1:0] _t_T_91 = 3'h4 == x_17 ? 2'h2 : 2'h0; // @[Mux.scala 81:58]
  wire [1:0] _t_T_93 = 3'h5 == x_17 ? 2'h1 : _t_T_91; // @[Mux.scala 81:58]
  wire [1:0] t_18 = 3'h6 == x_17 ? 2'h1 : _t_T_93; // @[Mux.scala 81:58]
  wire  _T_1079 = ~s_18; // @[Multiplier.scala 56:24]
  wire [58:0] pp_18 = {1'h1,_T_1079,pp_temp_18,t_18}; // @[Cat.scala 31:58]
  wire [2:0] x_19 = io_a[39:37]; // @[Multiplier.scala 34:90]
  wire [54:0] _pp_temp_T_210 = 3'h1 == x_19 ? b_sext : 55'h0; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_212 = 3'h2 == x_19 ? b_sext : _pp_temp_T_210; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_214 = 3'h3 == x_19 ? bx2 : _pp_temp_T_212; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_216 = 3'h4 == x_19 ? neg_bx2 : _pp_temp_T_214; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_218 = 3'h5 == x_19 ? neg_b : _pp_temp_T_216; // @[Mux.scala 81:58]
  wire [54:0] pp_temp_19 = 3'h6 == x_19 ? neg_b : _pp_temp_T_218; // @[Mux.scala 81:58]
  wire  s_19 = pp_temp_19[54]; // @[Multiplier.scala 43:20]
  wire [1:0] _t_T_96 = 3'h4 == x_18 ? 2'h2 : 2'h0; // @[Mux.scala 81:58]
  wire [1:0] _t_T_98 = 3'h5 == x_18 ? 2'h1 : _t_T_96; // @[Mux.scala 81:58]
  wire [1:0] t_19 = 3'h6 == x_18 ? 2'h1 : _t_T_98; // @[Mux.scala 81:58]
  wire  _T_1139 = ~s_19; // @[Multiplier.scala 56:24]
  wire [58:0] pp_19 = {1'h1,_T_1139,pp_temp_19,t_19}; // @[Cat.scala 31:58]
  wire [2:0] x_20 = io_a[41:39]; // @[Multiplier.scala 34:90]
  wire [54:0] _pp_temp_T_221 = 3'h1 == x_20 ? b_sext : 55'h0; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_223 = 3'h2 == x_20 ? b_sext : _pp_temp_T_221; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_225 = 3'h3 == x_20 ? bx2 : _pp_temp_T_223; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_227 = 3'h4 == x_20 ? neg_bx2 : _pp_temp_T_225; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_229 = 3'h5 == x_20 ? neg_b : _pp_temp_T_227; // @[Mux.scala 81:58]
  wire [54:0] pp_temp_20 = 3'h6 == x_20 ? neg_b : _pp_temp_T_229; // @[Mux.scala 81:58]
  wire  s_20 = pp_temp_20[54]; // @[Multiplier.scala 43:20]
  wire [1:0] _t_T_101 = 3'h4 == x_19 ? 2'h2 : 2'h0; // @[Mux.scala 81:58]
  wire [1:0] _t_T_103 = 3'h5 == x_19 ? 2'h1 : _t_T_101; // @[Mux.scala 81:58]
  wire [1:0] t_20 = 3'h6 == x_19 ? 2'h1 : _t_T_103; // @[Mux.scala 81:58]
  wire  _T_1199 = ~s_20; // @[Multiplier.scala 56:24]
  wire [58:0] pp_20 = {1'h1,_T_1199,pp_temp_20,t_20}; // @[Cat.scala 31:58]
  wire [2:0] x_21 = io_a[43:41]; // @[Multiplier.scala 34:90]
  wire [54:0] _pp_temp_T_232 = 3'h1 == x_21 ? b_sext : 55'h0; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_234 = 3'h2 == x_21 ? b_sext : _pp_temp_T_232; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_236 = 3'h3 == x_21 ? bx2 : _pp_temp_T_234; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_238 = 3'h4 == x_21 ? neg_bx2 : _pp_temp_T_236; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_240 = 3'h5 == x_21 ? neg_b : _pp_temp_T_238; // @[Mux.scala 81:58]
  wire [54:0] pp_temp_21 = 3'h6 == x_21 ? neg_b : _pp_temp_T_240; // @[Mux.scala 81:58]
  wire  s_21 = pp_temp_21[54]; // @[Multiplier.scala 43:20]
  wire [1:0] _t_T_106 = 3'h4 == x_20 ? 2'h2 : 2'h0; // @[Mux.scala 81:58]
  wire [1:0] _t_T_108 = 3'h5 == x_20 ? 2'h1 : _t_T_106; // @[Mux.scala 81:58]
  wire [1:0] t_21 = 3'h6 == x_20 ? 2'h1 : _t_T_108; // @[Mux.scala 81:58]
  wire  _T_1259 = ~s_21; // @[Multiplier.scala 56:24]
  wire [58:0] pp_21 = {1'h1,_T_1259,pp_temp_21,t_21}; // @[Cat.scala 31:58]
  wire [2:0] x_22 = io_a[45:43]; // @[Multiplier.scala 34:90]
  wire [54:0] _pp_temp_T_243 = 3'h1 == x_22 ? b_sext : 55'h0; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_245 = 3'h2 == x_22 ? b_sext : _pp_temp_T_243; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_247 = 3'h3 == x_22 ? bx2 : _pp_temp_T_245; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_249 = 3'h4 == x_22 ? neg_bx2 : _pp_temp_T_247; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_251 = 3'h5 == x_22 ? neg_b : _pp_temp_T_249; // @[Mux.scala 81:58]
  wire [54:0] pp_temp_22 = 3'h6 == x_22 ? neg_b : _pp_temp_T_251; // @[Mux.scala 81:58]
  wire  s_22 = pp_temp_22[54]; // @[Multiplier.scala 43:20]
  wire [1:0] _t_T_111 = 3'h4 == x_21 ? 2'h2 : 2'h0; // @[Mux.scala 81:58]
  wire [1:0] _t_T_113 = 3'h5 == x_21 ? 2'h1 : _t_T_111; // @[Mux.scala 81:58]
  wire [1:0] t_22 = 3'h6 == x_21 ? 2'h1 : _t_T_113; // @[Mux.scala 81:58]
  wire  _T_1319 = ~s_22; // @[Multiplier.scala 56:24]
  wire [58:0] pp_22 = {1'h1,_T_1319,pp_temp_22,t_22}; // @[Cat.scala 31:58]
  wire [2:0] x_23 = io_a[47:45]; // @[Multiplier.scala 34:90]
  wire [54:0] _pp_temp_T_254 = 3'h1 == x_23 ? b_sext : 55'h0; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_256 = 3'h2 == x_23 ? b_sext : _pp_temp_T_254; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_258 = 3'h3 == x_23 ? bx2 : _pp_temp_T_256; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_260 = 3'h4 == x_23 ? neg_bx2 : _pp_temp_T_258; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_262 = 3'h5 == x_23 ? neg_b : _pp_temp_T_260; // @[Mux.scala 81:58]
  wire [54:0] pp_temp_23 = 3'h6 == x_23 ? neg_b : _pp_temp_T_262; // @[Mux.scala 81:58]
  wire  s_23 = pp_temp_23[54]; // @[Multiplier.scala 43:20]
  wire [1:0] _t_T_116 = 3'h4 == x_22 ? 2'h2 : 2'h0; // @[Mux.scala 81:58]
  wire [1:0] _t_T_118 = 3'h5 == x_22 ? 2'h1 : _t_T_116; // @[Mux.scala 81:58]
  wire [1:0] t_23 = 3'h6 == x_22 ? 2'h1 : _t_T_118; // @[Mux.scala 81:58]
  wire  _T_1379 = ~s_23; // @[Multiplier.scala 56:24]
  wire [58:0] pp_23 = {1'h1,_T_1379,pp_temp_23,t_23}; // @[Cat.scala 31:58]
  wire [2:0] x_24 = io_a[49:47]; // @[Multiplier.scala 34:90]
  wire [54:0] _pp_temp_T_265 = 3'h1 == x_24 ? b_sext : 55'h0; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_267 = 3'h2 == x_24 ? b_sext : _pp_temp_T_265; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_269 = 3'h3 == x_24 ? bx2 : _pp_temp_T_267; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_271 = 3'h4 == x_24 ? neg_bx2 : _pp_temp_T_269; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_273 = 3'h5 == x_24 ? neg_b : _pp_temp_T_271; // @[Mux.scala 81:58]
  wire [54:0] pp_temp_24 = 3'h6 == x_24 ? neg_b : _pp_temp_T_273; // @[Mux.scala 81:58]
  wire  s_24 = pp_temp_24[54]; // @[Multiplier.scala 43:20]
  wire [1:0] _t_T_121 = 3'h4 == x_23 ? 2'h2 : 2'h0; // @[Mux.scala 81:58]
  wire [1:0] _t_T_123 = 3'h5 == x_23 ? 2'h1 : _t_T_121; // @[Mux.scala 81:58]
  wire [1:0] t_24 = 3'h6 == x_23 ? 2'h1 : _t_T_123; // @[Mux.scala 81:58]
  wire  _T_1439 = ~s_24; // @[Multiplier.scala 56:24]
  wire [58:0] pp_24 = {1'h1,_T_1439,pp_temp_24,t_24}; // @[Cat.scala 31:58]
  wire [2:0] x_25 = io_a[51:49]; // @[Multiplier.scala 34:90]
  wire [54:0] _pp_temp_T_276 = 3'h1 == x_25 ? b_sext : 55'h0; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_278 = 3'h2 == x_25 ? b_sext : _pp_temp_T_276; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_280 = 3'h3 == x_25 ? bx2 : _pp_temp_T_278; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_282 = 3'h4 == x_25 ? neg_bx2 : _pp_temp_T_280; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_284 = 3'h5 == x_25 ? neg_b : _pp_temp_T_282; // @[Mux.scala 81:58]
  wire [54:0] pp_temp_25 = 3'h6 == x_25 ? neg_b : _pp_temp_T_284; // @[Mux.scala 81:58]
  wire  s_25 = pp_temp_25[54]; // @[Multiplier.scala 43:20]
  wire [1:0] _t_T_126 = 3'h4 == x_24 ? 2'h2 : 2'h0; // @[Mux.scala 81:58]
  wire [1:0] _t_T_128 = 3'h5 == x_24 ? 2'h1 : _t_T_126; // @[Mux.scala 81:58]
  wire [1:0] t_25 = 3'h6 == x_24 ? 2'h1 : _t_T_128; // @[Mux.scala 81:58]
  wire  _T_1499 = ~s_25; // @[Multiplier.scala 56:24]
  wire [58:0] pp_25 = {1'h1,_T_1499,pp_temp_25,t_25}; // @[Cat.scala 31:58]
  wire [2:0] last_x_1 = io_a[53:51]; // @[Multiplier.scala 34:90]
  wire [54:0] _pp_temp_T_287 = 3'h1 == last_x_1 ? b_sext : 55'h0; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_289 = 3'h2 == last_x_1 ? b_sext : _pp_temp_T_287; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_291 = 3'h3 == last_x_1 ? bx2 : _pp_temp_T_289; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_293 = 3'h4 == last_x_1 ? neg_bx2 : _pp_temp_T_291; // @[Mux.scala 81:58]
  wire [54:0] _pp_temp_T_295 = 3'h5 == last_x_1 ? neg_b : _pp_temp_T_293; // @[Mux.scala 81:58]
  wire [54:0] pp_temp_26 = 3'h6 == last_x_1 ? neg_b : _pp_temp_T_295; // @[Mux.scala 81:58]
  wire  s_26 = pp_temp_26[54]; // @[Multiplier.scala 43:20]
  wire [1:0] _t_T_131 = 3'h4 == x_25 ? 2'h2 : 2'h0; // @[Mux.scala 81:58]
  wire [1:0] _t_T_133 = 3'h5 == x_25 ? 2'h1 : _t_T_131; // @[Mux.scala 81:58]
  wire [1:0] t_26 = 3'h6 == x_25 ? 2'h1 : _t_T_133; // @[Mux.scala 81:58]
  wire  _T_1559 = ~s_26; // @[Multiplier.scala 54:14]
  wire [57:0] pp_26 = {_T_1559,pp_temp_26,t_26}; // @[Cat.scala 31:58]
  wire  s_0 = c22_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_1_5 = c53_11_io_out_2; // @[Multiplier.scala 90:41]
  wire  c2_1_6 = c53_13_io_out_2; // @[Multiplier.scala 90:41]
  wire  c2_1_7 = c53_15_io_out_2; // @[Multiplier.scala 90:41]
  wire  c2_3_5 = c53_55_io_out_2; // @[Multiplier.scala 90:41]
  wire  c2_3_6 = c53_59_io_out_2; // @[Multiplier.scala 90:41]
  wire  c2_3_7 = c53_63_io_out_2; // @[Multiplier.scala 90:41]
  wire  c2_5_5 = c53_131_io_out_2; // @[Multiplier.scala 90:41]
  wire  c2_5_6 = c53_137_io_out_2; // @[Multiplier.scala 90:41]
  wire  c2_5_7 = c53_143_io_out_2; // @[Multiplier.scala 90:41]
  wire  c2_5_19 = c53_215_io_out_2; // @[Multiplier.scala 90:41]
  wire  c2_5_22 = c53_233_io_out_2; // @[Multiplier.scala 90:41]
  wire  c2_3_51 = c53_293_io_out_2; // @[Multiplier.scala 90:41]
  wire  c2_3_54 = c53_305_io_out_2; // @[Multiplier.scala 90:41]
  wire  c2_1_83 = c53_339_io_out_2; // @[Multiplier.scala 90:41]
  wire  c2_1_86 = c53_345_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_0_107 = c22_27_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_107 = c22_27_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_108 = c22_28_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_108 = c22_28_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_109 = c22_29_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_109 = c22_29_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_110 = c22_30_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_110 = c22_30_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_111 = c22_31_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_111 = c22_31_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_112 = c32_32_io_out_0; // @[Multiplier.scala 80:35]
  wire  c2_0_112 = c32_32_io_out_1; // @[Multiplier.scala 81:41]
  wire  s_0_113 = c32_33_io_out_0; // @[Multiplier.scala 80:35]
  wire  c2_0_113 = c32_33_io_out_1; // @[Multiplier.scala 81:41]
  wire  s_0_114 = c32_34_io_out_0; // @[Multiplier.scala 80:35]
  wire  c2_0_114 = c32_34_io_out_1; // @[Multiplier.scala 81:41]
  wire  s_0_115 = c53_354_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_115 = c53_354_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_0_116 = c53_355_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_116 = c53_355_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_0_117 = c53_356_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_117 = c53_356_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_0_118 = c53_357_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_118 = c53_357_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_0_119 = c53_358_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_119 = c53_358_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_0_120 = c53_359_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_120 = c53_359_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_0_121 = c53_360_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_121 = c53_360_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_0_122 = c53_361_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_122 = c53_361_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_0_123 = c53_362_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_123 = c53_362_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_1_92 = c22_32_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_1_91 = c22_32_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_124 = c53_363_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_124 = c53_363_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_1_93 = c22_33_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_1_92 = c22_33_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_125 = c53_364_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_125 = c53_364_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_1_94 = c22_34_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_1_93 = c22_34_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_126 = c53_365_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_126 = c53_365_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_1_95 = c22_35_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_1_94 = c22_35_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_127 = c53_366_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_127 = c53_366_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_1_96 = c22_36_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_1_95 = c22_36_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_128 = c53_367_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_128 = c53_367_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_1_97 = c32_35_io_out_0; // @[Multiplier.scala 80:35]
  wire  c2_1_96 = c32_35_io_out_1; // @[Multiplier.scala 81:41]
  wire  s_0_129 = c53_368_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_129 = c53_368_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_1_98 = c32_36_io_out_0; // @[Multiplier.scala 80:35]
  wire  c2_1_97 = c32_36_io_out_1; // @[Multiplier.scala 81:41]
  wire  s_0_130 = c53_369_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_130 = c53_369_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_1_99 = c32_37_io_out_0; // @[Multiplier.scala 80:35]
  wire  c2_1_98 = c32_37_io_out_1; // @[Multiplier.scala 81:41]
  wire  s_0_131 = c53_370_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_131 = c53_370_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_1_100 = c53_371_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_1_99 = c53_371_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_0_132 = c53_372_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_132 = c53_372_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_1_101 = c53_373_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_1_100 = c53_373_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_0_133 = c53_374_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_133 = c53_374_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_1_102 = c53_375_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_1_101 = c53_375_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_0_134 = c53_376_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_134 = c53_376_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_1_103 = c53_377_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_1_102 = c53_377_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_0_135 = c53_378_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_135 = c53_378_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_1_104 = c53_379_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_1_103 = c53_379_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_0_136 = c53_380_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_136 = c53_380_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_1_105 = c53_381_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_1_104 = c53_381_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_0_137 = c53_382_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_137 = c53_382_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_1_106 = c53_383_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_1_105 = c53_383_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_0_138 = c53_384_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_138 = c53_384_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_1_107 = c53_385_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_1_106 = c53_385_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_0_139 = c53_386_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_139 = c53_386_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_1_108 = c53_387_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_1_107 = c53_387_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_2_76 = c22_37_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_2_75 = c22_37_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_140 = c53_388_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_140 = c53_388_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_1_109 = c53_389_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_1_108 = c53_389_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_2_77 = c22_38_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_2_76 = c22_38_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_141 = c53_390_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_141 = c53_390_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_1_110 = c53_391_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_1_109 = c53_391_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_2_78 = c22_39_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_2_77 = c22_39_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_142 = c53_392_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_142 = c53_392_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_1_111 = c53_393_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_1_110 = c53_393_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_2_79 = c22_40_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_2_78 = c22_40_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_143 = c53_394_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_143 = c53_394_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_1_112 = c53_395_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_1_111 = c53_395_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_2_80 = c22_41_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_2_79 = c22_41_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_144 = c53_396_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_144 = c53_396_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_1_113 = c53_397_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_1_112 = c53_397_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_2_81 = c32_38_io_out_0; // @[Multiplier.scala 80:35]
  wire  c2_2_80 = c32_38_io_out_1; // @[Multiplier.scala 81:41]
  wire  s_0_145 = c53_398_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_145 = c53_398_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_1_114 = c53_399_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_1_113 = c53_399_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_2_82 = c32_39_io_out_0; // @[Multiplier.scala 80:35]
  wire  c2_2_81 = c32_39_io_out_1; // @[Multiplier.scala 81:41]
  wire  s_0_146 = c53_400_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_146 = c53_400_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_1_115 = c53_401_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_1_114 = c53_401_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_2_83 = c32_40_io_out_0; // @[Multiplier.scala 80:35]
  wire  c2_2_82 = c32_40_io_out_1; // @[Multiplier.scala 81:41]
  wire  s_0_147 = c53_402_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_147 = c53_402_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_1_116 = c53_403_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_1_115 = c53_403_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_2_84 = c53_404_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_2_83 = c53_404_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_0_148 = c53_405_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_148 = c53_405_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_1_117 = c53_406_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_1_116 = c53_406_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_2_85 = c53_407_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_2_84 = c53_407_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_0_149 = c53_408_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_149 = c53_408_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_1_118 = c53_409_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_1_117 = c53_409_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_2_86 = c53_410_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_2_85 = c53_410_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_0_150 = c53_411_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_150 = c53_411_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_1_119 = c53_412_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_1_118 = c53_412_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_2_87 = c53_413_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_2_86 = c53_413_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_0_151 = c53_414_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_151 = c53_414_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_1_120 = c53_415_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_1_119 = c53_415_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_2_88 = c53_416_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_2_87 = c53_416_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_0_152 = c53_417_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_152 = c53_417_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_1_121 = c53_418_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_1_120 = c53_418_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_2_89 = c53_419_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_2_88 = c53_419_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_0_153 = c53_420_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_153 = c53_420_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_1_122 = c53_421_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_1_121 = c53_421_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_2_90 = c53_422_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_2_89 = c53_422_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_0_154 = c53_423_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_154 = c53_423_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_1_123 = c53_424_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_1_122 = c53_424_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_2_91 = c53_425_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_2_90 = c53_425_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_0_155 = c53_426_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_155 = c53_426_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_1_124 = c53_427_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_1_123 = c53_427_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_2_92 = c53_428_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_2_91 = c53_428_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_3_60 = c22_42_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_3_59 = c22_42_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_156 = c53_429_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_156 = c53_429_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_1_125 = c53_430_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_1_124 = c53_430_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_2_93 = c53_431_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_2_92 = c53_431_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_3_61 = c22_43_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_3_60 = c22_43_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_157 = c53_432_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_157 = c53_432_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_1_126 = c53_433_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_1_125 = c53_433_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_2_94 = c53_434_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_2_93 = c53_434_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_3_62 = c22_44_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_3_61 = c22_44_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_158 = c53_435_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_158 = c53_435_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_1_127 = c53_436_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_1_126 = c53_436_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_2_95 = c53_437_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_2_94 = c53_437_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_3_63 = c22_45_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_3_62 = c22_45_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_159 = c53_438_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_159 = c53_438_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_1_128 = c53_439_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_1_127 = c53_439_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_2_96 = c53_440_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_2_95 = c53_440_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_3_64 = c22_46_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_3_63 = c22_46_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_160 = c53_441_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_160 = c53_441_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_1_129 = c53_442_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_1_128 = c53_442_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_2_97 = c53_443_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_2_96 = c53_443_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_3_65 = c22_47_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_3_64 = c22_47_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_161 = c53_444_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_161 = c53_444_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_1_130 = c53_445_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_1_129 = c53_445_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_2_98 = c53_446_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_2_97 = c53_446_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_3_66 = c22_48_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_3_65 = c22_48_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_162 = c53_447_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_162 = c53_447_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_1_131 = c53_448_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_1_130 = c53_448_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_2_99 = c53_449_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_2_98 = c53_449_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_3_67 = c22_49_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_3_66 = c22_49_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_163 = c53_450_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_163 = c53_450_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_1_132 = c53_451_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_1_131 = c53_451_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_2_100 = c53_452_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_2_99 = c53_452_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_3_68 = c22_50_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_3_67 = c22_50_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_164 = c53_453_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_164 = c53_453_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_1_133 = c53_454_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_1_132 = c53_454_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_2_101 = c53_455_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_2_100 = c53_455_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_3_69 = c22_51_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_3_68 = c22_51_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_165 = c53_456_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_165 = c53_456_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_1_134 = c53_457_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_1_133 = c53_457_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_2_102 = c53_458_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_2_101 = c53_458_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_3_70 = c22_52_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_3_69 = c22_52_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_166 = c53_459_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_166 = c53_459_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_1_135 = c53_460_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_1_134 = c53_460_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_2_103 = c53_461_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_2_102 = c53_461_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_0_167 = c53_462_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_167 = c53_462_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_1_136 = c53_463_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_1_135 = c53_463_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_2_104 = c53_464_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_2_103 = c53_464_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_0_168 = c53_465_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_168 = c53_465_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_1_137 = c53_466_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_1_136 = c53_466_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_2_105 = c53_467_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_2_104 = c53_467_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_0_169 = c53_468_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_169 = c53_468_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_1_138 = c53_469_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_1_137 = c53_469_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_2_106 = c53_470_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_2_105 = c53_470_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_0_170 = c53_471_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_170 = c53_471_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_1_139 = c53_472_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_1_138 = c53_472_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_2_107 = c53_473_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_2_106 = c53_473_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_0_171 = c53_474_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_171 = c53_474_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_1_140 = c53_475_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_1_139 = c53_475_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_2_108 = c53_476_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_2_107 = c53_476_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_0_172 = c53_477_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_172 = c53_477_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_1_141 = c53_478_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_1_140 = c53_478_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_2_109 = c53_479_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_2_108 = c53_479_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_0_173 = c53_480_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_173 = c53_480_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_1_142 = c53_481_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_1_141 = c53_481_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_2_110 = c53_482_io_out_0; // @[Multiplier.scala 88:39]
  wire  c1_2_93 = c53_482_io_out_1; // @[Multiplier.scala 89:41]
  wire  c2_2_109 = c53_482_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_0_174 = c53_483_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_174 = c53_483_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_1_143 = c53_484_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_1_142 = c53_484_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_2_111 = c32_41_io_out_0; // @[Multiplier.scala 80:35]
  wire  c2_2_110 = c32_41_io_out_1; // @[Multiplier.scala 81:41]
  wire  s_0_175 = c53_485_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_175 = c53_485_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_1_144 = c53_486_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_1_143 = c53_486_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_2_112 = c22_53_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_2_111 = c22_53_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_176 = c53_487_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_176 = c53_487_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_1_145 = c53_488_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_1_144 = c53_488_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_2_113 = c22_54_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_2_112 = c22_54_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_177 = c53_489_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_177 = c53_489_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_1_146 = c53_490_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_1_145 = c53_490_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_2_114 = c32_42_io_out_0; // @[Multiplier.scala 80:35]
  wire  c2_2_113 = c32_42_io_out_1; // @[Multiplier.scala 81:41]
  wire  s_0_178 = c53_491_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_178 = c53_491_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_1_147 = c53_492_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_1_146 = c53_492_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_2_115 = c22_55_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_2_114 = c22_55_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_179 = c53_493_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_179 = c53_493_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_1_148 = c53_494_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_1_147 = c53_494_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_2_116 = c22_56_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_2_115 = c22_56_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_180 = c53_495_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_180 = c53_495_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_1_149 = c53_496_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_1_148 = c53_496_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_2_117 = c22_57_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_2_116 = c22_57_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_181 = c53_497_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_181 = c53_497_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_1_150 = c53_498_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_1_149 = c53_498_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_2_118 = c22_58_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_2_117 = c22_58_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_182 = c53_499_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_182 = c53_499_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_1_151 = c53_500_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_1_150 = c53_500_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_0_183 = c53_501_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_183 = c53_501_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_1_152 = c53_502_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_1_151 = c53_502_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_0_184 = c53_503_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_184 = c53_503_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_1_153 = c53_504_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_1_152 = c53_504_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_0_185 = c53_505_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_185 = c53_505_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_1_154 = c53_506_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_1_153 = c53_506_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_0_186 = c53_507_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_186 = c53_507_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_1_155 = c53_508_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_1_154 = c53_508_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_0_187 = c53_509_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_187 = c53_509_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_1_156 = c53_510_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_1_155 = c53_510_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_0_188 = c53_511_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_188 = c53_511_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_1_157 = c53_512_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_1_156 = c53_512_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_0_189 = c53_513_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_189 = c53_513_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_1_158 = c53_514_io_out_0; // @[Multiplier.scala 88:39]
  wire  c1_1_141 = c53_514_io_out_1; // @[Multiplier.scala 89:41]
  wire  c2_1_157 = c53_514_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_0_190 = c53_515_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_190 = c53_515_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_1_159 = c32_43_io_out_0; // @[Multiplier.scala 80:35]
  wire  c2_1_158 = c32_43_io_out_1; // @[Multiplier.scala 81:41]
  wire  s_0_191 = c53_516_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_191 = c53_516_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_1_160 = c22_59_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_1_159 = c22_59_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_192 = c53_517_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_192 = c53_517_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_1_161 = c22_60_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_1_160 = c22_60_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_193 = c53_518_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_193 = c53_518_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_1_162 = c32_44_io_out_0; // @[Multiplier.scala 80:35]
  wire  c2_1_161 = c32_44_io_out_1; // @[Multiplier.scala 81:41]
  wire  s_0_194 = c53_519_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_194 = c53_519_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_1_163 = c22_61_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_1_162 = c22_61_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_195 = c53_520_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_195 = c53_520_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_1_164 = c22_62_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_1_163 = c22_62_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_196 = c53_521_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_196 = c53_521_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_1_165 = c22_63_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_1_164 = c22_63_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_197 = c53_522_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_197 = c53_522_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_1_166 = c22_64_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_1_165 = c22_64_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_198 = c53_523_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_198 = c53_523_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_0_199 = c53_524_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_199 = c53_524_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_0_200 = c53_525_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_200 = c53_525_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_0_201 = c53_526_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_201 = c53_526_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_0_202 = c53_527_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_202 = c53_527_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_0_203 = c53_528_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_203 = c53_528_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_0_204 = c53_529_io_out_0; // @[Multiplier.scala 88:39]
  wire  c2_0_204 = c53_529_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_0_205 = c53_530_io_out_0; // @[Multiplier.scala 88:39]
  wire  c1_0_189 = c53_530_io_out_1; // @[Multiplier.scala 89:41]
  wire  c2_0_205 = c53_530_io_out_2; // @[Multiplier.scala 90:41]
  wire  s_0_206 = c32_45_io_out_0; // @[Multiplier.scala 80:35]
  wire  c2_0_206 = c32_45_io_out_1; // @[Multiplier.scala 81:41]
  wire  s_0_207 = c22_65_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_207 = c22_65_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_208 = c22_66_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_208 = c22_66_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_209 = c32_46_io_out_0; // @[Multiplier.scala 80:35]
  wire  c2_0_209 = c32_46_io_out_1; // @[Multiplier.scala 81:41]
  wire  s_0_210 = c22_67_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_210 = c22_67_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_211 = c22_68_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_211 = c22_68_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_212 = c22_69_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_212 = c22_69_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_213 = c22_70_io_out_0; // @[Multiplier.scala 75:35]
  reg  r; // @[Reg.scala 16:16]
  reg  r_1; // @[Reg.scala 16:16]
  reg  r_2; // @[Reg.scala 16:16]
  reg  r_3; // @[Reg.scala 16:16]
  reg  r_4; // @[Reg.scala 16:16]
  reg  r_5; // @[Reg.scala 16:16]
  reg  r_6; // @[Reg.scala 16:16]
  reg  r_7; // @[Reg.scala 16:16]
  reg  r_8; // @[Reg.scala 16:16]
  reg  r_9; // @[Reg.scala 16:16]
  reg  r_10; // @[Reg.scala 16:16]
  reg  r_11; // @[Reg.scala 16:16]
  reg  r_12; // @[Reg.scala 16:16]
  reg  r_13; // @[Reg.scala 16:16]
  reg  r_14; // @[Reg.scala 16:16]
  reg  r_15; // @[Reg.scala 16:16]
  reg  r_16; // @[Reg.scala 16:16]
  reg  r_17; // @[Reg.scala 16:16]
  reg  r_18; // @[Reg.scala 16:16]
  reg  r_19; // @[Reg.scala 16:16]
  reg  r_20; // @[Reg.scala 16:16]
  reg  r_21; // @[Reg.scala 16:16]
  reg  r_22; // @[Reg.scala 16:16]
  reg  r_23; // @[Reg.scala 16:16]
  reg  r_24; // @[Reg.scala 16:16]
  reg  r_25; // @[Reg.scala 16:16]
  reg  r_26; // @[Reg.scala 16:16]
  reg  r_27; // @[Reg.scala 16:16]
  reg  r_28; // @[Reg.scala 16:16]
  reg  r_29; // @[Reg.scala 16:16]
  reg  r_30; // @[Reg.scala 16:16]
  reg  r_31; // @[Reg.scala 16:16]
  reg  r_32; // @[Reg.scala 16:16]
  reg  r_33; // @[Reg.scala 16:16]
  reg  r_34; // @[Reg.scala 16:16]
  reg  r_35; // @[Reg.scala 16:16]
  reg  r_36; // @[Reg.scala 16:16]
  reg  r_37; // @[Reg.scala 16:16]
  reg  r_38; // @[Reg.scala 16:16]
  reg  r_39; // @[Reg.scala 16:16]
  reg  r_40; // @[Reg.scala 16:16]
  reg  r_41; // @[Reg.scala 16:16]
  reg  r_42; // @[Reg.scala 16:16]
  reg  r_43; // @[Reg.scala 16:16]
  reg  r_44; // @[Reg.scala 16:16]
  reg  r_45; // @[Reg.scala 16:16]
  reg  r_46; // @[Reg.scala 16:16]
  reg  r_47; // @[Reg.scala 16:16]
  reg  r_48; // @[Reg.scala 16:16]
  reg  r_49; // @[Reg.scala 16:16]
  reg  r_50; // @[Reg.scala 16:16]
  reg  r_51; // @[Reg.scala 16:16]
  reg  r_52; // @[Reg.scala 16:16]
  reg  r_53; // @[Reg.scala 16:16]
  reg  r_54; // @[Reg.scala 16:16]
  reg  r_55; // @[Reg.scala 16:16]
  reg  r_56; // @[Reg.scala 16:16]
  reg  r_57; // @[Reg.scala 16:16]
  reg  r_58; // @[Reg.scala 16:16]
  reg  r_59; // @[Reg.scala 16:16]
  reg  r_60; // @[Reg.scala 16:16]
  reg  r_61; // @[Reg.scala 16:16]
  reg  r_62; // @[Reg.scala 16:16]
  reg  r_63; // @[Reg.scala 16:16]
  reg  r_64; // @[Reg.scala 16:16]
  reg  r_65; // @[Reg.scala 16:16]
  reg  r_66; // @[Reg.scala 16:16]
  reg  r_67; // @[Reg.scala 16:16]
  reg  r_68; // @[Reg.scala 16:16]
  reg  r_69; // @[Reg.scala 16:16]
  reg  r_70; // @[Reg.scala 16:16]
  reg  r_71; // @[Reg.scala 16:16]
  reg  r_72; // @[Reg.scala 16:16]
  reg  r_73; // @[Reg.scala 16:16]
  reg  r_74; // @[Reg.scala 16:16]
  reg  r_75; // @[Reg.scala 16:16]
  reg  r_76; // @[Reg.scala 16:16]
  reg  r_77; // @[Reg.scala 16:16]
  reg  r_78; // @[Reg.scala 16:16]
  reg  r_79; // @[Reg.scala 16:16]
  reg  r_80; // @[Reg.scala 16:16]
  reg  r_81; // @[Reg.scala 16:16]
  reg  r_82; // @[Reg.scala 16:16]
  reg  r_83; // @[Reg.scala 16:16]
  reg  r_84; // @[Reg.scala 16:16]
  reg  r_85; // @[Reg.scala 16:16]
  reg  r_86; // @[Reg.scala 16:16]
  reg  r_87; // @[Reg.scala 16:16]
  reg  r_88; // @[Reg.scala 16:16]
  reg  r_89; // @[Reg.scala 16:16]
  reg  r_90; // @[Reg.scala 16:16]
  reg  r_91; // @[Reg.scala 16:16]
  reg  r_92; // @[Reg.scala 16:16]
  reg  r_93; // @[Reg.scala 16:16]
  reg  r_94; // @[Reg.scala 16:16]
  reg  r_95; // @[Reg.scala 16:16]
  reg  r_96; // @[Reg.scala 16:16]
  reg  r_97; // @[Reg.scala 16:16]
  reg  r_98; // @[Reg.scala 16:16]
  reg  r_99; // @[Reg.scala 16:16]
  reg  r_100; // @[Reg.scala 16:16]
  reg  r_101; // @[Reg.scala 16:16]
  reg  r_102; // @[Reg.scala 16:16]
  reg  r_103; // @[Reg.scala 16:16]
  reg  r_104; // @[Reg.scala 16:16]
  reg  r_105; // @[Reg.scala 16:16]
  reg  r_106; // @[Reg.scala 16:16]
  reg  r_107; // @[Reg.scala 16:16]
  reg  r_108; // @[Reg.scala 16:16]
  reg  r_109; // @[Reg.scala 16:16]
  reg  r_110; // @[Reg.scala 16:16]
  reg  r_111; // @[Reg.scala 16:16]
  reg  r_112; // @[Reg.scala 16:16]
  reg  r_113; // @[Reg.scala 16:16]
  reg  r_114; // @[Reg.scala 16:16]
  reg  r_115; // @[Reg.scala 16:16]
  reg  r_116; // @[Reg.scala 16:16]
  reg  r_117; // @[Reg.scala 16:16]
  reg  r_118; // @[Reg.scala 16:16]
  reg  r_119; // @[Reg.scala 16:16]
  reg  r_120; // @[Reg.scala 16:16]
  reg  r_121; // @[Reg.scala 16:16]
  reg  r_122; // @[Reg.scala 16:16]
  reg  r_123; // @[Reg.scala 16:16]
  reg  r_124; // @[Reg.scala 16:16]
  reg  r_125; // @[Reg.scala 16:16]
  reg  r_126; // @[Reg.scala 16:16]
  reg  r_127; // @[Reg.scala 16:16]
  reg  r_128; // @[Reg.scala 16:16]
  reg  r_129; // @[Reg.scala 16:16]
  reg  r_130; // @[Reg.scala 16:16]
  reg  r_131; // @[Reg.scala 16:16]
  reg  r_132; // @[Reg.scala 16:16]
  reg  r_133; // @[Reg.scala 16:16]
  reg  r_134; // @[Reg.scala 16:16]
  reg  r_135; // @[Reg.scala 16:16]
  reg  r_136; // @[Reg.scala 16:16]
  reg  r_137; // @[Reg.scala 16:16]
  reg  r_138; // @[Reg.scala 16:16]
  reg  r_139; // @[Reg.scala 16:16]
  reg  r_140; // @[Reg.scala 16:16]
  reg  r_141; // @[Reg.scala 16:16]
  reg  r_142; // @[Reg.scala 16:16]
  reg  r_143; // @[Reg.scala 16:16]
  reg  r_144; // @[Reg.scala 16:16]
  reg  r_145; // @[Reg.scala 16:16]
  reg  r_146; // @[Reg.scala 16:16]
  reg  r_147; // @[Reg.scala 16:16]
  reg  r_148; // @[Reg.scala 16:16]
  reg  r_149; // @[Reg.scala 16:16]
  reg  r_150; // @[Reg.scala 16:16]
  reg  r_151; // @[Reg.scala 16:16]
  reg  r_152; // @[Reg.scala 16:16]
  reg  r_153; // @[Reg.scala 16:16]
  reg  r_154; // @[Reg.scala 16:16]
  reg  r_155; // @[Reg.scala 16:16]
  reg  r_156; // @[Reg.scala 16:16]
  reg  r_157; // @[Reg.scala 16:16]
  reg  r_158; // @[Reg.scala 16:16]
  reg  r_159; // @[Reg.scala 16:16]
  reg  r_160; // @[Reg.scala 16:16]
  reg  r_161; // @[Reg.scala 16:16]
  reg  r_162; // @[Reg.scala 16:16]
  reg  r_163; // @[Reg.scala 16:16]
  reg  r_164; // @[Reg.scala 16:16]
  reg  r_165; // @[Reg.scala 16:16]
  reg  r_166; // @[Reg.scala 16:16]
  reg  r_167; // @[Reg.scala 16:16]
  reg  r_168; // @[Reg.scala 16:16]
  reg  r_169; // @[Reg.scala 16:16]
  reg  r_170; // @[Reg.scala 16:16]
  reg  r_171; // @[Reg.scala 16:16]
  reg  r_172; // @[Reg.scala 16:16]
  reg  r_173; // @[Reg.scala 16:16]
  reg  r_174; // @[Reg.scala 16:16]
  reg  r_175; // @[Reg.scala 16:16]
  reg  r_176; // @[Reg.scala 16:16]
  reg  r_177; // @[Reg.scala 16:16]
  reg  r_178; // @[Reg.scala 16:16]
  reg  r_179; // @[Reg.scala 16:16]
  reg  r_180; // @[Reg.scala 16:16]
  reg  r_181; // @[Reg.scala 16:16]
  reg  r_182; // @[Reg.scala 16:16]
  reg  r_183; // @[Reg.scala 16:16]
  reg  r_184; // @[Reg.scala 16:16]
  reg  r_185; // @[Reg.scala 16:16]
  reg  r_186; // @[Reg.scala 16:16]
  reg  r_187; // @[Reg.scala 16:16]
  reg  r_188; // @[Reg.scala 16:16]
  reg  r_189; // @[Reg.scala 16:16]
  reg  r_190; // @[Reg.scala 16:16]
  reg  r_191; // @[Reg.scala 16:16]
  reg  r_192; // @[Reg.scala 16:16]
  reg  r_193; // @[Reg.scala 16:16]
  reg  r_194; // @[Reg.scala 16:16]
  reg  r_195; // @[Reg.scala 16:16]
  reg  r_196; // @[Reg.scala 16:16]
  reg  r_197; // @[Reg.scala 16:16]
  reg  r_198; // @[Reg.scala 16:16]
  reg  r_199; // @[Reg.scala 16:16]
  reg  r_200; // @[Reg.scala 16:16]
  reg  r_201; // @[Reg.scala 16:16]
  reg  r_202; // @[Reg.scala 16:16]
  reg  r_203; // @[Reg.scala 16:16]
  reg  r_204; // @[Reg.scala 16:16]
  reg  r_205; // @[Reg.scala 16:16]
  reg  r_206; // @[Reg.scala 16:16]
  reg  r_207; // @[Reg.scala 16:16]
  reg  r_208; // @[Reg.scala 16:16]
  reg  r_209; // @[Reg.scala 16:16]
  reg  r_210; // @[Reg.scala 16:16]
  reg  r_211; // @[Reg.scala 16:16]
  reg  r_212; // @[Reg.scala 16:16]
  reg  r_213; // @[Reg.scala 16:16]
  reg  r_214; // @[Reg.scala 16:16]
  reg  r_215; // @[Reg.scala 16:16]
  reg  r_216; // @[Reg.scala 16:16]
  reg  r_217; // @[Reg.scala 16:16]
  reg  r_218; // @[Reg.scala 16:16]
  reg  r_219; // @[Reg.scala 16:16]
  reg  r_220; // @[Reg.scala 16:16]
  reg  r_221; // @[Reg.scala 16:16]
  reg  r_222; // @[Reg.scala 16:16]
  reg  r_223; // @[Reg.scala 16:16]
  reg  r_224; // @[Reg.scala 16:16]
  reg  r_225; // @[Reg.scala 16:16]
  reg  r_226; // @[Reg.scala 16:16]
  reg  r_227; // @[Reg.scala 16:16]
  reg  r_228; // @[Reg.scala 16:16]
  reg  r_229; // @[Reg.scala 16:16]
  reg  r_230; // @[Reg.scala 16:16]
  reg  r_231; // @[Reg.scala 16:16]
  reg  r_232; // @[Reg.scala 16:16]
  reg  r_233; // @[Reg.scala 16:16]
  reg  r_234; // @[Reg.scala 16:16]
  reg  r_235; // @[Reg.scala 16:16]
  reg  r_236; // @[Reg.scala 16:16]
  reg  r_237; // @[Reg.scala 16:16]
  reg  r_238; // @[Reg.scala 16:16]
  reg  r_239; // @[Reg.scala 16:16]
  reg  r_240; // @[Reg.scala 16:16]
  reg  r_241; // @[Reg.scala 16:16]
  reg  r_242; // @[Reg.scala 16:16]
  reg  r_243; // @[Reg.scala 16:16]
  reg  r_244; // @[Reg.scala 16:16]
  reg  r_245; // @[Reg.scala 16:16]
  reg  r_246; // @[Reg.scala 16:16]
  reg  r_247; // @[Reg.scala 16:16]
  reg  r_248; // @[Reg.scala 16:16]
  reg  r_249; // @[Reg.scala 16:16]
  reg  r_250; // @[Reg.scala 16:16]
  reg  r_251; // @[Reg.scala 16:16]
  reg  r_252; // @[Reg.scala 16:16]
  reg  r_253; // @[Reg.scala 16:16]
  reg  r_254; // @[Reg.scala 16:16]
  reg  r_255; // @[Reg.scala 16:16]
  reg  r_256; // @[Reg.scala 16:16]
  reg  r_257; // @[Reg.scala 16:16]
  reg  r_258; // @[Reg.scala 16:16]
  reg  r_259; // @[Reg.scala 16:16]
  reg  r_260; // @[Reg.scala 16:16]
  reg  r_261; // @[Reg.scala 16:16]
  reg  r_262; // @[Reg.scala 16:16]
  reg  r_263; // @[Reg.scala 16:16]
  reg  r_264; // @[Reg.scala 16:16]
  reg  r_265; // @[Reg.scala 16:16]
  reg  r_266; // @[Reg.scala 16:16]
  reg  r_267; // @[Reg.scala 16:16]
  reg  r_268; // @[Reg.scala 16:16]
  reg  r_269; // @[Reg.scala 16:16]
  reg  r_270; // @[Reg.scala 16:16]
  reg  r_271; // @[Reg.scala 16:16]
  reg  r_272; // @[Reg.scala 16:16]
  reg  r_273; // @[Reg.scala 16:16]
  reg  r_274; // @[Reg.scala 16:16]
  reg  r_275; // @[Reg.scala 16:16]
  reg  r_276; // @[Reg.scala 16:16]
  reg  r_277; // @[Reg.scala 16:16]
  reg  r_278; // @[Reg.scala 16:16]
  reg  r_279; // @[Reg.scala 16:16]
  reg  r_280; // @[Reg.scala 16:16]
  reg  r_281; // @[Reg.scala 16:16]
  reg  r_282; // @[Reg.scala 16:16]
  reg  r_283; // @[Reg.scala 16:16]
  reg  r_284; // @[Reg.scala 16:16]
  reg  r_285; // @[Reg.scala 16:16]
  reg  r_286; // @[Reg.scala 16:16]
  reg  r_287; // @[Reg.scala 16:16]
  reg  r_288; // @[Reg.scala 16:16]
  reg  r_289; // @[Reg.scala 16:16]
  reg  r_290; // @[Reg.scala 16:16]
  reg  r_291; // @[Reg.scala 16:16]
  reg  r_292; // @[Reg.scala 16:16]
  reg  r_293; // @[Reg.scala 16:16]
  reg  r_294; // @[Reg.scala 16:16]
  reg  r_295; // @[Reg.scala 16:16]
  reg  r_296; // @[Reg.scala 16:16]
  reg  r_297; // @[Reg.scala 16:16]
  reg  r_298; // @[Reg.scala 16:16]
  reg  r_299; // @[Reg.scala 16:16]
  reg  r_300; // @[Reg.scala 16:16]
  reg  r_301; // @[Reg.scala 16:16]
  reg  r_302; // @[Reg.scala 16:16]
  reg  r_303; // @[Reg.scala 16:16]
  reg  r_304; // @[Reg.scala 16:16]
  reg  r_305; // @[Reg.scala 16:16]
  reg  r_306; // @[Reg.scala 16:16]
  reg  r_307; // @[Reg.scala 16:16]
  reg  r_308; // @[Reg.scala 16:16]
  reg  r_309; // @[Reg.scala 16:16]
  reg  r_310; // @[Reg.scala 16:16]
  reg  r_311; // @[Reg.scala 16:16]
  reg  r_312; // @[Reg.scala 16:16]
  reg  r_313; // @[Reg.scala 16:16]
  reg  r_314; // @[Reg.scala 16:16]
  reg  r_315; // @[Reg.scala 16:16]
  reg  r_316; // @[Reg.scala 16:16]
  reg  r_317; // @[Reg.scala 16:16]
  reg  r_318; // @[Reg.scala 16:16]
  reg  r_319; // @[Reg.scala 16:16]
  reg  r_320; // @[Reg.scala 16:16]
  reg  r_321; // @[Reg.scala 16:16]
  reg  r_322; // @[Reg.scala 16:16]
  reg  r_323; // @[Reg.scala 16:16]
  reg  r_324; // @[Reg.scala 16:16]
  reg  r_325; // @[Reg.scala 16:16]
  reg  r_326; // @[Reg.scala 16:16]
  reg  r_327; // @[Reg.scala 16:16]
  reg  r_328; // @[Reg.scala 16:16]
  reg  r_329; // @[Reg.scala 16:16]
  reg  r_330; // @[Reg.scala 16:16]
  reg  r_331; // @[Reg.scala 16:16]
  reg  r_332; // @[Reg.scala 16:16]
  reg  r_333; // @[Reg.scala 16:16]
  reg  r_334; // @[Reg.scala 16:16]
  reg  r_335; // @[Reg.scala 16:16]
  reg  r_336; // @[Reg.scala 16:16]
  reg  r_337; // @[Reg.scala 16:16]
  reg  r_338; // @[Reg.scala 16:16]
  reg  r_339; // @[Reg.scala 16:16]
  reg  r_340; // @[Reg.scala 16:16]
  reg  r_341; // @[Reg.scala 16:16]
  reg  r_342; // @[Reg.scala 16:16]
  reg  r_343; // @[Reg.scala 16:16]
  reg  r_344; // @[Reg.scala 16:16]
  reg  r_345; // @[Reg.scala 16:16]
  reg  r_346; // @[Reg.scala 16:16]
  reg  r_347; // @[Reg.scala 16:16]
  reg  r_348; // @[Reg.scala 16:16]
  reg  r_349; // @[Reg.scala 16:16]
  reg  r_350; // @[Reg.scala 16:16]
  reg  r_351; // @[Reg.scala 16:16]
  reg  r_352; // @[Reg.scala 16:16]
  reg  r_353; // @[Reg.scala 16:16]
  reg  r_354; // @[Reg.scala 16:16]
  reg  r_355; // @[Reg.scala 16:16]
  reg  r_356; // @[Reg.scala 16:16]
  reg  r_357; // @[Reg.scala 16:16]
  reg  r_358; // @[Reg.scala 16:16]
  reg  r_359; // @[Reg.scala 16:16]
  reg  r_360; // @[Reg.scala 16:16]
  reg  r_361; // @[Reg.scala 16:16]
  reg  r_362; // @[Reg.scala 16:16]
  reg  r_363; // @[Reg.scala 16:16]
  reg  r_364; // @[Reg.scala 16:16]
  reg  r_365; // @[Reg.scala 16:16]
  reg  r_366; // @[Reg.scala 16:16]
  reg  r_367; // @[Reg.scala 16:16]
  reg  r_368; // @[Reg.scala 16:16]
  reg  r_369; // @[Reg.scala 16:16]
  reg  r_370; // @[Reg.scala 16:16]
  reg  r_371; // @[Reg.scala 16:16]
  reg  r_372; // @[Reg.scala 16:16]
  reg  r_373; // @[Reg.scala 16:16]
  reg  r_374; // @[Reg.scala 16:16]
  reg  r_375; // @[Reg.scala 16:16]
  reg  r_376; // @[Reg.scala 16:16]
  reg  r_377; // @[Reg.scala 16:16]
  reg  r_378; // @[Reg.scala 16:16]
  reg  r_379; // @[Reg.scala 16:16]
  reg  r_380; // @[Reg.scala 16:16]
  reg  r_381; // @[Reg.scala 16:16]
  reg  r_382; // @[Reg.scala 16:16]
  reg  r_383; // @[Reg.scala 16:16]
  reg  r_384; // @[Reg.scala 16:16]
  reg  r_385; // @[Reg.scala 16:16]
  reg  r_386; // @[Reg.scala 16:16]
  reg  r_387; // @[Reg.scala 16:16]
  reg  r_388; // @[Reg.scala 16:16]
  reg  r_389; // @[Reg.scala 16:16]
  reg  r_390; // @[Reg.scala 16:16]
  reg  r_391; // @[Reg.scala 16:16]
  reg  r_392; // @[Reg.scala 16:16]
  reg  r_393; // @[Reg.scala 16:16]
  reg  r_394; // @[Reg.scala 16:16]
  reg  r_395; // @[Reg.scala 16:16]
  reg  r_396; // @[Reg.scala 16:16]
  reg  r_397; // @[Reg.scala 16:16]
  reg  r_398; // @[Reg.scala 16:16]
  reg  r_399; // @[Reg.scala 16:16]
  reg  r_400; // @[Reg.scala 16:16]
  reg  r_401; // @[Reg.scala 16:16]
  reg  r_402; // @[Reg.scala 16:16]
  reg  r_403; // @[Reg.scala 16:16]
  reg  r_404; // @[Reg.scala 16:16]
  reg  r_405; // @[Reg.scala 16:16]
  reg  r_406; // @[Reg.scala 16:16]
  reg  r_407; // @[Reg.scala 16:16]
  reg  r_408; // @[Reg.scala 16:16]
  reg  r_409; // @[Reg.scala 16:16]
  reg  r_410; // @[Reg.scala 16:16]
  reg  r_411; // @[Reg.scala 16:16]
  reg  r_412; // @[Reg.scala 16:16]
  reg  r_413; // @[Reg.scala 16:16]
  reg  r_414; // @[Reg.scala 16:16]
  reg  r_415; // @[Reg.scala 16:16]
  reg  r_416; // @[Reg.scala 16:16]
  reg  r_417; // @[Reg.scala 16:16]
  reg  r_418; // @[Reg.scala 16:16]
  reg  r_419; // @[Reg.scala 16:16]
  reg  r_420; // @[Reg.scala 16:16]
  reg  r_421; // @[Reg.scala 16:16]
  reg  r_422; // @[Reg.scala 16:16]
  reg  r_423; // @[Reg.scala 16:16]
  reg  r_424; // @[Reg.scala 16:16]
  reg  r_425; // @[Reg.scala 16:16]
  reg  r_426; // @[Reg.scala 16:16]
  reg  r_427; // @[Reg.scala 16:16]
  reg  r_428; // @[Reg.scala 16:16]
  reg  r_429; // @[Reg.scala 16:16]
  reg  r_430; // @[Reg.scala 16:16]
  reg  r_431; // @[Reg.scala 16:16]
  reg  r_432; // @[Reg.scala 16:16]
  reg  r_433; // @[Reg.scala 16:16]
  reg  r_434; // @[Reg.scala 16:16]
  reg  r_435; // @[Reg.scala 16:16]
  reg  r_436; // @[Reg.scala 16:16]
  reg  r_437; // @[Reg.scala 16:16]
  reg  r_438; // @[Reg.scala 16:16]
  reg  r_439; // @[Reg.scala 16:16]
  reg  r_440; // @[Reg.scala 16:16]
  reg  r_441; // @[Reg.scala 16:16]
  reg  r_442; // @[Reg.scala 16:16]
  reg  r_443; // @[Reg.scala 16:16]
  reg  r_444; // @[Reg.scala 16:16]
  reg  r_445; // @[Reg.scala 16:16]
  reg  r_446; // @[Reg.scala 16:16]
  reg  r_447; // @[Reg.scala 16:16]
  reg  r_448; // @[Reg.scala 16:16]
  reg  r_449; // @[Reg.scala 16:16]
  reg  r_450; // @[Reg.scala 16:16]
  reg  r_451; // @[Reg.scala 16:16]
  reg  r_452; // @[Reg.scala 16:16]
  reg  r_453; // @[Reg.scala 16:16]
  reg  r_454; // @[Reg.scala 16:16]
  reg  r_455; // @[Reg.scala 16:16]
  reg  r_456; // @[Reg.scala 16:16]
  reg  r_457; // @[Reg.scala 16:16]
  reg  r_458; // @[Reg.scala 16:16]
  reg  r_459; // @[Reg.scala 16:16]
  reg  r_460; // @[Reg.scala 16:16]
  reg  r_461; // @[Reg.scala 16:16]
  reg  r_462; // @[Reg.scala 16:16]
  reg  r_463; // @[Reg.scala 16:16]
  reg  r_464; // @[Reg.scala 16:16]
  reg  r_465; // @[Reg.scala 16:16]
  reg  r_466; // @[Reg.scala 16:16]
  reg  r_467; // @[Reg.scala 16:16]
  reg  r_468; // @[Reg.scala 16:16]
  reg  r_469; // @[Reg.scala 16:16]
  reg  r_470; // @[Reg.scala 16:16]
  reg  r_471; // @[Reg.scala 16:16]
  reg  r_472; // @[Reg.scala 16:16]
  reg  r_473; // @[Reg.scala 16:16]
  reg  r_474; // @[Reg.scala 16:16]
  reg  r_475; // @[Reg.scala 16:16]
  reg  r_476; // @[Reg.scala 16:16]
  reg  r_477; // @[Reg.scala 16:16]
  reg  r_478; // @[Reg.scala 16:16]
  reg  r_479; // @[Reg.scala 16:16]
  reg  r_480; // @[Reg.scala 16:16]
  reg  r_481; // @[Reg.scala 16:16]
  reg  r_482; // @[Reg.scala 16:16]
  reg  r_483; // @[Reg.scala 16:16]
  reg  r_484; // @[Reg.scala 16:16]
  reg  r_485; // @[Reg.scala 16:16]
  reg  r_486; // @[Reg.scala 16:16]
  reg  r_487; // @[Reg.scala 16:16]
  reg  r_488; // @[Reg.scala 16:16]
  reg  r_489; // @[Reg.scala 16:16]
  wire  s_0_214 = c22_71_io_out_0; // @[Multiplier.scala 75:35]
  wire  s_0_320 = c22_122_io_out_0; // @[Multiplier.scala 75:35]
  wire  s_0_425 = c22_176_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_425 = c22_176_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_426 = c22_177_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_426 = c22_177_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_427 = c22_178_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_427 = c22_178_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_428 = c22_179_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_428 = c22_179_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_429 = c22_180_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_429 = c22_180_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_430 = c22_181_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_430 = c22_181_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_431 = c22_182_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_431 = c22_182_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_432 = c22_183_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_432 = c22_183_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_433 = c22_184_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_433 = c22_184_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_434 = c22_185_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_434 = c22_185_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_435 = c22_186_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_435 = c22_186_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_436 = c22_187_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_436 = c22_187_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_437 = c22_188_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_437 = c22_188_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_438 = c22_189_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_438 = c22_189_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_439 = c22_190_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_439 = c22_190_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_440 = c22_191_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_440 = c22_191_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_441 = c22_192_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_441 = c22_192_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_442 = c22_193_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_442 = c22_193_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_443 = c22_194_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_443 = c22_194_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_444 = c22_195_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_444 = c22_195_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_445 = c22_196_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_445 = c22_196_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_446 = c22_197_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_446 = c22_197_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_447 = c22_198_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_447 = c22_198_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_448 = c22_199_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_448 = c22_199_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_449 = c22_200_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_449 = c22_200_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_450 = c22_201_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_450 = c22_201_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_451 = c22_202_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_451 = c22_202_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_452 = c22_203_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_452 = c22_203_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_453 = c22_204_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_453 = c22_204_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_454 = c22_205_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_454 = c22_205_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_455 = c22_206_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_455 = c22_206_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_456 = c22_207_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_456 = c22_207_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_457 = c22_208_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_457 = c22_208_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_458 = c22_209_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_458 = c22_209_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_459 = c22_210_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_459 = c22_210_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_460 = c22_211_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_460 = c22_211_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_461 = c22_212_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_461 = c22_212_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_462 = c22_213_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_462 = c22_213_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_463 = c22_214_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_463 = c22_214_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_464 = c22_215_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_464 = c22_215_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_465 = c22_216_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_465 = c22_216_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_466 = c22_217_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_466 = c22_217_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_467 = c22_218_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_467 = c22_218_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_468 = c22_219_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_468 = c22_219_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_469 = c22_220_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_469 = c22_220_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_470 = c22_221_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_470 = c22_221_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_471 = c22_222_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_471 = c22_222_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_472 = c22_223_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_472 = c22_223_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_473 = c22_224_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_473 = c22_224_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_474 = c22_225_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_474 = c22_225_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_475 = c22_226_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_475 = c22_226_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_476 = c22_227_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_476 = c22_227_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_477 = c22_228_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_477 = c22_228_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_478 = c22_229_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_478 = c22_229_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_479 = c22_230_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_479 = c22_230_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_480 = c22_231_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_480 = c22_231_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_481 = c22_232_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_481 = c22_232_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_482 = c32_68_io_out_0; // @[Multiplier.scala 80:35]
  wire  c2_0_482 = c32_68_io_out_1; // @[Multiplier.scala 81:41]
  wire  s_0_483 = c22_233_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_483 = c22_233_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_484 = c22_234_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_484 = c22_234_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_485 = c22_235_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_485 = c22_235_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_486 = c22_236_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_486 = c22_236_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_487 = c22_237_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_487 = c22_237_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_488 = c22_238_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_488 = c22_238_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_489 = c22_239_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_489 = c22_239_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_490 = c22_240_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_490 = c22_240_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_491 = c22_241_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_491 = c22_241_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_492 = c22_242_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_492 = c22_242_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_493 = c22_243_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_493 = c22_243_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_494 = c22_244_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_494 = c22_244_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_495 = c22_245_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_495 = c22_245_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_496 = c22_246_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_496 = c22_246_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_497 = c22_247_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_497 = c22_247_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_498 = c32_69_io_out_0; // @[Multiplier.scala 80:35]
  wire  c2_0_498 = c32_69_io_out_1; // @[Multiplier.scala 81:41]
  wire  s_0_499 = c22_248_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_499 = c22_248_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_500 = c22_249_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_500 = c22_249_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_501 = c22_250_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_501 = c22_250_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_502 = c22_251_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_502 = c22_251_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_503 = c22_252_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_503 = c22_252_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_504 = c22_253_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_504 = c22_253_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_505 = c22_254_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_505 = c22_254_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_506 = c22_255_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_506 = c22_255_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_507 = c22_256_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_507 = c22_256_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_508 = c22_257_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_508 = c22_257_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_509 = c22_258_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_509 = c22_258_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_510 = c22_259_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_510 = c22_259_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_511 = c22_260_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_511 = c22_260_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_512 = c22_261_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_512 = c22_261_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_513 = c22_262_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_513 = c22_262_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_514 = c22_263_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_514 = c22_263_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_515 = c22_264_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_515 = c22_264_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_516 = c22_265_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_516 = c22_265_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_517 = c22_266_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_517 = c22_266_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_518 = c22_267_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_518 = c22_267_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_519 = c22_268_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_519 = c22_268_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_520 = c22_269_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_520 = c22_269_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_521 = c22_270_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_521 = c22_270_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_522 = c22_271_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_522 = c22_271_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_523 = c22_272_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_523 = c22_272_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_524 = c22_273_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_524 = c22_273_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_525 = c22_274_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_525 = c22_274_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_526 = c22_275_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_526 = c22_275_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_527 = c22_276_io_out_0; // @[Multiplier.scala 75:35]
  wire  c2_0_527 = c22_276_io_out_1; // @[Multiplier.scala 76:41]
  wire  s_0_528 = c22_277_io_out_0; // @[Multiplier.scala 75:35]
  wire [5:0] sum_lo_lo_lo_lo = {s_0_426,s_0_425,s_0_320,s_0_214,r_1,r}; // @[Cat.scala 31:58]
  wire [12:0] sum_lo_lo_lo = {s_0_433,s_0_432,s_0_431,s_0_430,s_0_429,s_0_428,s_0_427,sum_lo_lo_lo_lo}; // @[Cat.scala 31:58]
  wire [6:0] sum_lo_lo_hi_lo = {s_0_440,s_0_439,s_0_438,s_0_437,s_0_436,s_0_435,s_0_434}; // @[Cat.scala 31:58]
  wire [26:0] sum_lo_lo = {s_0_447,s_0_446,s_0_445,s_0_444,s_0_443,s_0_442,s_0_441,sum_lo_lo_hi_lo,sum_lo_lo_lo}; // @[Cat.scala 31:58]
  wire [5:0] sum_lo_hi_lo_lo = {s_0_453,s_0_452,s_0_451,s_0_450,s_0_449,s_0_448}; // @[Cat.scala 31:58]
  wire [12:0] sum_lo_hi_lo = {s_0_460,s_0_459,s_0_458,s_0_457,s_0_456,s_0_455,s_0_454,sum_lo_hi_lo_lo}; // @[Cat.scala 31:58]
  wire [6:0] sum_lo_hi_hi_lo = {s_0_467,s_0_466,s_0_465,s_0_464,s_0_463,s_0_462,s_0_461}; // @[Cat.scala 31:58]
  wire [53:0] sum_lo = {s_0_474,s_0_473,s_0_472,s_0_471,s_0_470,s_0_469,s_0_468,sum_lo_hi_hi_lo,sum_lo_hi_lo,sum_lo_lo}; // @[Cat.scala 31:58]
  wire [5:0] sum_hi_lo_lo_lo = {s_0_480,s_0_479,s_0_478,s_0_477,s_0_476,s_0_475}; // @[Cat.scala 31:58]
  wire [12:0] sum_hi_lo_lo = {s_0_487,s_0_486,s_0_485,s_0_484,s_0_483,s_0_482,s_0_481,sum_hi_lo_lo_lo}; // @[Cat.scala 31:58]
  wire [6:0] sum_hi_lo_hi_lo = {s_0_494,s_0_493,s_0_492,s_0_491,s_0_490,s_0_489,s_0_488}; // @[Cat.scala 31:58]
  wire [26:0] sum_hi_lo = {s_0_501,s_0_500,s_0_499,s_0_498,s_0_497,s_0_496,s_0_495,sum_hi_lo_hi_lo,sum_hi_lo_lo}; // @[Cat.scala 31:58]
  wire [5:0] sum_hi_hi_lo_lo = {s_0_507,s_0_506,s_0_505,s_0_504,s_0_503,s_0_502}; // @[Cat.scala 31:58]
  wire [12:0] sum_hi_hi_lo = {s_0_514,s_0_513,s_0_512,s_0_511,s_0_510,s_0_509,s_0_508,sum_hi_hi_lo_lo}; // @[Cat.scala 31:58]
  wire [6:0] sum_hi_hi_hi_lo = {s_0_521,s_0_520,s_0_519,s_0_518,s_0_517,s_0_516,s_0_515}; // @[Cat.scala 31:58]
  wire [53:0] sum_hi = {s_0_528,s_0_527,s_0_526,s_0_525,s_0_524,s_0_523,s_0_522,sum_hi_hi_hi_lo,sum_hi_hi_lo,sum_hi_lo}; // @[Cat.scala 31:58]
  wire [107:0] sum = {sum_hi,sum_lo}; // @[Cat.scala 31:58]
  wire [5:0] carry_lo_lo_lo_lo = {c2_0_430,c2_0_429,c2_0_428,c2_0_427,c2_0_426,c2_0_425}; // @[Cat.scala 31:58]
  wire [11:0] carry_lo_lo_lo = {c2_0_436,c2_0_435,c2_0_434,c2_0_433,c2_0_432,c2_0_431,carry_lo_lo_lo_lo}; // @[Cat.scala 31:58]
  wire [5:0] carry_lo_lo_hi_lo = {c2_0_442,c2_0_441,c2_0_440,c2_0_439,c2_0_438,c2_0_437}; // @[Cat.scala 31:58]
  wire [24:0] carry_lo_lo = {c2_0_449,c2_0_448,c2_0_447,c2_0_446,c2_0_445,c2_0_444,c2_0_443,carry_lo_lo_hi_lo,
    carry_lo_lo_lo}; // @[Cat.scala 31:58]
  wire [5:0] carry_lo_hi_lo_lo = {c2_0_455,c2_0_454,c2_0_453,c2_0_452,c2_0_451,c2_0_450}; // @[Cat.scala 31:58]
  wire [12:0] carry_lo_hi_lo = {c2_0_462,c2_0_461,c2_0_460,c2_0_459,c2_0_458,c2_0_457,c2_0_456,carry_lo_hi_lo_lo}; // @[Cat.scala 31:58]
  wire [5:0] carry_lo_hi_hi_lo = {c2_0_468,c2_0_467,c2_0_466,c2_0_465,c2_0_464,c2_0_463}; // @[Cat.scala 31:58]
  wire [50:0] carry_lo = {c2_0_475,c2_0_474,c2_0_473,c2_0_472,c2_0_471,c2_0_470,c2_0_469,carry_lo_hi_hi_lo,
    carry_lo_hi_lo,carry_lo_lo}; // @[Cat.scala 31:58]
  wire [5:0] carry_hi_lo_lo_lo = {c2_0_481,c2_0_480,c2_0_479,c2_0_478,c2_0_477,c2_0_476}; // @[Cat.scala 31:58]
  wire [12:0] carry_hi_lo_lo = {c2_0_488,c2_0_487,c2_0_486,c2_0_485,c2_0_484,c2_0_483,c2_0_482,carry_hi_lo_lo_lo}; // @[Cat.scala 31:58]
  wire [5:0] carry_hi_lo_hi_lo = {c2_0_494,c2_0_493,c2_0_492,c2_0_491,c2_0_490,c2_0_489}; // @[Cat.scala 31:58]
  wire [25:0] carry_hi_lo = {c2_0_501,c2_0_500,c2_0_499,c2_0_498,c2_0_497,c2_0_496,c2_0_495,carry_hi_lo_hi_lo,
    carry_hi_lo_lo}; // @[Cat.scala 31:58]
  wire [5:0] carry_hi_hi_lo_lo = {c2_0_507,c2_0_506,c2_0_505,c2_0_504,c2_0_503,c2_0_502}; // @[Cat.scala 31:58]
  wire [12:0] carry_hi_hi_lo = {c2_0_514,c2_0_513,c2_0_512,c2_0_511,c2_0_510,c2_0_509,c2_0_508,carry_hi_hi_lo_lo}; // @[Cat.scala 31:58]
  wire [5:0] carry_hi_hi_hi_lo = {c2_0_520,c2_0_519,c2_0_518,c2_0_517,c2_0_516,c2_0_515}; // @[Cat.scala 31:58]
  wire [51:0] carry_hi = {c2_0_527,c2_0_526,c2_0_525,c2_0_524,c2_0_523,c2_0_522,c2_0_521,carry_hi_hi_hi_lo,
    carry_hi_hi_lo,carry_hi_lo}; // @[Cat.scala 31:58]
  wire [107:0] carry_1 = {carry_hi,carry_lo,5'h0}; // @[Cat.scala 31:58]
  C22 c22 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_io_in_0),
    .io_in_1(c22_io_in_1),
    .io_out_0(c22_io_out_0),
    .io_out_1(c22_io_out_1)
  );
  C22 c22_1 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_1_io_in_0),
    .io_in_1(c22_1_io_in_1),
    .io_out_0(c22_1_io_out_0),
    .io_out_1(c22_1_io_out_1)
  );
  C32 c32 ( // @[Multiplier.scala 78:25]
    .io_in_0(c32_io_in_0),
    .io_in_1(c32_io_in_1),
    .io_in_2(c32_io_in_2),
    .io_out_0(c32_io_out_0),
    .io_out_1(c32_io_out_1)
  );
  C32 c32_1 ( // @[Multiplier.scala 78:25]
    .io_in_0(c32_1_io_in_0),
    .io_in_1(c32_1_io_in_1),
    .io_in_2(c32_1_io_in_2),
    .io_out_0(c32_1_io_out_0),
    .io_out_1(c32_1_io_out_1)
  );
  C53 c53 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_io_in_0),
    .io_in_1(c53_io_in_1),
    .io_in_2(c53_io_in_2),
    .io_in_3(c53_io_in_3),
    .io_in_4(c53_io_in_4),
    .io_out_0(c53_io_out_0),
    .io_out_1(c53_io_out_1),
    .io_out_2(c53_io_out_2)
  );
  C53 c53_1 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_1_io_in_0),
    .io_in_1(c53_1_io_in_1),
    .io_in_2(c53_1_io_in_2),
    .io_in_3(c53_1_io_in_3),
    .io_in_4(c53_1_io_in_4),
    .io_out_0(c53_1_io_out_0),
    .io_out_1(c53_1_io_out_1),
    .io_out_2(c53_1_io_out_2)
  );
  C53 c53_2 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_2_io_in_0),
    .io_in_1(c53_2_io_in_1),
    .io_in_2(c53_2_io_in_2),
    .io_in_3(c53_2_io_in_3),
    .io_in_4(c53_2_io_in_4),
    .io_out_0(c53_2_io_out_0),
    .io_out_1(c53_2_io_out_1),
    .io_out_2(c53_2_io_out_2)
  );
  C53 c53_3 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_3_io_in_0),
    .io_in_1(c53_3_io_in_1),
    .io_in_2(c53_3_io_in_2),
    .io_in_3(c53_3_io_in_3),
    .io_in_4(c53_3_io_in_4),
    .io_out_0(c53_3_io_out_0),
    .io_out_1(c53_3_io_out_1),
    .io_out_2(c53_3_io_out_2)
  );
  C53 c53_4 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_4_io_in_0),
    .io_in_1(c53_4_io_in_1),
    .io_in_2(c53_4_io_in_2),
    .io_in_3(c53_4_io_in_3),
    .io_in_4(c53_4_io_in_4),
    .io_out_0(c53_4_io_out_0),
    .io_out_1(c53_4_io_out_1),
    .io_out_2(c53_4_io_out_2)
  );
  C22 c22_2 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_2_io_in_0),
    .io_in_1(c22_2_io_in_1),
    .io_out_0(c22_2_io_out_0),
    .io_out_1(c22_2_io_out_1)
  );
  C53 c53_5 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_5_io_in_0),
    .io_in_1(c53_5_io_in_1),
    .io_in_2(c53_5_io_in_2),
    .io_in_3(c53_5_io_in_3),
    .io_in_4(c53_5_io_in_4),
    .io_out_0(c53_5_io_out_0),
    .io_out_1(c53_5_io_out_1),
    .io_out_2(c53_5_io_out_2)
  );
  C22 c22_3 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_3_io_in_0),
    .io_in_1(c22_3_io_in_1),
    .io_out_0(c22_3_io_out_0),
    .io_out_1(c22_3_io_out_1)
  );
  C53 c53_6 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_6_io_in_0),
    .io_in_1(c53_6_io_in_1),
    .io_in_2(c53_6_io_in_2),
    .io_in_3(c53_6_io_in_3),
    .io_in_4(c53_6_io_in_4),
    .io_out_0(c53_6_io_out_0),
    .io_out_1(c53_6_io_out_1),
    .io_out_2(c53_6_io_out_2)
  );
  C32 c32_2 ( // @[Multiplier.scala 78:25]
    .io_in_0(c32_2_io_in_0),
    .io_in_1(c32_2_io_in_1),
    .io_in_2(c32_2_io_in_2),
    .io_out_0(c32_2_io_out_0),
    .io_out_1(c32_2_io_out_1)
  );
  C53 c53_7 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_7_io_in_0),
    .io_in_1(c53_7_io_in_1),
    .io_in_2(c53_7_io_in_2),
    .io_in_3(c53_7_io_in_3),
    .io_in_4(c53_7_io_in_4),
    .io_out_0(c53_7_io_out_0),
    .io_out_1(c53_7_io_out_1),
    .io_out_2(c53_7_io_out_2)
  );
  C32 c32_3 ( // @[Multiplier.scala 78:25]
    .io_in_0(c32_3_io_in_0),
    .io_in_1(c32_3_io_in_1),
    .io_in_2(c32_3_io_in_2),
    .io_out_0(c32_3_io_out_0),
    .io_out_1(c32_3_io_out_1)
  );
  C53 c53_8 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_8_io_in_0),
    .io_in_1(c53_8_io_in_1),
    .io_in_2(c53_8_io_in_2),
    .io_in_3(c53_8_io_in_3),
    .io_in_4(c53_8_io_in_4),
    .io_out_0(c53_8_io_out_0),
    .io_out_1(c53_8_io_out_1),
    .io_out_2(c53_8_io_out_2)
  );
  C53 c53_9 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_9_io_in_0),
    .io_in_1(c53_9_io_in_1),
    .io_in_2(c53_9_io_in_2),
    .io_in_3(c53_9_io_in_3),
    .io_in_4(c53_9_io_in_4),
    .io_out_0(c53_9_io_out_0),
    .io_out_1(c53_9_io_out_1),
    .io_out_2(c53_9_io_out_2)
  );
  C53 c53_10 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_10_io_in_0),
    .io_in_1(c53_10_io_in_1),
    .io_in_2(c53_10_io_in_2),
    .io_in_3(c53_10_io_in_3),
    .io_in_4(c53_10_io_in_4),
    .io_out_0(c53_10_io_out_0),
    .io_out_1(c53_10_io_out_1),
    .io_out_2(c53_10_io_out_2)
  );
  C53 c53_11 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_11_io_in_0),
    .io_in_1(c53_11_io_in_1),
    .io_in_2(c53_11_io_in_2),
    .io_in_3(c53_11_io_in_3),
    .io_in_4(c53_11_io_in_4),
    .io_out_0(c53_11_io_out_0),
    .io_out_1(c53_11_io_out_1),
    .io_out_2(c53_11_io_out_2)
  );
  C53 c53_12 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_12_io_in_0),
    .io_in_1(c53_12_io_in_1),
    .io_in_2(c53_12_io_in_2),
    .io_in_3(c53_12_io_in_3),
    .io_in_4(c53_12_io_in_4),
    .io_out_0(c53_12_io_out_0),
    .io_out_1(c53_12_io_out_1),
    .io_out_2(c53_12_io_out_2)
  );
  C53 c53_13 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_13_io_in_0),
    .io_in_1(c53_13_io_in_1),
    .io_in_2(c53_13_io_in_2),
    .io_in_3(c53_13_io_in_3),
    .io_in_4(c53_13_io_in_4),
    .io_out_0(c53_13_io_out_0),
    .io_out_1(c53_13_io_out_1),
    .io_out_2(c53_13_io_out_2)
  );
  C53 c53_14 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_14_io_in_0),
    .io_in_1(c53_14_io_in_1),
    .io_in_2(c53_14_io_in_2),
    .io_in_3(c53_14_io_in_3),
    .io_in_4(c53_14_io_in_4),
    .io_out_0(c53_14_io_out_0),
    .io_out_1(c53_14_io_out_1),
    .io_out_2(c53_14_io_out_2)
  );
  C53 c53_15 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_15_io_in_0),
    .io_in_1(c53_15_io_in_1),
    .io_in_2(c53_15_io_in_2),
    .io_in_3(c53_15_io_in_3),
    .io_in_4(c53_15_io_in_4),
    .io_out_0(c53_15_io_out_0),
    .io_out_1(c53_15_io_out_1),
    .io_out_2(c53_15_io_out_2)
  );
  C53 c53_16 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_16_io_in_0),
    .io_in_1(c53_16_io_in_1),
    .io_in_2(c53_16_io_in_2),
    .io_in_3(c53_16_io_in_3),
    .io_in_4(c53_16_io_in_4),
    .io_out_0(c53_16_io_out_0),
    .io_out_1(c53_16_io_out_1),
    .io_out_2(c53_16_io_out_2)
  );
  C53 c53_17 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_17_io_in_0),
    .io_in_1(c53_17_io_in_1),
    .io_in_2(c53_17_io_in_2),
    .io_in_3(c53_17_io_in_3),
    .io_in_4(c53_17_io_in_4),
    .io_out_0(c53_17_io_out_0),
    .io_out_1(c53_17_io_out_1),
    .io_out_2(c53_17_io_out_2)
  );
  C22 c22_4 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_4_io_in_0),
    .io_in_1(c22_4_io_in_1),
    .io_out_0(c22_4_io_out_0),
    .io_out_1(c22_4_io_out_1)
  );
  C53 c53_18 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_18_io_in_0),
    .io_in_1(c53_18_io_in_1),
    .io_in_2(c53_18_io_in_2),
    .io_in_3(c53_18_io_in_3),
    .io_in_4(c53_18_io_in_4),
    .io_out_0(c53_18_io_out_0),
    .io_out_1(c53_18_io_out_1),
    .io_out_2(c53_18_io_out_2)
  );
  C53 c53_19 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_19_io_in_0),
    .io_in_1(c53_19_io_in_1),
    .io_in_2(c53_19_io_in_2),
    .io_in_3(c53_19_io_in_3),
    .io_in_4(c53_19_io_in_4),
    .io_out_0(c53_19_io_out_0),
    .io_out_1(c53_19_io_out_1),
    .io_out_2(c53_19_io_out_2)
  );
  C22 c22_5 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_5_io_in_0),
    .io_in_1(c22_5_io_in_1),
    .io_out_0(c22_5_io_out_0),
    .io_out_1(c22_5_io_out_1)
  );
  C53 c53_20 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_20_io_in_0),
    .io_in_1(c53_20_io_in_1),
    .io_in_2(c53_20_io_in_2),
    .io_in_3(c53_20_io_in_3),
    .io_in_4(c53_20_io_in_4),
    .io_out_0(c53_20_io_out_0),
    .io_out_1(c53_20_io_out_1),
    .io_out_2(c53_20_io_out_2)
  );
  C53 c53_21 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_21_io_in_0),
    .io_in_1(c53_21_io_in_1),
    .io_in_2(c53_21_io_in_2),
    .io_in_3(c53_21_io_in_3),
    .io_in_4(c53_21_io_in_4),
    .io_out_0(c53_21_io_out_0),
    .io_out_1(c53_21_io_out_1),
    .io_out_2(c53_21_io_out_2)
  );
  C32 c32_4 ( // @[Multiplier.scala 78:25]
    .io_in_0(c32_4_io_in_0),
    .io_in_1(c32_4_io_in_1),
    .io_in_2(c32_4_io_in_2),
    .io_out_0(c32_4_io_out_0),
    .io_out_1(c32_4_io_out_1)
  );
  C53 c53_22 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_22_io_in_0),
    .io_in_1(c53_22_io_in_1),
    .io_in_2(c53_22_io_in_2),
    .io_in_3(c53_22_io_in_3),
    .io_in_4(c53_22_io_in_4),
    .io_out_0(c53_22_io_out_0),
    .io_out_1(c53_22_io_out_1),
    .io_out_2(c53_22_io_out_2)
  );
  C53 c53_23 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_23_io_in_0),
    .io_in_1(c53_23_io_in_1),
    .io_in_2(c53_23_io_in_2),
    .io_in_3(c53_23_io_in_3),
    .io_in_4(c53_23_io_in_4),
    .io_out_0(c53_23_io_out_0),
    .io_out_1(c53_23_io_out_1),
    .io_out_2(c53_23_io_out_2)
  );
  C32 c32_5 ( // @[Multiplier.scala 78:25]
    .io_in_0(c32_5_io_in_0),
    .io_in_1(c32_5_io_in_1),
    .io_in_2(c32_5_io_in_2),
    .io_out_0(c32_5_io_out_0),
    .io_out_1(c32_5_io_out_1)
  );
  C53 c53_24 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_24_io_in_0),
    .io_in_1(c53_24_io_in_1),
    .io_in_2(c53_24_io_in_2),
    .io_in_3(c53_24_io_in_3),
    .io_in_4(c53_24_io_in_4),
    .io_out_0(c53_24_io_out_0),
    .io_out_1(c53_24_io_out_1),
    .io_out_2(c53_24_io_out_2)
  );
  C53 c53_25 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_25_io_in_0),
    .io_in_1(c53_25_io_in_1),
    .io_in_2(c53_25_io_in_2),
    .io_in_3(c53_25_io_in_3),
    .io_in_4(c53_25_io_in_4),
    .io_out_0(c53_25_io_out_0),
    .io_out_1(c53_25_io_out_1),
    .io_out_2(c53_25_io_out_2)
  );
  C53 c53_26 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_26_io_in_0),
    .io_in_1(c53_26_io_in_1),
    .io_in_2(c53_26_io_in_2),
    .io_in_3(c53_26_io_in_3),
    .io_in_4(c53_26_io_in_4),
    .io_out_0(c53_26_io_out_0),
    .io_out_1(c53_26_io_out_1),
    .io_out_2(c53_26_io_out_2)
  );
  C53 c53_27 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_27_io_in_0),
    .io_in_1(c53_27_io_in_1),
    .io_in_2(c53_27_io_in_2),
    .io_in_3(c53_27_io_in_3),
    .io_in_4(c53_27_io_in_4),
    .io_out_0(c53_27_io_out_0),
    .io_out_1(c53_27_io_out_1),
    .io_out_2(c53_27_io_out_2)
  );
  C53 c53_28 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_28_io_in_0),
    .io_in_1(c53_28_io_in_1),
    .io_in_2(c53_28_io_in_2),
    .io_in_3(c53_28_io_in_3),
    .io_in_4(c53_28_io_in_4),
    .io_out_0(c53_28_io_out_0),
    .io_out_1(c53_28_io_out_1),
    .io_out_2(c53_28_io_out_2)
  );
  C53 c53_29 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_29_io_in_0),
    .io_in_1(c53_29_io_in_1),
    .io_in_2(c53_29_io_in_2),
    .io_in_3(c53_29_io_in_3),
    .io_in_4(c53_29_io_in_4),
    .io_out_0(c53_29_io_out_0),
    .io_out_1(c53_29_io_out_1),
    .io_out_2(c53_29_io_out_2)
  );
  C53 c53_30 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_30_io_in_0),
    .io_in_1(c53_30_io_in_1),
    .io_in_2(c53_30_io_in_2),
    .io_in_3(c53_30_io_in_3),
    .io_in_4(c53_30_io_in_4),
    .io_out_0(c53_30_io_out_0),
    .io_out_1(c53_30_io_out_1),
    .io_out_2(c53_30_io_out_2)
  );
  C53 c53_31 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_31_io_in_0),
    .io_in_1(c53_31_io_in_1),
    .io_in_2(c53_31_io_in_2),
    .io_in_3(c53_31_io_in_3),
    .io_in_4(c53_31_io_in_4),
    .io_out_0(c53_31_io_out_0),
    .io_out_1(c53_31_io_out_1),
    .io_out_2(c53_31_io_out_2)
  );
  C53 c53_32 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_32_io_in_0),
    .io_in_1(c53_32_io_in_1),
    .io_in_2(c53_32_io_in_2),
    .io_in_3(c53_32_io_in_3),
    .io_in_4(c53_32_io_in_4),
    .io_out_0(c53_32_io_out_0),
    .io_out_1(c53_32_io_out_1),
    .io_out_2(c53_32_io_out_2)
  );
  C53 c53_33 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_33_io_in_0),
    .io_in_1(c53_33_io_in_1),
    .io_in_2(c53_33_io_in_2),
    .io_in_3(c53_33_io_in_3),
    .io_in_4(c53_33_io_in_4),
    .io_out_0(c53_33_io_out_0),
    .io_out_1(c53_33_io_out_1),
    .io_out_2(c53_33_io_out_2)
  );
  C53 c53_34 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_34_io_in_0),
    .io_in_1(c53_34_io_in_1),
    .io_in_2(c53_34_io_in_2),
    .io_in_3(c53_34_io_in_3),
    .io_in_4(c53_34_io_in_4),
    .io_out_0(c53_34_io_out_0),
    .io_out_1(c53_34_io_out_1),
    .io_out_2(c53_34_io_out_2)
  );
  C53 c53_35 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_35_io_in_0),
    .io_in_1(c53_35_io_in_1),
    .io_in_2(c53_35_io_in_2),
    .io_in_3(c53_35_io_in_3),
    .io_in_4(c53_35_io_in_4),
    .io_out_0(c53_35_io_out_0),
    .io_out_1(c53_35_io_out_1),
    .io_out_2(c53_35_io_out_2)
  );
  C53 c53_36 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_36_io_in_0),
    .io_in_1(c53_36_io_in_1),
    .io_in_2(c53_36_io_in_2),
    .io_in_3(c53_36_io_in_3),
    .io_in_4(c53_36_io_in_4),
    .io_out_0(c53_36_io_out_0),
    .io_out_1(c53_36_io_out_1),
    .io_out_2(c53_36_io_out_2)
  );
  C53 c53_37 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_37_io_in_0),
    .io_in_1(c53_37_io_in_1),
    .io_in_2(c53_37_io_in_2),
    .io_in_3(c53_37_io_in_3),
    .io_in_4(c53_37_io_in_4),
    .io_out_0(c53_37_io_out_0),
    .io_out_1(c53_37_io_out_1),
    .io_out_2(c53_37_io_out_2)
  );
  C53 c53_38 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_38_io_in_0),
    .io_in_1(c53_38_io_in_1),
    .io_in_2(c53_38_io_in_2),
    .io_in_3(c53_38_io_in_3),
    .io_in_4(c53_38_io_in_4),
    .io_out_0(c53_38_io_out_0),
    .io_out_1(c53_38_io_out_1),
    .io_out_2(c53_38_io_out_2)
  );
  C22 c22_6 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_6_io_in_0),
    .io_in_1(c22_6_io_in_1),
    .io_out_0(c22_6_io_out_0),
    .io_out_1(c22_6_io_out_1)
  );
  C53 c53_39 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_39_io_in_0),
    .io_in_1(c53_39_io_in_1),
    .io_in_2(c53_39_io_in_2),
    .io_in_3(c53_39_io_in_3),
    .io_in_4(c53_39_io_in_4),
    .io_out_0(c53_39_io_out_0),
    .io_out_1(c53_39_io_out_1),
    .io_out_2(c53_39_io_out_2)
  );
  C53 c53_40 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_40_io_in_0),
    .io_in_1(c53_40_io_in_1),
    .io_in_2(c53_40_io_in_2),
    .io_in_3(c53_40_io_in_3),
    .io_in_4(c53_40_io_in_4),
    .io_out_0(c53_40_io_out_0),
    .io_out_1(c53_40_io_out_1),
    .io_out_2(c53_40_io_out_2)
  );
  C53 c53_41 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_41_io_in_0),
    .io_in_1(c53_41_io_in_1),
    .io_in_2(c53_41_io_in_2),
    .io_in_3(c53_41_io_in_3),
    .io_in_4(c53_41_io_in_4),
    .io_out_0(c53_41_io_out_0),
    .io_out_1(c53_41_io_out_1),
    .io_out_2(c53_41_io_out_2)
  );
  C22 c22_7 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_7_io_in_0),
    .io_in_1(c22_7_io_in_1),
    .io_out_0(c22_7_io_out_0),
    .io_out_1(c22_7_io_out_1)
  );
  C53 c53_42 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_42_io_in_0),
    .io_in_1(c53_42_io_in_1),
    .io_in_2(c53_42_io_in_2),
    .io_in_3(c53_42_io_in_3),
    .io_in_4(c53_42_io_in_4),
    .io_out_0(c53_42_io_out_0),
    .io_out_1(c53_42_io_out_1),
    .io_out_2(c53_42_io_out_2)
  );
  C53 c53_43 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_43_io_in_0),
    .io_in_1(c53_43_io_in_1),
    .io_in_2(c53_43_io_in_2),
    .io_in_3(c53_43_io_in_3),
    .io_in_4(c53_43_io_in_4),
    .io_out_0(c53_43_io_out_0),
    .io_out_1(c53_43_io_out_1),
    .io_out_2(c53_43_io_out_2)
  );
  C53 c53_44 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_44_io_in_0),
    .io_in_1(c53_44_io_in_1),
    .io_in_2(c53_44_io_in_2),
    .io_in_3(c53_44_io_in_3),
    .io_in_4(c53_44_io_in_4),
    .io_out_0(c53_44_io_out_0),
    .io_out_1(c53_44_io_out_1),
    .io_out_2(c53_44_io_out_2)
  );
  C32 c32_6 ( // @[Multiplier.scala 78:25]
    .io_in_0(c32_6_io_in_0),
    .io_in_1(c32_6_io_in_1),
    .io_in_2(c32_6_io_in_2),
    .io_out_0(c32_6_io_out_0),
    .io_out_1(c32_6_io_out_1)
  );
  C53 c53_45 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_45_io_in_0),
    .io_in_1(c53_45_io_in_1),
    .io_in_2(c53_45_io_in_2),
    .io_in_3(c53_45_io_in_3),
    .io_in_4(c53_45_io_in_4),
    .io_out_0(c53_45_io_out_0),
    .io_out_1(c53_45_io_out_1),
    .io_out_2(c53_45_io_out_2)
  );
  C53 c53_46 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_46_io_in_0),
    .io_in_1(c53_46_io_in_1),
    .io_in_2(c53_46_io_in_2),
    .io_in_3(c53_46_io_in_3),
    .io_in_4(c53_46_io_in_4),
    .io_out_0(c53_46_io_out_0),
    .io_out_1(c53_46_io_out_1),
    .io_out_2(c53_46_io_out_2)
  );
  C53 c53_47 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_47_io_in_0),
    .io_in_1(c53_47_io_in_1),
    .io_in_2(c53_47_io_in_2),
    .io_in_3(c53_47_io_in_3),
    .io_in_4(c53_47_io_in_4),
    .io_out_0(c53_47_io_out_0),
    .io_out_1(c53_47_io_out_1),
    .io_out_2(c53_47_io_out_2)
  );
  C32 c32_7 ( // @[Multiplier.scala 78:25]
    .io_in_0(c32_7_io_in_0),
    .io_in_1(c32_7_io_in_1),
    .io_in_2(c32_7_io_in_2),
    .io_out_0(c32_7_io_out_0),
    .io_out_1(c32_7_io_out_1)
  );
  C53 c53_48 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_48_io_in_0),
    .io_in_1(c53_48_io_in_1),
    .io_in_2(c53_48_io_in_2),
    .io_in_3(c53_48_io_in_3),
    .io_in_4(c53_48_io_in_4),
    .io_out_0(c53_48_io_out_0),
    .io_out_1(c53_48_io_out_1),
    .io_out_2(c53_48_io_out_2)
  );
  C53 c53_49 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_49_io_in_0),
    .io_in_1(c53_49_io_in_1),
    .io_in_2(c53_49_io_in_2),
    .io_in_3(c53_49_io_in_3),
    .io_in_4(c53_49_io_in_4),
    .io_out_0(c53_49_io_out_0),
    .io_out_1(c53_49_io_out_1),
    .io_out_2(c53_49_io_out_2)
  );
  C53 c53_50 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_50_io_in_0),
    .io_in_1(c53_50_io_in_1),
    .io_in_2(c53_50_io_in_2),
    .io_in_3(c53_50_io_in_3),
    .io_in_4(c53_50_io_in_4),
    .io_out_0(c53_50_io_out_0),
    .io_out_1(c53_50_io_out_1),
    .io_out_2(c53_50_io_out_2)
  );
  C53 c53_51 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_51_io_in_0),
    .io_in_1(c53_51_io_in_1),
    .io_in_2(c53_51_io_in_2),
    .io_in_3(c53_51_io_in_3),
    .io_in_4(c53_51_io_in_4),
    .io_out_0(c53_51_io_out_0),
    .io_out_1(c53_51_io_out_1),
    .io_out_2(c53_51_io_out_2)
  );
  C53 c53_52 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_52_io_in_0),
    .io_in_1(c53_52_io_in_1),
    .io_in_2(c53_52_io_in_2),
    .io_in_3(c53_52_io_in_3),
    .io_in_4(c53_52_io_in_4),
    .io_out_0(c53_52_io_out_0),
    .io_out_1(c53_52_io_out_1),
    .io_out_2(c53_52_io_out_2)
  );
  C53 c53_53 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_53_io_in_0),
    .io_in_1(c53_53_io_in_1),
    .io_in_2(c53_53_io_in_2),
    .io_in_3(c53_53_io_in_3),
    .io_in_4(c53_53_io_in_4),
    .io_out_0(c53_53_io_out_0),
    .io_out_1(c53_53_io_out_1),
    .io_out_2(c53_53_io_out_2)
  );
  C53 c53_54 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_54_io_in_0),
    .io_in_1(c53_54_io_in_1),
    .io_in_2(c53_54_io_in_2),
    .io_in_3(c53_54_io_in_3),
    .io_in_4(c53_54_io_in_4),
    .io_out_0(c53_54_io_out_0),
    .io_out_1(c53_54_io_out_1),
    .io_out_2(c53_54_io_out_2)
  );
  C53 c53_55 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_55_io_in_0),
    .io_in_1(c53_55_io_in_1),
    .io_in_2(c53_55_io_in_2),
    .io_in_3(c53_55_io_in_3),
    .io_in_4(c53_55_io_in_4),
    .io_out_0(c53_55_io_out_0),
    .io_out_1(c53_55_io_out_1),
    .io_out_2(c53_55_io_out_2)
  );
  C53 c53_56 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_56_io_in_0),
    .io_in_1(c53_56_io_in_1),
    .io_in_2(c53_56_io_in_2),
    .io_in_3(c53_56_io_in_3),
    .io_in_4(c53_56_io_in_4),
    .io_out_0(c53_56_io_out_0),
    .io_out_1(c53_56_io_out_1),
    .io_out_2(c53_56_io_out_2)
  );
  C53 c53_57 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_57_io_in_0),
    .io_in_1(c53_57_io_in_1),
    .io_in_2(c53_57_io_in_2),
    .io_in_3(c53_57_io_in_3),
    .io_in_4(c53_57_io_in_4),
    .io_out_0(c53_57_io_out_0),
    .io_out_1(c53_57_io_out_1),
    .io_out_2(c53_57_io_out_2)
  );
  C53 c53_58 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_58_io_in_0),
    .io_in_1(c53_58_io_in_1),
    .io_in_2(c53_58_io_in_2),
    .io_in_3(c53_58_io_in_3),
    .io_in_4(c53_58_io_in_4),
    .io_out_0(c53_58_io_out_0),
    .io_out_1(c53_58_io_out_1),
    .io_out_2(c53_58_io_out_2)
  );
  C53 c53_59 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_59_io_in_0),
    .io_in_1(c53_59_io_in_1),
    .io_in_2(c53_59_io_in_2),
    .io_in_3(c53_59_io_in_3),
    .io_in_4(c53_59_io_in_4),
    .io_out_0(c53_59_io_out_0),
    .io_out_1(c53_59_io_out_1),
    .io_out_2(c53_59_io_out_2)
  );
  C53 c53_60 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_60_io_in_0),
    .io_in_1(c53_60_io_in_1),
    .io_in_2(c53_60_io_in_2),
    .io_in_3(c53_60_io_in_3),
    .io_in_4(c53_60_io_in_4),
    .io_out_0(c53_60_io_out_0),
    .io_out_1(c53_60_io_out_1),
    .io_out_2(c53_60_io_out_2)
  );
  C53 c53_61 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_61_io_in_0),
    .io_in_1(c53_61_io_in_1),
    .io_in_2(c53_61_io_in_2),
    .io_in_3(c53_61_io_in_3),
    .io_in_4(c53_61_io_in_4),
    .io_out_0(c53_61_io_out_0),
    .io_out_1(c53_61_io_out_1),
    .io_out_2(c53_61_io_out_2)
  );
  C53 c53_62 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_62_io_in_0),
    .io_in_1(c53_62_io_in_1),
    .io_in_2(c53_62_io_in_2),
    .io_in_3(c53_62_io_in_3),
    .io_in_4(c53_62_io_in_4),
    .io_out_0(c53_62_io_out_0),
    .io_out_1(c53_62_io_out_1),
    .io_out_2(c53_62_io_out_2)
  );
  C53 c53_63 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_63_io_in_0),
    .io_in_1(c53_63_io_in_1),
    .io_in_2(c53_63_io_in_2),
    .io_in_3(c53_63_io_in_3),
    .io_in_4(c53_63_io_in_4),
    .io_out_0(c53_63_io_out_0),
    .io_out_1(c53_63_io_out_1),
    .io_out_2(c53_63_io_out_2)
  );
  C53 c53_64 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_64_io_in_0),
    .io_in_1(c53_64_io_in_1),
    .io_in_2(c53_64_io_in_2),
    .io_in_3(c53_64_io_in_3),
    .io_in_4(c53_64_io_in_4),
    .io_out_0(c53_64_io_out_0),
    .io_out_1(c53_64_io_out_1),
    .io_out_2(c53_64_io_out_2)
  );
  C53 c53_65 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_65_io_in_0),
    .io_in_1(c53_65_io_in_1),
    .io_in_2(c53_65_io_in_2),
    .io_in_3(c53_65_io_in_3),
    .io_in_4(c53_65_io_in_4),
    .io_out_0(c53_65_io_out_0),
    .io_out_1(c53_65_io_out_1),
    .io_out_2(c53_65_io_out_2)
  );
  C53 c53_66 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_66_io_in_0),
    .io_in_1(c53_66_io_in_1),
    .io_in_2(c53_66_io_in_2),
    .io_in_3(c53_66_io_in_3),
    .io_in_4(c53_66_io_in_4),
    .io_out_0(c53_66_io_out_0),
    .io_out_1(c53_66_io_out_1),
    .io_out_2(c53_66_io_out_2)
  );
  C53 c53_67 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_67_io_in_0),
    .io_in_1(c53_67_io_in_1),
    .io_in_2(c53_67_io_in_2),
    .io_in_3(c53_67_io_in_3),
    .io_in_4(c53_67_io_in_4),
    .io_out_0(c53_67_io_out_0),
    .io_out_1(c53_67_io_out_1),
    .io_out_2(c53_67_io_out_2)
  );
  C22 c22_8 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_8_io_in_0),
    .io_in_1(c22_8_io_in_1),
    .io_out_0(c22_8_io_out_0),
    .io_out_1(c22_8_io_out_1)
  );
  C53 c53_68 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_68_io_in_0),
    .io_in_1(c53_68_io_in_1),
    .io_in_2(c53_68_io_in_2),
    .io_in_3(c53_68_io_in_3),
    .io_in_4(c53_68_io_in_4),
    .io_out_0(c53_68_io_out_0),
    .io_out_1(c53_68_io_out_1),
    .io_out_2(c53_68_io_out_2)
  );
  C53 c53_69 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_69_io_in_0),
    .io_in_1(c53_69_io_in_1),
    .io_in_2(c53_69_io_in_2),
    .io_in_3(c53_69_io_in_3),
    .io_in_4(c53_69_io_in_4),
    .io_out_0(c53_69_io_out_0),
    .io_out_1(c53_69_io_out_1),
    .io_out_2(c53_69_io_out_2)
  );
  C53 c53_70 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_70_io_in_0),
    .io_in_1(c53_70_io_in_1),
    .io_in_2(c53_70_io_in_2),
    .io_in_3(c53_70_io_in_3),
    .io_in_4(c53_70_io_in_4),
    .io_out_0(c53_70_io_out_0),
    .io_out_1(c53_70_io_out_1),
    .io_out_2(c53_70_io_out_2)
  );
  C53 c53_71 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_71_io_in_0),
    .io_in_1(c53_71_io_in_1),
    .io_in_2(c53_71_io_in_2),
    .io_in_3(c53_71_io_in_3),
    .io_in_4(c53_71_io_in_4),
    .io_out_0(c53_71_io_out_0),
    .io_out_1(c53_71_io_out_1),
    .io_out_2(c53_71_io_out_2)
  );
  C22 c22_9 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_9_io_in_0),
    .io_in_1(c22_9_io_in_1),
    .io_out_0(c22_9_io_out_0),
    .io_out_1(c22_9_io_out_1)
  );
  C53 c53_72 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_72_io_in_0),
    .io_in_1(c53_72_io_in_1),
    .io_in_2(c53_72_io_in_2),
    .io_in_3(c53_72_io_in_3),
    .io_in_4(c53_72_io_in_4),
    .io_out_0(c53_72_io_out_0),
    .io_out_1(c53_72_io_out_1),
    .io_out_2(c53_72_io_out_2)
  );
  C53 c53_73 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_73_io_in_0),
    .io_in_1(c53_73_io_in_1),
    .io_in_2(c53_73_io_in_2),
    .io_in_3(c53_73_io_in_3),
    .io_in_4(c53_73_io_in_4),
    .io_out_0(c53_73_io_out_0),
    .io_out_1(c53_73_io_out_1),
    .io_out_2(c53_73_io_out_2)
  );
  C53 c53_74 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_74_io_in_0),
    .io_in_1(c53_74_io_in_1),
    .io_in_2(c53_74_io_in_2),
    .io_in_3(c53_74_io_in_3),
    .io_in_4(c53_74_io_in_4),
    .io_out_0(c53_74_io_out_0),
    .io_out_1(c53_74_io_out_1),
    .io_out_2(c53_74_io_out_2)
  );
  C53 c53_75 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_75_io_in_0),
    .io_in_1(c53_75_io_in_1),
    .io_in_2(c53_75_io_in_2),
    .io_in_3(c53_75_io_in_3),
    .io_in_4(c53_75_io_in_4),
    .io_out_0(c53_75_io_out_0),
    .io_out_1(c53_75_io_out_1),
    .io_out_2(c53_75_io_out_2)
  );
  C32 c32_8 ( // @[Multiplier.scala 78:25]
    .io_in_0(c32_8_io_in_0),
    .io_in_1(c32_8_io_in_1),
    .io_in_2(c32_8_io_in_2),
    .io_out_0(c32_8_io_out_0),
    .io_out_1(c32_8_io_out_1)
  );
  C53 c53_76 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_76_io_in_0),
    .io_in_1(c53_76_io_in_1),
    .io_in_2(c53_76_io_in_2),
    .io_in_3(c53_76_io_in_3),
    .io_in_4(c53_76_io_in_4),
    .io_out_0(c53_76_io_out_0),
    .io_out_1(c53_76_io_out_1),
    .io_out_2(c53_76_io_out_2)
  );
  C53 c53_77 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_77_io_in_0),
    .io_in_1(c53_77_io_in_1),
    .io_in_2(c53_77_io_in_2),
    .io_in_3(c53_77_io_in_3),
    .io_in_4(c53_77_io_in_4),
    .io_out_0(c53_77_io_out_0),
    .io_out_1(c53_77_io_out_1),
    .io_out_2(c53_77_io_out_2)
  );
  C53 c53_78 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_78_io_in_0),
    .io_in_1(c53_78_io_in_1),
    .io_in_2(c53_78_io_in_2),
    .io_in_3(c53_78_io_in_3),
    .io_in_4(c53_78_io_in_4),
    .io_out_0(c53_78_io_out_0),
    .io_out_1(c53_78_io_out_1),
    .io_out_2(c53_78_io_out_2)
  );
  C53 c53_79 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_79_io_in_0),
    .io_in_1(c53_79_io_in_1),
    .io_in_2(c53_79_io_in_2),
    .io_in_3(c53_79_io_in_3),
    .io_in_4(c53_79_io_in_4),
    .io_out_0(c53_79_io_out_0),
    .io_out_1(c53_79_io_out_1),
    .io_out_2(c53_79_io_out_2)
  );
  C32 c32_9 ( // @[Multiplier.scala 78:25]
    .io_in_0(c32_9_io_in_0),
    .io_in_1(c32_9_io_in_1),
    .io_in_2(c32_9_io_in_2),
    .io_out_0(c32_9_io_out_0),
    .io_out_1(c32_9_io_out_1)
  );
  C53 c53_80 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_80_io_in_0),
    .io_in_1(c53_80_io_in_1),
    .io_in_2(c53_80_io_in_2),
    .io_in_3(c53_80_io_in_3),
    .io_in_4(c53_80_io_in_4),
    .io_out_0(c53_80_io_out_0),
    .io_out_1(c53_80_io_out_1),
    .io_out_2(c53_80_io_out_2)
  );
  C53 c53_81 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_81_io_in_0),
    .io_in_1(c53_81_io_in_1),
    .io_in_2(c53_81_io_in_2),
    .io_in_3(c53_81_io_in_3),
    .io_in_4(c53_81_io_in_4),
    .io_out_0(c53_81_io_out_0),
    .io_out_1(c53_81_io_out_1),
    .io_out_2(c53_81_io_out_2)
  );
  C53 c53_82 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_82_io_in_0),
    .io_in_1(c53_82_io_in_1),
    .io_in_2(c53_82_io_in_2),
    .io_in_3(c53_82_io_in_3),
    .io_in_4(c53_82_io_in_4),
    .io_out_0(c53_82_io_out_0),
    .io_out_1(c53_82_io_out_1),
    .io_out_2(c53_82_io_out_2)
  );
  C53 c53_83 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_83_io_in_0),
    .io_in_1(c53_83_io_in_1),
    .io_in_2(c53_83_io_in_2),
    .io_in_3(c53_83_io_in_3),
    .io_in_4(c53_83_io_in_4),
    .io_out_0(c53_83_io_out_0),
    .io_out_1(c53_83_io_out_1),
    .io_out_2(c53_83_io_out_2)
  );
  C53 c53_84 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_84_io_in_0),
    .io_in_1(c53_84_io_in_1),
    .io_in_2(c53_84_io_in_2),
    .io_in_3(c53_84_io_in_3),
    .io_in_4(c53_84_io_in_4),
    .io_out_0(c53_84_io_out_0),
    .io_out_1(c53_84_io_out_1),
    .io_out_2(c53_84_io_out_2)
  );
  C53 c53_85 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_85_io_in_0),
    .io_in_1(c53_85_io_in_1),
    .io_in_2(c53_85_io_in_2),
    .io_in_3(c53_85_io_in_3),
    .io_in_4(c53_85_io_in_4),
    .io_out_0(c53_85_io_out_0),
    .io_out_1(c53_85_io_out_1),
    .io_out_2(c53_85_io_out_2)
  );
  C53 c53_86 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_86_io_in_0),
    .io_in_1(c53_86_io_in_1),
    .io_in_2(c53_86_io_in_2),
    .io_in_3(c53_86_io_in_3),
    .io_in_4(c53_86_io_in_4),
    .io_out_0(c53_86_io_out_0),
    .io_out_1(c53_86_io_out_1),
    .io_out_2(c53_86_io_out_2)
  );
  C53 c53_87 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_87_io_in_0),
    .io_in_1(c53_87_io_in_1),
    .io_in_2(c53_87_io_in_2),
    .io_in_3(c53_87_io_in_3),
    .io_in_4(c53_87_io_in_4),
    .io_out_0(c53_87_io_out_0),
    .io_out_1(c53_87_io_out_1),
    .io_out_2(c53_87_io_out_2)
  );
  C53 c53_88 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_88_io_in_0),
    .io_in_1(c53_88_io_in_1),
    .io_in_2(c53_88_io_in_2),
    .io_in_3(c53_88_io_in_3),
    .io_in_4(c53_88_io_in_4),
    .io_out_0(c53_88_io_out_0),
    .io_out_1(c53_88_io_out_1),
    .io_out_2(c53_88_io_out_2)
  );
  C53 c53_89 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_89_io_in_0),
    .io_in_1(c53_89_io_in_1),
    .io_in_2(c53_89_io_in_2),
    .io_in_3(c53_89_io_in_3),
    .io_in_4(c53_89_io_in_4),
    .io_out_0(c53_89_io_out_0),
    .io_out_1(c53_89_io_out_1),
    .io_out_2(c53_89_io_out_2)
  );
  C53 c53_90 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_90_io_in_0),
    .io_in_1(c53_90_io_in_1),
    .io_in_2(c53_90_io_in_2),
    .io_in_3(c53_90_io_in_3),
    .io_in_4(c53_90_io_in_4),
    .io_out_0(c53_90_io_out_0),
    .io_out_1(c53_90_io_out_1),
    .io_out_2(c53_90_io_out_2)
  );
  C53 c53_91 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_91_io_in_0),
    .io_in_1(c53_91_io_in_1),
    .io_in_2(c53_91_io_in_2),
    .io_in_3(c53_91_io_in_3),
    .io_in_4(c53_91_io_in_4),
    .io_out_0(c53_91_io_out_0),
    .io_out_1(c53_91_io_out_1),
    .io_out_2(c53_91_io_out_2)
  );
  C53 c53_92 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_92_io_in_0),
    .io_in_1(c53_92_io_in_1),
    .io_in_2(c53_92_io_in_2),
    .io_in_3(c53_92_io_in_3),
    .io_in_4(c53_92_io_in_4),
    .io_out_0(c53_92_io_out_0),
    .io_out_1(c53_92_io_out_1),
    .io_out_2(c53_92_io_out_2)
  );
  C53 c53_93 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_93_io_in_0),
    .io_in_1(c53_93_io_in_1),
    .io_in_2(c53_93_io_in_2),
    .io_in_3(c53_93_io_in_3),
    .io_in_4(c53_93_io_in_4),
    .io_out_0(c53_93_io_out_0),
    .io_out_1(c53_93_io_out_1),
    .io_out_2(c53_93_io_out_2)
  );
  C53 c53_94 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_94_io_in_0),
    .io_in_1(c53_94_io_in_1),
    .io_in_2(c53_94_io_in_2),
    .io_in_3(c53_94_io_in_3),
    .io_in_4(c53_94_io_in_4),
    .io_out_0(c53_94_io_out_0),
    .io_out_1(c53_94_io_out_1),
    .io_out_2(c53_94_io_out_2)
  );
  C53 c53_95 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_95_io_in_0),
    .io_in_1(c53_95_io_in_1),
    .io_in_2(c53_95_io_in_2),
    .io_in_3(c53_95_io_in_3),
    .io_in_4(c53_95_io_in_4),
    .io_out_0(c53_95_io_out_0),
    .io_out_1(c53_95_io_out_1),
    .io_out_2(c53_95_io_out_2)
  );
  C53 c53_96 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_96_io_in_0),
    .io_in_1(c53_96_io_in_1),
    .io_in_2(c53_96_io_in_2),
    .io_in_3(c53_96_io_in_3),
    .io_in_4(c53_96_io_in_4),
    .io_out_0(c53_96_io_out_0),
    .io_out_1(c53_96_io_out_1),
    .io_out_2(c53_96_io_out_2)
  );
  C53 c53_97 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_97_io_in_0),
    .io_in_1(c53_97_io_in_1),
    .io_in_2(c53_97_io_in_2),
    .io_in_3(c53_97_io_in_3),
    .io_in_4(c53_97_io_in_4),
    .io_out_0(c53_97_io_out_0),
    .io_out_1(c53_97_io_out_1),
    .io_out_2(c53_97_io_out_2)
  );
  C53 c53_98 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_98_io_in_0),
    .io_in_1(c53_98_io_in_1),
    .io_in_2(c53_98_io_in_2),
    .io_in_3(c53_98_io_in_3),
    .io_in_4(c53_98_io_in_4),
    .io_out_0(c53_98_io_out_0),
    .io_out_1(c53_98_io_out_1),
    .io_out_2(c53_98_io_out_2)
  );
  C53 c53_99 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_99_io_in_0),
    .io_in_1(c53_99_io_in_1),
    .io_in_2(c53_99_io_in_2),
    .io_in_3(c53_99_io_in_3),
    .io_in_4(c53_99_io_in_4),
    .io_out_0(c53_99_io_out_0),
    .io_out_1(c53_99_io_out_1),
    .io_out_2(c53_99_io_out_2)
  );
  C53 c53_100 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_100_io_in_0),
    .io_in_1(c53_100_io_in_1),
    .io_in_2(c53_100_io_in_2),
    .io_in_3(c53_100_io_in_3),
    .io_in_4(c53_100_io_in_4),
    .io_out_0(c53_100_io_out_0),
    .io_out_1(c53_100_io_out_1),
    .io_out_2(c53_100_io_out_2)
  );
  C53 c53_101 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_101_io_in_0),
    .io_in_1(c53_101_io_in_1),
    .io_in_2(c53_101_io_in_2),
    .io_in_3(c53_101_io_in_3),
    .io_in_4(c53_101_io_in_4),
    .io_out_0(c53_101_io_out_0),
    .io_out_1(c53_101_io_out_1),
    .io_out_2(c53_101_io_out_2)
  );
  C53 c53_102 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_102_io_in_0),
    .io_in_1(c53_102_io_in_1),
    .io_in_2(c53_102_io_in_2),
    .io_in_3(c53_102_io_in_3),
    .io_in_4(c53_102_io_in_4),
    .io_out_0(c53_102_io_out_0),
    .io_out_1(c53_102_io_out_1),
    .io_out_2(c53_102_io_out_2)
  );
  C53 c53_103 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_103_io_in_0),
    .io_in_1(c53_103_io_in_1),
    .io_in_2(c53_103_io_in_2),
    .io_in_3(c53_103_io_in_3),
    .io_in_4(c53_103_io_in_4),
    .io_out_0(c53_103_io_out_0),
    .io_out_1(c53_103_io_out_1),
    .io_out_2(c53_103_io_out_2)
  );
  C53 c53_104 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_104_io_in_0),
    .io_in_1(c53_104_io_in_1),
    .io_in_2(c53_104_io_in_2),
    .io_in_3(c53_104_io_in_3),
    .io_in_4(c53_104_io_in_4),
    .io_out_0(c53_104_io_out_0),
    .io_out_1(c53_104_io_out_1),
    .io_out_2(c53_104_io_out_2)
  );
  C22 c22_10 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_10_io_in_0),
    .io_in_1(c22_10_io_in_1),
    .io_out_0(c22_10_io_out_0),
    .io_out_1(c22_10_io_out_1)
  );
  C53 c53_105 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_105_io_in_0),
    .io_in_1(c53_105_io_in_1),
    .io_in_2(c53_105_io_in_2),
    .io_in_3(c53_105_io_in_3),
    .io_in_4(c53_105_io_in_4),
    .io_out_0(c53_105_io_out_0),
    .io_out_1(c53_105_io_out_1),
    .io_out_2(c53_105_io_out_2)
  );
  C53 c53_106 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_106_io_in_0),
    .io_in_1(c53_106_io_in_1),
    .io_in_2(c53_106_io_in_2),
    .io_in_3(c53_106_io_in_3),
    .io_in_4(c53_106_io_in_4),
    .io_out_0(c53_106_io_out_0),
    .io_out_1(c53_106_io_out_1),
    .io_out_2(c53_106_io_out_2)
  );
  C53 c53_107 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_107_io_in_0),
    .io_in_1(c53_107_io_in_1),
    .io_in_2(c53_107_io_in_2),
    .io_in_3(c53_107_io_in_3),
    .io_in_4(c53_107_io_in_4),
    .io_out_0(c53_107_io_out_0),
    .io_out_1(c53_107_io_out_1),
    .io_out_2(c53_107_io_out_2)
  );
  C53 c53_108 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_108_io_in_0),
    .io_in_1(c53_108_io_in_1),
    .io_in_2(c53_108_io_in_2),
    .io_in_3(c53_108_io_in_3),
    .io_in_4(c53_108_io_in_4),
    .io_out_0(c53_108_io_out_0),
    .io_out_1(c53_108_io_out_1),
    .io_out_2(c53_108_io_out_2)
  );
  C53 c53_109 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_109_io_in_0),
    .io_in_1(c53_109_io_in_1),
    .io_in_2(c53_109_io_in_2),
    .io_in_3(c53_109_io_in_3),
    .io_in_4(c53_109_io_in_4),
    .io_out_0(c53_109_io_out_0),
    .io_out_1(c53_109_io_out_1),
    .io_out_2(c53_109_io_out_2)
  );
  C22 c22_11 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_11_io_in_0),
    .io_in_1(c22_11_io_in_1),
    .io_out_0(c22_11_io_out_0),
    .io_out_1(c22_11_io_out_1)
  );
  C53 c53_110 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_110_io_in_0),
    .io_in_1(c53_110_io_in_1),
    .io_in_2(c53_110_io_in_2),
    .io_in_3(c53_110_io_in_3),
    .io_in_4(c53_110_io_in_4),
    .io_out_0(c53_110_io_out_0),
    .io_out_1(c53_110_io_out_1),
    .io_out_2(c53_110_io_out_2)
  );
  C53 c53_111 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_111_io_in_0),
    .io_in_1(c53_111_io_in_1),
    .io_in_2(c53_111_io_in_2),
    .io_in_3(c53_111_io_in_3),
    .io_in_4(c53_111_io_in_4),
    .io_out_0(c53_111_io_out_0),
    .io_out_1(c53_111_io_out_1),
    .io_out_2(c53_111_io_out_2)
  );
  C53 c53_112 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_112_io_in_0),
    .io_in_1(c53_112_io_in_1),
    .io_in_2(c53_112_io_in_2),
    .io_in_3(c53_112_io_in_3),
    .io_in_4(c53_112_io_in_4),
    .io_out_0(c53_112_io_out_0),
    .io_out_1(c53_112_io_out_1),
    .io_out_2(c53_112_io_out_2)
  );
  C53 c53_113 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_113_io_in_0),
    .io_in_1(c53_113_io_in_1),
    .io_in_2(c53_113_io_in_2),
    .io_in_3(c53_113_io_in_3),
    .io_in_4(c53_113_io_in_4),
    .io_out_0(c53_113_io_out_0),
    .io_out_1(c53_113_io_out_1),
    .io_out_2(c53_113_io_out_2)
  );
  C53 c53_114 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_114_io_in_0),
    .io_in_1(c53_114_io_in_1),
    .io_in_2(c53_114_io_in_2),
    .io_in_3(c53_114_io_in_3),
    .io_in_4(c53_114_io_in_4),
    .io_out_0(c53_114_io_out_0),
    .io_out_1(c53_114_io_out_1),
    .io_out_2(c53_114_io_out_2)
  );
  C32 c32_10 ( // @[Multiplier.scala 78:25]
    .io_in_0(c32_10_io_in_0),
    .io_in_1(c32_10_io_in_1),
    .io_in_2(c32_10_io_in_2),
    .io_out_0(c32_10_io_out_0),
    .io_out_1(c32_10_io_out_1)
  );
  C53 c53_115 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_115_io_in_0),
    .io_in_1(c53_115_io_in_1),
    .io_in_2(c53_115_io_in_2),
    .io_in_3(c53_115_io_in_3),
    .io_in_4(c53_115_io_in_4),
    .io_out_0(c53_115_io_out_0),
    .io_out_1(c53_115_io_out_1),
    .io_out_2(c53_115_io_out_2)
  );
  C53 c53_116 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_116_io_in_0),
    .io_in_1(c53_116_io_in_1),
    .io_in_2(c53_116_io_in_2),
    .io_in_3(c53_116_io_in_3),
    .io_in_4(c53_116_io_in_4),
    .io_out_0(c53_116_io_out_0),
    .io_out_1(c53_116_io_out_1),
    .io_out_2(c53_116_io_out_2)
  );
  C53 c53_117 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_117_io_in_0),
    .io_in_1(c53_117_io_in_1),
    .io_in_2(c53_117_io_in_2),
    .io_in_3(c53_117_io_in_3),
    .io_in_4(c53_117_io_in_4),
    .io_out_0(c53_117_io_out_0),
    .io_out_1(c53_117_io_out_1),
    .io_out_2(c53_117_io_out_2)
  );
  C53 c53_118 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_118_io_in_0),
    .io_in_1(c53_118_io_in_1),
    .io_in_2(c53_118_io_in_2),
    .io_in_3(c53_118_io_in_3),
    .io_in_4(c53_118_io_in_4),
    .io_out_0(c53_118_io_out_0),
    .io_out_1(c53_118_io_out_1),
    .io_out_2(c53_118_io_out_2)
  );
  C53 c53_119 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_119_io_in_0),
    .io_in_1(c53_119_io_in_1),
    .io_in_2(c53_119_io_in_2),
    .io_in_3(c53_119_io_in_3),
    .io_in_4(c53_119_io_in_4),
    .io_out_0(c53_119_io_out_0),
    .io_out_1(c53_119_io_out_1),
    .io_out_2(c53_119_io_out_2)
  );
  C32 c32_11 ( // @[Multiplier.scala 78:25]
    .io_in_0(c32_11_io_in_0),
    .io_in_1(c32_11_io_in_1),
    .io_in_2(c32_11_io_in_2),
    .io_out_0(c32_11_io_out_0),
    .io_out_1(c32_11_io_out_1)
  );
  C53 c53_120 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_120_io_in_0),
    .io_in_1(c53_120_io_in_1),
    .io_in_2(c53_120_io_in_2),
    .io_in_3(c53_120_io_in_3),
    .io_in_4(c53_120_io_in_4),
    .io_out_0(c53_120_io_out_0),
    .io_out_1(c53_120_io_out_1),
    .io_out_2(c53_120_io_out_2)
  );
  C53 c53_121 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_121_io_in_0),
    .io_in_1(c53_121_io_in_1),
    .io_in_2(c53_121_io_in_2),
    .io_in_3(c53_121_io_in_3),
    .io_in_4(c53_121_io_in_4),
    .io_out_0(c53_121_io_out_0),
    .io_out_1(c53_121_io_out_1),
    .io_out_2(c53_121_io_out_2)
  );
  C53 c53_122 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_122_io_in_0),
    .io_in_1(c53_122_io_in_1),
    .io_in_2(c53_122_io_in_2),
    .io_in_3(c53_122_io_in_3),
    .io_in_4(c53_122_io_in_4),
    .io_out_0(c53_122_io_out_0),
    .io_out_1(c53_122_io_out_1),
    .io_out_2(c53_122_io_out_2)
  );
  C53 c53_123 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_123_io_in_0),
    .io_in_1(c53_123_io_in_1),
    .io_in_2(c53_123_io_in_2),
    .io_in_3(c53_123_io_in_3),
    .io_in_4(c53_123_io_in_4),
    .io_out_0(c53_123_io_out_0),
    .io_out_1(c53_123_io_out_1),
    .io_out_2(c53_123_io_out_2)
  );
  C53 c53_124 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_124_io_in_0),
    .io_in_1(c53_124_io_in_1),
    .io_in_2(c53_124_io_in_2),
    .io_in_3(c53_124_io_in_3),
    .io_in_4(c53_124_io_in_4),
    .io_out_0(c53_124_io_out_0),
    .io_out_1(c53_124_io_out_1),
    .io_out_2(c53_124_io_out_2)
  );
  C53 c53_125 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_125_io_in_0),
    .io_in_1(c53_125_io_in_1),
    .io_in_2(c53_125_io_in_2),
    .io_in_3(c53_125_io_in_3),
    .io_in_4(c53_125_io_in_4),
    .io_out_0(c53_125_io_out_0),
    .io_out_1(c53_125_io_out_1),
    .io_out_2(c53_125_io_out_2)
  );
  C53 c53_126 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_126_io_in_0),
    .io_in_1(c53_126_io_in_1),
    .io_in_2(c53_126_io_in_2),
    .io_in_3(c53_126_io_in_3),
    .io_in_4(c53_126_io_in_4),
    .io_out_0(c53_126_io_out_0),
    .io_out_1(c53_126_io_out_1),
    .io_out_2(c53_126_io_out_2)
  );
  C53 c53_127 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_127_io_in_0),
    .io_in_1(c53_127_io_in_1),
    .io_in_2(c53_127_io_in_2),
    .io_in_3(c53_127_io_in_3),
    .io_in_4(c53_127_io_in_4),
    .io_out_0(c53_127_io_out_0),
    .io_out_1(c53_127_io_out_1),
    .io_out_2(c53_127_io_out_2)
  );
  C53 c53_128 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_128_io_in_0),
    .io_in_1(c53_128_io_in_1),
    .io_in_2(c53_128_io_in_2),
    .io_in_3(c53_128_io_in_3),
    .io_in_4(c53_128_io_in_4),
    .io_out_0(c53_128_io_out_0),
    .io_out_1(c53_128_io_out_1),
    .io_out_2(c53_128_io_out_2)
  );
  C53 c53_129 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_129_io_in_0),
    .io_in_1(c53_129_io_in_1),
    .io_in_2(c53_129_io_in_2),
    .io_in_3(c53_129_io_in_3),
    .io_in_4(c53_129_io_in_4),
    .io_out_0(c53_129_io_out_0),
    .io_out_1(c53_129_io_out_1),
    .io_out_2(c53_129_io_out_2)
  );
  C53 c53_130 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_130_io_in_0),
    .io_in_1(c53_130_io_in_1),
    .io_in_2(c53_130_io_in_2),
    .io_in_3(c53_130_io_in_3),
    .io_in_4(c53_130_io_in_4),
    .io_out_0(c53_130_io_out_0),
    .io_out_1(c53_130_io_out_1),
    .io_out_2(c53_130_io_out_2)
  );
  C53 c53_131 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_131_io_in_0),
    .io_in_1(c53_131_io_in_1),
    .io_in_2(c53_131_io_in_2),
    .io_in_3(c53_131_io_in_3),
    .io_in_4(c53_131_io_in_4),
    .io_out_0(c53_131_io_out_0),
    .io_out_1(c53_131_io_out_1),
    .io_out_2(c53_131_io_out_2)
  );
  C53 c53_132 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_132_io_in_0),
    .io_in_1(c53_132_io_in_1),
    .io_in_2(c53_132_io_in_2),
    .io_in_3(c53_132_io_in_3),
    .io_in_4(c53_132_io_in_4),
    .io_out_0(c53_132_io_out_0),
    .io_out_1(c53_132_io_out_1),
    .io_out_2(c53_132_io_out_2)
  );
  C53 c53_133 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_133_io_in_0),
    .io_in_1(c53_133_io_in_1),
    .io_in_2(c53_133_io_in_2),
    .io_in_3(c53_133_io_in_3),
    .io_in_4(c53_133_io_in_4),
    .io_out_0(c53_133_io_out_0),
    .io_out_1(c53_133_io_out_1),
    .io_out_2(c53_133_io_out_2)
  );
  C53 c53_134 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_134_io_in_0),
    .io_in_1(c53_134_io_in_1),
    .io_in_2(c53_134_io_in_2),
    .io_in_3(c53_134_io_in_3),
    .io_in_4(c53_134_io_in_4),
    .io_out_0(c53_134_io_out_0),
    .io_out_1(c53_134_io_out_1),
    .io_out_2(c53_134_io_out_2)
  );
  C53 c53_135 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_135_io_in_0),
    .io_in_1(c53_135_io_in_1),
    .io_in_2(c53_135_io_in_2),
    .io_in_3(c53_135_io_in_3),
    .io_in_4(c53_135_io_in_4),
    .io_out_0(c53_135_io_out_0),
    .io_out_1(c53_135_io_out_1),
    .io_out_2(c53_135_io_out_2)
  );
  C53 c53_136 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_136_io_in_0),
    .io_in_1(c53_136_io_in_1),
    .io_in_2(c53_136_io_in_2),
    .io_in_3(c53_136_io_in_3),
    .io_in_4(c53_136_io_in_4),
    .io_out_0(c53_136_io_out_0),
    .io_out_1(c53_136_io_out_1),
    .io_out_2(c53_136_io_out_2)
  );
  C53 c53_137 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_137_io_in_0),
    .io_in_1(c53_137_io_in_1),
    .io_in_2(c53_137_io_in_2),
    .io_in_3(c53_137_io_in_3),
    .io_in_4(c53_137_io_in_4),
    .io_out_0(c53_137_io_out_0),
    .io_out_1(c53_137_io_out_1),
    .io_out_2(c53_137_io_out_2)
  );
  C53 c53_138 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_138_io_in_0),
    .io_in_1(c53_138_io_in_1),
    .io_in_2(c53_138_io_in_2),
    .io_in_3(c53_138_io_in_3),
    .io_in_4(c53_138_io_in_4),
    .io_out_0(c53_138_io_out_0),
    .io_out_1(c53_138_io_out_1),
    .io_out_2(c53_138_io_out_2)
  );
  C53 c53_139 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_139_io_in_0),
    .io_in_1(c53_139_io_in_1),
    .io_in_2(c53_139_io_in_2),
    .io_in_3(c53_139_io_in_3),
    .io_in_4(c53_139_io_in_4),
    .io_out_0(c53_139_io_out_0),
    .io_out_1(c53_139_io_out_1),
    .io_out_2(c53_139_io_out_2)
  );
  C53 c53_140 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_140_io_in_0),
    .io_in_1(c53_140_io_in_1),
    .io_in_2(c53_140_io_in_2),
    .io_in_3(c53_140_io_in_3),
    .io_in_4(c53_140_io_in_4),
    .io_out_0(c53_140_io_out_0),
    .io_out_1(c53_140_io_out_1),
    .io_out_2(c53_140_io_out_2)
  );
  C53 c53_141 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_141_io_in_0),
    .io_in_1(c53_141_io_in_1),
    .io_in_2(c53_141_io_in_2),
    .io_in_3(c53_141_io_in_3),
    .io_in_4(c53_141_io_in_4),
    .io_out_0(c53_141_io_out_0),
    .io_out_1(c53_141_io_out_1),
    .io_out_2(c53_141_io_out_2)
  );
  C53 c53_142 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_142_io_in_0),
    .io_in_1(c53_142_io_in_1),
    .io_in_2(c53_142_io_in_2),
    .io_in_3(c53_142_io_in_3),
    .io_in_4(c53_142_io_in_4),
    .io_out_0(c53_142_io_out_0),
    .io_out_1(c53_142_io_out_1),
    .io_out_2(c53_142_io_out_2)
  );
  C53 c53_143 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_143_io_in_0),
    .io_in_1(c53_143_io_in_1),
    .io_in_2(c53_143_io_in_2),
    .io_in_3(c53_143_io_in_3),
    .io_in_4(c53_143_io_in_4),
    .io_out_0(c53_143_io_out_0),
    .io_out_1(c53_143_io_out_1),
    .io_out_2(c53_143_io_out_2)
  );
  C53 c53_144 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_144_io_in_0),
    .io_in_1(c53_144_io_in_1),
    .io_in_2(c53_144_io_in_2),
    .io_in_3(c53_144_io_in_3),
    .io_in_4(c53_144_io_in_4),
    .io_out_0(c53_144_io_out_0),
    .io_out_1(c53_144_io_out_1),
    .io_out_2(c53_144_io_out_2)
  );
  C53 c53_145 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_145_io_in_0),
    .io_in_1(c53_145_io_in_1),
    .io_in_2(c53_145_io_in_2),
    .io_in_3(c53_145_io_in_3),
    .io_in_4(c53_145_io_in_4),
    .io_out_0(c53_145_io_out_0),
    .io_out_1(c53_145_io_out_1),
    .io_out_2(c53_145_io_out_2)
  );
  C53 c53_146 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_146_io_in_0),
    .io_in_1(c53_146_io_in_1),
    .io_in_2(c53_146_io_in_2),
    .io_in_3(c53_146_io_in_3),
    .io_in_4(c53_146_io_in_4),
    .io_out_0(c53_146_io_out_0),
    .io_out_1(c53_146_io_out_1),
    .io_out_2(c53_146_io_out_2)
  );
  C53 c53_147 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_147_io_in_0),
    .io_in_1(c53_147_io_in_1),
    .io_in_2(c53_147_io_in_2),
    .io_in_3(c53_147_io_in_3),
    .io_in_4(c53_147_io_in_4),
    .io_out_0(c53_147_io_out_0),
    .io_out_1(c53_147_io_out_1),
    .io_out_2(c53_147_io_out_2)
  );
  C53 c53_148 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_148_io_in_0),
    .io_in_1(c53_148_io_in_1),
    .io_in_2(c53_148_io_in_2),
    .io_in_3(c53_148_io_in_3),
    .io_in_4(c53_148_io_in_4),
    .io_out_0(c53_148_io_out_0),
    .io_out_1(c53_148_io_out_1),
    .io_out_2(c53_148_io_out_2)
  );
  C53 c53_149 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_149_io_in_0),
    .io_in_1(c53_149_io_in_1),
    .io_in_2(c53_149_io_in_2),
    .io_in_3(c53_149_io_in_3),
    .io_in_4(c53_149_io_in_4),
    .io_out_0(c53_149_io_out_0),
    .io_out_1(c53_149_io_out_1),
    .io_out_2(c53_149_io_out_2)
  );
  C22 c22_12 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_12_io_in_0),
    .io_in_1(c22_12_io_in_1),
    .io_out_0(c22_12_io_out_0),
    .io_out_1(c22_12_io_out_1)
  );
  C53 c53_150 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_150_io_in_0),
    .io_in_1(c53_150_io_in_1),
    .io_in_2(c53_150_io_in_2),
    .io_in_3(c53_150_io_in_3),
    .io_in_4(c53_150_io_in_4),
    .io_out_0(c53_150_io_out_0),
    .io_out_1(c53_150_io_out_1),
    .io_out_2(c53_150_io_out_2)
  );
  C53 c53_151 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_151_io_in_0),
    .io_in_1(c53_151_io_in_1),
    .io_in_2(c53_151_io_in_2),
    .io_in_3(c53_151_io_in_3),
    .io_in_4(c53_151_io_in_4),
    .io_out_0(c53_151_io_out_0),
    .io_out_1(c53_151_io_out_1),
    .io_out_2(c53_151_io_out_2)
  );
  C53 c53_152 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_152_io_in_0),
    .io_in_1(c53_152_io_in_1),
    .io_in_2(c53_152_io_in_2),
    .io_in_3(c53_152_io_in_3),
    .io_in_4(c53_152_io_in_4),
    .io_out_0(c53_152_io_out_0),
    .io_out_1(c53_152_io_out_1),
    .io_out_2(c53_152_io_out_2)
  );
  C53 c53_153 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_153_io_in_0),
    .io_in_1(c53_153_io_in_1),
    .io_in_2(c53_153_io_in_2),
    .io_in_3(c53_153_io_in_3),
    .io_in_4(c53_153_io_in_4),
    .io_out_0(c53_153_io_out_0),
    .io_out_1(c53_153_io_out_1),
    .io_out_2(c53_153_io_out_2)
  );
  C53 c53_154 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_154_io_in_0),
    .io_in_1(c53_154_io_in_1),
    .io_in_2(c53_154_io_in_2),
    .io_in_3(c53_154_io_in_3),
    .io_in_4(c53_154_io_in_4),
    .io_out_0(c53_154_io_out_0),
    .io_out_1(c53_154_io_out_1),
    .io_out_2(c53_154_io_out_2)
  );
  C53 c53_155 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_155_io_in_0),
    .io_in_1(c53_155_io_in_1),
    .io_in_2(c53_155_io_in_2),
    .io_in_3(c53_155_io_in_3),
    .io_in_4(c53_155_io_in_4),
    .io_out_0(c53_155_io_out_0),
    .io_out_1(c53_155_io_out_1),
    .io_out_2(c53_155_io_out_2)
  );
  C22 c22_13 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_13_io_in_0),
    .io_in_1(c22_13_io_in_1),
    .io_out_0(c22_13_io_out_0),
    .io_out_1(c22_13_io_out_1)
  );
  C53 c53_156 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_156_io_in_0),
    .io_in_1(c53_156_io_in_1),
    .io_in_2(c53_156_io_in_2),
    .io_in_3(c53_156_io_in_3),
    .io_in_4(c53_156_io_in_4),
    .io_out_0(c53_156_io_out_0),
    .io_out_1(c53_156_io_out_1),
    .io_out_2(c53_156_io_out_2)
  );
  C53 c53_157 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_157_io_in_0),
    .io_in_1(c53_157_io_in_1),
    .io_in_2(c53_157_io_in_2),
    .io_in_3(c53_157_io_in_3),
    .io_in_4(c53_157_io_in_4),
    .io_out_0(c53_157_io_out_0),
    .io_out_1(c53_157_io_out_1),
    .io_out_2(c53_157_io_out_2)
  );
  C53 c53_158 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_158_io_in_0),
    .io_in_1(c53_158_io_in_1),
    .io_in_2(c53_158_io_in_2),
    .io_in_3(c53_158_io_in_3),
    .io_in_4(c53_158_io_in_4),
    .io_out_0(c53_158_io_out_0),
    .io_out_1(c53_158_io_out_1),
    .io_out_2(c53_158_io_out_2)
  );
  C53 c53_159 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_159_io_in_0),
    .io_in_1(c53_159_io_in_1),
    .io_in_2(c53_159_io_in_2),
    .io_in_3(c53_159_io_in_3),
    .io_in_4(c53_159_io_in_4),
    .io_out_0(c53_159_io_out_0),
    .io_out_1(c53_159_io_out_1),
    .io_out_2(c53_159_io_out_2)
  );
  C53 c53_160 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_160_io_in_0),
    .io_in_1(c53_160_io_in_1),
    .io_in_2(c53_160_io_in_2),
    .io_in_3(c53_160_io_in_3),
    .io_in_4(c53_160_io_in_4),
    .io_out_0(c53_160_io_out_0),
    .io_out_1(c53_160_io_out_1),
    .io_out_2(c53_160_io_out_2)
  );
  C53 c53_161 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_161_io_in_0),
    .io_in_1(c53_161_io_in_1),
    .io_in_2(c53_161_io_in_2),
    .io_in_3(c53_161_io_in_3),
    .io_in_4(c53_161_io_in_4),
    .io_out_0(c53_161_io_out_0),
    .io_out_1(c53_161_io_out_1),
    .io_out_2(c53_161_io_out_2)
  );
  C32 c32_12 ( // @[Multiplier.scala 78:25]
    .io_in_0(c32_12_io_in_0),
    .io_in_1(c32_12_io_in_1),
    .io_in_2(c32_12_io_in_2),
    .io_out_0(c32_12_io_out_0),
    .io_out_1(c32_12_io_out_1)
  );
  C53 c53_162 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_162_io_in_0),
    .io_in_1(c53_162_io_in_1),
    .io_in_2(c53_162_io_in_2),
    .io_in_3(c53_162_io_in_3),
    .io_in_4(c53_162_io_in_4),
    .io_out_0(c53_162_io_out_0),
    .io_out_1(c53_162_io_out_1),
    .io_out_2(c53_162_io_out_2)
  );
  C53 c53_163 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_163_io_in_0),
    .io_in_1(c53_163_io_in_1),
    .io_in_2(c53_163_io_in_2),
    .io_in_3(c53_163_io_in_3),
    .io_in_4(c53_163_io_in_4),
    .io_out_0(c53_163_io_out_0),
    .io_out_1(c53_163_io_out_1),
    .io_out_2(c53_163_io_out_2)
  );
  C53 c53_164 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_164_io_in_0),
    .io_in_1(c53_164_io_in_1),
    .io_in_2(c53_164_io_in_2),
    .io_in_3(c53_164_io_in_3),
    .io_in_4(c53_164_io_in_4),
    .io_out_0(c53_164_io_out_0),
    .io_out_1(c53_164_io_out_1),
    .io_out_2(c53_164_io_out_2)
  );
  C53 c53_165 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_165_io_in_0),
    .io_in_1(c53_165_io_in_1),
    .io_in_2(c53_165_io_in_2),
    .io_in_3(c53_165_io_in_3),
    .io_in_4(c53_165_io_in_4),
    .io_out_0(c53_165_io_out_0),
    .io_out_1(c53_165_io_out_1),
    .io_out_2(c53_165_io_out_2)
  );
  C53 c53_166 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_166_io_in_0),
    .io_in_1(c53_166_io_in_1),
    .io_in_2(c53_166_io_in_2),
    .io_in_3(c53_166_io_in_3),
    .io_in_4(c53_166_io_in_4),
    .io_out_0(c53_166_io_out_0),
    .io_out_1(c53_166_io_out_1),
    .io_out_2(c53_166_io_out_2)
  );
  C53 c53_167 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_167_io_in_0),
    .io_in_1(c53_167_io_in_1),
    .io_in_2(c53_167_io_in_2),
    .io_in_3(c53_167_io_in_3),
    .io_in_4(c53_167_io_in_4),
    .io_out_0(c53_167_io_out_0),
    .io_out_1(c53_167_io_out_1),
    .io_out_2(c53_167_io_out_2)
  );
  C32 c32_13 ( // @[Multiplier.scala 78:25]
    .io_in_0(c32_13_io_in_0),
    .io_in_1(c32_13_io_in_1),
    .io_in_2(c32_13_io_in_2),
    .io_out_0(c32_13_io_out_0),
    .io_out_1(c32_13_io_out_1)
  );
  C53 c53_168 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_168_io_in_0),
    .io_in_1(c53_168_io_in_1),
    .io_in_2(c53_168_io_in_2),
    .io_in_3(c53_168_io_in_3),
    .io_in_4(c53_168_io_in_4),
    .io_out_0(c53_168_io_out_0),
    .io_out_1(c53_168_io_out_1),
    .io_out_2(c53_168_io_out_2)
  );
  C53 c53_169 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_169_io_in_0),
    .io_in_1(c53_169_io_in_1),
    .io_in_2(c53_169_io_in_2),
    .io_in_3(c53_169_io_in_3),
    .io_in_4(c53_169_io_in_4),
    .io_out_0(c53_169_io_out_0),
    .io_out_1(c53_169_io_out_1),
    .io_out_2(c53_169_io_out_2)
  );
  C53 c53_170 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_170_io_in_0),
    .io_in_1(c53_170_io_in_1),
    .io_in_2(c53_170_io_in_2),
    .io_in_3(c53_170_io_in_3),
    .io_in_4(c53_170_io_in_4),
    .io_out_0(c53_170_io_out_0),
    .io_out_1(c53_170_io_out_1),
    .io_out_2(c53_170_io_out_2)
  );
  C53 c53_171 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_171_io_in_0),
    .io_in_1(c53_171_io_in_1),
    .io_in_2(c53_171_io_in_2),
    .io_in_3(c53_171_io_in_3),
    .io_in_4(c53_171_io_in_4),
    .io_out_0(c53_171_io_out_0),
    .io_out_1(c53_171_io_out_1),
    .io_out_2(c53_171_io_out_2)
  );
  C53 c53_172 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_172_io_in_0),
    .io_in_1(c53_172_io_in_1),
    .io_in_2(c53_172_io_in_2),
    .io_in_3(c53_172_io_in_3),
    .io_in_4(c53_172_io_in_4),
    .io_out_0(c53_172_io_out_0),
    .io_out_1(c53_172_io_out_1),
    .io_out_2(c53_172_io_out_2)
  );
  C53 c53_173 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_173_io_in_0),
    .io_in_1(c53_173_io_in_1),
    .io_in_2(c53_173_io_in_2),
    .io_in_3(c53_173_io_in_3),
    .io_in_4(c53_173_io_in_4),
    .io_out_0(c53_173_io_out_0),
    .io_out_1(c53_173_io_out_1),
    .io_out_2(c53_173_io_out_2)
  );
  C32 c32_14 ( // @[Multiplier.scala 78:25]
    .io_in_0(c32_14_io_in_0),
    .io_in_1(c32_14_io_in_1),
    .io_in_2(c32_14_io_in_2),
    .io_out_0(c32_14_io_out_0),
    .io_out_1(c32_14_io_out_1)
  );
  C53 c53_174 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_174_io_in_0),
    .io_in_1(c53_174_io_in_1),
    .io_in_2(c53_174_io_in_2),
    .io_in_3(c53_174_io_in_3),
    .io_in_4(c53_174_io_in_4),
    .io_out_0(c53_174_io_out_0),
    .io_out_1(c53_174_io_out_1),
    .io_out_2(c53_174_io_out_2)
  );
  C53 c53_175 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_175_io_in_0),
    .io_in_1(c53_175_io_in_1),
    .io_in_2(c53_175_io_in_2),
    .io_in_3(c53_175_io_in_3),
    .io_in_4(c53_175_io_in_4),
    .io_out_0(c53_175_io_out_0),
    .io_out_1(c53_175_io_out_1),
    .io_out_2(c53_175_io_out_2)
  );
  C53 c53_176 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_176_io_in_0),
    .io_in_1(c53_176_io_in_1),
    .io_in_2(c53_176_io_in_2),
    .io_in_3(c53_176_io_in_3),
    .io_in_4(c53_176_io_in_4),
    .io_out_0(c53_176_io_out_0),
    .io_out_1(c53_176_io_out_1),
    .io_out_2(c53_176_io_out_2)
  );
  C53 c53_177 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_177_io_in_0),
    .io_in_1(c53_177_io_in_1),
    .io_in_2(c53_177_io_in_2),
    .io_in_3(c53_177_io_in_3),
    .io_in_4(c53_177_io_in_4),
    .io_out_0(c53_177_io_out_0),
    .io_out_1(c53_177_io_out_1),
    .io_out_2(c53_177_io_out_2)
  );
  C53 c53_178 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_178_io_in_0),
    .io_in_1(c53_178_io_in_1),
    .io_in_2(c53_178_io_in_2),
    .io_in_3(c53_178_io_in_3),
    .io_in_4(c53_178_io_in_4),
    .io_out_0(c53_178_io_out_0),
    .io_out_1(c53_178_io_out_1),
    .io_out_2(c53_178_io_out_2)
  );
  C53 c53_179 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_179_io_in_0),
    .io_in_1(c53_179_io_in_1),
    .io_in_2(c53_179_io_in_2),
    .io_in_3(c53_179_io_in_3),
    .io_in_4(c53_179_io_in_4),
    .io_out_0(c53_179_io_out_0),
    .io_out_1(c53_179_io_out_1),
    .io_out_2(c53_179_io_out_2)
  );
  C32 c32_15 ( // @[Multiplier.scala 78:25]
    .io_in_0(c32_15_io_in_0),
    .io_in_1(c32_15_io_in_1),
    .io_in_2(c32_15_io_in_2),
    .io_out_0(c32_15_io_out_0),
    .io_out_1(c32_15_io_out_1)
  );
  C53 c53_180 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_180_io_in_0),
    .io_in_1(c53_180_io_in_1),
    .io_in_2(c53_180_io_in_2),
    .io_in_3(c53_180_io_in_3),
    .io_in_4(c53_180_io_in_4),
    .io_out_0(c53_180_io_out_0),
    .io_out_1(c53_180_io_out_1),
    .io_out_2(c53_180_io_out_2)
  );
  C53 c53_181 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_181_io_in_0),
    .io_in_1(c53_181_io_in_1),
    .io_in_2(c53_181_io_in_2),
    .io_in_3(c53_181_io_in_3),
    .io_in_4(c53_181_io_in_4),
    .io_out_0(c53_181_io_out_0),
    .io_out_1(c53_181_io_out_1),
    .io_out_2(c53_181_io_out_2)
  );
  C53 c53_182 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_182_io_in_0),
    .io_in_1(c53_182_io_in_1),
    .io_in_2(c53_182_io_in_2),
    .io_in_3(c53_182_io_in_3),
    .io_in_4(c53_182_io_in_4),
    .io_out_0(c53_182_io_out_0),
    .io_out_1(c53_182_io_out_1),
    .io_out_2(c53_182_io_out_2)
  );
  C53 c53_183 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_183_io_in_0),
    .io_in_1(c53_183_io_in_1),
    .io_in_2(c53_183_io_in_2),
    .io_in_3(c53_183_io_in_3),
    .io_in_4(c53_183_io_in_4),
    .io_out_0(c53_183_io_out_0),
    .io_out_1(c53_183_io_out_1),
    .io_out_2(c53_183_io_out_2)
  );
  C53 c53_184 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_184_io_in_0),
    .io_in_1(c53_184_io_in_1),
    .io_in_2(c53_184_io_in_2),
    .io_in_3(c53_184_io_in_3),
    .io_in_4(c53_184_io_in_4),
    .io_out_0(c53_184_io_out_0),
    .io_out_1(c53_184_io_out_1),
    .io_out_2(c53_184_io_out_2)
  );
  C53 c53_185 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_185_io_in_0),
    .io_in_1(c53_185_io_in_1),
    .io_in_2(c53_185_io_in_2),
    .io_in_3(c53_185_io_in_3),
    .io_in_4(c53_185_io_in_4),
    .io_out_0(c53_185_io_out_0),
    .io_out_1(c53_185_io_out_1),
    .io_out_2(c53_185_io_out_2)
  );
  C32 c32_16 ( // @[Multiplier.scala 78:25]
    .io_in_0(c32_16_io_in_0),
    .io_in_1(c32_16_io_in_1),
    .io_in_2(c32_16_io_in_2),
    .io_out_0(c32_16_io_out_0),
    .io_out_1(c32_16_io_out_1)
  );
  C53 c53_186 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_186_io_in_0),
    .io_in_1(c53_186_io_in_1),
    .io_in_2(c53_186_io_in_2),
    .io_in_3(c53_186_io_in_3),
    .io_in_4(c53_186_io_in_4),
    .io_out_0(c53_186_io_out_0),
    .io_out_1(c53_186_io_out_1),
    .io_out_2(c53_186_io_out_2)
  );
  C53 c53_187 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_187_io_in_0),
    .io_in_1(c53_187_io_in_1),
    .io_in_2(c53_187_io_in_2),
    .io_in_3(c53_187_io_in_3),
    .io_in_4(c53_187_io_in_4),
    .io_out_0(c53_187_io_out_0),
    .io_out_1(c53_187_io_out_1),
    .io_out_2(c53_187_io_out_2)
  );
  C53 c53_188 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_188_io_in_0),
    .io_in_1(c53_188_io_in_1),
    .io_in_2(c53_188_io_in_2),
    .io_in_3(c53_188_io_in_3),
    .io_in_4(c53_188_io_in_4),
    .io_out_0(c53_188_io_out_0),
    .io_out_1(c53_188_io_out_1),
    .io_out_2(c53_188_io_out_2)
  );
  C53 c53_189 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_189_io_in_0),
    .io_in_1(c53_189_io_in_1),
    .io_in_2(c53_189_io_in_2),
    .io_in_3(c53_189_io_in_3),
    .io_in_4(c53_189_io_in_4),
    .io_out_0(c53_189_io_out_0),
    .io_out_1(c53_189_io_out_1),
    .io_out_2(c53_189_io_out_2)
  );
  C53 c53_190 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_190_io_in_0),
    .io_in_1(c53_190_io_in_1),
    .io_in_2(c53_190_io_in_2),
    .io_in_3(c53_190_io_in_3),
    .io_in_4(c53_190_io_in_4),
    .io_out_0(c53_190_io_out_0),
    .io_out_1(c53_190_io_out_1),
    .io_out_2(c53_190_io_out_2)
  );
  C53 c53_191 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_191_io_in_0),
    .io_in_1(c53_191_io_in_1),
    .io_in_2(c53_191_io_in_2),
    .io_in_3(c53_191_io_in_3),
    .io_in_4(c53_191_io_in_4),
    .io_out_0(c53_191_io_out_0),
    .io_out_1(c53_191_io_out_1),
    .io_out_2(c53_191_io_out_2)
  );
  C32 c32_17 ( // @[Multiplier.scala 78:25]
    .io_in_0(c32_17_io_in_0),
    .io_in_1(c32_17_io_in_1),
    .io_in_2(c32_17_io_in_2),
    .io_out_0(c32_17_io_out_0),
    .io_out_1(c32_17_io_out_1)
  );
  C53 c53_192 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_192_io_in_0),
    .io_in_1(c53_192_io_in_1),
    .io_in_2(c53_192_io_in_2),
    .io_in_3(c53_192_io_in_3),
    .io_in_4(c53_192_io_in_4),
    .io_out_0(c53_192_io_out_0),
    .io_out_1(c53_192_io_out_1),
    .io_out_2(c53_192_io_out_2)
  );
  C53 c53_193 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_193_io_in_0),
    .io_in_1(c53_193_io_in_1),
    .io_in_2(c53_193_io_in_2),
    .io_in_3(c53_193_io_in_3),
    .io_in_4(c53_193_io_in_4),
    .io_out_0(c53_193_io_out_0),
    .io_out_1(c53_193_io_out_1),
    .io_out_2(c53_193_io_out_2)
  );
  C53 c53_194 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_194_io_in_0),
    .io_in_1(c53_194_io_in_1),
    .io_in_2(c53_194_io_in_2),
    .io_in_3(c53_194_io_in_3),
    .io_in_4(c53_194_io_in_4),
    .io_out_0(c53_194_io_out_0),
    .io_out_1(c53_194_io_out_1),
    .io_out_2(c53_194_io_out_2)
  );
  C53 c53_195 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_195_io_in_0),
    .io_in_1(c53_195_io_in_1),
    .io_in_2(c53_195_io_in_2),
    .io_in_3(c53_195_io_in_3),
    .io_in_4(c53_195_io_in_4),
    .io_out_0(c53_195_io_out_0),
    .io_out_1(c53_195_io_out_1),
    .io_out_2(c53_195_io_out_2)
  );
  C53 c53_196 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_196_io_in_0),
    .io_in_1(c53_196_io_in_1),
    .io_in_2(c53_196_io_in_2),
    .io_in_3(c53_196_io_in_3),
    .io_in_4(c53_196_io_in_4),
    .io_out_0(c53_196_io_out_0),
    .io_out_1(c53_196_io_out_1),
    .io_out_2(c53_196_io_out_2)
  );
  C53 c53_197 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_197_io_in_0),
    .io_in_1(c53_197_io_in_1),
    .io_in_2(c53_197_io_in_2),
    .io_in_3(c53_197_io_in_3),
    .io_in_4(c53_197_io_in_4),
    .io_out_0(c53_197_io_out_0),
    .io_out_1(c53_197_io_out_1),
    .io_out_2(c53_197_io_out_2)
  );
  C32 c32_18 ( // @[Multiplier.scala 78:25]
    .io_in_0(c32_18_io_in_0),
    .io_in_1(c32_18_io_in_1),
    .io_in_2(c32_18_io_in_2),
    .io_out_0(c32_18_io_out_0),
    .io_out_1(c32_18_io_out_1)
  );
  C53 c53_198 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_198_io_in_0),
    .io_in_1(c53_198_io_in_1),
    .io_in_2(c53_198_io_in_2),
    .io_in_3(c53_198_io_in_3),
    .io_in_4(c53_198_io_in_4),
    .io_out_0(c53_198_io_out_0),
    .io_out_1(c53_198_io_out_1),
    .io_out_2(c53_198_io_out_2)
  );
  C53 c53_199 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_199_io_in_0),
    .io_in_1(c53_199_io_in_1),
    .io_in_2(c53_199_io_in_2),
    .io_in_3(c53_199_io_in_3),
    .io_in_4(c53_199_io_in_4),
    .io_out_0(c53_199_io_out_0),
    .io_out_1(c53_199_io_out_1),
    .io_out_2(c53_199_io_out_2)
  );
  C53 c53_200 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_200_io_in_0),
    .io_in_1(c53_200_io_in_1),
    .io_in_2(c53_200_io_in_2),
    .io_in_3(c53_200_io_in_3),
    .io_in_4(c53_200_io_in_4),
    .io_out_0(c53_200_io_out_0),
    .io_out_1(c53_200_io_out_1),
    .io_out_2(c53_200_io_out_2)
  );
  C53 c53_201 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_201_io_in_0),
    .io_in_1(c53_201_io_in_1),
    .io_in_2(c53_201_io_in_2),
    .io_in_3(c53_201_io_in_3),
    .io_in_4(c53_201_io_in_4),
    .io_out_0(c53_201_io_out_0),
    .io_out_1(c53_201_io_out_1),
    .io_out_2(c53_201_io_out_2)
  );
  C53 c53_202 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_202_io_in_0),
    .io_in_1(c53_202_io_in_1),
    .io_in_2(c53_202_io_in_2),
    .io_in_3(c53_202_io_in_3),
    .io_in_4(c53_202_io_in_4),
    .io_out_0(c53_202_io_out_0),
    .io_out_1(c53_202_io_out_1),
    .io_out_2(c53_202_io_out_2)
  );
  C53 c53_203 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_203_io_in_0),
    .io_in_1(c53_203_io_in_1),
    .io_in_2(c53_203_io_in_2),
    .io_in_3(c53_203_io_in_3),
    .io_in_4(c53_203_io_in_4),
    .io_out_0(c53_203_io_out_0),
    .io_out_1(c53_203_io_out_1),
    .io_out_2(c53_203_io_out_2)
  );
  C32 c32_19 ( // @[Multiplier.scala 78:25]
    .io_in_0(c32_19_io_in_0),
    .io_in_1(c32_19_io_in_1),
    .io_in_2(c32_19_io_in_2),
    .io_out_0(c32_19_io_out_0),
    .io_out_1(c32_19_io_out_1)
  );
  C53 c53_204 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_204_io_in_0),
    .io_in_1(c53_204_io_in_1),
    .io_in_2(c53_204_io_in_2),
    .io_in_3(c53_204_io_in_3),
    .io_in_4(c53_204_io_in_4),
    .io_out_0(c53_204_io_out_0),
    .io_out_1(c53_204_io_out_1),
    .io_out_2(c53_204_io_out_2)
  );
  C53 c53_205 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_205_io_in_0),
    .io_in_1(c53_205_io_in_1),
    .io_in_2(c53_205_io_in_2),
    .io_in_3(c53_205_io_in_3),
    .io_in_4(c53_205_io_in_4),
    .io_out_0(c53_205_io_out_0),
    .io_out_1(c53_205_io_out_1),
    .io_out_2(c53_205_io_out_2)
  );
  C53 c53_206 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_206_io_in_0),
    .io_in_1(c53_206_io_in_1),
    .io_in_2(c53_206_io_in_2),
    .io_in_3(c53_206_io_in_3),
    .io_in_4(c53_206_io_in_4),
    .io_out_0(c53_206_io_out_0),
    .io_out_1(c53_206_io_out_1),
    .io_out_2(c53_206_io_out_2)
  );
  C53 c53_207 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_207_io_in_0),
    .io_in_1(c53_207_io_in_1),
    .io_in_2(c53_207_io_in_2),
    .io_in_3(c53_207_io_in_3),
    .io_in_4(c53_207_io_in_4),
    .io_out_0(c53_207_io_out_0),
    .io_out_1(c53_207_io_out_1),
    .io_out_2(c53_207_io_out_2)
  );
  C53 c53_208 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_208_io_in_0),
    .io_in_1(c53_208_io_in_1),
    .io_in_2(c53_208_io_in_2),
    .io_in_3(c53_208_io_in_3),
    .io_in_4(c53_208_io_in_4),
    .io_out_0(c53_208_io_out_0),
    .io_out_1(c53_208_io_out_1),
    .io_out_2(c53_208_io_out_2)
  );
  C53 c53_209 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_209_io_in_0),
    .io_in_1(c53_209_io_in_1),
    .io_in_2(c53_209_io_in_2),
    .io_in_3(c53_209_io_in_3),
    .io_in_4(c53_209_io_in_4),
    .io_out_0(c53_209_io_out_0),
    .io_out_1(c53_209_io_out_1),
    .io_out_2(c53_209_io_out_2)
  );
  C22 c22_14 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_14_io_in_0),
    .io_in_1(c22_14_io_in_1),
    .io_out_0(c22_14_io_out_0),
    .io_out_1(c22_14_io_out_1)
  );
  C53 c53_210 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_210_io_in_0),
    .io_in_1(c53_210_io_in_1),
    .io_in_2(c53_210_io_in_2),
    .io_in_3(c53_210_io_in_3),
    .io_in_4(c53_210_io_in_4),
    .io_out_0(c53_210_io_out_0),
    .io_out_1(c53_210_io_out_1),
    .io_out_2(c53_210_io_out_2)
  );
  C53 c53_211 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_211_io_in_0),
    .io_in_1(c53_211_io_in_1),
    .io_in_2(c53_211_io_in_2),
    .io_in_3(c53_211_io_in_3),
    .io_in_4(c53_211_io_in_4),
    .io_out_0(c53_211_io_out_0),
    .io_out_1(c53_211_io_out_1),
    .io_out_2(c53_211_io_out_2)
  );
  C53 c53_212 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_212_io_in_0),
    .io_in_1(c53_212_io_in_1),
    .io_in_2(c53_212_io_in_2),
    .io_in_3(c53_212_io_in_3),
    .io_in_4(c53_212_io_in_4),
    .io_out_0(c53_212_io_out_0),
    .io_out_1(c53_212_io_out_1),
    .io_out_2(c53_212_io_out_2)
  );
  C53 c53_213 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_213_io_in_0),
    .io_in_1(c53_213_io_in_1),
    .io_in_2(c53_213_io_in_2),
    .io_in_3(c53_213_io_in_3),
    .io_in_4(c53_213_io_in_4),
    .io_out_0(c53_213_io_out_0),
    .io_out_1(c53_213_io_out_1),
    .io_out_2(c53_213_io_out_2)
  );
  C53 c53_214 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_214_io_in_0),
    .io_in_1(c53_214_io_in_1),
    .io_in_2(c53_214_io_in_2),
    .io_in_3(c53_214_io_in_3),
    .io_in_4(c53_214_io_in_4),
    .io_out_0(c53_214_io_out_0),
    .io_out_1(c53_214_io_out_1),
    .io_out_2(c53_214_io_out_2)
  );
  C53 c53_215 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_215_io_in_0),
    .io_in_1(c53_215_io_in_1),
    .io_in_2(c53_215_io_in_2),
    .io_in_3(c53_215_io_in_3),
    .io_in_4(c53_215_io_in_4),
    .io_out_0(c53_215_io_out_0),
    .io_out_1(c53_215_io_out_1),
    .io_out_2(c53_215_io_out_2)
  );
  C53 c53_216 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_216_io_in_0),
    .io_in_1(c53_216_io_in_1),
    .io_in_2(c53_216_io_in_2),
    .io_in_3(c53_216_io_in_3),
    .io_in_4(c53_216_io_in_4),
    .io_out_0(c53_216_io_out_0),
    .io_out_1(c53_216_io_out_1),
    .io_out_2(c53_216_io_out_2)
  );
  C53 c53_217 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_217_io_in_0),
    .io_in_1(c53_217_io_in_1),
    .io_in_2(c53_217_io_in_2),
    .io_in_3(c53_217_io_in_3),
    .io_in_4(c53_217_io_in_4),
    .io_out_0(c53_217_io_out_0),
    .io_out_1(c53_217_io_out_1),
    .io_out_2(c53_217_io_out_2)
  );
  C53 c53_218 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_218_io_in_0),
    .io_in_1(c53_218_io_in_1),
    .io_in_2(c53_218_io_in_2),
    .io_in_3(c53_218_io_in_3),
    .io_in_4(c53_218_io_in_4),
    .io_out_0(c53_218_io_out_0),
    .io_out_1(c53_218_io_out_1),
    .io_out_2(c53_218_io_out_2)
  );
  C53 c53_219 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_219_io_in_0),
    .io_in_1(c53_219_io_in_1),
    .io_in_2(c53_219_io_in_2),
    .io_in_3(c53_219_io_in_3),
    .io_in_4(c53_219_io_in_4),
    .io_out_0(c53_219_io_out_0),
    .io_out_1(c53_219_io_out_1),
    .io_out_2(c53_219_io_out_2)
  );
  C53 c53_220 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_220_io_in_0),
    .io_in_1(c53_220_io_in_1),
    .io_in_2(c53_220_io_in_2),
    .io_in_3(c53_220_io_in_3),
    .io_in_4(c53_220_io_in_4),
    .io_out_0(c53_220_io_out_0),
    .io_out_1(c53_220_io_out_1),
    .io_out_2(c53_220_io_out_2)
  );
  C53 c53_221 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_221_io_in_0),
    .io_in_1(c53_221_io_in_1),
    .io_in_2(c53_221_io_in_2),
    .io_in_3(c53_221_io_in_3),
    .io_in_4(c53_221_io_in_4),
    .io_out_0(c53_221_io_out_0),
    .io_out_1(c53_221_io_out_1),
    .io_out_2(c53_221_io_out_2)
  );
  C53 c53_222 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_222_io_in_0),
    .io_in_1(c53_222_io_in_1),
    .io_in_2(c53_222_io_in_2),
    .io_in_3(c53_222_io_in_3),
    .io_in_4(c53_222_io_in_4),
    .io_out_0(c53_222_io_out_0),
    .io_out_1(c53_222_io_out_1),
    .io_out_2(c53_222_io_out_2)
  );
  C53 c53_223 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_223_io_in_0),
    .io_in_1(c53_223_io_in_1),
    .io_in_2(c53_223_io_in_2),
    .io_in_3(c53_223_io_in_3),
    .io_in_4(c53_223_io_in_4),
    .io_out_0(c53_223_io_out_0),
    .io_out_1(c53_223_io_out_1),
    .io_out_2(c53_223_io_out_2)
  );
  C53 c53_224 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_224_io_in_0),
    .io_in_1(c53_224_io_in_1),
    .io_in_2(c53_224_io_in_2),
    .io_in_3(c53_224_io_in_3),
    .io_in_4(c53_224_io_in_4),
    .io_out_0(c53_224_io_out_0),
    .io_out_1(c53_224_io_out_1),
    .io_out_2(c53_224_io_out_2)
  );
  C53 c53_225 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_225_io_in_0),
    .io_in_1(c53_225_io_in_1),
    .io_in_2(c53_225_io_in_2),
    .io_in_3(c53_225_io_in_3),
    .io_in_4(c53_225_io_in_4),
    .io_out_0(c53_225_io_out_0),
    .io_out_1(c53_225_io_out_1),
    .io_out_2(c53_225_io_out_2)
  );
  C53 c53_226 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_226_io_in_0),
    .io_in_1(c53_226_io_in_1),
    .io_in_2(c53_226_io_in_2),
    .io_in_3(c53_226_io_in_3),
    .io_in_4(c53_226_io_in_4),
    .io_out_0(c53_226_io_out_0),
    .io_out_1(c53_226_io_out_1),
    .io_out_2(c53_226_io_out_2)
  );
  C53 c53_227 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_227_io_in_0),
    .io_in_1(c53_227_io_in_1),
    .io_in_2(c53_227_io_in_2),
    .io_in_3(c53_227_io_in_3),
    .io_in_4(c53_227_io_in_4),
    .io_out_0(c53_227_io_out_0),
    .io_out_1(c53_227_io_out_1),
    .io_out_2(c53_227_io_out_2)
  );
  C53 c53_228 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_228_io_in_0),
    .io_in_1(c53_228_io_in_1),
    .io_in_2(c53_228_io_in_2),
    .io_in_3(c53_228_io_in_3),
    .io_in_4(c53_228_io_in_4),
    .io_out_0(c53_228_io_out_0),
    .io_out_1(c53_228_io_out_1),
    .io_out_2(c53_228_io_out_2)
  );
  C53 c53_229 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_229_io_in_0),
    .io_in_1(c53_229_io_in_1),
    .io_in_2(c53_229_io_in_2),
    .io_in_3(c53_229_io_in_3),
    .io_in_4(c53_229_io_in_4),
    .io_out_0(c53_229_io_out_0),
    .io_out_1(c53_229_io_out_1),
    .io_out_2(c53_229_io_out_2)
  );
  C53 c53_230 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_230_io_in_0),
    .io_in_1(c53_230_io_in_1),
    .io_in_2(c53_230_io_in_2),
    .io_in_3(c53_230_io_in_3),
    .io_in_4(c53_230_io_in_4),
    .io_out_0(c53_230_io_out_0),
    .io_out_1(c53_230_io_out_1),
    .io_out_2(c53_230_io_out_2)
  );
  C53 c53_231 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_231_io_in_0),
    .io_in_1(c53_231_io_in_1),
    .io_in_2(c53_231_io_in_2),
    .io_in_3(c53_231_io_in_3),
    .io_in_4(c53_231_io_in_4),
    .io_out_0(c53_231_io_out_0),
    .io_out_1(c53_231_io_out_1),
    .io_out_2(c53_231_io_out_2)
  );
  C53 c53_232 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_232_io_in_0),
    .io_in_1(c53_232_io_in_1),
    .io_in_2(c53_232_io_in_2),
    .io_in_3(c53_232_io_in_3),
    .io_in_4(c53_232_io_in_4),
    .io_out_0(c53_232_io_out_0),
    .io_out_1(c53_232_io_out_1),
    .io_out_2(c53_232_io_out_2)
  );
  C53 c53_233 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_233_io_in_0),
    .io_in_1(c53_233_io_in_1),
    .io_in_2(c53_233_io_in_2),
    .io_in_3(c53_233_io_in_3),
    .io_in_4(c53_233_io_in_4),
    .io_out_0(c53_233_io_out_0),
    .io_out_1(c53_233_io_out_1),
    .io_out_2(c53_233_io_out_2)
  );
  C53 c53_234 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_234_io_in_0),
    .io_in_1(c53_234_io_in_1),
    .io_in_2(c53_234_io_in_2),
    .io_in_3(c53_234_io_in_3),
    .io_in_4(c53_234_io_in_4),
    .io_out_0(c53_234_io_out_0),
    .io_out_1(c53_234_io_out_1),
    .io_out_2(c53_234_io_out_2)
  );
  C53 c53_235 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_235_io_in_0),
    .io_in_1(c53_235_io_in_1),
    .io_in_2(c53_235_io_in_2),
    .io_in_3(c53_235_io_in_3),
    .io_in_4(c53_235_io_in_4),
    .io_out_0(c53_235_io_out_0),
    .io_out_1(c53_235_io_out_1),
    .io_out_2(c53_235_io_out_2)
  );
  C53 c53_236 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_236_io_in_0),
    .io_in_1(c53_236_io_in_1),
    .io_in_2(c53_236_io_in_2),
    .io_in_3(c53_236_io_in_3),
    .io_in_4(c53_236_io_in_4),
    .io_out_0(c53_236_io_out_0),
    .io_out_1(c53_236_io_out_1),
    .io_out_2(c53_236_io_out_2)
  );
  C53 c53_237 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_237_io_in_0),
    .io_in_1(c53_237_io_in_1),
    .io_in_2(c53_237_io_in_2),
    .io_in_3(c53_237_io_in_3),
    .io_in_4(c53_237_io_in_4),
    .io_out_0(c53_237_io_out_0),
    .io_out_1(c53_237_io_out_1),
    .io_out_2(c53_237_io_out_2)
  );
  C53 c53_238 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_238_io_in_0),
    .io_in_1(c53_238_io_in_1),
    .io_in_2(c53_238_io_in_2),
    .io_in_3(c53_238_io_in_3),
    .io_in_4(c53_238_io_in_4),
    .io_out_0(c53_238_io_out_0),
    .io_out_1(c53_238_io_out_1),
    .io_out_2(c53_238_io_out_2)
  );
  C32 c32_20 ( // @[Multiplier.scala 78:25]
    .io_in_0(c32_20_io_in_0),
    .io_in_1(c32_20_io_in_1),
    .io_in_2(c32_20_io_in_2),
    .io_out_0(c32_20_io_out_0),
    .io_out_1(c32_20_io_out_1)
  );
  C53 c53_239 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_239_io_in_0),
    .io_in_1(c53_239_io_in_1),
    .io_in_2(c53_239_io_in_2),
    .io_in_3(c53_239_io_in_3),
    .io_in_4(c53_239_io_in_4),
    .io_out_0(c53_239_io_out_0),
    .io_out_1(c53_239_io_out_1),
    .io_out_2(c53_239_io_out_2)
  );
  C53 c53_240 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_240_io_in_0),
    .io_in_1(c53_240_io_in_1),
    .io_in_2(c53_240_io_in_2),
    .io_in_3(c53_240_io_in_3),
    .io_in_4(c53_240_io_in_4),
    .io_out_0(c53_240_io_out_0),
    .io_out_1(c53_240_io_out_1),
    .io_out_2(c53_240_io_out_2)
  );
  C53 c53_241 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_241_io_in_0),
    .io_in_1(c53_241_io_in_1),
    .io_in_2(c53_241_io_in_2),
    .io_in_3(c53_241_io_in_3),
    .io_in_4(c53_241_io_in_4),
    .io_out_0(c53_241_io_out_0),
    .io_out_1(c53_241_io_out_1),
    .io_out_2(c53_241_io_out_2)
  );
  C53 c53_242 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_242_io_in_0),
    .io_in_1(c53_242_io_in_1),
    .io_in_2(c53_242_io_in_2),
    .io_in_3(c53_242_io_in_3),
    .io_in_4(c53_242_io_in_4),
    .io_out_0(c53_242_io_out_0),
    .io_out_1(c53_242_io_out_1),
    .io_out_2(c53_242_io_out_2)
  );
  C53 c53_243 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_243_io_in_0),
    .io_in_1(c53_243_io_in_1),
    .io_in_2(c53_243_io_in_2),
    .io_in_3(c53_243_io_in_3),
    .io_in_4(c53_243_io_in_4),
    .io_out_0(c53_243_io_out_0),
    .io_out_1(c53_243_io_out_1),
    .io_out_2(c53_243_io_out_2)
  );
  C32 c32_21 ( // @[Multiplier.scala 78:25]
    .io_in_0(c32_21_io_in_0),
    .io_in_1(c32_21_io_in_1),
    .io_in_2(c32_21_io_in_2),
    .io_out_0(c32_21_io_out_0),
    .io_out_1(c32_21_io_out_1)
  );
  C53 c53_244 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_244_io_in_0),
    .io_in_1(c53_244_io_in_1),
    .io_in_2(c53_244_io_in_2),
    .io_in_3(c53_244_io_in_3),
    .io_in_4(c53_244_io_in_4),
    .io_out_0(c53_244_io_out_0),
    .io_out_1(c53_244_io_out_1),
    .io_out_2(c53_244_io_out_2)
  );
  C53 c53_245 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_245_io_in_0),
    .io_in_1(c53_245_io_in_1),
    .io_in_2(c53_245_io_in_2),
    .io_in_3(c53_245_io_in_3),
    .io_in_4(c53_245_io_in_4),
    .io_out_0(c53_245_io_out_0),
    .io_out_1(c53_245_io_out_1),
    .io_out_2(c53_245_io_out_2)
  );
  C53 c53_246 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_246_io_in_0),
    .io_in_1(c53_246_io_in_1),
    .io_in_2(c53_246_io_in_2),
    .io_in_3(c53_246_io_in_3),
    .io_in_4(c53_246_io_in_4),
    .io_out_0(c53_246_io_out_0),
    .io_out_1(c53_246_io_out_1),
    .io_out_2(c53_246_io_out_2)
  );
  C53 c53_247 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_247_io_in_0),
    .io_in_1(c53_247_io_in_1),
    .io_in_2(c53_247_io_in_2),
    .io_in_3(c53_247_io_in_3),
    .io_in_4(c53_247_io_in_4),
    .io_out_0(c53_247_io_out_0),
    .io_out_1(c53_247_io_out_1),
    .io_out_2(c53_247_io_out_2)
  );
  C53 c53_248 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_248_io_in_0),
    .io_in_1(c53_248_io_in_1),
    .io_in_2(c53_248_io_in_2),
    .io_in_3(c53_248_io_in_3),
    .io_in_4(c53_248_io_in_4),
    .io_out_0(c53_248_io_out_0),
    .io_out_1(c53_248_io_out_1),
    .io_out_2(c53_248_io_out_2)
  );
  C22 c22_15 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_15_io_in_0),
    .io_in_1(c22_15_io_in_1),
    .io_out_0(c22_15_io_out_0),
    .io_out_1(c22_15_io_out_1)
  );
  C53 c53_249 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_249_io_in_0),
    .io_in_1(c53_249_io_in_1),
    .io_in_2(c53_249_io_in_2),
    .io_in_3(c53_249_io_in_3),
    .io_in_4(c53_249_io_in_4),
    .io_out_0(c53_249_io_out_0),
    .io_out_1(c53_249_io_out_1),
    .io_out_2(c53_249_io_out_2)
  );
  C53 c53_250 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_250_io_in_0),
    .io_in_1(c53_250_io_in_1),
    .io_in_2(c53_250_io_in_2),
    .io_in_3(c53_250_io_in_3),
    .io_in_4(c53_250_io_in_4),
    .io_out_0(c53_250_io_out_0),
    .io_out_1(c53_250_io_out_1),
    .io_out_2(c53_250_io_out_2)
  );
  C53 c53_251 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_251_io_in_0),
    .io_in_1(c53_251_io_in_1),
    .io_in_2(c53_251_io_in_2),
    .io_in_3(c53_251_io_in_3),
    .io_in_4(c53_251_io_in_4),
    .io_out_0(c53_251_io_out_0),
    .io_out_1(c53_251_io_out_1),
    .io_out_2(c53_251_io_out_2)
  );
  C53 c53_252 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_252_io_in_0),
    .io_in_1(c53_252_io_in_1),
    .io_in_2(c53_252_io_in_2),
    .io_in_3(c53_252_io_in_3),
    .io_in_4(c53_252_io_in_4),
    .io_out_0(c53_252_io_out_0),
    .io_out_1(c53_252_io_out_1),
    .io_out_2(c53_252_io_out_2)
  );
  C53 c53_253 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_253_io_in_0),
    .io_in_1(c53_253_io_in_1),
    .io_in_2(c53_253_io_in_2),
    .io_in_3(c53_253_io_in_3),
    .io_in_4(c53_253_io_in_4),
    .io_out_0(c53_253_io_out_0),
    .io_out_1(c53_253_io_out_1),
    .io_out_2(c53_253_io_out_2)
  );
  C22 c22_16 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_16_io_in_0),
    .io_in_1(c22_16_io_in_1),
    .io_out_0(c22_16_io_out_0),
    .io_out_1(c22_16_io_out_1)
  );
  C53 c53_254 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_254_io_in_0),
    .io_in_1(c53_254_io_in_1),
    .io_in_2(c53_254_io_in_2),
    .io_in_3(c53_254_io_in_3),
    .io_in_4(c53_254_io_in_4),
    .io_out_0(c53_254_io_out_0),
    .io_out_1(c53_254_io_out_1),
    .io_out_2(c53_254_io_out_2)
  );
  C53 c53_255 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_255_io_in_0),
    .io_in_1(c53_255_io_in_1),
    .io_in_2(c53_255_io_in_2),
    .io_in_3(c53_255_io_in_3),
    .io_in_4(c53_255_io_in_4),
    .io_out_0(c53_255_io_out_0),
    .io_out_1(c53_255_io_out_1),
    .io_out_2(c53_255_io_out_2)
  );
  C53 c53_256 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_256_io_in_0),
    .io_in_1(c53_256_io_in_1),
    .io_in_2(c53_256_io_in_2),
    .io_in_3(c53_256_io_in_3),
    .io_in_4(c53_256_io_in_4),
    .io_out_0(c53_256_io_out_0),
    .io_out_1(c53_256_io_out_1),
    .io_out_2(c53_256_io_out_2)
  );
  C53 c53_257 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_257_io_in_0),
    .io_in_1(c53_257_io_in_1),
    .io_in_2(c53_257_io_in_2),
    .io_in_3(c53_257_io_in_3),
    .io_in_4(c53_257_io_in_4),
    .io_out_0(c53_257_io_out_0),
    .io_out_1(c53_257_io_out_1),
    .io_out_2(c53_257_io_out_2)
  );
  C53 c53_258 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_258_io_in_0),
    .io_in_1(c53_258_io_in_1),
    .io_in_2(c53_258_io_in_2),
    .io_in_3(c53_258_io_in_3),
    .io_in_4(c53_258_io_in_4),
    .io_out_0(c53_258_io_out_0),
    .io_out_1(c53_258_io_out_1),
    .io_out_2(c53_258_io_out_2)
  );
  C53 c53_259 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_259_io_in_0),
    .io_in_1(c53_259_io_in_1),
    .io_in_2(c53_259_io_in_2),
    .io_in_3(c53_259_io_in_3),
    .io_in_4(c53_259_io_in_4),
    .io_out_0(c53_259_io_out_0),
    .io_out_1(c53_259_io_out_1),
    .io_out_2(c53_259_io_out_2)
  );
  C53 c53_260 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_260_io_in_0),
    .io_in_1(c53_260_io_in_1),
    .io_in_2(c53_260_io_in_2),
    .io_in_3(c53_260_io_in_3),
    .io_in_4(c53_260_io_in_4),
    .io_out_0(c53_260_io_out_0),
    .io_out_1(c53_260_io_out_1),
    .io_out_2(c53_260_io_out_2)
  );
  C53 c53_261 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_261_io_in_0),
    .io_in_1(c53_261_io_in_1),
    .io_in_2(c53_261_io_in_2),
    .io_in_3(c53_261_io_in_3),
    .io_in_4(c53_261_io_in_4),
    .io_out_0(c53_261_io_out_0),
    .io_out_1(c53_261_io_out_1),
    .io_out_2(c53_261_io_out_2)
  );
  C53 c53_262 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_262_io_in_0),
    .io_in_1(c53_262_io_in_1),
    .io_in_2(c53_262_io_in_2),
    .io_in_3(c53_262_io_in_3),
    .io_in_4(c53_262_io_in_4),
    .io_out_0(c53_262_io_out_0),
    .io_out_1(c53_262_io_out_1),
    .io_out_2(c53_262_io_out_2)
  );
  C53 c53_263 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_263_io_in_0),
    .io_in_1(c53_263_io_in_1),
    .io_in_2(c53_263_io_in_2),
    .io_in_3(c53_263_io_in_3),
    .io_in_4(c53_263_io_in_4),
    .io_out_0(c53_263_io_out_0),
    .io_out_1(c53_263_io_out_1),
    .io_out_2(c53_263_io_out_2)
  );
  C53 c53_264 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_264_io_in_0),
    .io_in_1(c53_264_io_in_1),
    .io_in_2(c53_264_io_in_2),
    .io_in_3(c53_264_io_in_3),
    .io_in_4(c53_264_io_in_4),
    .io_out_0(c53_264_io_out_0),
    .io_out_1(c53_264_io_out_1),
    .io_out_2(c53_264_io_out_2)
  );
  C53 c53_265 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_265_io_in_0),
    .io_in_1(c53_265_io_in_1),
    .io_in_2(c53_265_io_in_2),
    .io_in_3(c53_265_io_in_3),
    .io_in_4(c53_265_io_in_4),
    .io_out_0(c53_265_io_out_0),
    .io_out_1(c53_265_io_out_1),
    .io_out_2(c53_265_io_out_2)
  );
  C53 c53_266 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_266_io_in_0),
    .io_in_1(c53_266_io_in_1),
    .io_in_2(c53_266_io_in_2),
    .io_in_3(c53_266_io_in_3),
    .io_in_4(c53_266_io_in_4),
    .io_out_0(c53_266_io_out_0),
    .io_out_1(c53_266_io_out_1),
    .io_out_2(c53_266_io_out_2)
  );
  C53 c53_267 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_267_io_in_0),
    .io_in_1(c53_267_io_in_1),
    .io_in_2(c53_267_io_in_2),
    .io_in_3(c53_267_io_in_3),
    .io_in_4(c53_267_io_in_4),
    .io_out_0(c53_267_io_out_0),
    .io_out_1(c53_267_io_out_1),
    .io_out_2(c53_267_io_out_2)
  );
  C53 c53_268 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_268_io_in_0),
    .io_in_1(c53_268_io_in_1),
    .io_in_2(c53_268_io_in_2),
    .io_in_3(c53_268_io_in_3),
    .io_in_4(c53_268_io_in_4),
    .io_out_0(c53_268_io_out_0),
    .io_out_1(c53_268_io_out_1),
    .io_out_2(c53_268_io_out_2)
  );
  C53 c53_269 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_269_io_in_0),
    .io_in_1(c53_269_io_in_1),
    .io_in_2(c53_269_io_in_2),
    .io_in_3(c53_269_io_in_3),
    .io_in_4(c53_269_io_in_4),
    .io_out_0(c53_269_io_out_0),
    .io_out_1(c53_269_io_out_1),
    .io_out_2(c53_269_io_out_2)
  );
  C53 c53_270 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_270_io_in_0),
    .io_in_1(c53_270_io_in_1),
    .io_in_2(c53_270_io_in_2),
    .io_in_3(c53_270_io_in_3),
    .io_in_4(c53_270_io_in_4),
    .io_out_0(c53_270_io_out_0),
    .io_out_1(c53_270_io_out_1),
    .io_out_2(c53_270_io_out_2)
  );
  C53 c53_271 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_271_io_in_0),
    .io_in_1(c53_271_io_in_1),
    .io_in_2(c53_271_io_in_2),
    .io_in_3(c53_271_io_in_3),
    .io_in_4(c53_271_io_in_4),
    .io_out_0(c53_271_io_out_0),
    .io_out_1(c53_271_io_out_1),
    .io_out_2(c53_271_io_out_2)
  );
  C53 c53_272 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_272_io_in_0),
    .io_in_1(c53_272_io_in_1),
    .io_in_2(c53_272_io_in_2),
    .io_in_3(c53_272_io_in_3),
    .io_in_4(c53_272_io_in_4),
    .io_out_0(c53_272_io_out_0),
    .io_out_1(c53_272_io_out_1),
    .io_out_2(c53_272_io_out_2)
  );
  C53 c53_273 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_273_io_in_0),
    .io_in_1(c53_273_io_in_1),
    .io_in_2(c53_273_io_in_2),
    .io_in_3(c53_273_io_in_3),
    .io_in_4(c53_273_io_in_4),
    .io_out_0(c53_273_io_out_0),
    .io_out_1(c53_273_io_out_1),
    .io_out_2(c53_273_io_out_2)
  );
  C53 c53_274 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_274_io_in_0),
    .io_in_1(c53_274_io_in_1),
    .io_in_2(c53_274_io_in_2),
    .io_in_3(c53_274_io_in_3),
    .io_in_4(c53_274_io_in_4),
    .io_out_0(c53_274_io_out_0),
    .io_out_1(c53_274_io_out_1),
    .io_out_2(c53_274_io_out_2)
  );
  C53 c53_275 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_275_io_in_0),
    .io_in_1(c53_275_io_in_1),
    .io_in_2(c53_275_io_in_2),
    .io_in_3(c53_275_io_in_3),
    .io_in_4(c53_275_io_in_4),
    .io_out_0(c53_275_io_out_0),
    .io_out_1(c53_275_io_out_1),
    .io_out_2(c53_275_io_out_2)
  );
  C53 c53_276 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_276_io_in_0),
    .io_in_1(c53_276_io_in_1),
    .io_in_2(c53_276_io_in_2),
    .io_in_3(c53_276_io_in_3),
    .io_in_4(c53_276_io_in_4),
    .io_out_0(c53_276_io_out_0),
    .io_out_1(c53_276_io_out_1),
    .io_out_2(c53_276_io_out_2)
  );
  C53 c53_277 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_277_io_in_0),
    .io_in_1(c53_277_io_in_1),
    .io_in_2(c53_277_io_in_2),
    .io_in_3(c53_277_io_in_3),
    .io_in_4(c53_277_io_in_4),
    .io_out_0(c53_277_io_out_0),
    .io_out_1(c53_277_io_out_1),
    .io_out_2(c53_277_io_out_2)
  );
  C32 c32_22 ( // @[Multiplier.scala 78:25]
    .io_in_0(c32_22_io_in_0),
    .io_in_1(c32_22_io_in_1),
    .io_in_2(c32_22_io_in_2),
    .io_out_0(c32_22_io_out_0),
    .io_out_1(c32_22_io_out_1)
  );
  C53 c53_278 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_278_io_in_0),
    .io_in_1(c53_278_io_in_1),
    .io_in_2(c53_278_io_in_2),
    .io_in_3(c53_278_io_in_3),
    .io_in_4(c53_278_io_in_4),
    .io_out_0(c53_278_io_out_0),
    .io_out_1(c53_278_io_out_1),
    .io_out_2(c53_278_io_out_2)
  );
  C53 c53_279 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_279_io_in_0),
    .io_in_1(c53_279_io_in_1),
    .io_in_2(c53_279_io_in_2),
    .io_in_3(c53_279_io_in_3),
    .io_in_4(c53_279_io_in_4),
    .io_out_0(c53_279_io_out_0),
    .io_out_1(c53_279_io_out_1),
    .io_out_2(c53_279_io_out_2)
  );
  C53 c53_280 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_280_io_in_0),
    .io_in_1(c53_280_io_in_1),
    .io_in_2(c53_280_io_in_2),
    .io_in_3(c53_280_io_in_3),
    .io_in_4(c53_280_io_in_4),
    .io_out_0(c53_280_io_out_0),
    .io_out_1(c53_280_io_out_1),
    .io_out_2(c53_280_io_out_2)
  );
  C53 c53_281 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_281_io_in_0),
    .io_in_1(c53_281_io_in_1),
    .io_in_2(c53_281_io_in_2),
    .io_in_3(c53_281_io_in_3),
    .io_in_4(c53_281_io_in_4),
    .io_out_0(c53_281_io_out_0),
    .io_out_1(c53_281_io_out_1),
    .io_out_2(c53_281_io_out_2)
  );
  C32 c32_23 ( // @[Multiplier.scala 78:25]
    .io_in_0(c32_23_io_in_0),
    .io_in_1(c32_23_io_in_1),
    .io_in_2(c32_23_io_in_2),
    .io_out_0(c32_23_io_out_0),
    .io_out_1(c32_23_io_out_1)
  );
  C53 c53_282 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_282_io_in_0),
    .io_in_1(c53_282_io_in_1),
    .io_in_2(c53_282_io_in_2),
    .io_in_3(c53_282_io_in_3),
    .io_in_4(c53_282_io_in_4),
    .io_out_0(c53_282_io_out_0),
    .io_out_1(c53_282_io_out_1),
    .io_out_2(c53_282_io_out_2)
  );
  C53 c53_283 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_283_io_in_0),
    .io_in_1(c53_283_io_in_1),
    .io_in_2(c53_283_io_in_2),
    .io_in_3(c53_283_io_in_3),
    .io_in_4(c53_283_io_in_4),
    .io_out_0(c53_283_io_out_0),
    .io_out_1(c53_283_io_out_1),
    .io_out_2(c53_283_io_out_2)
  );
  C53 c53_284 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_284_io_in_0),
    .io_in_1(c53_284_io_in_1),
    .io_in_2(c53_284_io_in_2),
    .io_in_3(c53_284_io_in_3),
    .io_in_4(c53_284_io_in_4),
    .io_out_0(c53_284_io_out_0),
    .io_out_1(c53_284_io_out_1),
    .io_out_2(c53_284_io_out_2)
  );
  C53 c53_285 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_285_io_in_0),
    .io_in_1(c53_285_io_in_1),
    .io_in_2(c53_285_io_in_2),
    .io_in_3(c53_285_io_in_3),
    .io_in_4(c53_285_io_in_4),
    .io_out_0(c53_285_io_out_0),
    .io_out_1(c53_285_io_out_1),
    .io_out_2(c53_285_io_out_2)
  );
  C22 c22_17 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_17_io_in_0),
    .io_in_1(c22_17_io_in_1),
    .io_out_0(c22_17_io_out_0),
    .io_out_1(c22_17_io_out_1)
  );
  C53 c53_286 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_286_io_in_0),
    .io_in_1(c53_286_io_in_1),
    .io_in_2(c53_286_io_in_2),
    .io_in_3(c53_286_io_in_3),
    .io_in_4(c53_286_io_in_4),
    .io_out_0(c53_286_io_out_0),
    .io_out_1(c53_286_io_out_1),
    .io_out_2(c53_286_io_out_2)
  );
  C53 c53_287 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_287_io_in_0),
    .io_in_1(c53_287_io_in_1),
    .io_in_2(c53_287_io_in_2),
    .io_in_3(c53_287_io_in_3),
    .io_in_4(c53_287_io_in_4),
    .io_out_0(c53_287_io_out_0),
    .io_out_1(c53_287_io_out_1),
    .io_out_2(c53_287_io_out_2)
  );
  C53 c53_288 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_288_io_in_0),
    .io_in_1(c53_288_io_in_1),
    .io_in_2(c53_288_io_in_2),
    .io_in_3(c53_288_io_in_3),
    .io_in_4(c53_288_io_in_4),
    .io_out_0(c53_288_io_out_0),
    .io_out_1(c53_288_io_out_1),
    .io_out_2(c53_288_io_out_2)
  );
  C53 c53_289 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_289_io_in_0),
    .io_in_1(c53_289_io_in_1),
    .io_in_2(c53_289_io_in_2),
    .io_in_3(c53_289_io_in_3),
    .io_in_4(c53_289_io_in_4),
    .io_out_0(c53_289_io_out_0),
    .io_out_1(c53_289_io_out_1),
    .io_out_2(c53_289_io_out_2)
  );
  C22 c22_18 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_18_io_in_0),
    .io_in_1(c22_18_io_in_1),
    .io_out_0(c22_18_io_out_0),
    .io_out_1(c22_18_io_out_1)
  );
  C53 c53_290 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_290_io_in_0),
    .io_in_1(c53_290_io_in_1),
    .io_in_2(c53_290_io_in_2),
    .io_in_3(c53_290_io_in_3),
    .io_in_4(c53_290_io_in_4),
    .io_out_0(c53_290_io_out_0),
    .io_out_1(c53_290_io_out_1),
    .io_out_2(c53_290_io_out_2)
  );
  C53 c53_291 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_291_io_in_0),
    .io_in_1(c53_291_io_in_1),
    .io_in_2(c53_291_io_in_2),
    .io_in_3(c53_291_io_in_3),
    .io_in_4(c53_291_io_in_4),
    .io_out_0(c53_291_io_out_0),
    .io_out_1(c53_291_io_out_1),
    .io_out_2(c53_291_io_out_2)
  );
  C53 c53_292 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_292_io_in_0),
    .io_in_1(c53_292_io_in_1),
    .io_in_2(c53_292_io_in_2),
    .io_in_3(c53_292_io_in_3),
    .io_in_4(c53_292_io_in_4),
    .io_out_0(c53_292_io_out_0),
    .io_out_1(c53_292_io_out_1),
    .io_out_2(c53_292_io_out_2)
  );
  C53 c53_293 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_293_io_in_0),
    .io_in_1(c53_293_io_in_1),
    .io_in_2(c53_293_io_in_2),
    .io_in_3(c53_293_io_in_3),
    .io_in_4(c53_293_io_in_4),
    .io_out_0(c53_293_io_out_0),
    .io_out_1(c53_293_io_out_1),
    .io_out_2(c53_293_io_out_2)
  );
  C53 c53_294 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_294_io_in_0),
    .io_in_1(c53_294_io_in_1),
    .io_in_2(c53_294_io_in_2),
    .io_in_3(c53_294_io_in_3),
    .io_in_4(c53_294_io_in_4),
    .io_out_0(c53_294_io_out_0),
    .io_out_1(c53_294_io_out_1),
    .io_out_2(c53_294_io_out_2)
  );
  C53 c53_295 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_295_io_in_0),
    .io_in_1(c53_295_io_in_1),
    .io_in_2(c53_295_io_in_2),
    .io_in_3(c53_295_io_in_3),
    .io_in_4(c53_295_io_in_4),
    .io_out_0(c53_295_io_out_0),
    .io_out_1(c53_295_io_out_1),
    .io_out_2(c53_295_io_out_2)
  );
  C53 c53_296 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_296_io_in_0),
    .io_in_1(c53_296_io_in_1),
    .io_in_2(c53_296_io_in_2),
    .io_in_3(c53_296_io_in_3),
    .io_in_4(c53_296_io_in_4),
    .io_out_0(c53_296_io_out_0),
    .io_out_1(c53_296_io_out_1),
    .io_out_2(c53_296_io_out_2)
  );
  C53 c53_297 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_297_io_in_0),
    .io_in_1(c53_297_io_in_1),
    .io_in_2(c53_297_io_in_2),
    .io_in_3(c53_297_io_in_3),
    .io_in_4(c53_297_io_in_4),
    .io_out_0(c53_297_io_out_0),
    .io_out_1(c53_297_io_out_1),
    .io_out_2(c53_297_io_out_2)
  );
  C53 c53_298 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_298_io_in_0),
    .io_in_1(c53_298_io_in_1),
    .io_in_2(c53_298_io_in_2),
    .io_in_3(c53_298_io_in_3),
    .io_in_4(c53_298_io_in_4),
    .io_out_0(c53_298_io_out_0),
    .io_out_1(c53_298_io_out_1),
    .io_out_2(c53_298_io_out_2)
  );
  C53 c53_299 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_299_io_in_0),
    .io_in_1(c53_299_io_in_1),
    .io_in_2(c53_299_io_in_2),
    .io_in_3(c53_299_io_in_3),
    .io_in_4(c53_299_io_in_4),
    .io_out_0(c53_299_io_out_0),
    .io_out_1(c53_299_io_out_1),
    .io_out_2(c53_299_io_out_2)
  );
  C53 c53_300 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_300_io_in_0),
    .io_in_1(c53_300_io_in_1),
    .io_in_2(c53_300_io_in_2),
    .io_in_3(c53_300_io_in_3),
    .io_in_4(c53_300_io_in_4),
    .io_out_0(c53_300_io_out_0),
    .io_out_1(c53_300_io_out_1),
    .io_out_2(c53_300_io_out_2)
  );
  C53 c53_301 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_301_io_in_0),
    .io_in_1(c53_301_io_in_1),
    .io_in_2(c53_301_io_in_2),
    .io_in_3(c53_301_io_in_3),
    .io_in_4(c53_301_io_in_4),
    .io_out_0(c53_301_io_out_0),
    .io_out_1(c53_301_io_out_1),
    .io_out_2(c53_301_io_out_2)
  );
  C53 c53_302 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_302_io_in_0),
    .io_in_1(c53_302_io_in_1),
    .io_in_2(c53_302_io_in_2),
    .io_in_3(c53_302_io_in_3),
    .io_in_4(c53_302_io_in_4),
    .io_out_0(c53_302_io_out_0),
    .io_out_1(c53_302_io_out_1),
    .io_out_2(c53_302_io_out_2)
  );
  C53 c53_303 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_303_io_in_0),
    .io_in_1(c53_303_io_in_1),
    .io_in_2(c53_303_io_in_2),
    .io_in_3(c53_303_io_in_3),
    .io_in_4(c53_303_io_in_4),
    .io_out_0(c53_303_io_out_0),
    .io_out_1(c53_303_io_out_1),
    .io_out_2(c53_303_io_out_2)
  );
  C53 c53_304 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_304_io_in_0),
    .io_in_1(c53_304_io_in_1),
    .io_in_2(c53_304_io_in_2),
    .io_in_3(c53_304_io_in_3),
    .io_in_4(c53_304_io_in_4),
    .io_out_0(c53_304_io_out_0),
    .io_out_1(c53_304_io_out_1),
    .io_out_2(c53_304_io_out_2)
  );
  C53 c53_305 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_305_io_in_0),
    .io_in_1(c53_305_io_in_1),
    .io_in_2(c53_305_io_in_2),
    .io_in_3(c53_305_io_in_3),
    .io_in_4(c53_305_io_in_4),
    .io_out_0(c53_305_io_out_0),
    .io_out_1(c53_305_io_out_1),
    .io_out_2(c53_305_io_out_2)
  );
  C53 c53_306 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_306_io_in_0),
    .io_in_1(c53_306_io_in_1),
    .io_in_2(c53_306_io_in_2),
    .io_in_3(c53_306_io_in_3),
    .io_in_4(c53_306_io_in_4),
    .io_out_0(c53_306_io_out_0),
    .io_out_1(c53_306_io_out_1),
    .io_out_2(c53_306_io_out_2)
  );
  C53 c53_307 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_307_io_in_0),
    .io_in_1(c53_307_io_in_1),
    .io_in_2(c53_307_io_in_2),
    .io_in_3(c53_307_io_in_3),
    .io_in_4(c53_307_io_in_4),
    .io_out_0(c53_307_io_out_0),
    .io_out_1(c53_307_io_out_1),
    .io_out_2(c53_307_io_out_2)
  );
  C53 c53_308 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_308_io_in_0),
    .io_in_1(c53_308_io_in_1),
    .io_in_2(c53_308_io_in_2),
    .io_in_3(c53_308_io_in_3),
    .io_in_4(c53_308_io_in_4),
    .io_out_0(c53_308_io_out_0),
    .io_out_1(c53_308_io_out_1),
    .io_out_2(c53_308_io_out_2)
  );
  C32 c32_24 ( // @[Multiplier.scala 78:25]
    .io_in_0(c32_24_io_in_0),
    .io_in_1(c32_24_io_in_1),
    .io_in_2(c32_24_io_in_2),
    .io_out_0(c32_24_io_out_0),
    .io_out_1(c32_24_io_out_1)
  );
  C53 c53_309 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_309_io_in_0),
    .io_in_1(c53_309_io_in_1),
    .io_in_2(c53_309_io_in_2),
    .io_in_3(c53_309_io_in_3),
    .io_in_4(c53_309_io_in_4),
    .io_out_0(c53_309_io_out_0),
    .io_out_1(c53_309_io_out_1),
    .io_out_2(c53_309_io_out_2)
  );
  C53 c53_310 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_310_io_in_0),
    .io_in_1(c53_310_io_in_1),
    .io_in_2(c53_310_io_in_2),
    .io_in_3(c53_310_io_in_3),
    .io_in_4(c53_310_io_in_4),
    .io_out_0(c53_310_io_out_0),
    .io_out_1(c53_310_io_out_1),
    .io_out_2(c53_310_io_out_2)
  );
  C53 c53_311 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_311_io_in_0),
    .io_in_1(c53_311_io_in_1),
    .io_in_2(c53_311_io_in_2),
    .io_in_3(c53_311_io_in_3),
    .io_in_4(c53_311_io_in_4),
    .io_out_0(c53_311_io_out_0),
    .io_out_1(c53_311_io_out_1),
    .io_out_2(c53_311_io_out_2)
  );
  C32 c32_25 ( // @[Multiplier.scala 78:25]
    .io_in_0(c32_25_io_in_0),
    .io_in_1(c32_25_io_in_1),
    .io_in_2(c32_25_io_in_2),
    .io_out_0(c32_25_io_out_0),
    .io_out_1(c32_25_io_out_1)
  );
  C53 c53_312 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_312_io_in_0),
    .io_in_1(c53_312_io_in_1),
    .io_in_2(c53_312_io_in_2),
    .io_in_3(c53_312_io_in_3),
    .io_in_4(c53_312_io_in_4),
    .io_out_0(c53_312_io_out_0),
    .io_out_1(c53_312_io_out_1),
    .io_out_2(c53_312_io_out_2)
  );
  C53 c53_313 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_313_io_in_0),
    .io_in_1(c53_313_io_in_1),
    .io_in_2(c53_313_io_in_2),
    .io_in_3(c53_313_io_in_3),
    .io_in_4(c53_313_io_in_4),
    .io_out_0(c53_313_io_out_0),
    .io_out_1(c53_313_io_out_1),
    .io_out_2(c53_313_io_out_2)
  );
  C53 c53_314 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_314_io_in_0),
    .io_in_1(c53_314_io_in_1),
    .io_in_2(c53_314_io_in_2),
    .io_in_3(c53_314_io_in_3),
    .io_in_4(c53_314_io_in_4),
    .io_out_0(c53_314_io_out_0),
    .io_out_1(c53_314_io_out_1),
    .io_out_2(c53_314_io_out_2)
  );
  C22 c22_19 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_19_io_in_0),
    .io_in_1(c22_19_io_in_1),
    .io_out_0(c22_19_io_out_0),
    .io_out_1(c22_19_io_out_1)
  );
  C53 c53_315 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_315_io_in_0),
    .io_in_1(c53_315_io_in_1),
    .io_in_2(c53_315_io_in_2),
    .io_in_3(c53_315_io_in_3),
    .io_in_4(c53_315_io_in_4),
    .io_out_0(c53_315_io_out_0),
    .io_out_1(c53_315_io_out_1),
    .io_out_2(c53_315_io_out_2)
  );
  C53 c53_316 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_316_io_in_0),
    .io_in_1(c53_316_io_in_1),
    .io_in_2(c53_316_io_in_2),
    .io_in_3(c53_316_io_in_3),
    .io_in_4(c53_316_io_in_4),
    .io_out_0(c53_316_io_out_0),
    .io_out_1(c53_316_io_out_1),
    .io_out_2(c53_316_io_out_2)
  );
  C53 c53_317 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_317_io_in_0),
    .io_in_1(c53_317_io_in_1),
    .io_in_2(c53_317_io_in_2),
    .io_in_3(c53_317_io_in_3),
    .io_in_4(c53_317_io_in_4),
    .io_out_0(c53_317_io_out_0),
    .io_out_1(c53_317_io_out_1),
    .io_out_2(c53_317_io_out_2)
  );
  C22 c22_20 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_20_io_in_0),
    .io_in_1(c22_20_io_in_1),
    .io_out_0(c22_20_io_out_0),
    .io_out_1(c22_20_io_out_1)
  );
  C53 c53_318 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_318_io_in_0),
    .io_in_1(c53_318_io_in_1),
    .io_in_2(c53_318_io_in_2),
    .io_in_3(c53_318_io_in_3),
    .io_in_4(c53_318_io_in_4),
    .io_out_0(c53_318_io_out_0),
    .io_out_1(c53_318_io_out_1),
    .io_out_2(c53_318_io_out_2)
  );
  C53 c53_319 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_319_io_in_0),
    .io_in_1(c53_319_io_in_1),
    .io_in_2(c53_319_io_in_2),
    .io_in_3(c53_319_io_in_3),
    .io_in_4(c53_319_io_in_4),
    .io_out_0(c53_319_io_out_0),
    .io_out_1(c53_319_io_out_1),
    .io_out_2(c53_319_io_out_2)
  );
  C53 c53_320 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_320_io_in_0),
    .io_in_1(c53_320_io_in_1),
    .io_in_2(c53_320_io_in_2),
    .io_in_3(c53_320_io_in_3),
    .io_in_4(c53_320_io_in_4),
    .io_out_0(c53_320_io_out_0),
    .io_out_1(c53_320_io_out_1),
    .io_out_2(c53_320_io_out_2)
  );
  C53 c53_321 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_321_io_in_0),
    .io_in_1(c53_321_io_in_1),
    .io_in_2(c53_321_io_in_2),
    .io_in_3(c53_321_io_in_3),
    .io_in_4(c53_321_io_in_4),
    .io_out_0(c53_321_io_out_0),
    .io_out_1(c53_321_io_out_1),
    .io_out_2(c53_321_io_out_2)
  );
  C53 c53_322 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_322_io_in_0),
    .io_in_1(c53_322_io_in_1),
    .io_in_2(c53_322_io_in_2),
    .io_in_3(c53_322_io_in_3),
    .io_in_4(c53_322_io_in_4),
    .io_out_0(c53_322_io_out_0),
    .io_out_1(c53_322_io_out_1),
    .io_out_2(c53_322_io_out_2)
  );
  C53 c53_323 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_323_io_in_0),
    .io_in_1(c53_323_io_in_1),
    .io_in_2(c53_323_io_in_2),
    .io_in_3(c53_323_io_in_3),
    .io_in_4(c53_323_io_in_4),
    .io_out_0(c53_323_io_out_0),
    .io_out_1(c53_323_io_out_1),
    .io_out_2(c53_323_io_out_2)
  );
  C53 c53_324 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_324_io_in_0),
    .io_in_1(c53_324_io_in_1),
    .io_in_2(c53_324_io_in_2),
    .io_in_3(c53_324_io_in_3),
    .io_in_4(c53_324_io_in_4),
    .io_out_0(c53_324_io_out_0),
    .io_out_1(c53_324_io_out_1),
    .io_out_2(c53_324_io_out_2)
  );
  C53 c53_325 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_325_io_in_0),
    .io_in_1(c53_325_io_in_1),
    .io_in_2(c53_325_io_in_2),
    .io_in_3(c53_325_io_in_3),
    .io_in_4(c53_325_io_in_4),
    .io_out_0(c53_325_io_out_0),
    .io_out_1(c53_325_io_out_1),
    .io_out_2(c53_325_io_out_2)
  );
  C53 c53_326 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_326_io_in_0),
    .io_in_1(c53_326_io_in_1),
    .io_in_2(c53_326_io_in_2),
    .io_in_3(c53_326_io_in_3),
    .io_in_4(c53_326_io_in_4),
    .io_out_0(c53_326_io_out_0),
    .io_out_1(c53_326_io_out_1),
    .io_out_2(c53_326_io_out_2)
  );
  C53 c53_327 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_327_io_in_0),
    .io_in_1(c53_327_io_in_1),
    .io_in_2(c53_327_io_in_2),
    .io_in_3(c53_327_io_in_3),
    .io_in_4(c53_327_io_in_4),
    .io_out_0(c53_327_io_out_0),
    .io_out_1(c53_327_io_out_1),
    .io_out_2(c53_327_io_out_2)
  );
  C53 c53_328 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_328_io_in_0),
    .io_in_1(c53_328_io_in_1),
    .io_in_2(c53_328_io_in_2),
    .io_in_3(c53_328_io_in_3),
    .io_in_4(c53_328_io_in_4),
    .io_out_0(c53_328_io_out_0),
    .io_out_1(c53_328_io_out_1),
    .io_out_2(c53_328_io_out_2)
  );
  C53 c53_329 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_329_io_in_0),
    .io_in_1(c53_329_io_in_1),
    .io_in_2(c53_329_io_in_2),
    .io_in_3(c53_329_io_in_3),
    .io_in_4(c53_329_io_in_4),
    .io_out_0(c53_329_io_out_0),
    .io_out_1(c53_329_io_out_1),
    .io_out_2(c53_329_io_out_2)
  );
  C53 c53_330 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_330_io_in_0),
    .io_in_1(c53_330_io_in_1),
    .io_in_2(c53_330_io_in_2),
    .io_in_3(c53_330_io_in_3),
    .io_in_4(c53_330_io_in_4),
    .io_out_0(c53_330_io_out_0),
    .io_out_1(c53_330_io_out_1),
    .io_out_2(c53_330_io_out_2)
  );
  C53 c53_331 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_331_io_in_0),
    .io_in_1(c53_331_io_in_1),
    .io_in_2(c53_331_io_in_2),
    .io_in_3(c53_331_io_in_3),
    .io_in_4(c53_331_io_in_4),
    .io_out_0(c53_331_io_out_0),
    .io_out_1(c53_331_io_out_1),
    .io_out_2(c53_331_io_out_2)
  );
  C32 c32_26 ( // @[Multiplier.scala 78:25]
    .io_in_0(c32_26_io_in_0),
    .io_in_1(c32_26_io_in_1),
    .io_in_2(c32_26_io_in_2),
    .io_out_0(c32_26_io_out_0),
    .io_out_1(c32_26_io_out_1)
  );
  C53 c53_332 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_332_io_in_0),
    .io_in_1(c53_332_io_in_1),
    .io_in_2(c53_332_io_in_2),
    .io_in_3(c53_332_io_in_3),
    .io_in_4(c53_332_io_in_4),
    .io_out_0(c53_332_io_out_0),
    .io_out_1(c53_332_io_out_1),
    .io_out_2(c53_332_io_out_2)
  );
  C53 c53_333 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_333_io_in_0),
    .io_in_1(c53_333_io_in_1),
    .io_in_2(c53_333_io_in_2),
    .io_in_3(c53_333_io_in_3),
    .io_in_4(c53_333_io_in_4),
    .io_out_0(c53_333_io_out_0),
    .io_out_1(c53_333_io_out_1),
    .io_out_2(c53_333_io_out_2)
  );
  C32 c32_27 ( // @[Multiplier.scala 78:25]
    .io_in_0(c32_27_io_in_0),
    .io_in_1(c32_27_io_in_1),
    .io_in_2(c32_27_io_in_2),
    .io_out_0(c32_27_io_out_0),
    .io_out_1(c32_27_io_out_1)
  );
  C53 c53_334 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_334_io_in_0),
    .io_in_1(c53_334_io_in_1),
    .io_in_2(c53_334_io_in_2),
    .io_in_3(c53_334_io_in_3),
    .io_in_4(c53_334_io_in_4),
    .io_out_0(c53_334_io_out_0),
    .io_out_1(c53_334_io_out_1),
    .io_out_2(c53_334_io_out_2)
  );
  C53 c53_335 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_335_io_in_0),
    .io_in_1(c53_335_io_in_1),
    .io_in_2(c53_335_io_in_2),
    .io_in_3(c53_335_io_in_3),
    .io_in_4(c53_335_io_in_4),
    .io_out_0(c53_335_io_out_0),
    .io_out_1(c53_335_io_out_1),
    .io_out_2(c53_335_io_out_2)
  );
  C22 c22_21 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_21_io_in_0),
    .io_in_1(c22_21_io_in_1),
    .io_out_0(c22_21_io_out_0),
    .io_out_1(c22_21_io_out_1)
  );
  C53 c53_336 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_336_io_in_0),
    .io_in_1(c53_336_io_in_1),
    .io_in_2(c53_336_io_in_2),
    .io_in_3(c53_336_io_in_3),
    .io_in_4(c53_336_io_in_4),
    .io_out_0(c53_336_io_out_0),
    .io_out_1(c53_336_io_out_1),
    .io_out_2(c53_336_io_out_2)
  );
  C53 c53_337 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_337_io_in_0),
    .io_in_1(c53_337_io_in_1),
    .io_in_2(c53_337_io_in_2),
    .io_in_3(c53_337_io_in_3),
    .io_in_4(c53_337_io_in_4),
    .io_out_0(c53_337_io_out_0),
    .io_out_1(c53_337_io_out_1),
    .io_out_2(c53_337_io_out_2)
  );
  C22 c22_22 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_22_io_in_0),
    .io_in_1(c22_22_io_in_1),
    .io_out_0(c22_22_io_out_0),
    .io_out_1(c22_22_io_out_1)
  );
  C53 c53_338 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_338_io_in_0),
    .io_in_1(c53_338_io_in_1),
    .io_in_2(c53_338_io_in_2),
    .io_in_3(c53_338_io_in_3),
    .io_in_4(c53_338_io_in_4),
    .io_out_0(c53_338_io_out_0),
    .io_out_1(c53_338_io_out_1),
    .io_out_2(c53_338_io_out_2)
  );
  C53 c53_339 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_339_io_in_0),
    .io_in_1(c53_339_io_in_1),
    .io_in_2(c53_339_io_in_2),
    .io_in_3(c53_339_io_in_3),
    .io_in_4(c53_339_io_in_4),
    .io_out_0(c53_339_io_out_0),
    .io_out_1(c53_339_io_out_1),
    .io_out_2(c53_339_io_out_2)
  );
  C53 c53_340 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_340_io_in_0),
    .io_in_1(c53_340_io_in_1),
    .io_in_2(c53_340_io_in_2),
    .io_in_3(c53_340_io_in_3),
    .io_in_4(c53_340_io_in_4),
    .io_out_0(c53_340_io_out_0),
    .io_out_1(c53_340_io_out_1),
    .io_out_2(c53_340_io_out_2)
  );
  C53 c53_341 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_341_io_in_0),
    .io_in_1(c53_341_io_in_1),
    .io_in_2(c53_341_io_in_2),
    .io_in_3(c53_341_io_in_3),
    .io_in_4(c53_341_io_in_4),
    .io_out_0(c53_341_io_out_0),
    .io_out_1(c53_341_io_out_1),
    .io_out_2(c53_341_io_out_2)
  );
  C53 c53_342 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_342_io_in_0),
    .io_in_1(c53_342_io_in_1),
    .io_in_2(c53_342_io_in_2),
    .io_in_3(c53_342_io_in_3),
    .io_in_4(c53_342_io_in_4),
    .io_out_0(c53_342_io_out_0),
    .io_out_1(c53_342_io_out_1),
    .io_out_2(c53_342_io_out_2)
  );
  C53 c53_343 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_343_io_in_0),
    .io_in_1(c53_343_io_in_1),
    .io_in_2(c53_343_io_in_2),
    .io_in_3(c53_343_io_in_3),
    .io_in_4(c53_343_io_in_4),
    .io_out_0(c53_343_io_out_0),
    .io_out_1(c53_343_io_out_1),
    .io_out_2(c53_343_io_out_2)
  );
  C53 c53_344 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_344_io_in_0),
    .io_in_1(c53_344_io_in_1),
    .io_in_2(c53_344_io_in_2),
    .io_in_3(c53_344_io_in_3),
    .io_in_4(c53_344_io_in_4),
    .io_out_0(c53_344_io_out_0),
    .io_out_1(c53_344_io_out_1),
    .io_out_2(c53_344_io_out_2)
  );
  C53 c53_345 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_345_io_in_0),
    .io_in_1(c53_345_io_in_1),
    .io_in_2(c53_345_io_in_2),
    .io_in_3(c53_345_io_in_3),
    .io_in_4(c53_345_io_in_4),
    .io_out_0(c53_345_io_out_0),
    .io_out_1(c53_345_io_out_1),
    .io_out_2(c53_345_io_out_2)
  );
  C53 c53_346 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_346_io_in_0),
    .io_in_1(c53_346_io_in_1),
    .io_in_2(c53_346_io_in_2),
    .io_in_3(c53_346_io_in_3),
    .io_in_4(c53_346_io_in_4),
    .io_out_0(c53_346_io_out_0),
    .io_out_1(c53_346_io_out_1),
    .io_out_2(c53_346_io_out_2)
  );
  C32 c32_28 ( // @[Multiplier.scala 78:25]
    .io_in_0(c32_28_io_in_0),
    .io_in_1(c32_28_io_in_1),
    .io_in_2(c32_28_io_in_2),
    .io_out_0(c32_28_io_out_0),
    .io_out_1(c32_28_io_out_1)
  );
  C53 c53_347 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_347_io_in_0),
    .io_in_1(c53_347_io_in_1),
    .io_in_2(c53_347_io_in_2),
    .io_in_3(c53_347_io_in_3),
    .io_in_4(c53_347_io_in_4),
    .io_out_0(c53_347_io_out_0),
    .io_out_1(c53_347_io_out_1),
    .io_out_2(c53_347_io_out_2)
  );
  C32 c32_29 ( // @[Multiplier.scala 78:25]
    .io_in_0(c32_29_io_in_0),
    .io_in_1(c32_29_io_in_1),
    .io_in_2(c32_29_io_in_2),
    .io_out_0(c32_29_io_out_0),
    .io_out_1(c32_29_io_out_1)
  );
  C53 c53_348 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_348_io_in_0),
    .io_in_1(c53_348_io_in_1),
    .io_in_2(c53_348_io_in_2),
    .io_in_3(c53_348_io_in_3),
    .io_in_4(c53_348_io_in_4),
    .io_out_0(c53_348_io_out_0),
    .io_out_1(c53_348_io_out_1),
    .io_out_2(c53_348_io_out_2)
  );
  C22 c22_23 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_23_io_in_0),
    .io_in_1(c22_23_io_in_1),
    .io_out_0(c22_23_io_out_0),
    .io_out_1(c22_23_io_out_1)
  );
  C53 c53_349 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_349_io_in_0),
    .io_in_1(c53_349_io_in_1),
    .io_in_2(c53_349_io_in_2),
    .io_in_3(c53_349_io_in_3),
    .io_in_4(c53_349_io_in_4),
    .io_out_0(c53_349_io_out_0),
    .io_out_1(c53_349_io_out_1),
    .io_out_2(c53_349_io_out_2)
  );
  C22 c22_24 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_24_io_in_0),
    .io_in_1(c22_24_io_in_1),
    .io_out_0(c22_24_io_out_0),
    .io_out_1(c22_24_io_out_1)
  );
  C53 c53_350 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_350_io_in_0),
    .io_in_1(c53_350_io_in_1),
    .io_in_2(c53_350_io_in_2),
    .io_in_3(c53_350_io_in_3),
    .io_in_4(c53_350_io_in_4),
    .io_out_0(c53_350_io_out_0),
    .io_out_1(c53_350_io_out_1),
    .io_out_2(c53_350_io_out_2)
  );
  C53 c53_351 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_351_io_in_0),
    .io_in_1(c53_351_io_in_1),
    .io_in_2(c53_351_io_in_2),
    .io_in_3(c53_351_io_in_3),
    .io_in_4(c53_351_io_in_4),
    .io_out_0(c53_351_io_out_0),
    .io_out_1(c53_351_io_out_1),
    .io_out_2(c53_351_io_out_2)
  );
  C53 c53_352 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_352_io_in_0),
    .io_in_1(c53_352_io_in_1),
    .io_in_2(c53_352_io_in_2),
    .io_in_3(c53_352_io_in_3),
    .io_in_4(c53_352_io_in_4),
    .io_out_0(c53_352_io_out_0),
    .io_out_1(c53_352_io_out_1),
    .io_out_2(c53_352_io_out_2)
  );
  C53 c53_353 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_353_io_in_0),
    .io_in_1(c53_353_io_in_1),
    .io_in_2(c53_353_io_in_2),
    .io_in_3(c53_353_io_in_3),
    .io_in_4(c53_353_io_in_4),
    .io_out_0(c53_353_io_out_0),
    .io_out_1(c53_353_io_out_1),
    .io_out_2(c53_353_io_out_2)
  );
  C32 c32_30 ( // @[Multiplier.scala 78:25]
    .io_in_0(c32_30_io_in_0),
    .io_in_1(c32_30_io_in_1),
    .io_in_2(c32_30_io_in_2),
    .io_out_0(c32_30_io_out_0),
    .io_out_1(c32_30_io_out_1)
  );
  C32 c32_31 ( // @[Multiplier.scala 78:25]
    .io_in_0(c32_31_io_in_0),
    .io_in_1(c32_31_io_in_1),
    .io_in_2(c32_31_io_in_2),
    .io_out_0(c32_31_io_out_0),
    .io_out_1(c32_31_io_out_1)
  );
  C22 c22_25 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_25_io_in_0),
    .io_in_1(c22_25_io_in_1),
    .io_out_0(c22_25_io_out_0),
    .io_out_1(c22_25_io_out_1)
  );
  C22 c22_26 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_26_io_in_0),
    .io_in_1(c22_26_io_in_1),
    .io_out_0(c22_26_io_out_0),
    .io_out_1(c22_26_io_out_1)
  );
  C22 c22_27 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_27_io_in_0),
    .io_in_1(c22_27_io_in_1),
    .io_out_0(c22_27_io_out_0),
    .io_out_1(c22_27_io_out_1)
  );
  C22 c22_28 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_28_io_in_0),
    .io_in_1(c22_28_io_in_1),
    .io_out_0(c22_28_io_out_0),
    .io_out_1(c22_28_io_out_1)
  );
  C22 c22_29 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_29_io_in_0),
    .io_in_1(c22_29_io_in_1),
    .io_out_0(c22_29_io_out_0),
    .io_out_1(c22_29_io_out_1)
  );
  C22 c22_30 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_30_io_in_0),
    .io_in_1(c22_30_io_in_1),
    .io_out_0(c22_30_io_out_0),
    .io_out_1(c22_30_io_out_1)
  );
  C22 c22_31 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_31_io_in_0),
    .io_in_1(c22_31_io_in_1),
    .io_out_0(c22_31_io_out_0),
    .io_out_1(c22_31_io_out_1)
  );
  C32 c32_32 ( // @[Multiplier.scala 78:25]
    .io_in_0(c32_32_io_in_0),
    .io_in_1(c32_32_io_in_1),
    .io_in_2(c32_32_io_in_2),
    .io_out_0(c32_32_io_out_0),
    .io_out_1(c32_32_io_out_1)
  );
  C32 c32_33 ( // @[Multiplier.scala 78:25]
    .io_in_0(c32_33_io_in_0),
    .io_in_1(c32_33_io_in_1),
    .io_in_2(c32_33_io_in_2),
    .io_out_0(c32_33_io_out_0),
    .io_out_1(c32_33_io_out_1)
  );
  C32 c32_34 ( // @[Multiplier.scala 78:25]
    .io_in_0(c32_34_io_in_0),
    .io_in_1(c32_34_io_in_1),
    .io_in_2(c32_34_io_in_2),
    .io_out_0(c32_34_io_out_0),
    .io_out_1(c32_34_io_out_1)
  );
  C53 c53_354 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_354_io_in_0),
    .io_in_1(c53_354_io_in_1),
    .io_in_2(c53_354_io_in_2),
    .io_in_3(c53_354_io_in_3),
    .io_in_4(c53_354_io_in_4),
    .io_out_0(c53_354_io_out_0),
    .io_out_1(c53_354_io_out_1),
    .io_out_2(c53_354_io_out_2)
  );
  C53 c53_355 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_355_io_in_0),
    .io_in_1(c53_355_io_in_1),
    .io_in_2(c53_355_io_in_2),
    .io_in_3(c53_355_io_in_3),
    .io_in_4(c53_355_io_in_4),
    .io_out_0(c53_355_io_out_0),
    .io_out_1(c53_355_io_out_1),
    .io_out_2(c53_355_io_out_2)
  );
  C53 c53_356 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_356_io_in_0),
    .io_in_1(c53_356_io_in_1),
    .io_in_2(c53_356_io_in_2),
    .io_in_3(c53_356_io_in_3),
    .io_in_4(c53_356_io_in_4),
    .io_out_0(c53_356_io_out_0),
    .io_out_1(c53_356_io_out_1),
    .io_out_2(c53_356_io_out_2)
  );
  C53 c53_357 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_357_io_in_0),
    .io_in_1(c53_357_io_in_1),
    .io_in_2(c53_357_io_in_2),
    .io_in_3(c53_357_io_in_3),
    .io_in_4(c53_357_io_in_4),
    .io_out_0(c53_357_io_out_0),
    .io_out_1(c53_357_io_out_1),
    .io_out_2(c53_357_io_out_2)
  );
  C53 c53_358 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_358_io_in_0),
    .io_in_1(c53_358_io_in_1),
    .io_in_2(c53_358_io_in_2),
    .io_in_3(c53_358_io_in_3),
    .io_in_4(c53_358_io_in_4),
    .io_out_0(c53_358_io_out_0),
    .io_out_1(c53_358_io_out_1),
    .io_out_2(c53_358_io_out_2)
  );
  C53 c53_359 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_359_io_in_0),
    .io_in_1(c53_359_io_in_1),
    .io_in_2(c53_359_io_in_2),
    .io_in_3(c53_359_io_in_3),
    .io_in_4(c53_359_io_in_4),
    .io_out_0(c53_359_io_out_0),
    .io_out_1(c53_359_io_out_1),
    .io_out_2(c53_359_io_out_2)
  );
  C53 c53_360 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_360_io_in_0),
    .io_in_1(c53_360_io_in_1),
    .io_in_2(c53_360_io_in_2),
    .io_in_3(c53_360_io_in_3),
    .io_in_4(c53_360_io_in_4),
    .io_out_0(c53_360_io_out_0),
    .io_out_1(c53_360_io_out_1),
    .io_out_2(c53_360_io_out_2)
  );
  C53 c53_361 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_361_io_in_0),
    .io_in_1(c53_361_io_in_1),
    .io_in_2(c53_361_io_in_2),
    .io_in_3(c53_361_io_in_3),
    .io_in_4(c53_361_io_in_4),
    .io_out_0(c53_361_io_out_0),
    .io_out_1(c53_361_io_out_1),
    .io_out_2(c53_361_io_out_2)
  );
  C53 c53_362 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_362_io_in_0),
    .io_in_1(c53_362_io_in_1),
    .io_in_2(c53_362_io_in_2),
    .io_in_3(c53_362_io_in_3),
    .io_in_4(c53_362_io_in_4),
    .io_out_0(c53_362_io_out_0),
    .io_out_1(c53_362_io_out_1),
    .io_out_2(c53_362_io_out_2)
  );
  C22 c22_32 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_32_io_in_0),
    .io_in_1(c22_32_io_in_1),
    .io_out_0(c22_32_io_out_0),
    .io_out_1(c22_32_io_out_1)
  );
  C53 c53_363 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_363_io_in_0),
    .io_in_1(c53_363_io_in_1),
    .io_in_2(c53_363_io_in_2),
    .io_in_3(c53_363_io_in_3),
    .io_in_4(c53_363_io_in_4),
    .io_out_0(c53_363_io_out_0),
    .io_out_1(c53_363_io_out_1),
    .io_out_2(c53_363_io_out_2)
  );
  C22 c22_33 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_33_io_in_0),
    .io_in_1(c22_33_io_in_1),
    .io_out_0(c22_33_io_out_0),
    .io_out_1(c22_33_io_out_1)
  );
  C53 c53_364 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_364_io_in_0),
    .io_in_1(c53_364_io_in_1),
    .io_in_2(c53_364_io_in_2),
    .io_in_3(c53_364_io_in_3),
    .io_in_4(c53_364_io_in_4),
    .io_out_0(c53_364_io_out_0),
    .io_out_1(c53_364_io_out_1),
    .io_out_2(c53_364_io_out_2)
  );
  C22 c22_34 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_34_io_in_0),
    .io_in_1(c22_34_io_in_1),
    .io_out_0(c22_34_io_out_0),
    .io_out_1(c22_34_io_out_1)
  );
  C53 c53_365 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_365_io_in_0),
    .io_in_1(c53_365_io_in_1),
    .io_in_2(c53_365_io_in_2),
    .io_in_3(c53_365_io_in_3),
    .io_in_4(c53_365_io_in_4),
    .io_out_0(c53_365_io_out_0),
    .io_out_1(c53_365_io_out_1),
    .io_out_2(c53_365_io_out_2)
  );
  C22 c22_35 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_35_io_in_0),
    .io_in_1(c22_35_io_in_1),
    .io_out_0(c22_35_io_out_0),
    .io_out_1(c22_35_io_out_1)
  );
  C53 c53_366 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_366_io_in_0),
    .io_in_1(c53_366_io_in_1),
    .io_in_2(c53_366_io_in_2),
    .io_in_3(c53_366_io_in_3),
    .io_in_4(c53_366_io_in_4),
    .io_out_0(c53_366_io_out_0),
    .io_out_1(c53_366_io_out_1),
    .io_out_2(c53_366_io_out_2)
  );
  C22 c22_36 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_36_io_in_0),
    .io_in_1(c22_36_io_in_1),
    .io_out_0(c22_36_io_out_0),
    .io_out_1(c22_36_io_out_1)
  );
  C53 c53_367 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_367_io_in_0),
    .io_in_1(c53_367_io_in_1),
    .io_in_2(c53_367_io_in_2),
    .io_in_3(c53_367_io_in_3),
    .io_in_4(c53_367_io_in_4),
    .io_out_0(c53_367_io_out_0),
    .io_out_1(c53_367_io_out_1),
    .io_out_2(c53_367_io_out_2)
  );
  C32 c32_35 ( // @[Multiplier.scala 78:25]
    .io_in_0(c32_35_io_in_0),
    .io_in_1(c32_35_io_in_1),
    .io_in_2(c32_35_io_in_2),
    .io_out_0(c32_35_io_out_0),
    .io_out_1(c32_35_io_out_1)
  );
  C53 c53_368 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_368_io_in_0),
    .io_in_1(c53_368_io_in_1),
    .io_in_2(c53_368_io_in_2),
    .io_in_3(c53_368_io_in_3),
    .io_in_4(c53_368_io_in_4),
    .io_out_0(c53_368_io_out_0),
    .io_out_1(c53_368_io_out_1),
    .io_out_2(c53_368_io_out_2)
  );
  C32 c32_36 ( // @[Multiplier.scala 78:25]
    .io_in_0(c32_36_io_in_0),
    .io_in_1(c32_36_io_in_1),
    .io_in_2(c32_36_io_in_2),
    .io_out_0(c32_36_io_out_0),
    .io_out_1(c32_36_io_out_1)
  );
  C53 c53_369 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_369_io_in_0),
    .io_in_1(c53_369_io_in_1),
    .io_in_2(c53_369_io_in_2),
    .io_in_3(c53_369_io_in_3),
    .io_in_4(c53_369_io_in_4),
    .io_out_0(c53_369_io_out_0),
    .io_out_1(c53_369_io_out_1),
    .io_out_2(c53_369_io_out_2)
  );
  C32 c32_37 ( // @[Multiplier.scala 78:25]
    .io_in_0(c32_37_io_in_0),
    .io_in_1(c32_37_io_in_1),
    .io_in_2(c32_37_io_in_2),
    .io_out_0(c32_37_io_out_0),
    .io_out_1(c32_37_io_out_1)
  );
  C53 c53_370 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_370_io_in_0),
    .io_in_1(c53_370_io_in_1),
    .io_in_2(c53_370_io_in_2),
    .io_in_3(c53_370_io_in_3),
    .io_in_4(c53_370_io_in_4),
    .io_out_0(c53_370_io_out_0),
    .io_out_1(c53_370_io_out_1),
    .io_out_2(c53_370_io_out_2)
  );
  C53 c53_371 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_371_io_in_0),
    .io_in_1(c53_371_io_in_1),
    .io_in_2(c53_371_io_in_2),
    .io_in_3(c53_371_io_in_3),
    .io_in_4(c53_371_io_in_4),
    .io_out_0(c53_371_io_out_0),
    .io_out_1(c53_371_io_out_1),
    .io_out_2(c53_371_io_out_2)
  );
  C53 c53_372 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_372_io_in_0),
    .io_in_1(c53_372_io_in_1),
    .io_in_2(c53_372_io_in_2),
    .io_in_3(c53_372_io_in_3),
    .io_in_4(c53_372_io_in_4),
    .io_out_0(c53_372_io_out_0),
    .io_out_1(c53_372_io_out_1),
    .io_out_2(c53_372_io_out_2)
  );
  C53 c53_373 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_373_io_in_0),
    .io_in_1(c53_373_io_in_1),
    .io_in_2(c53_373_io_in_2),
    .io_in_3(c53_373_io_in_3),
    .io_in_4(c53_373_io_in_4),
    .io_out_0(c53_373_io_out_0),
    .io_out_1(c53_373_io_out_1),
    .io_out_2(c53_373_io_out_2)
  );
  C53 c53_374 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_374_io_in_0),
    .io_in_1(c53_374_io_in_1),
    .io_in_2(c53_374_io_in_2),
    .io_in_3(c53_374_io_in_3),
    .io_in_4(c53_374_io_in_4),
    .io_out_0(c53_374_io_out_0),
    .io_out_1(c53_374_io_out_1),
    .io_out_2(c53_374_io_out_2)
  );
  C53 c53_375 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_375_io_in_0),
    .io_in_1(c53_375_io_in_1),
    .io_in_2(c53_375_io_in_2),
    .io_in_3(c53_375_io_in_3),
    .io_in_4(c53_375_io_in_4),
    .io_out_0(c53_375_io_out_0),
    .io_out_1(c53_375_io_out_1),
    .io_out_2(c53_375_io_out_2)
  );
  C53 c53_376 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_376_io_in_0),
    .io_in_1(c53_376_io_in_1),
    .io_in_2(c53_376_io_in_2),
    .io_in_3(c53_376_io_in_3),
    .io_in_4(c53_376_io_in_4),
    .io_out_0(c53_376_io_out_0),
    .io_out_1(c53_376_io_out_1),
    .io_out_2(c53_376_io_out_2)
  );
  C53 c53_377 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_377_io_in_0),
    .io_in_1(c53_377_io_in_1),
    .io_in_2(c53_377_io_in_2),
    .io_in_3(c53_377_io_in_3),
    .io_in_4(c53_377_io_in_4),
    .io_out_0(c53_377_io_out_0),
    .io_out_1(c53_377_io_out_1),
    .io_out_2(c53_377_io_out_2)
  );
  C53 c53_378 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_378_io_in_0),
    .io_in_1(c53_378_io_in_1),
    .io_in_2(c53_378_io_in_2),
    .io_in_3(c53_378_io_in_3),
    .io_in_4(c53_378_io_in_4),
    .io_out_0(c53_378_io_out_0),
    .io_out_1(c53_378_io_out_1),
    .io_out_2(c53_378_io_out_2)
  );
  C53 c53_379 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_379_io_in_0),
    .io_in_1(c53_379_io_in_1),
    .io_in_2(c53_379_io_in_2),
    .io_in_3(c53_379_io_in_3),
    .io_in_4(c53_379_io_in_4),
    .io_out_0(c53_379_io_out_0),
    .io_out_1(c53_379_io_out_1),
    .io_out_2(c53_379_io_out_2)
  );
  C53 c53_380 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_380_io_in_0),
    .io_in_1(c53_380_io_in_1),
    .io_in_2(c53_380_io_in_2),
    .io_in_3(c53_380_io_in_3),
    .io_in_4(c53_380_io_in_4),
    .io_out_0(c53_380_io_out_0),
    .io_out_1(c53_380_io_out_1),
    .io_out_2(c53_380_io_out_2)
  );
  C53 c53_381 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_381_io_in_0),
    .io_in_1(c53_381_io_in_1),
    .io_in_2(c53_381_io_in_2),
    .io_in_3(c53_381_io_in_3),
    .io_in_4(c53_381_io_in_4),
    .io_out_0(c53_381_io_out_0),
    .io_out_1(c53_381_io_out_1),
    .io_out_2(c53_381_io_out_2)
  );
  C53 c53_382 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_382_io_in_0),
    .io_in_1(c53_382_io_in_1),
    .io_in_2(c53_382_io_in_2),
    .io_in_3(c53_382_io_in_3),
    .io_in_4(c53_382_io_in_4),
    .io_out_0(c53_382_io_out_0),
    .io_out_1(c53_382_io_out_1),
    .io_out_2(c53_382_io_out_2)
  );
  C53 c53_383 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_383_io_in_0),
    .io_in_1(c53_383_io_in_1),
    .io_in_2(c53_383_io_in_2),
    .io_in_3(c53_383_io_in_3),
    .io_in_4(c53_383_io_in_4),
    .io_out_0(c53_383_io_out_0),
    .io_out_1(c53_383_io_out_1),
    .io_out_2(c53_383_io_out_2)
  );
  C53 c53_384 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_384_io_in_0),
    .io_in_1(c53_384_io_in_1),
    .io_in_2(c53_384_io_in_2),
    .io_in_3(c53_384_io_in_3),
    .io_in_4(c53_384_io_in_4),
    .io_out_0(c53_384_io_out_0),
    .io_out_1(c53_384_io_out_1),
    .io_out_2(c53_384_io_out_2)
  );
  C53 c53_385 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_385_io_in_0),
    .io_in_1(c53_385_io_in_1),
    .io_in_2(c53_385_io_in_2),
    .io_in_3(c53_385_io_in_3),
    .io_in_4(c53_385_io_in_4),
    .io_out_0(c53_385_io_out_0),
    .io_out_1(c53_385_io_out_1),
    .io_out_2(c53_385_io_out_2)
  );
  C53 c53_386 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_386_io_in_0),
    .io_in_1(c53_386_io_in_1),
    .io_in_2(c53_386_io_in_2),
    .io_in_3(c53_386_io_in_3),
    .io_in_4(c53_386_io_in_4),
    .io_out_0(c53_386_io_out_0),
    .io_out_1(c53_386_io_out_1),
    .io_out_2(c53_386_io_out_2)
  );
  C53 c53_387 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_387_io_in_0),
    .io_in_1(c53_387_io_in_1),
    .io_in_2(c53_387_io_in_2),
    .io_in_3(c53_387_io_in_3),
    .io_in_4(c53_387_io_in_4),
    .io_out_0(c53_387_io_out_0),
    .io_out_1(c53_387_io_out_1),
    .io_out_2(c53_387_io_out_2)
  );
  C22 c22_37 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_37_io_in_0),
    .io_in_1(c22_37_io_in_1),
    .io_out_0(c22_37_io_out_0),
    .io_out_1(c22_37_io_out_1)
  );
  C53 c53_388 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_388_io_in_0),
    .io_in_1(c53_388_io_in_1),
    .io_in_2(c53_388_io_in_2),
    .io_in_3(c53_388_io_in_3),
    .io_in_4(c53_388_io_in_4),
    .io_out_0(c53_388_io_out_0),
    .io_out_1(c53_388_io_out_1),
    .io_out_2(c53_388_io_out_2)
  );
  C53 c53_389 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_389_io_in_0),
    .io_in_1(c53_389_io_in_1),
    .io_in_2(c53_389_io_in_2),
    .io_in_3(c53_389_io_in_3),
    .io_in_4(c53_389_io_in_4),
    .io_out_0(c53_389_io_out_0),
    .io_out_1(c53_389_io_out_1),
    .io_out_2(c53_389_io_out_2)
  );
  C22 c22_38 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_38_io_in_0),
    .io_in_1(c22_38_io_in_1),
    .io_out_0(c22_38_io_out_0),
    .io_out_1(c22_38_io_out_1)
  );
  C53 c53_390 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_390_io_in_0),
    .io_in_1(c53_390_io_in_1),
    .io_in_2(c53_390_io_in_2),
    .io_in_3(c53_390_io_in_3),
    .io_in_4(c53_390_io_in_4),
    .io_out_0(c53_390_io_out_0),
    .io_out_1(c53_390_io_out_1),
    .io_out_2(c53_390_io_out_2)
  );
  C53 c53_391 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_391_io_in_0),
    .io_in_1(c53_391_io_in_1),
    .io_in_2(c53_391_io_in_2),
    .io_in_3(c53_391_io_in_3),
    .io_in_4(c53_391_io_in_4),
    .io_out_0(c53_391_io_out_0),
    .io_out_1(c53_391_io_out_1),
    .io_out_2(c53_391_io_out_2)
  );
  C22 c22_39 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_39_io_in_0),
    .io_in_1(c22_39_io_in_1),
    .io_out_0(c22_39_io_out_0),
    .io_out_1(c22_39_io_out_1)
  );
  C53 c53_392 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_392_io_in_0),
    .io_in_1(c53_392_io_in_1),
    .io_in_2(c53_392_io_in_2),
    .io_in_3(c53_392_io_in_3),
    .io_in_4(c53_392_io_in_4),
    .io_out_0(c53_392_io_out_0),
    .io_out_1(c53_392_io_out_1),
    .io_out_2(c53_392_io_out_2)
  );
  C53 c53_393 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_393_io_in_0),
    .io_in_1(c53_393_io_in_1),
    .io_in_2(c53_393_io_in_2),
    .io_in_3(c53_393_io_in_3),
    .io_in_4(c53_393_io_in_4),
    .io_out_0(c53_393_io_out_0),
    .io_out_1(c53_393_io_out_1),
    .io_out_2(c53_393_io_out_2)
  );
  C22 c22_40 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_40_io_in_0),
    .io_in_1(c22_40_io_in_1),
    .io_out_0(c22_40_io_out_0),
    .io_out_1(c22_40_io_out_1)
  );
  C53 c53_394 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_394_io_in_0),
    .io_in_1(c53_394_io_in_1),
    .io_in_2(c53_394_io_in_2),
    .io_in_3(c53_394_io_in_3),
    .io_in_4(c53_394_io_in_4),
    .io_out_0(c53_394_io_out_0),
    .io_out_1(c53_394_io_out_1),
    .io_out_2(c53_394_io_out_2)
  );
  C53 c53_395 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_395_io_in_0),
    .io_in_1(c53_395_io_in_1),
    .io_in_2(c53_395_io_in_2),
    .io_in_3(c53_395_io_in_3),
    .io_in_4(c53_395_io_in_4),
    .io_out_0(c53_395_io_out_0),
    .io_out_1(c53_395_io_out_1),
    .io_out_2(c53_395_io_out_2)
  );
  C22 c22_41 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_41_io_in_0),
    .io_in_1(c22_41_io_in_1),
    .io_out_0(c22_41_io_out_0),
    .io_out_1(c22_41_io_out_1)
  );
  C53 c53_396 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_396_io_in_0),
    .io_in_1(c53_396_io_in_1),
    .io_in_2(c53_396_io_in_2),
    .io_in_3(c53_396_io_in_3),
    .io_in_4(c53_396_io_in_4),
    .io_out_0(c53_396_io_out_0),
    .io_out_1(c53_396_io_out_1),
    .io_out_2(c53_396_io_out_2)
  );
  C53 c53_397 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_397_io_in_0),
    .io_in_1(c53_397_io_in_1),
    .io_in_2(c53_397_io_in_2),
    .io_in_3(c53_397_io_in_3),
    .io_in_4(c53_397_io_in_4),
    .io_out_0(c53_397_io_out_0),
    .io_out_1(c53_397_io_out_1),
    .io_out_2(c53_397_io_out_2)
  );
  C32 c32_38 ( // @[Multiplier.scala 78:25]
    .io_in_0(c32_38_io_in_0),
    .io_in_1(c32_38_io_in_1),
    .io_in_2(c32_38_io_in_2),
    .io_out_0(c32_38_io_out_0),
    .io_out_1(c32_38_io_out_1)
  );
  C53 c53_398 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_398_io_in_0),
    .io_in_1(c53_398_io_in_1),
    .io_in_2(c53_398_io_in_2),
    .io_in_3(c53_398_io_in_3),
    .io_in_4(c53_398_io_in_4),
    .io_out_0(c53_398_io_out_0),
    .io_out_1(c53_398_io_out_1),
    .io_out_2(c53_398_io_out_2)
  );
  C53 c53_399 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_399_io_in_0),
    .io_in_1(c53_399_io_in_1),
    .io_in_2(c53_399_io_in_2),
    .io_in_3(c53_399_io_in_3),
    .io_in_4(c53_399_io_in_4),
    .io_out_0(c53_399_io_out_0),
    .io_out_1(c53_399_io_out_1),
    .io_out_2(c53_399_io_out_2)
  );
  C32 c32_39 ( // @[Multiplier.scala 78:25]
    .io_in_0(c32_39_io_in_0),
    .io_in_1(c32_39_io_in_1),
    .io_in_2(c32_39_io_in_2),
    .io_out_0(c32_39_io_out_0),
    .io_out_1(c32_39_io_out_1)
  );
  C53 c53_400 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_400_io_in_0),
    .io_in_1(c53_400_io_in_1),
    .io_in_2(c53_400_io_in_2),
    .io_in_3(c53_400_io_in_3),
    .io_in_4(c53_400_io_in_4),
    .io_out_0(c53_400_io_out_0),
    .io_out_1(c53_400_io_out_1),
    .io_out_2(c53_400_io_out_2)
  );
  C53 c53_401 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_401_io_in_0),
    .io_in_1(c53_401_io_in_1),
    .io_in_2(c53_401_io_in_2),
    .io_in_3(c53_401_io_in_3),
    .io_in_4(c53_401_io_in_4),
    .io_out_0(c53_401_io_out_0),
    .io_out_1(c53_401_io_out_1),
    .io_out_2(c53_401_io_out_2)
  );
  C32 c32_40 ( // @[Multiplier.scala 78:25]
    .io_in_0(c32_40_io_in_0),
    .io_in_1(c32_40_io_in_1),
    .io_in_2(c32_40_io_in_2),
    .io_out_0(c32_40_io_out_0),
    .io_out_1(c32_40_io_out_1)
  );
  C53 c53_402 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_402_io_in_0),
    .io_in_1(c53_402_io_in_1),
    .io_in_2(c53_402_io_in_2),
    .io_in_3(c53_402_io_in_3),
    .io_in_4(c53_402_io_in_4),
    .io_out_0(c53_402_io_out_0),
    .io_out_1(c53_402_io_out_1),
    .io_out_2(c53_402_io_out_2)
  );
  C53 c53_403 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_403_io_in_0),
    .io_in_1(c53_403_io_in_1),
    .io_in_2(c53_403_io_in_2),
    .io_in_3(c53_403_io_in_3),
    .io_in_4(c53_403_io_in_4),
    .io_out_0(c53_403_io_out_0),
    .io_out_1(c53_403_io_out_1),
    .io_out_2(c53_403_io_out_2)
  );
  C53 c53_404 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_404_io_in_0),
    .io_in_1(c53_404_io_in_1),
    .io_in_2(c53_404_io_in_2),
    .io_in_3(c53_404_io_in_3),
    .io_in_4(c53_404_io_in_4),
    .io_out_0(c53_404_io_out_0),
    .io_out_1(c53_404_io_out_1),
    .io_out_2(c53_404_io_out_2)
  );
  C53 c53_405 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_405_io_in_0),
    .io_in_1(c53_405_io_in_1),
    .io_in_2(c53_405_io_in_2),
    .io_in_3(c53_405_io_in_3),
    .io_in_4(c53_405_io_in_4),
    .io_out_0(c53_405_io_out_0),
    .io_out_1(c53_405_io_out_1),
    .io_out_2(c53_405_io_out_2)
  );
  C53 c53_406 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_406_io_in_0),
    .io_in_1(c53_406_io_in_1),
    .io_in_2(c53_406_io_in_2),
    .io_in_3(c53_406_io_in_3),
    .io_in_4(c53_406_io_in_4),
    .io_out_0(c53_406_io_out_0),
    .io_out_1(c53_406_io_out_1),
    .io_out_2(c53_406_io_out_2)
  );
  C53 c53_407 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_407_io_in_0),
    .io_in_1(c53_407_io_in_1),
    .io_in_2(c53_407_io_in_2),
    .io_in_3(c53_407_io_in_3),
    .io_in_4(c53_407_io_in_4),
    .io_out_0(c53_407_io_out_0),
    .io_out_1(c53_407_io_out_1),
    .io_out_2(c53_407_io_out_2)
  );
  C53 c53_408 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_408_io_in_0),
    .io_in_1(c53_408_io_in_1),
    .io_in_2(c53_408_io_in_2),
    .io_in_3(c53_408_io_in_3),
    .io_in_4(c53_408_io_in_4),
    .io_out_0(c53_408_io_out_0),
    .io_out_1(c53_408_io_out_1),
    .io_out_2(c53_408_io_out_2)
  );
  C53 c53_409 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_409_io_in_0),
    .io_in_1(c53_409_io_in_1),
    .io_in_2(c53_409_io_in_2),
    .io_in_3(c53_409_io_in_3),
    .io_in_4(c53_409_io_in_4),
    .io_out_0(c53_409_io_out_0),
    .io_out_1(c53_409_io_out_1),
    .io_out_2(c53_409_io_out_2)
  );
  C53 c53_410 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_410_io_in_0),
    .io_in_1(c53_410_io_in_1),
    .io_in_2(c53_410_io_in_2),
    .io_in_3(c53_410_io_in_3),
    .io_in_4(c53_410_io_in_4),
    .io_out_0(c53_410_io_out_0),
    .io_out_1(c53_410_io_out_1),
    .io_out_2(c53_410_io_out_2)
  );
  C53 c53_411 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_411_io_in_0),
    .io_in_1(c53_411_io_in_1),
    .io_in_2(c53_411_io_in_2),
    .io_in_3(c53_411_io_in_3),
    .io_in_4(c53_411_io_in_4),
    .io_out_0(c53_411_io_out_0),
    .io_out_1(c53_411_io_out_1),
    .io_out_2(c53_411_io_out_2)
  );
  C53 c53_412 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_412_io_in_0),
    .io_in_1(c53_412_io_in_1),
    .io_in_2(c53_412_io_in_2),
    .io_in_3(c53_412_io_in_3),
    .io_in_4(c53_412_io_in_4),
    .io_out_0(c53_412_io_out_0),
    .io_out_1(c53_412_io_out_1),
    .io_out_2(c53_412_io_out_2)
  );
  C53 c53_413 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_413_io_in_0),
    .io_in_1(c53_413_io_in_1),
    .io_in_2(c53_413_io_in_2),
    .io_in_3(c53_413_io_in_3),
    .io_in_4(c53_413_io_in_4),
    .io_out_0(c53_413_io_out_0),
    .io_out_1(c53_413_io_out_1),
    .io_out_2(c53_413_io_out_2)
  );
  C53 c53_414 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_414_io_in_0),
    .io_in_1(c53_414_io_in_1),
    .io_in_2(c53_414_io_in_2),
    .io_in_3(c53_414_io_in_3),
    .io_in_4(c53_414_io_in_4),
    .io_out_0(c53_414_io_out_0),
    .io_out_1(c53_414_io_out_1),
    .io_out_2(c53_414_io_out_2)
  );
  C53 c53_415 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_415_io_in_0),
    .io_in_1(c53_415_io_in_1),
    .io_in_2(c53_415_io_in_2),
    .io_in_3(c53_415_io_in_3),
    .io_in_4(c53_415_io_in_4),
    .io_out_0(c53_415_io_out_0),
    .io_out_1(c53_415_io_out_1),
    .io_out_2(c53_415_io_out_2)
  );
  C53 c53_416 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_416_io_in_0),
    .io_in_1(c53_416_io_in_1),
    .io_in_2(c53_416_io_in_2),
    .io_in_3(c53_416_io_in_3),
    .io_in_4(c53_416_io_in_4),
    .io_out_0(c53_416_io_out_0),
    .io_out_1(c53_416_io_out_1),
    .io_out_2(c53_416_io_out_2)
  );
  C53 c53_417 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_417_io_in_0),
    .io_in_1(c53_417_io_in_1),
    .io_in_2(c53_417_io_in_2),
    .io_in_3(c53_417_io_in_3),
    .io_in_4(c53_417_io_in_4),
    .io_out_0(c53_417_io_out_0),
    .io_out_1(c53_417_io_out_1),
    .io_out_2(c53_417_io_out_2)
  );
  C53 c53_418 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_418_io_in_0),
    .io_in_1(c53_418_io_in_1),
    .io_in_2(c53_418_io_in_2),
    .io_in_3(c53_418_io_in_3),
    .io_in_4(c53_418_io_in_4),
    .io_out_0(c53_418_io_out_0),
    .io_out_1(c53_418_io_out_1),
    .io_out_2(c53_418_io_out_2)
  );
  C53 c53_419 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_419_io_in_0),
    .io_in_1(c53_419_io_in_1),
    .io_in_2(c53_419_io_in_2),
    .io_in_3(c53_419_io_in_3),
    .io_in_4(c53_419_io_in_4),
    .io_out_0(c53_419_io_out_0),
    .io_out_1(c53_419_io_out_1),
    .io_out_2(c53_419_io_out_2)
  );
  C53 c53_420 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_420_io_in_0),
    .io_in_1(c53_420_io_in_1),
    .io_in_2(c53_420_io_in_2),
    .io_in_3(c53_420_io_in_3),
    .io_in_4(c53_420_io_in_4),
    .io_out_0(c53_420_io_out_0),
    .io_out_1(c53_420_io_out_1),
    .io_out_2(c53_420_io_out_2)
  );
  C53 c53_421 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_421_io_in_0),
    .io_in_1(c53_421_io_in_1),
    .io_in_2(c53_421_io_in_2),
    .io_in_3(c53_421_io_in_3),
    .io_in_4(c53_421_io_in_4),
    .io_out_0(c53_421_io_out_0),
    .io_out_1(c53_421_io_out_1),
    .io_out_2(c53_421_io_out_2)
  );
  C53 c53_422 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_422_io_in_0),
    .io_in_1(c53_422_io_in_1),
    .io_in_2(c53_422_io_in_2),
    .io_in_3(c53_422_io_in_3),
    .io_in_4(c53_422_io_in_4),
    .io_out_0(c53_422_io_out_0),
    .io_out_1(c53_422_io_out_1),
    .io_out_2(c53_422_io_out_2)
  );
  C53 c53_423 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_423_io_in_0),
    .io_in_1(c53_423_io_in_1),
    .io_in_2(c53_423_io_in_2),
    .io_in_3(c53_423_io_in_3),
    .io_in_4(c53_423_io_in_4),
    .io_out_0(c53_423_io_out_0),
    .io_out_1(c53_423_io_out_1),
    .io_out_2(c53_423_io_out_2)
  );
  C53 c53_424 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_424_io_in_0),
    .io_in_1(c53_424_io_in_1),
    .io_in_2(c53_424_io_in_2),
    .io_in_3(c53_424_io_in_3),
    .io_in_4(c53_424_io_in_4),
    .io_out_0(c53_424_io_out_0),
    .io_out_1(c53_424_io_out_1),
    .io_out_2(c53_424_io_out_2)
  );
  C53 c53_425 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_425_io_in_0),
    .io_in_1(c53_425_io_in_1),
    .io_in_2(c53_425_io_in_2),
    .io_in_3(c53_425_io_in_3),
    .io_in_4(c53_425_io_in_4),
    .io_out_0(c53_425_io_out_0),
    .io_out_1(c53_425_io_out_1),
    .io_out_2(c53_425_io_out_2)
  );
  C53 c53_426 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_426_io_in_0),
    .io_in_1(c53_426_io_in_1),
    .io_in_2(c53_426_io_in_2),
    .io_in_3(c53_426_io_in_3),
    .io_in_4(c53_426_io_in_4),
    .io_out_0(c53_426_io_out_0),
    .io_out_1(c53_426_io_out_1),
    .io_out_2(c53_426_io_out_2)
  );
  C53 c53_427 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_427_io_in_0),
    .io_in_1(c53_427_io_in_1),
    .io_in_2(c53_427_io_in_2),
    .io_in_3(c53_427_io_in_3),
    .io_in_4(c53_427_io_in_4),
    .io_out_0(c53_427_io_out_0),
    .io_out_1(c53_427_io_out_1),
    .io_out_2(c53_427_io_out_2)
  );
  C53 c53_428 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_428_io_in_0),
    .io_in_1(c53_428_io_in_1),
    .io_in_2(c53_428_io_in_2),
    .io_in_3(c53_428_io_in_3),
    .io_in_4(c53_428_io_in_4),
    .io_out_0(c53_428_io_out_0),
    .io_out_1(c53_428_io_out_1),
    .io_out_2(c53_428_io_out_2)
  );
  C22 c22_42 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_42_io_in_0),
    .io_in_1(c22_42_io_in_1),
    .io_out_0(c22_42_io_out_0),
    .io_out_1(c22_42_io_out_1)
  );
  C53 c53_429 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_429_io_in_0),
    .io_in_1(c53_429_io_in_1),
    .io_in_2(c53_429_io_in_2),
    .io_in_3(c53_429_io_in_3),
    .io_in_4(c53_429_io_in_4),
    .io_out_0(c53_429_io_out_0),
    .io_out_1(c53_429_io_out_1),
    .io_out_2(c53_429_io_out_2)
  );
  C53 c53_430 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_430_io_in_0),
    .io_in_1(c53_430_io_in_1),
    .io_in_2(c53_430_io_in_2),
    .io_in_3(c53_430_io_in_3),
    .io_in_4(c53_430_io_in_4),
    .io_out_0(c53_430_io_out_0),
    .io_out_1(c53_430_io_out_1),
    .io_out_2(c53_430_io_out_2)
  );
  C53 c53_431 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_431_io_in_0),
    .io_in_1(c53_431_io_in_1),
    .io_in_2(c53_431_io_in_2),
    .io_in_3(c53_431_io_in_3),
    .io_in_4(c53_431_io_in_4),
    .io_out_0(c53_431_io_out_0),
    .io_out_1(c53_431_io_out_1),
    .io_out_2(c53_431_io_out_2)
  );
  C22 c22_43 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_43_io_in_0),
    .io_in_1(c22_43_io_in_1),
    .io_out_0(c22_43_io_out_0),
    .io_out_1(c22_43_io_out_1)
  );
  C53 c53_432 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_432_io_in_0),
    .io_in_1(c53_432_io_in_1),
    .io_in_2(c53_432_io_in_2),
    .io_in_3(c53_432_io_in_3),
    .io_in_4(c53_432_io_in_4),
    .io_out_0(c53_432_io_out_0),
    .io_out_1(c53_432_io_out_1),
    .io_out_2(c53_432_io_out_2)
  );
  C53 c53_433 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_433_io_in_0),
    .io_in_1(c53_433_io_in_1),
    .io_in_2(c53_433_io_in_2),
    .io_in_3(c53_433_io_in_3),
    .io_in_4(c53_433_io_in_4),
    .io_out_0(c53_433_io_out_0),
    .io_out_1(c53_433_io_out_1),
    .io_out_2(c53_433_io_out_2)
  );
  C53 c53_434 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_434_io_in_0),
    .io_in_1(c53_434_io_in_1),
    .io_in_2(c53_434_io_in_2),
    .io_in_3(c53_434_io_in_3),
    .io_in_4(c53_434_io_in_4),
    .io_out_0(c53_434_io_out_0),
    .io_out_1(c53_434_io_out_1),
    .io_out_2(c53_434_io_out_2)
  );
  C22 c22_44 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_44_io_in_0),
    .io_in_1(c22_44_io_in_1),
    .io_out_0(c22_44_io_out_0),
    .io_out_1(c22_44_io_out_1)
  );
  C53 c53_435 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_435_io_in_0),
    .io_in_1(c53_435_io_in_1),
    .io_in_2(c53_435_io_in_2),
    .io_in_3(c53_435_io_in_3),
    .io_in_4(c53_435_io_in_4),
    .io_out_0(c53_435_io_out_0),
    .io_out_1(c53_435_io_out_1),
    .io_out_2(c53_435_io_out_2)
  );
  C53 c53_436 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_436_io_in_0),
    .io_in_1(c53_436_io_in_1),
    .io_in_2(c53_436_io_in_2),
    .io_in_3(c53_436_io_in_3),
    .io_in_4(c53_436_io_in_4),
    .io_out_0(c53_436_io_out_0),
    .io_out_1(c53_436_io_out_1),
    .io_out_2(c53_436_io_out_2)
  );
  C53 c53_437 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_437_io_in_0),
    .io_in_1(c53_437_io_in_1),
    .io_in_2(c53_437_io_in_2),
    .io_in_3(c53_437_io_in_3),
    .io_in_4(c53_437_io_in_4),
    .io_out_0(c53_437_io_out_0),
    .io_out_1(c53_437_io_out_1),
    .io_out_2(c53_437_io_out_2)
  );
  C22 c22_45 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_45_io_in_0),
    .io_in_1(c22_45_io_in_1),
    .io_out_0(c22_45_io_out_0),
    .io_out_1(c22_45_io_out_1)
  );
  C53 c53_438 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_438_io_in_0),
    .io_in_1(c53_438_io_in_1),
    .io_in_2(c53_438_io_in_2),
    .io_in_3(c53_438_io_in_3),
    .io_in_4(c53_438_io_in_4),
    .io_out_0(c53_438_io_out_0),
    .io_out_1(c53_438_io_out_1),
    .io_out_2(c53_438_io_out_2)
  );
  C53 c53_439 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_439_io_in_0),
    .io_in_1(c53_439_io_in_1),
    .io_in_2(c53_439_io_in_2),
    .io_in_3(c53_439_io_in_3),
    .io_in_4(c53_439_io_in_4),
    .io_out_0(c53_439_io_out_0),
    .io_out_1(c53_439_io_out_1),
    .io_out_2(c53_439_io_out_2)
  );
  C53 c53_440 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_440_io_in_0),
    .io_in_1(c53_440_io_in_1),
    .io_in_2(c53_440_io_in_2),
    .io_in_3(c53_440_io_in_3),
    .io_in_4(c53_440_io_in_4),
    .io_out_0(c53_440_io_out_0),
    .io_out_1(c53_440_io_out_1),
    .io_out_2(c53_440_io_out_2)
  );
  C22 c22_46 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_46_io_in_0),
    .io_in_1(c22_46_io_in_1),
    .io_out_0(c22_46_io_out_0),
    .io_out_1(c22_46_io_out_1)
  );
  C53 c53_441 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_441_io_in_0),
    .io_in_1(c53_441_io_in_1),
    .io_in_2(c53_441_io_in_2),
    .io_in_3(c53_441_io_in_3),
    .io_in_4(c53_441_io_in_4),
    .io_out_0(c53_441_io_out_0),
    .io_out_1(c53_441_io_out_1),
    .io_out_2(c53_441_io_out_2)
  );
  C53 c53_442 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_442_io_in_0),
    .io_in_1(c53_442_io_in_1),
    .io_in_2(c53_442_io_in_2),
    .io_in_3(c53_442_io_in_3),
    .io_in_4(c53_442_io_in_4),
    .io_out_0(c53_442_io_out_0),
    .io_out_1(c53_442_io_out_1),
    .io_out_2(c53_442_io_out_2)
  );
  C53 c53_443 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_443_io_in_0),
    .io_in_1(c53_443_io_in_1),
    .io_in_2(c53_443_io_in_2),
    .io_in_3(c53_443_io_in_3),
    .io_in_4(c53_443_io_in_4),
    .io_out_0(c53_443_io_out_0),
    .io_out_1(c53_443_io_out_1),
    .io_out_2(c53_443_io_out_2)
  );
  C22 c22_47 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_47_io_in_0),
    .io_in_1(c22_47_io_in_1),
    .io_out_0(c22_47_io_out_0),
    .io_out_1(c22_47_io_out_1)
  );
  C53 c53_444 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_444_io_in_0),
    .io_in_1(c53_444_io_in_1),
    .io_in_2(c53_444_io_in_2),
    .io_in_3(c53_444_io_in_3),
    .io_in_4(c53_444_io_in_4),
    .io_out_0(c53_444_io_out_0),
    .io_out_1(c53_444_io_out_1),
    .io_out_2(c53_444_io_out_2)
  );
  C53 c53_445 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_445_io_in_0),
    .io_in_1(c53_445_io_in_1),
    .io_in_2(c53_445_io_in_2),
    .io_in_3(c53_445_io_in_3),
    .io_in_4(c53_445_io_in_4),
    .io_out_0(c53_445_io_out_0),
    .io_out_1(c53_445_io_out_1),
    .io_out_2(c53_445_io_out_2)
  );
  C53 c53_446 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_446_io_in_0),
    .io_in_1(c53_446_io_in_1),
    .io_in_2(c53_446_io_in_2),
    .io_in_3(c53_446_io_in_3),
    .io_in_4(c53_446_io_in_4),
    .io_out_0(c53_446_io_out_0),
    .io_out_1(c53_446_io_out_1),
    .io_out_2(c53_446_io_out_2)
  );
  C22 c22_48 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_48_io_in_0),
    .io_in_1(c22_48_io_in_1),
    .io_out_0(c22_48_io_out_0),
    .io_out_1(c22_48_io_out_1)
  );
  C53 c53_447 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_447_io_in_0),
    .io_in_1(c53_447_io_in_1),
    .io_in_2(c53_447_io_in_2),
    .io_in_3(c53_447_io_in_3),
    .io_in_4(c53_447_io_in_4),
    .io_out_0(c53_447_io_out_0),
    .io_out_1(c53_447_io_out_1),
    .io_out_2(c53_447_io_out_2)
  );
  C53 c53_448 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_448_io_in_0),
    .io_in_1(c53_448_io_in_1),
    .io_in_2(c53_448_io_in_2),
    .io_in_3(c53_448_io_in_3),
    .io_in_4(c53_448_io_in_4),
    .io_out_0(c53_448_io_out_0),
    .io_out_1(c53_448_io_out_1),
    .io_out_2(c53_448_io_out_2)
  );
  C53 c53_449 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_449_io_in_0),
    .io_in_1(c53_449_io_in_1),
    .io_in_2(c53_449_io_in_2),
    .io_in_3(c53_449_io_in_3),
    .io_in_4(c53_449_io_in_4),
    .io_out_0(c53_449_io_out_0),
    .io_out_1(c53_449_io_out_1),
    .io_out_2(c53_449_io_out_2)
  );
  C22 c22_49 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_49_io_in_0),
    .io_in_1(c22_49_io_in_1),
    .io_out_0(c22_49_io_out_0),
    .io_out_1(c22_49_io_out_1)
  );
  C53 c53_450 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_450_io_in_0),
    .io_in_1(c53_450_io_in_1),
    .io_in_2(c53_450_io_in_2),
    .io_in_3(c53_450_io_in_3),
    .io_in_4(c53_450_io_in_4),
    .io_out_0(c53_450_io_out_0),
    .io_out_1(c53_450_io_out_1),
    .io_out_2(c53_450_io_out_2)
  );
  C53 c53_451 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_451_io_in_0),
    .io_in_1(c53_451_io_in_1),
    .io_in_2(c53_451_io_in_2),
    .io_in_3(c53_451_io_in_3),
    .io_in_4(c53_451_io_in_4),
    .io_out_0(c53_451_io_out_0),
    .io_out_1(c53_451_io_out_1),
    .io_out_2(c53_451_io_out_2)
  );
  C53 c53_452 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_452_io_in_0),
    .io_in_1(c53_452_io_in_1),
    .io_in_2(c53_452_io_in_2),
    .io_in_3(c53_452_io_in_3),
    .io_in_4(c53_452_io_in_4),
    .io_out_0(c53_452_io_out_0),
    .io_out_1(c53_452_io_out_1),
    .io_out_2(c53_452_io_out_2)
  );
  C22 c22_50 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_50_io_in_0),
    .io_in_1(c22_50_io_in_1),
    .io_out_0(c22_50_io_out_0),
    .io_out_1(c22_50_io_out_1)
  );
  C53 c53_453 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_453_io_in_0),
    .io_in_1(c53_453_io_in_1),
    .io_in_2(c53_453_io_in_2),
    .io_in_3(c53_453_io_in_3),
    .io_in_4(c53_453_io_in_4),
    .io_out_0(c53_453_io_out_0),
    .io_out_1(c53_453_io_out_1),
    .io_out_2(c53_453_io_out_2)
  );
  C53 c53_454 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_454_io_in_0),
    .io_in_1(c53_454_io_in_1),
    .io_in_2(c53_454_io_in_2),
    .io_in_3(c53_454_io_in_3),
    .io_in_4(c53_454_io_in_4),
    .io_out_0(c53_454_io_out_0),
    .io_out_1(c53_454_io_out_1),
    .io_out_2(c53_454_io_out_2)
  );
  C53 c53_455 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_455_io_in_0),
    .io_in_1(c53_455_io_in_1),
    .io_in_2(c53_455_io_in_2),
    .io_in_3(c53_455_io_in_3),
    .io_in_4(c53_455_io_in_4),
    .io_out_0(c53_455_io_out_0),
    .io_out_1(c53_455_io_out_1),
    .io_out_2(c53_455_io_out_2)
  );
  C22 c22_51 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_51_io_in_0),
    .io_in_1(c22_51_io_in_1),
    .io_out_0(c22_51_io_out_0),
    .io_out_1(c22_51_io_out_1)
  );
  C53 c53_456 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_456_io_in_0),
    .io_in_1(c53_456_io_in_1),
    .io_in_2(c53_456_io_in_2),
    .io_in_3(c53_456_io_in_3),
    .io_in_4(c53_456_io_in_4),
    .io_out_0(c53_456_io_out_0),
    .io_out_1(c53_456_io_out_1),
    .io_out_2(c53_456_io_out_2)
  );
  C53 c53_457 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_457_io_in_0),
    .io_in_1(c53_457_io_in_1),
    .io_in_2(c53_457_io_in_2),
    .io_in_3(c53_457_io_in_3),
    .io_in_4(c53_457_io_in_4),
    .io_out_0(c53_457_io_out_0),
    .io_out_1(c53_457_io_out_1),
    .io_out_2(c53_457_io_out_2)
  );
  C53 c53_458 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_458_io_in_0),
    .io_in_1(c53_458_io_in_1),
    .io_in_2(c53_458_io_in_2),
    .io_in_3(c53_458_io_in_3),
    .io_in_4(c53_458_io_in_4),
    .io_out_0(c53_458_io_out_0),
    .io_out_1(c53_458_io_out_1),
    .io_out_2(c53_458_io_out_2)
  );
  C22 c22_52 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_52_io_in_0),
    .io_in_1(c22_52_io_in_1),
    .io_out_0(c22_52_io_out_0),
    .io_out_1(c22_52_io_out_1)
  );
  C53 c53_459 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_459_io_in_0),
    .io_in_1(c53_459_io_in_1),
    .io_in_2(c53_459_io_in_2),
    .io_in_3(c53_459_io_in_3),
    .io_in_4(c53_459_io_in_4),
    .io_out_0(c53_459_io_out_0),
    .io_out_1(c53_459_io_out_1),
    .io_out_2(c53_459_io_out_2)
  );
  C53 c53_460 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_460_io_in_0),
    .io_in_1(c53_460_io_in_1),
    .io_in_2(c53_460_io_in_2),
    .io_in_3(c53_460_io_in_3),
    .io_in_4(c53_460_io_in_4),
    .io_out_0(c53_460_io_out_0),
    .io_out_1(c53_460_io_out_1),
    .io_out_2(c53_460_io_out_2)
  );
  C53 c53_461 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_461_io_in_0),
    .io_in_1(c53_461_io_in_1),
    .io_in_2(c53_461_io_in_2),
    .io_in_3(c53_461_io_in_3),
    .io_in_4(c53_461_io_in_4),
    .io_out_0(c53_461_io_out_0),
    .io_out_1(c53_461_io_out_1),
    .io_out_2(c53_461_io_out_2)
  );
  C53 c53_462 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_462_io_in_0),
    .io_in_1(c53_462_io_in_1),
    .io_in_2(c53_462_io_in_2),
    .io_in_3(c53_462_io_in_3),
    .io_in_4(c53_462_io_in_4),
    .io_out_0(c53_462_io_out_0),
    .io_out_1(c53_462_io_out_1),
    .io_out_2(c53_462_io_out_2)
  );
  C53 c53_463 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_463_io_in_0),
    .io_in_1(c53_463_io_in_1),
    .io_in_2(c53_463_io_in_2),
    .io_in_3(c53_463_io_in_3),
    .io_in_4(c53_463_io_in_4),
    .io_out_0(c53_463_io_out_0),
    .io_out_1(c53_463_io_out_1),
    .io_out_2(c53_463_io_out_2)
  );
  C53 c53_464 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_464_io_in_0),
    .io_in_1(c53_464_io_in_1),
    .io_in_2(c53_464_io_in_2),
    .io_in_3(c53_464_io_in_3),
    .io_in_4(c53_464_io_in_4),
    .io_out_0(c53_464_io_out_0),
    .io_out_1(c53_464_io_out_1),
    .io_out_2(c53_464_io_out_2)
  );
  C53 c53_465 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_465_io_in_0),
    .io_in_1(c53_465_io_in_1),
    .io_in_2(c53_465_io_in_2),
    .io_in_3(c53_465_io_in_3),
    .io_in_4(c53_465_io_in_4),
    .io_out_0(c53_465_io_out_0),
    .io_out_1(c53_465_io_out_1),
    .io_out_2(c53_465_io_out_2)
  );
  C53 c53_466 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_466_io_in_0),
    .io_in_1(c53_466_io_in_1),
    .io_in_2(c53_466_io_in_2),
    .io_in_3(c53_466_io_in_3),
    .io_in_4(c53_466_io_in_4),
    .io_out_0(c53_466_io_out_0),
    .io_out_1(c53_466_io_out_1),
    .io_out_2(c53_466_io_out_2)
  );
  C53 c53_467 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_467_io_in_0),
    .io_in_1(c53_467_io_in_1),
    .io_in_2(c53_467_io_in_2),
    .io_in_3(c53_467_io_in_3),
    .io_in_4(c53_467_io_in_4),
    .io_out_0(c53_467_io_out_0),
    .io_out_1(c53_467_io_out_1),
    .io_out_2(c53_467_io_out_2)
  );
  C53 c53_468 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_468_io_in_0),
    .io_in_1(c53_468_io_in_1),
    .io_in_2(c53_468_io_in_2),
    .io_in_3(c53_468_io_in_3),
    .io_in_4(c53_468_io_in_4),
    .io_out_0(c53_468_io_out_0),
    .io_out_1(c53_468_io_out_1),
    .io_out_2(c53_468_io_out_2)
  );
  C53 c53_469 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_469_io_in_0),
    .io_in_1(c53_469_io_in_1),
    .io_in_2(c53_469_io_in_2),
    .io_in_3(c53_469_io_in_3),
    .io_in_4(c53_469_io_in_4),
    .io_out_0(c53_469_io_out_0),
    .io_out_1(c53_469_io_out_1),
    .io_out_2(c53_469_io_out_2)
  );
  C53 c53_470 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_470_io_in_0),
    .io_in_1(c53_470_io_in_1),
    .io_in_2(c53_470_io_in_2),
    .io_in_3(c53_470_io_in_3),
    .io_in_4(c53_470_io_in_4),
    .io_out_0(c53_470_io_out_0),
    .io_out_1(c53_470_io_out_1),
    .io_out_2(c53_470_io_out_2)
  );
  C53 c53_471 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_471_io_in_0),
    .io_in_1(c53_471_io_in_1),
    .io_in_2(c53_471_io_in_2),
    .io_in_3(c53_471_io_in_3),
    .io_in_4(c53_471_io_in_4),
    .io_out_0(c53_471_io_out_0),
    .io_out_1(c53_471_io_out_1),
    .io_out_2(c53_471_io_out_2)
  );
  C53 c53_472 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_472_io_in_0),
    .io_in_1(c53_472_io_in_1),
    .io_in_2(c53_472_io_in_2),
    .io_in_3(c53_472_io_in_3),
    .io_in_4(c53_472_io_in_4),
    .io_out_0(c53_472_io_out_0),
    .io_out_1(c53_472_io_out_1),
    .io_out_2(c53_472_io_out_2)
  );
  C53 c53_473 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_473_io_in_0),
    .io_in_1(c53_473_io_in_1),
    .io_in_2(c53_473_io_in_2),
    .io_in_3(c53_473_io_in_3),
    .io_in_4(c53_473_io_in_4),
    .io_out_0(c53_473_io_out_0),
    .io_out_1(c53_473_io_out_1),
    .io_out_2(c53_473_io_out_2)
  );
  C53 c53_474 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_474_io_in_0),
    .io_in_1(c53_474_io_in_1),
    .io_in_2(c53_474_io_in_2),
    .io_in_3(c53_474_io_in_3),
    .io_in_4(c53_474_io_in_4),
    .io_out_0(c53_474_io_out_0),
    .io_out_1(c53_474_io_out_1),
    .io_out_2(c53_474_io_out_2)
  );
  C53 c53_475 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_475_io_in_0),
    .io_in_1(c53_475_io_in_1),
    .io_in_2(c53_475_io_in_2),
    .io_in_3(c53_475_io_in_3),
    .io_in_4(c53_475_io_in_4),
    .io_out_0(c53_475_io_out_0),
    .io_out_1(c53_475_io_out_1),
    .io_out_2(c53_475_io_out_2)
  );
  C53 c53_476 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_476_io_in_0),
    .io_in_1(c53_476_io_in_1),
    .io_in_2(c53_476_io_in_2),
    .io_in_3(c53_476_io_in_3),
    .io_in_4(c53_476_io_in_4),
    .io_out_0(c53_476_io_out_0),
    .io_out_1(c53_476_io_out_1),
    .io_out_2(c53_476_io_out_2)
  );
  C53 c53_477 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_477_io_in_0),
    .io_in_1(c53_477_io_in_1),
    .io_in_2(c53_477_io_in_2),
    .io_in_3(c53_477_io_in_3),
    .io_in_4(c53_477_io_in_4),
    .io_out_0(c53_477_io_out_0),
    .io_out_1(c53_477_io_out_1),
    .io_out_2(c53_477_io_out_2)
  );
  C53 c53_478 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_478_io_in_0),
    .io_in_1(c53_478_io_in_1),
    .io_in_2(c53_478_io_in_2),
    .io_in_3(c53_478_io_in_3),
    .io_in_4(c53_478_io_in_4),
    .io_out_0(c53_478_io_out_0),
    .io_out_1(c53_478_io_out_1),
    .io_out_2(c53_478_io_out_2)
  );
  C53 c53_479 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_479_io_in_0),
    .io_in_1(c53_479_io_in_1),
    .io_in_2(c53_479_io_in_2),
    .io_in_3(c53_479_io_in_3),
    .io_in_4(c53_479_io_in_4),
    .io_out_0(c53_479_io_out_0),
    .io_out_1(c53_479_io_out_1),
    .io_out_2(c53_479_io_out_2)
  );
  C53 c53_480 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_480_io_in_0),
    .io_in_1(c53_480_io_in_1),
    .io_in_2(c53_480_io_in_2),
    .io_in_3(c53_480_io_in_3),
    .io_in_4(c53_480_io_in_4),
    .io_out_0(c53_480_io_out_0),
    .io_out_1(c53_480_io_out_1),
    .io_out_2(c53_480_io_out_2)
  );
  C53 c53_481 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_481_io_in_0),
    .io_in_1(c53_481_io_in_1),
    .io_in_2(c53_481_io_in_2),
    .io_in_3(c53_481_io_in_3),
    .io_in_4(c53_481_io_in_4),
    .io_out_0(c53_481_io_out_0),
    .io_out_1(c53_481_io_out_1),
    .io_out_2(c53_481_io_out_2)
  );
  C53 c53_482 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_482_io_in_0),
    .io_in_1(c53_482_io_in_1),
    .io_in_2(c53_482_io_in_2),
    .io_in_3(c53_482_io_in_3),
    .io_in_4(c53_482_io_in_4),
    .io_out_0(c53_482_io_out_0),
    .io_out_1(c53_482_io_out_1),
    .io_out_2(c53_482_io_out_2)
  );
  C53 c53_483 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_483_io_in_0),
    .io_in_1(c53_483_io_in_1),
    .io_in_2(c53_483_io_in_2),
    .io_in_3(c53_483_io_in_3),
    .io_in_4(c53_483_io_in_4),
    .io_out_0(c53_483_io_out_0),
    .io_out_1(c53_483_io_out_1),
    .io_out_2(c53_483_io_out_2)
  );
  C53 c53_484 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_484_io_in_0),
    .io_in_1(c53_484_io_in_1),
    .io_in_2(c53_484_io_in_2),
    .io_in_3(c53_484_io_in_3),
    .io_in_4(c53_484_io_in_4),
    .io_out_0(c53_484_io_out_0),
    .io_out_1(c53_484_io_out_1),
    .io_out_2(c53_484_io_out_2)
  );
  C32 c32_41 ( // @[Multiplier.scala 78:25]
    .io_in_0(c32_41_io_in_0),
    .io_in_1(c32_41_io_in_1),
    .io_in_2(c32_41_io_in_2),
    .io_out_0(c32_41_io_out_0),
    .io_out_1(c32_41_io_out_1)
  );
  C53 c53_485 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_485_io_in_0),
    .io_in_1(c53_485_io_in_1),
    .io_in_2(c53_485_io_in_2),
    .io_in_3(c53_485_io_in_3),
    .io_in_4(c53_485_io_in_4),
    .io_out_0(c53_485_io_out_0),
    .io_out_1(c53_485_io_out_1),
    .io_out_2(c53_485_io_out_2)
  );
  C53 c53_486 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_486_io_in_0),
    .io_in_1(c53_486_io_in_1),
    .io_in_2(c53_486_io_in_2),
    .io_in_3(c53_486_io_in_3),
    .io_in_4(c53_486_io_in_4),
    .io_out_0(c53_486_io_out_0),
    .io_out_1(c53_486_io_out_1),
    .io_out_2(c53_486_io_out_2)
  );
  C22 c22_53 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_53_io_in_0),
    .io_in_1(c22_53_io_in_1),
    .io_out_0(c22_53_io_out_0),
    .io_out_1(c22_53_io_out_1)
  );
  C53 c53_487 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_487_io_in_0),
    .io_in_1(c53_487_io_in_1),
    .io_in_2(c53_487_io_in_2),
    .io_in_3(c53_487_io_in_3),
    .io_in_4(c53_487_io_in_4),
    .io_out_0(c53_487_io_out_0),
    .io_out_1(c53_487_io_out_1),
    .io_out_2(c53_487_io_out_2)
  );
  C53 c53_488 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_488_io_in_0),
    .io_in_1(c53_488_io_in_1),
    .io_in_2(c53_488_io_in_2),
    .io_in_3(c53_488_io_in_3),
    .io_in_4(c53_488_io_in_4),
    .io_out_0(c53_488_io_out_0),
    .io_out_1(c53_488_io_out_1),
    .io_out_2(c53_488_io_out_2)
  );
  C22 c22_54 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_54_io_in_0),
    .io_in_1(c22_54_io_in_1),
    .io_out_0(c22_54_io_out_0),
    .io_out_1(c22_54_io_out_1)
  );
  C53 c53_489 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_489_io_in_0),
    .io_in_1(c53_489_io_in_1),
    .io_in_2(c53_489_io_in_2),
    .io_in_3(c53_489_io_in_3),
    .io_in_4(c53_489_io_in_4),
    .io_out_0(c53_489_io_out_0),
    .io_out_1(c53_489_io_out_1),
    .io_out_2(c53_489_io_out_2)
  );
  C53 c53_490 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_490_io_in_0),
    .io_in_1(c53_490_io_in_1),
    .io_in_2(c53_490_io_in_2),
    .io_in_3(c53_490_io_in_3),
    .io_in_4(c53_490_io_in_4),
    .io_out_0(c53_490_io_out_0),
    .io_out_1(c53_490_io_out_1),
    .io_out_2(c53_490_io_out_2)
  );
  C32 c32_42 ( // @[Multiplier.scala 78:25]
    .io_in_0(c32_42_io_in_0),
    .io_in_1(c32_42_io_in_1),
    .io_in_2(c32_42_io_in_2),
    .io_out_0(c32_42_io_out_0),
    .io_out_1(c32_42_io_out_1)
  );
  C53 c53_491 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_491_io_in_0),
    .io_in_1(c53_491_io_in_1),
    .io_in_2(c53_491_io_in_2),
    .io_in_3(c53_491_io_in_3),
    .io_in_4(c53_491_io_in_4),
    .io_out_0(c53_491_io_out_0),
    .io_out_1(c53_491_io_out_1),
    .io_out_2(c53_491_io_out_2)
  );
  C53 c53_492 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_492_io_in_0),
    .io_in_1(c53_492_io_in_1),
    .io_in_2(c53_492_io_in_2),
    .io_in_3(c53_492_io_in_3),
    .io_in_4(c53_492_io_in_4),
    .io_out_0(c53_492_io_out_0),
    .io_out_1(c53_492_io_out_1),
    .io_out_2(c53_492_io_out_2)
  );
  C22 c22_55 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_55_io_in_0),
    .io_in_1(c22_55_io_in_1),
    .io_out_0(c22_55_io_out_0),
    .io_out_1(c22_55_io_out_1)
  );
  C53 c53_493 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_493_io_in_0),
    .io_in_1(c53_493_io_in_1),
    .io_in_2(c53_493_io_in_2),
    .io_in_3(c53_493_io_in_3),
    .io_in_4(c53_493_io_in_4),
    .io_out_0(c53_493_io_out_0),
    .io_out_1(c53_493_io_out_1),
    .io_out_2(c53_493_io_out_2)
  );
  C53 c53_494 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_494_io_in_0),
    .io_in_1(c53_494_io_in_1),
    .io_in_2(c53_494_io_in_2),
    .io_in_3(c53_494_io_in_3),
    .io_in_4(c53_494_io_in_4),
    .io_out_0(c53_494_io_out_0),
    .io_out_1(c53_494_io_out_1),
    .io_out_2(c53_494_io_out_2)
  );
  C22 c22_56 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_56_io_in_0),
    .io_in_1(c22_56_io_in_1),
    .io_out_0(c22_56_io_out_0),
    .io_out_1(c22_56_io_out_1)
  );
  C53 c53_495 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_495_io_in_0),
    .io_in_1(c53_495_io_in_1),
    .io_in_2(c53_495_io_in_2),
    .io_in_3(c53_495_io_in_3),
    .io_in_4(c53_495_io_in_4),
    .io_out_0(c53_495_io_out_0),
    .io_out_1(c53_495_io_out_1),
    .io_out_2(c53_495_io_out_2)
  );
  C53 c53_496 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_496_io_in_0),
    .io_in_1(c53_496_io_in_1),
    .io_in_2(c53_496_io_in_2),
    .io_in_3(c53_496_io_in_3),
    .io_in_4(c53_496_io_in_4),
    .io_out_0(c53_496_io_out_0),
    .io_out_1(c53_496_io_out_1),
    .io_out_2(c53_496_io_out_2)
  );
  C22 c22_57 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_57_io_in_0),
    .io_in_1(c22_57_io_in_1),
    .io_out_0(c22_57_io_out_0),
    .io_out_1(c22_57_io_out_1)
  );
  C53 c53_497 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_497_io_in_0),
    .io_in_1(c53_497_io_in_1),
    .io_in_2(c53_497_io_in_2),
    .io_in_3(c53_497_io_in_3),
    .io_in_4(c53_497_io_in_4),
    .io_out_0(c53_497_io_out_0),
    .io_out_1(c53_497_io_out_1),
    .io_out_2(c53_497_io_out_2)
  );
  C53 c53_498 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_498_io_in_0),
    .io_in_1(c53_498_io_in_1),
    .io_in_2(c53_498_io_in_2),
    .io_in_3(c53_498_io_in_3),
    .io_in_4(c53_498_io_in_4),
    .io_out_0(c53_498_io_out_0),
    .io_out_1(c53_498_io_out_1),
    .io_out_2(c53_498_io_out_2)
  );
  C22 c22_58 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_58_io_in_0),
    .io_in_1(c22_58_io_in_1),
    .io_out_0(c22_58_io_out_0),
    .io_out_1(c22_58_io_out_1)
  );
  C53 c53_499 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_499_io_in_0),
    .io_in_1(c53_499_io_in_1),
    .io_in_2(c53_499_io_in_2),
    .io_in_3(c53_499_io_in_3),
    .io_in_4(c53_499_io_in_4),
    .io_out_0(c53_499_io_out_0),
    .io_out_1(c53_499_io_out_1),
    .io_out_2(c53_499_io_out_2)
  );
  C53 c53_500 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_500_io_in_0),
    .io_in_1(c53_500_io_in_1),
    .io_in_2(c53_500_io_in_2),
    .io_in_3(c53_500_io_in_3),
    .io_in_4(c53_500_io_in_4),
    .io_out_0(c53_500_io_out_0),
    .io_out_1(c53_500_io_out_1),
    .io_out_2(c53_500_io_out_2)
  );
  C53 c53_501 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_501_io_in_0),
    .io_in_1(c53_501_io_in_1),
    .io_in_2(c53_501_io_in_2),
    .io_in_3(c53_501_io_in_3),
    .io_in_4(c53_501_io_in_4),
    .io_out_0(c53_501_io_out_0),
    .io_out_1(c53_501_io_out_1),
    .io_out_2(c53_501_io_out_2)
  );
  C53 c53_502 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_502_io_in_0),
    .io_in_1(c53_502_io_in_1),
    .io_in_2(c53_502_io_in_2),
    .io_in_3(c53_502_io_in_3),
    .io_in_4(c53_502_io_in_4),
    .io_out_0(c53_502_io_out_0),
    .io_out_1(c53_502_io_out_1),
    .io_out_2(c53_502_io_out_2)
  );
  C53 c53_503 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_503_io_in_0),
    .io_in_1(c53_503_io_in_1),
    .io_in_2(c53_503_io_in_2),
    .io_in_3(c53_503_io_in_3),
    .io_in_4(c53_503_io_in_4),
    .io_out_0(c53_503_io_out_0),
    .io_out_1(c53_503_io_out_1),
    .io_out_2(c53_503_io_out_2)
  );
  C53 c53_504 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_504_io_in_0),
    .io_in_1(c53_504_io_in_1),
    .io_in_2(c53_504_io_in_2),
    .io_in_3(c53_504_io_in_3),
    .io_in_4(c53_504_io_in_4),
    .io_out_0(c53_504_io_out_0),
    .io_out_1(c53_504_io_out_1),
    .io_out_2(c53_504_io_out_2)
  );
  C53 c53_505 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_505_io_in_0),
    .io_in_1(c53_505_io_in_1),
    .io_in_2(c53_505_io_in_2),
    .io_in_3(c53_505_io_in_3),
    .io_in_4(c53_505_io_in_4),
    .io_out_0(c53_505_io_out_0),
    .io_out_1(c53_505_io_out_1),
    .io_out_2(c53_505_io_out_2)
  );
  C53 c53_506 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_506_io_in_0),
    .io_in_1(c53_506_io_in_1),
    .io_in_2(c53_506_io_in_2),
    .io_in_3(c53_506_io_in_3),
    .io_in_4(c53_506_io_in_4),
    .io_out_0(c53_506_io_out_0),
    .io_out_1(c53_506_io_out_1),
    .io_out_2(c53_506_io_out_2)
  );
  C53 c53_507 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_507_io_in_0),
    .io_in_1(c53_507_io_in_1),
    .io_in_2(c53_507_io_in_2),
    .io_in_3(c53_507_io_in_3),
    .io_in_4(c53_507_io_in_4),
    .io_out_0(c53_507_io_out_0),
    .io_out_1(c53_507_io_out_1),
    .io_out_2(c53_507_io_out_2)
  );
  C53 c53_508 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_508_io_in_0),
    .io_in_1(c53_508_io_in_1),
    .io_in_2(c53_508_io_in_2),
    .io_in_3(c53_508_io_in_3),
    .io_in_4(c53_508_io_in_4),
    .io_out_0(c53_508_io_out_0),
    .io_out_1(c53_508_io_out_1),
    .io_out_2(c53_508_io_out_2)
  );
  C53 c53_509 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_509_io_in_0),
    .io_in_1(c53_509_io_in_1),
    .io_in_2(c53_509_io_in_2),
    .io_in_3(c53_509_io_in_3),
    .io_in_4(c53_509_io_in_4),
    .io_out_0(c53_509_io_out_0),
    .io_out_1(c53_509_io_out_1),
    .io_out_2(c53_509_io_out_2)
  );
  C53 c53_510 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_510_io_in_0),
    .io_in_1(c53_510_io_in_1),
    .io_in_2(c53_510_io_in_2),
    .io_in_3(c53_510_io_in_3),
    .io_in_4(c53_510_io_in_4),
    .io_out_0(c53_510_io_out_0),
    .io_out_1(c53_510_io_out_1),
    .io_out_2(c53_510_io_out_2)
  );
  C53 c53_511 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_511_io_in_0),
    .io_in_1(c53_511_io_in_1),
    .io_in_2(c53_511_io_in_2),
    .io_in_3(c53_511_io_in_3),
    .io_in_4(c53_511_io_in_4),
    .io_out_0(c53_511_io_out_0),
    .io_out_1(c53_511_io_out_1),
    .io_out_2(c53_511_io_out_2)
  );
  C53 c53_512 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_512_io_in_0),
    .io_in_1(c53_512_io_in_1),
    .io_in_2(c53_512_io_in_2),
    .io_in_3(c53_512_io_in_3),
    .io_in_4(c53_512_io_in_4),
    .io_out_0(c53_512_io_out_0),
    .io_out_1(c53_512_io_out_1),
    .io_out_2(c53_512_io_out_2)
  );
  C53 c53_513 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_513_io_in_0),
    .io_in_1(c53_513_io_in_1),
    .io_in_2(c53_513_io_in_2),
    .io_in_3(c53_513_io_in_3),
    .io_in_4(c53_513_io_in_4),
    .io_out_0(c53_513_io_out_0),
    .io_out_1(c53_513_io_out_1),
    .io_out_2(c53_513_io_out_2)
  );
  C53 c53_514 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_514_io_in_0),
    .io_in_1(c53_514_io_in_1),
    .io_in_2(c53_514_io_in_2),
    .io_in_3(c53_514_io_in_3),
    .io_in_4(c53_514_io_in_4),
    .io_out_0(c53_514_io_out_0),
    .io_out_1(c53_514_io_out_1),
    .io_out_2(c53_514_io_out_2)
  );
  C53 c53_515 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_515_io_in_0),
    .io_in_1(c53_515_io_in_1),
    .io_in_2(c53_515_io_in_2),
    .io_in_3(c53_515_io_in_3),
    .io_in_4(c53_515_io_in_4),
    .io_out_0(c53_515_io_out_0),
    .io_out_1(c53_515_io_out_1),
    .io_out_2(c53_515_io_out_2)
  );
  C32 c32_43 ( // @[Multiplier.scala 78:25]
    .io_in_0(c32_43_io_in_0),
    .io_in_1(c32_43_io_in_1),
    .io_in_2(c32_43_io_in_2),
    .io_out_0(c32_43_io_out_0),
    .io_out_1(c32_43_io_out_1)
  );
  C53 c53_516 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_516_io_in_0),
    .io_in_1(c53_516_io_in_1),
    .io_in_2(c53_516_io_in_2),
    .io_in_3(c53_516_io_in_3),
    .io_in_4(c53_516_io_in_4),
    .io_out_0(c53_516_io_out_0),
    .io_out_1(c53_516_io_out_1),
    .io_out_2(c53_516_io_out_2)
  );
  C22 c22_59 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_59_io_in_0),
    .io_in_1(c22_59_io_in_1),
    .io_out_0(c22_59_io_out_0),
    .io_out_1(c22_59_io_out_1)
  );
  C53 c53_517 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_517_io_in_0),
    .io_in_1(c53_517_io_in_1),
    .io_in_2(c53_517_io_in_2),
    .io_in_3(c53_517_io_in_3),
    .io_in_4(c53_517_io_in_4),
    .io_out_0(c53_517_io_out_0),
    .io_out_1(c53_517_io_out_1),
    .io_out_2(c53_517_io_out_2)
  );
  C22 c22_60 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_60_io_in_0),
    .io_in_1(c22_60_io_in_1),
    .io_out_0(c22_60_io_out_0),
    .io_out_1(c22_60_io_out_1)
  );
  C53 c53_518 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_518_io_in_0),
    .io_in_1(c53_518_io_in_1),
    .io_in_2(c53_518_io_in_2),
    .io_in_3(c53_518_io_in_3),
    .io_in_4(c53_518_io_in_4),
    .io_out_0(c53_518_io_out_0),
    .io_out_1(c53_518_io_out_1),
    .io_out_2(c53_518_io_out_2)
  );
  C32 c32_44 ( // @[Multiplier.scala 78:25]
    .io_in_0(c32_44_io_in_0),
    .io_in_1(c32_44_io_in_1),
    .io_in_2(c32_44_io_in_2),
    .io_out_0(c32_44_io_out_0),
    .io_out_1(c32_44_io_out_1)
  );
  C53 c53_519 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_519_io_in_0),
    .io_in_1(c53_519_io_in_1),
    .io_in_2(c53_519_io_in_2),
    .io_in_3(c53_519_io_in_3),
    .io_in_4(c53_519_io_in_4),
    .io_out_0(c53_519_io_out_0),
    .io_out_1(c53_519_io_out_1),
    .io_out_2(c53_519_io_out_2)
  );
  C22 c22_61 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_61_io_in_0),
    .io_in_1(c22_61_io_in_1),
    .io_out_0(c22_61_io_out_0),
    .io_out_1(c22_61_io_out_1)
  );
  C53 c53_520 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_520_io_in_0),
    .io_in_1(c53_520_io_in_1),
    .io_in_2(c53_520_io_in_2),
    .io_in_3(c53_520_io_in_3),
    .io_in_4(c53_520_io_in_4),
    .io_out_0(c53_520_io_out_0),
    .io_out_1(c53_520_io_out_1),
    .io_out_2(c53_520_io_out_2)
  );
  C22 c22_62 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_62_io_in_0),
    .io_in_1(c22_62_io_in_1),
    .io_out_0(c22_62_io_out_0),
    .io_out_1(c22_62_io_out_1)
  );
  C53 c53_521 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_521_io_in_0),
    .io_in_1(c53_521_io_in_1),
    .io_in_2(c53_521_io_in_2),
    .io_in_3(c53_521_io_in_3),
    .io_in_4(c53_521_io_in_4),
    .io_out_0(c53_521_io_out_0),
    .io_out_1(c53_521_io_out_1),
    .io_out_2(c53_521_io_out_2)
  );
  C22 c22_63 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_63_io_in_0),
    .io_in_1(c22_63_io_in_1),
    .io_out_0(c22_63_io_out_0),
    .io_out_1(c22_63_io_out_1)
  );
  C53 c53_522 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_522_io_in_0),
    .io_in_1(c53_522_io_in_1),
    .io_in_2(c53_522_io_in_2),
    .io_in_3(c53_522_io_in_3),
    .io_in_4(c53_522_io_in_4),
    .io_out_0(c53_522_io_out_0),
    .io_out_1(c53_522_io_out_1),
    .io_out_2(c53_522_io_out_2)
  );
  C22 c22_64 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_64_io_in_0),
    .io_in_1(c22_64_io_in_1),
    .io_out_0(c22_64_io_out_0),
    .io_out_1(c22_64_io_out_1)
  );
  C53 c53_523 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_523_io_in_0),
    .io_in_1(c53_523_io_in_1),
    .io_in_2(c53_523_io_in_2),
    .io_in_3(c53_523_io_in_3),
    .io_in_4(c53_523_io_in_4),
    .io_out_0(c53_523_io_out_0),
    .io_out_1(c53_523_io_out_1),
    .io_out_2(c53_523_io_out_2)
  );
  C53 c53_524 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_524_io_in_0),
    .io_in_1(c53_524_io_in_1),
    .io_in_2(c53_524_io_in_2),
    .io_in_3(c53_524_io_in_3),
    .io_in_4(c53_524_io_in_4),
    .io_out_0(c53_524_io_out_0),
    .io_out_1(c53_524_io_out_1),
    .io_out_2(c53_524_io_out_2)
  );
  C53 c53_525 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_525_io_in_0),
    .io_in_1(c53_525_io_in_1),
    .io_in_2(c53_525_io_in_2),
    .io_in_3(c53_525_io_in_3),
    .io_in_4(c53_525_io_in_4),
    .io_out_0(c53_525_io_out_0),
    .io_out_1(c53_525_io_out_1),
    .io_out_2(c53_525_io_out_2)
  );
  C53 c53_526 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_526_io_in_0),
    .io_in_1(c53_526_io_in_1),
    .io_in_2(c53_526_io_in_2),
    .io_in_3(c53_526_io_in_3),
    .io_in_4(c53_526_io_in_4),
    .io_out_0(c53_526_io_out_0),
    .io_out_1(c53_526_io_out_1),
    .io_out_2(c53_526_io_out_2)
  );
  C53 c53_527 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_527_io_in_0),
    .io_in_1(c53_527_io_in_1),
    .io_in_2(c53_527_io_in_2),
    .io_in_3(c53_527_io_in_3),
    .io_in_4(c53_527_io_in_4),
    .io_out_0(c53_527_io_out_0),
    .io_out_1(c53_527_io_out_1),
    .io_out_2(c53_527_io_out_2)
  );
  C53 c53_528 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_528_io_in_0),
    .io_in_1(c53_528_io_in_1),
    .io_in_2(c53_528_io_in_2),
    .io_in_3(c53_528_io_in_3),
    .io_in_4(c53_528_io_in_4),
    .io_out_0(c53_528_io_out_0),
    .io_out_1(c53_528_io_out_1),
    .io_out_2(c53_528_io_out_2)
  );
  C53 c53_529 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_529_io_in_0),
    .io_in_1(c53_529_io_in_1),
    .io_in_2(c53_529_io_in_2),
    .io_in_3(c53_529_io_in_3),
    .io_in_4(c53_529_io_in_4),
    .io_out_0(c53_529_io_out_0),
    .io_out_1(c53_529_io_out_1),
    .io_out_2(c53_529_io_out_2)
  );
  C53 c53_530 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_530_io_in_0),
    .io_in_1(c53_530_io_in_1),
    .io_in_2(c53_530_io_in_2),
    .io_in_3(c53_530_io_in_3),
    .io_in_4(c53_530_io_in_4),
    .io_out_0(c53_530_io_out_0),
    .io_out_1(c53_530_io_out_1),
    .io_out_2(c53_530_io_out_2)
  );
  C32 c32_45 ( // @[Multiplier.scala 78:25]
    .io_in_0(c32_45_io_in_0),
    .io_in_1(c32_45_io_in_1),
    .io_in_2(c32_45_io_in_2),
    .io_out_0(c32_45_io_out_0),
    .io_out_1(c32_45_io_out_1)
  );
  C22 c22_65 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_65_io_in_0),
    .io_in_1(c22_65_io_in_1),
    .io_out_0(c22_65_io_out_0),
    .io_out_1(c22_65_io_out_1)
  );
  C22 c22_66 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_66_io_in_0),
    .io_in_1(c22_66_io_in_1),
    .io_out_0(c22_66_io_out_0),
    .io_out_1(c22_66_io_out_1)
  );
  C32 c32_46 ( // @[Multiplier.scala 78:25]
    .io_in_0(c32_46_io_in_0),
    .io_in_1(c32_46_io_in_1),
    .io_in_2(c32_46_io_in_2),
    .io_out_0(c32_46_io_out_0),
    .io_out_1(c32_46_io_out_1)
  );
  C22 c22_67 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_67_io_in_0),
    .io_in_1(c22_67_io_in_1),
    .io_out_0(c22_67_io_out_0),
    .io_out_1(c22_67_io_out_1)
  );
  C22 c22_68 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_68_io_in_0),
    .io_in_1(c22_68_io_in_1),
    .io_out_0(c22_68_io_out_0),
    .io_out_1(c22_68_io_out_1)
  );
  C22 c22_69 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_69_io_in_0),
    .io_in_1(c22_69_io_in_1),
    .io_out_0(c22_69_io_out_0),
    .io_out_1(c22_69_io_out_1)
  );
  C22 c22_70 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_70_io_in_0),
    .io_in_1(c22_70_io_in_1),
    .io_out_0(c22_70_io_out_0),
    .io_out_1(c22_70_io_out_1)
  );
  C22 c22_71 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_71_io_in_0),
    .io_in_1(c22_71_io_in_1),
    .io_out_0(c22_71_io_out_0),
    .io_out_1(c22_71_io_out_1)
  );
  C22 c22_72 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_72_io_in_0),
    .io_in_1(c22_72_io_in_1),
    .io_out_0(c22_72_io_out_0),
    .io_out_1(c22_72_io_out_1)
  );
  C22 c22_73 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_73_io_in_0),
    .io_in_1(c22_73_io_in_1),
    .io_out_0(c22_73_io_out_0),
    .io_out_1(c22_73_io_out_1)
  );
  C22 c22_74 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_74_io_in_0),
    .io_in_1(c22_74_io_in_1),
    .io_out_0(c22_74_io_out_0),
    .io_out_1(c22_74_io_out_1)
  );
  C22 c22_75 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_75_io_in_0),
    .io_in_1(c22_75_io_in_1),
    .io_out_0(c22_75_io_out_0),
    .io_out_1(c22_75_io_out_1)
  );
  C22 c22_76 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_76_io_in_0),
    .io_in_1(c22_76_io_in_1),
    .io_out_0(c22_76_io_out_0),
    .io_out_1(c22_76_io_out_1)
  );
  C22 c22_77 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_77_io_in_0),
    .io_in_1(c22_77_io_in_1),
    .io_out_0(c22_77_io_out_0),
    .io_out_1(c22_77_io_out_1)
  );
  C22 c22_78 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_78_io_in_0),
    .io_in_1(c22_78_io_in_1),
    .io_out_0(c22_78_io_out_0),
    .io_out_1(c22_78_io_out_1)
  );
  C22 c22_79 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_79_io_in_0),
    .io_in_1(c22_79_io_in_1),
    .io_out_0(c22_79_io_out_0),
    .io_out_1(c22_79_io_out_1)
  );
  C22 c22_80 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_80_io_in_0),
    .io_in_1(c22_80_io_in_1),
    .io_out_0(c22_80_io_out_0),
    .io_out_1(c22_80_io_out_1)
  );
  C22 c22_81 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_81_io_in_0),
    .io_in_1(c22_81_io_in_1),
    .io_out_0(c22_81_io_out_0),
    .io_out_1(c22_81_io_out_1)
  );
  C22 c22_82 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_82_io_in_0),
    .io_in_1(c22_82_io_in_1),
    .io_out_0(c22_82_io_out_0),
    .io_out_1(c22_82_io_out_1)
  );
  C32 c32_47 ( // @[Multiplier.scala 78:25]
    .io_in_0(c32_47_io_in_0),
    .io_in_1(c32_47_io_in_1),
    .io_in_2(c32_47_io_in_2),
    .io_out_0(c32_47_io_out_0),
    .io_out_1(c32_47_io_out_1)
  );
  C32 c32_48 ( // @[Multiplier.scala 78:25]
    .io_in_0(c32_48_io_in_0),
    .io_in_1(c32_48_io_in_1),
    .io_in_2(c32_48_io_in_2),
    .io_out_0(c32_48_io_out_0),
    .io_out_1(c32_48_io_out_1)
  );
  C32 c32_49 ( // @[Multiplier.scala 78:25]
    .io_in_0(c32_49_io_in_0),
    .io_in_1(c32_49_io_in_1),
    .io_in_2(c32_49_io_in_2),
    .io_out_0(c32_49_io_out_0),
    .io_out_1(c32_49_io_out_1)
  );
  C32 c32_50 ( // @[Multiplier.scala 78:25]
    .io_in_0(c32_50_io_in_0),
    .io_in_1(c32_50_io_in_1),
    .io_in_2(c32_50_io_in_2),
    .io_out_0(c32_50_io_out_0),
    .io_out_1(c32_50_io_out_1)
  );
  C53 c53_531 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_531_io_in_0),
    .io_in_1(c53_531_io_in_1),
    .io_in_2(c53_531_io_in_2),
    .io_in_3(c53_531_io_in_3),
    .io_in_4(c53_531_io_in_4),
    .io_out_0(c53_531_io_out_0),
    .io_out_1(c53_531_io_out_1),
    .io_out_2(c53_531_io_out_2)
  );
  C53 c53_532 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_532_io_in_0),
    .io_in_1(c53_532_io_in_1),
    .io_in_2(c53_532_io_in_2),
    .io_in_3(c53_532_io_in_3),
    .io_in_4(c53_532_io_in_4),
    .io_out_0(c53_532_io_out_0),
    .io_out_1(c53_532_io_out_1),
    .io_out_2(c53_532_io_out_2)
  );
  C53 c53_533 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_533_io_in_0),
    .io_in_1(c53_533_io_in_1),
    .io_in_2(c53_533_io_in_2),
    .io_in_3(c53_533_io_in_3),
    .io_in_4(c53_533_io_in_4),
    .io_out_0(c53_533_io_out_0),
    .io_out_1(c53_533_io_out_1),
    .io_out_2(c53_533_io_out_2)
  );
  C53 c53_534 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_534_io_in_0),
    .io_in_1(c53_534_io_in_1),
    .io_in_2(c53_534_io_in_2),
    .io_in_3(c53_534_io_in_3),
    .io_in_4(c53_534_io_in_4),
    .io_out_0(c53_534_io_out_0),
    .io_out_1(c53_534_io_out_1),
    .io_out_2(c53_534_io_out_2)
  );
  C53 c53_535 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_535_io_in_0),
    .io_in_1(c53_535_io_in_1),
    .io_in_2(c53_535_io_in_2),
    .io_in_3(c53_535_io_in_3),
    .io_in_4(c53_535_io_in_4),
    .io_out_0(c53_535_io_out_0),
    .io_out_1(c53_535_io_out_1),
    .io_out_2(c53_535_io_out_2)
  );
  C53 c53_536 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_536_io_in_0),
    .io_in_1(c53_536_io_in_1),
    .io_in_2(c53_536_io_in_2),
    .io_in_3(c53_536_io_in_3),
    .io_in_4(c53_536_io_in_4),
    .io_out_0(c53_536_io_out_0),
    .io_out_1(c53_536_io_out_1),
    .io_out_2(c53_536_io_out_2)
  );
  C53 c53_537 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_537_io_in_0),
    .io_in_1(c53_537_io_in_1),
    .io_in_2(c53_537_io_in_2),
    .io_in_3(c53_537_io_in_3),
    .io_in_4(c53_537_io_in_4),
    .io_out_0(c53_537_io_out_0),
    .io_out_1(c53_537_io_out_1),
    .io_out_2(c53_537_io_out_2)
  );
  C53 c53_538 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_538_io_in_0),
    .io_in_1(c53_538_io_in_1),
    .io_in_2(c53_538_io_in_2),
    .io_in_3(c53_538_io_in_3),
    .io_in_4(c53_538_io_in_4),
    .io_out_0(c53_538_io_out_0),
    .io_out_1(c53_538_io_out_1),
    .io_out_2(c53_538_io_out_2)
  );
  C53 c53_539 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_539_io_in_0),
    .io_in_1(c53_539_io_in_1),
    .io_in_2(c53_539_io_in_2),
    .io_in_3(c53_539_io_in_3),
    .io_in_4(c53_539_io_in_4),
    .io_out_0(c53_539_io_out_0),
    .io_out_1(c53_539_io_out_1),
    .io_out_2(c53_539_io_out_2)
  );
  C53 c53_540 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_540_io_in_0),
    .io_in_1(c53_540_io_in_1),
    .io_in_2(c53_540_io_in_2),
    .io_in_3(c53_540_io_in_3),
    .io_in_4(c53_540_io_in_4),
    .io_out_0(c53_540_io_out_0),
    .io_out_1(c53_540_io_out_1),
    .io_out_2(c53_540_io_out_2)
  );
  C53 c53_541 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_541_io_in_0),
    .io_in_1(c53_541_io_in_1),
    .io_in_2(c53_541_io_in_2),
    .io_in_3(c53_541_io_in_3),
    .io_in_4(c53_541_io_in_4),
    .io_out_0(c53_541_io_out_0),
    .io_out_1(c53_541_io_out_1),
    .io_out_2(c53_541_io_out_2)
  );
  C53 c53_542 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_542_io_in_0),
    .io_in_1(c53_542_io_in_1),
    .io_in_2(c53_542_io_in_2),
    .io_in_3(c53_542_io_in_3),
    .io_in_4(c53_542_io_in_4),
    .io_out_0(c53_542_io_out_0),
    .io_out_1(c53_542_io_out_1),
    .io_out_2(c53_542_io_out_2)
  );
  C53 c53_543 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_543_io_in_0),
    .io_in_1(c53_543_io_in_1),
    .io_in_2(c53_543_io_in_2),
    .io_in_3(c53_543_io_in_3),
    .io_in_4(c53_543_io_in_4),
    .io_out_0(c53_543_io_out_0),
    .io_out_1(c53_543_io_out_1),
    .io_out_2(c53_543_io_out_2)
  );
  C53 c53_544 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_544_io_in_0),
    .io_in_1(c53_544_io_in_1),
    .io_in_2(c53_544_io_in_2),
    .io_in_3(c53_544_io_in_3),
    .io_in_4(c53_544_io_in_4),
    .io_out_0(c53_544_io_out_0),
    .io_out_1(c53_544_io_out_1),
    .io_out_2(c53_544_io_out_2)
  );
  C53 c53_545 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_545_io_in_0),
    .io_in_1(c53_545_io_in_1),
    .io_in_2(c53_545_io_in_2),
    .io_in_3(c53_545_io_in_3),
    .io_in_4(c53_545_io_in_4),
    .io_out_0(c53_545_io_out_0),
    .io_out_1(c53_545_io_out_1),
    .io_out_2(c53_545_io_out_2)
  );
  C53 c53_546 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_546_io_in_0),
    .io_in_1(c53_546_io_in_1),
    .io_in_2(c53_546_io_in_2),
    .io_in_3(c53_546_io_in_3),
    .io_in_4(c53_546_io_in_4),
    .io_out_0(c53_546_io_out_0),
    .io_out_1(c53_546_io_out_1),
    .io_out_2(c53_546_io_out_2)
  );
  C53 c53_547 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_547_io_in_0),
    .io_in_1(c53_547_io_in_1),
    .io_in_2(c53_547_io_in_2),
    .io_in_3(c53_547_io_in_3),
    .io_in_4(c53_547_io_in_4),
    .io_out_0(c53_547_io_out_0),
    .io_out_1(c53_547_io_out_1),
    .io_out_2(c53_547_io_out_2)
  );
  C22 c22_83 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_83_io_in_0),
    .io_in_1(c22_83_io_in_1),
    .io_out_0(c22_83_io_out_0),
    .io_out_1(c22_83_io_out_1)
  );
  C53 c53_548 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_548_io_in_0),
    .io_in_1(c53_548_io_in_1),
    .io_in_2(c53_548_io_in_2),
    .io_in_3(c53_548_io_in_3),
    .io_in_4(c53_548_io_in_4),
    .io_out_0(c53_548_io_out_0),
    .io_out_1(c53_548_io_out_1),
    .io_out_2(c53_548_io_out_2)
  );
  C22 c22_84 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_84_io_in_0),
    .io_in_1(c22_84_io_in_1),
    .io_out_0(c22_84_io_out_0),
    .io_out_1(c22_84_io_out_1)
  );
  C53 c53_549 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_549_io_in_0),
    .io_in_1(c53_549_io_in_1),
    .io_in_2(c53_549_io_in_2),
    .io_in_3(c53_549_io_in_3),
    .io_in_4(c53_549_io_in_4),
    .io_out_0(c53_549_io_out_0),
    .io_out_1(c53_549_io_out_1),
    .io_out_2(c53_549_io_out_2)
  );
  C22 c22_85 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_85_io_in_0),
    .io_in_1(c22_85_io_in_1),
    .io_out_0(c22_85_io_out_0),
    .io_out_1(c22_85_io_out_1)
  );
  C53 c53_550 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_550_io_in_0),
    .io_in_1(c53_550_io_in_1),
    .io_in_2(c53_550_io_in_2),
    .io_in_3(c53_550_io_in_3),
    .io_in_4(c53_550_io_in_4),
    .io_out_0(c53_550_io_out_0),
    .io_out_1(c53_550_io_out_1),
    .io_out_2(c53_550_io_out_2)
  );
  C22 c22_86 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_86_io_in_0),
    .io_in_1(c22_86_io_in_1),
    .io_out_0(c22_86_io_out_0),
    .io_out_1(c22_86_io_out_1)
  );
  C53 c53_551 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_551_io_in_0),
    .io_in_1(c53_551_io_in_1),
    .io_in_2(c53_551_io_in_2),
    .io_in_3(c53_551_io_in_3),
    .io_in_4(c53_551_io_in_4),
    .io_out_0(c53_551_io_out_0),
    .io_out_1(c53_551_io_out_1),
    .io_out_2(c53_551_io_out_2)
  );
  C22 c22_87 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_87_io_in_0),
    .io_in_1(c22_87_io_in_1),
    .io_out_0(c22_87_io_out_0),
    .io_out_1(c22_87_io_out_1)
  );
  C53 c53_552 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_552_io_in_0),
    .io_in_1(c53_552_io_in_1),
    .io_in_2(c53_552_io_in_2),
    .io_in_3(c53_552_io_in_3),
    .io_in_4(c53_552_io_in_4),
    .io_out_0(c53_552_io_out_0),
    .io_out_1(c53_552_io_out_1),
    .io_out_2(c53_552_io_out_2)
  );
  C22 c22_88 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_88_io_in_0),
    .io_in_1(c22_88_io_in_1),
    .io_out_0(c22_88_io_out_0),
    .io_out_1(c22_88_io_out_1)
  );
  C53 c53_553 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_553_io_in_0),
    .io_in_1(c53_553_io_in_1),
    .io_in_2(c53_553_io_in_2),
    .io_in_3(c53_553_io_in_3),
    .io_in_4(c53_553_io_in_4),
    .io_out_0(c53_553_io_out_0),
    .io_out_1(c53_553_io_out_1),
    .io_out_2(c53_553_io_out_2)
  );
  C22 c22_89 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_89_io_in_0),
    .io_in_1(c22_89_io_in_1),
    .io_out_0(c22_89_io_out_0),
    .io_out_1(c22_89_io_out_1)
  );
  C53 c53_554 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_554_io_in_0),
    .io_in_1(c53_554_io_in_1),
    .io_in_2(c53_554_io_in_2),
    .io_in_3(c53_554_io_in_3),
    .io_in_4(c53_554_io_in_4),
    .io_out_0(c53_554_io_out_0),
    .io_out_1(c53_554_io_out_1),
    .io_out_2(c53_554_io_out_2)
  );
  C22 c22_90 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_90_io_in_0),
    .io_in_1(c22_90_io_in_1),
    .io_out_0(c22_90_io_out_0),
    .io_out_1(c22_90_io_out_1)
  );
  C53 c53_555 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_555_io_in_0),
    .io_in_1(c53_555_io_in_1),
    .io_in_2(c53_555_io_in_2),
    .io_in_3(c53_555_io_in_3),
    .io_in_4(c53_555_io_in_4),
    .io_out_0(c53_555_io_out_0),
    .io_out_1(c53_555_io_out_1),
    .io_out_2(c53_555_io_out_2)
  );
  C22 c22_91 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_91_io_in_0),
    .io_in_1(c22_91_io_in_1),
    .io_out_0(c22_91_io_out_0),
    .io_out_1(c22_91_io_out_1)
  );
  C53 c53_556 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_556_io_in_0),
    .io_in_1(c53_556_io_in_1),
    .io_in_2(c53_556_io_in_2),
    .io_in_3(c53_556_io_in_3),
    .io_in_4(c53_556_io_in_4),
    .io_out_0(c53_556_io_out_0),
    .io_out_1(c53_556_io_out_1),
    .io_out_2(c53_556_io_out_2)
  );
  C22 c22_92 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_92_io_in_0),
    .io_in_1(c22_92_io_in_1),
    .io_out_0(c22_92_io_out_0),
    .io_out_1(c22_92_io_out_1)
  );
  C53 c53_557 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_557_io_in_0),
    .io_in_1(c53_557_io_in_1),
    .io_in_2(c53_557_io_in_2),
    .io_in_3(c53_557_io_in_3),
    .io_in_4(c53_557_io_in_4),
    .io_out_0(c53_557_io_out_0),
    .io_out_1(c53_557_io_out_1),
    .io_out_2(c53_557_io_out_2)
  );
  C22 c22_93 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_93_io_in_0),
    .io_in_1(c22_93_io_in_1),
    .io_out_0(c22_93_io_out_0),
    .io_out_1(c22_93_io_out_1)
  );
  C53 c53_558 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_558_io_in_0),
    .io_in_1(c53_558_io_in_1),
    .io_in_2(c53_558_io_in_2),
    .io_in_3(c53_558_io_in_3),
    .io_in_4(c53_558_io_in_4),
    .io_out_0(c53_558_io_out_0),
    .io_out_1(c53_558_io_out_1),
    .io_out_2(c53_558_io_out_2)
  );
  C22 c22_94 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_94_io_in_0),
    .io_in_1(c22_94_io_in_1),
    .io_out_0(c22_94_io_out_0),
    .io_out_1(c22_94_io_out_1)
  );
  C53 c53_559 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_559_io_in_0),
    .io_in_1(c53_559_io_in_1),
    .io_in_2(c53_559_io_in_2),
    .io_in_3(c53_559_io_in_3),
    .io_in_4(c53_559_io_in_4),
    .io_out_0(c53_559_io_out_0),
    .io_out_1(c53_559_io_out_1),
    .io_out_2(c53_559_io_out_2)
  );
  C32 c32_51 ( // @[Multiplier.scala 78:25]
    .io_in_0(c32_51_io_in_0),
    .io_in_1(c32_51_io_in_1),
    .io_in_2(c32_51_io_in_2),
    .io_out_0(c32_51_io_out_0),
    .io_out_1(c32_51_io_out_1)
  );
  C53 c53_560 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_560_io_in_0),
    .io_in_1(c53_560_io_in_1),
    .io_in_2(c53_560_io_in_2),
    .io_in_3(c53_560_io_in_3),
    .io_in_4(c53_560_io_in_4),
    .io_out_0(c53_560_io_out_0),
    .io_out_1(c53_560_io_out_1),
    .io_out_2(c53_560_io_out_2)
  );
  C32 c32_52 ( // @[Multiplier.scala 78:25]
    .io_in_0(c32_52_io_in_0),
    .io_in_1(c32_52_io_in_1),
    .io_in_2(c32_52_io_in_2),
    .io_out_0(c32_52_io_out_0),
    .io_out_1(c32_52_io_out_1)
  );
  C53 c53_561 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_561_io_in_0),
    .io_in_1(c53_561_io_in_1),
    .io_in_2(c53_561_io_in_2),
    .io_in_3(c53_561_io_in_3),
    .io_in_4(c53_561_io_in_4),
    .io_out_0(c53_561_io_out_0),
    .io_out_1(c53_561_io_out_1),
    .io_out_2(c53_561_io_out_2)
  );
  C32 c32_53 ( // @[Multiplier.scala 78:25]
    .io_in_0(c32_53_io_in_0),
    .io_in_1(c32_53_io_in_1),
    .io_in_2(c32_53_io_in_2),
    .io_out_0(c32_53_io_out_0),
    .io_out_1(c32_53_io_out_1)
  );
  C53 c53_562 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_562_io_in_0),
    .io_in_1(c53_562_io_in_1),
    .io_in_2(c53_562_io_in_2),
    .io_in_3(c53_562_io_in_3),
    .io_in_4(c53_562_io_in_4),
    .io_out_0(c53_562_io_out_0),
    .io_out_1(c53_562_io_out_1),
    .io_out_2(c53_562_io_out_2)
  );
  C32 c32_54 ( // @[Multiplier.scala 78:25]
    .io_in_0(c32_54_io_in_0),
    .io_in_1(c32_54_io_in_1),
    .io_in_2(c32_54_io_in_2),
    .io_out_0(c32_54_io_out_0),
    .io_out_1(c32_54_io_out_1)
  );
  C53 c53_563 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_563_io_in_0),
    .io_in_1(c53_563_io_in_1),
    .io_in_2(c53_563_io_in_2),
    .io_in_3(c53_563_io_in_3),
    .io_in_4(c53_563_io_in_4),
    .io_out_0(c53_563_io_out_0),
    .io_out_1(c53_563_io_out_1),
    .io_out_2(c53_563_io_out_2)
  );
  C53 c53_564 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_564_io_in_0),
    .io_in_1(c53_564_io_in_1),
    .io_in_2(c53_564_io_in_2),
    .io_in_3(c53_564_io_in_3),
    .io_in_4(c53_564_io_in_4),
    .io_out_0(c53_564_io_out_0),
    .io_out_1(c53_564_io_out_1),
    .io_out_2(c53_564_io_out_2)
  );
  C53 c53_565 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_565_io_in_0),
    .io_in_1(c53_565_io_in_1),
    .io_in_2(c53_565_io_in_2),
    .io_in_3(c53_565_io_in_3),
    .io_in_4(c53_565_io_in_4),
    .io_out_0(c53_565_io_out_0),
    .io_out_1(c53_565_io_out_1),
    .io_out_2(c53_565_io_out_2)
  );
  C53 c53_566 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_566_io_in_0),
    .io_in_1(c53_566_io_in_1),
    .io_in_2(c53_566_io_in_2),
    .io_in_3(c53_566_io_in_3),
    .io_in_4(c53_566_io_in_4),
    .io_out_0(c53_566_io_out_0),
    .io_out_1(c53_566_io_out_1),
    .io_out_2(c53_566_io_out_2)
  );
  C53 c53_567 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_567_io_in_0),
    .io_in_1(c53_567_io_in_1),
    .io_in_2(c53_567_io_in_2),
    .io_in_3(c53_567_io_in_3),
    .io_in_4(c53_567_io_in_4),
    .io_out_0(c53_567_io_out_0),
    .io_out_1(c53_567_io_out_1),
    .io_out_2(c53_567_io_out_2)
  );
  C53 c53_568 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_568_io_in_0),
    .io_in_1(c53_568_io_in_1),
    .io_in_2(c53_568_io_in_2),
    .io_in_3(c53_568_io_in_3),
    .io_in_4(c53_568_io_in_4),
    .io_out_0(c53_568_io_out_0),
    .io_out_1(c53_568_io_out_1),
    .io_out_2(c53_568_io_out_2)
  );
  C53 c53_569 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_569_io_in_0),
    .io_in_1(c53_569_io_in_1),
    .io_in_2(c53_569_io_in_2),
    .io_in_3(c53_569_io_in_3),
    .io_in_4(c53_569_io_in_4),
    .io_out_0(c53_569_io_out_0),
    .io_out_1(c53_569_io_out_1),
    .io_out_2(c53_569_io_out_2)
  );
  C53 c53_570 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_570_io_in_0),
    .io_in_1(c53_570_io_in_1),
    .io_in_2(c53_570_io_in_2),
    .io_in_3(c53_570_io_in_3),
    .io_in_4(c53_570_io_in_4),
    .io_out_0(c53_570_io_out_0),
    .io_out_1(c53_570_io_out_1),
    .io_out_2(c53_570_io_out_2)
  );
  C53 c53_571 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_571_io_in_0),
    .io_in_1(c53_571_io_in_1),
    .io_in_2(c53_571_io_in_2),
    .io_in_3(c53_571_io_in_3),
    .io_in_4(c53_571_io_in_4),
    .io_out_0(c53_571_io_out_0),
    .io_out_1(c53_571_io_out_1),
    .io_out_2(c53_571_io_out_2)
  );
  C53 c53_572 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_572_io_in_0),
    .io_in_1(c53_572_io_in_1),
    .io_in_2(c53_572_io_in_2),
    .io_in_3(c53_572_io_in_3),
    .io_in_4(c53_572_io_in_4),
    .io_out_0(c53_572_io_out_0),
    .io_out_1(c53_572_io_out_1),
    .io_out_2(c53_572_io_out_2)
  );
  C53 c53_573 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_573_io_in_0),
    .io_in_1(c53_573_io_in_1),
    .io_in_2(c53_573_io_in_2),
    .io_in_3(c53_573_io_in_3),
    .io_in_4(c53_573_io_in_4),
    .io_out_0(c53_573_io_out_0),
    .io_out_1(c53_573_io_out_1),
    .io_out_2(c53_573_io_out_2)
  );
  C53 c53_574 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_574_io_in_0),
    .io_in_1(c53_574_io_in_1),
    .io_in_2(c53_574_io_in_2),
    .io_in_3(c53_574_io_in_3),
    .io_in_4(c53_574_io_in_4),
    .io_out_0(c53_574_io_out_0),
    .io_out_1(c53_574_io_out_1),
    .io_out_2(c53_574_io_out_2)
  );
  C53 c53_575 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_575_io_in_0),
    .io_in_1(c53_575_io_in_1),
    .io_in_2(c53_575_io_in_2),
    .io_in_3(c53_575_io_in_3),
    .io_in_4(c53_575_io_in_4),
    .io_out_0(c53_575_io_out_0),
    .io_out_1(c53_575_io_out_1),
    .io_out_2(c53_575_io_out_2)
  );
  C53 c53_576 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_576_io_in_0),
    .io_in_1(c53_576_io_in_1),
    .io_in_2(c53_576_io_in_2),
    .io_in_3(c53_576_io_in_3),
    .io_in_4(c53_576_io_in_4),
    .io_out_0(c53_576_io_out_0),
    .io_out_1(c53_576_io_out_1),
    .io_out_2(c53_576_io_out_2)
  );
  C53 c53_577 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_577_io_in_0),
    .io_in_1(c53_577_io_in_1),
    .io_in_2(c53_577_io_in_2),
    .io_in_3(c53_577_io_in_3),
    .io_in_4(c53_577_io_in_4),
    .io_out_0(c53_577_io_out_0),
    .io_out_1(c53_577_io_out_1),
    .io_out_2(c53_577_io_out_2)
  );
  C53 c53_578 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_578_io_in_0),
    .io_in_1(c53_578_io_in_1),
    .io_in_2(c53_578_io_in_2),
    .io_in_3(c53_578_io_in_3),
    .io_in_4(c53_578_io_in_4),
    .io_out_0(c53_578_io_out_0),
    .io_out_1(c53_578_io_out_1),
    .io_out_2(c53_578_io_out_2)
  );
  C53 c53_579 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_579_io_in_0),
    .io_in_1(c53_579_io_in_1),
    .io_in_2(c53_579_io_in_2),
    .io_in_3(c53_579_io_in_3),
    .io_in_4(c53_579_io_in_4),
    .io_out_0(c53_579_io_out_0),
    .io_out_1(c53_579_io_out_1),
    .io_out_2(c53_579_io_out_2)
  );
  C53 c53_580 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_580_io_in_0),
    .io_in_1(c53_580_io_in_1),
    .io_in_2(c53_580_io_in_2),
    .io_in_3(c53_580_io_in_3),
    .io_in_4(c53_580_io_in_4),
    .io_out_0(c53_580_io_out_0),
    .io_out_1(c53_580_io_out_1),
    .io_out_2(c53_580_io_out_2)
  );
  C53 c53_581 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_581_io_in_0),
    .io_in_1(c53_581_io_in_1),
    .io_in_2(c53_581_io_in_2),
    .io_in_3(c53_581_io_in_3),
    .io_in_4(c53_581_io_in_4),
    .io_out_0(c53_581_io_out_0),
    .io_out_1(c53_581_io_out_1),
    .io_out_2(c53_581_io_out_2)
  );
  C53 c53_582 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_582_io_in_0),
    .io_in_1(c53_582_io_in_1),
    .io_in_2(c53_582_io_in_2),
    .io_in_3(c53_582_io_in_3),
    .io_in_4(c53_582_io_in_4),
    .io_out_0(c53_582_io_out_0),
    .io_out_1(c53_582_io_out_1),
    .io_out_2(c53_582_io_out_2)
  );
  C53 c53_583 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_583_io_in_0),
    .io_in_1(c53_583_io_in_1),
    .io_in_2(c53_583_io_in_2),
    .io_in_3(c53_583_io_in_3),
    .io_in_4(c53_583_io_in_4),
    .io_out_0(c53_583_io_out_0),
    .io_out_1(c53_583_io_out_1),
    .io_out_2(c53_583_io_out_2)
  );
  C53 c53_584 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_584_io_in_0),
    .io_in_1(c53_584_io_in_1),
    .io_in_2(c53_584_io_in_2),
    .io_in_3(c53_584_io_in_3),
    .io_in_4(c53_584_io_in_4),
    .io_out_0(c53_584_io_out_0),
    .io_out_1(c53_584_io_out_1),
    .io_out_2(c53_584_io_out_2)
  );
  C53 c53_585 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_585_io_in_0),
    .io_in_1(c53_585_io_in_1),
    .io_in_2(c53_585_io_in_2),
    .io_in_3(c53_585_io_in_3),
    .io_in_4(c53_585_io_in_4),
    .io_out_0(c53_585_io_out_0),
    .io_out_1(c53_585_io_out_1),
    .io_out_2(c53_585_io_out_2)
  );
  C22 c22_95 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_95_io_in_0),
    .io_in_1(c22_95_io_in_1),
    .io_out_0(c22_95_io_out_0),
    .io_out_1(c22_95_io_out_1)
  );
  C53 c53_586 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_586_io_in_0),
    .io_in_1(c53_586_io_in_1),
    .io_in_2(c53_586_io_in_2),
    .io_in_3(c53_586_io_in_3),
    .io_in_4(c53_586_io_in_4),
    .io_out_0(c53_586_io_out_0),
    .io_out_1(c53_586_io_out_1),
    .io_out_2(c53_586_io_out_2)
  );
  C22 c22_96 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_96_io_in_0),
    .io_in_1(c22_96_io_in_1),
    .io_out_0(c22_96_io_out_0),
    .io_out_1(c22_96_io_out_1)
  );
  C53 c53_587 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_587_io_in_0),
    .io_in_1(c53_587_io_in_1),
    .io_in_2(c53_587_io_in_2),
    .io_in_3(c53_587_io_in_3),
    .io_in_4(c53_587_io_in_4),
    .io_out_0(c53_587_io_out_0),
    .io_out_1(c53_587_io_out_1),
    .io_out_2(c53_587_io_out_2)
  );
  C32 c32_55 ( // @[Multiplier.scala 78:25]
    .io_in_0(c32_55_io_in_0),
    .io_in_1(c32_55_io_in_1),
    .io_in_2(c32_55_io_in_2),
    .io_out_0(c32_55_io_out_0),
    .io_out_1(c32_55_io_out_1)
  );
  C53 c53_588 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_588_io_in_0),
    .io_in_1(c53_588_io_in_1),
    .io_in_2(c53_588_io_in_2),
    .io_in_3(c53_588_io_in_3),
    .io_in_4(c53_588_io_in_4),
    .io_out_0(c53_588_io_out_0),
    .io_out_1(c53_588_io_out_1),
    .io_out_2(c53_588_io_out_2)
  );
  C22 c22_97 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_97_io_in_0),
    .io_in_1(c22_97_io_in_1),
    .io_out_0(c22_97_io_out_0),
    .io_out_1(c22_97_io_out_1)
  );
  C53 c53_589 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_589_io_in_0),
    .io_in_1(c53_589_io_in_1),
    .io_in_2(c53_589_io_in_2),
    .io_in_3(c53_589_io_in_3),
    .io_in_4(c53_589_io_in_4),
    .io_out_0(c53_589_io_out_0),
    .io_out_1(c53_589_io_out_1),
    .io_out_2(c53_589_io_out_2)
  );
  C22 c22_98 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_98_io_in_0),
    .io_in_1(c22_98_io_in_1),
    .io_out_0(c22_98_io_out_0),
    .io_out_1(c22_98_io_out_1)
  );
  C53 c53_590 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_590_io_in_0),
    .io_in_1(c53_590_io_in_1),
    .io_in_2(c53_590_io_in_2),
    .io_in_3(c53_590_io_in_3),
    .io_in_4(c53_590_io_in_4),
    .io_out_0(c53_590_io_out_0),
    .io_out_1(c53_590_io_out_1),
    .io_out_2(c53_590_io_out_2)
  );
  C22 c22_99 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_99_io_in_0),
    .io_in_1(c22_99_io_in_1),
    .io_out_0(c22_99_io_out_0),
    .io_out_1(c22_99_io_out_1)
  );
  C53 c53_591 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_591_io_in_0),
    .io_in_1(c53_591_io_in_1),
    .io_in_2(c53_591_io_in_2),
    .io_in_3(c53_591_io_in_3),
    .io_in_4(c53_591_io_in_4),
    .io_out_0(c53_591_io_out_0),
    .io_out_1(c53_591_io_out_1),
    .io_out_2(c53_591_io_out_2)
  );
  C22 c22_100 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_100_io_in_0),
    .io_in_1(c22_100_io_in_1),
    .io_out_0(c22_100_io_out_0),
    .io_out_1(c22_100_io_out_1)
  );
  C53 c53_592 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_592_io_in_0),
    .io_in_1(c53_592_io_in_1),
    .io_in_2(c53_592_io_in_2),
    .io_in_3(c53_592_io_in_3),
    .io_in_4(c53_592_io_in_4),
    .io_out_0(c53_592_io_out_0),
    .io_out_1(c53_592_io_out_1),
    .io_out_2(c53_592_io_out_2)
  );
  C32 c32_56 ( // @[Multiplier.scala 78:25]
    .io_in_0(c32_56_io_in_0),
    .io_in_1(c32_56_io_in_1),
    .io_in_2(c32_56_io_in_2),
    .io_out_0(c32_56_io_out_0),
    .io_out_1(c32_56_io_out_1)
  );
  C53 c53_593 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_593_io_in_0),
    .io_in_1(c53_593_io_in_1),
    .io_in_2(c53_593_io_in_2),
    .io_in_3(c53_593_io_in_3),
    .io_in_4(c53_593_io_in_4),
    .io_out_0(c53_593_io_out_0),
    .io_out_1(c53_593_io_out_1),
    .io_out_2(c53_593_io_out_2)
  );
  C22 c22_101 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_101_io_in_0),
    .io_in_1(c22_101_io_in_1),
    .io_out_0(c22_101_io_out_0),
    .io_out_1(c22_101_io_out_1)
  );
  C53 c53_594 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_594_io_in_0),
    .io_in_1(c53_594_io_in_1),
    .io_in_2(c53_594_io_in_2),
    .io_in_3(c53_594_io_in_3),
    .io_in_4(c53_594_io_in_4),
    .io_out_0(c53_594_io_out_0),
    .io_out_1(c53_594_io_out_1),
    .io_out_2(c53_594_io_out_2)
  );
  C22 c22_102 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_102_io_in_0),
    .io_in_1(c22_102_io_in_1),
    .io_out_0(c22_102_io_out_0),
    .io_out_1(c22_102_io_out_1)
  );
  C53 c53_595 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_595_io_in_0),
    .io_in_1(c53_595_io_in_1),
    .io_in_2(c53_595_io_in_2),
    .io_in_3(c53_595_io_in_3),
    .io_in_4(c53_595_io_in_4),
    .io_out_0(c53_595_io_out_0),
    .io_out_1(c53_595_io_out_1),
    .io_out_2(c53_595_io_out_2)
  );
  C22 c22_103 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_103_io_in_0),
    .io_in_1(c22_103_io_in_1),
    .io_out_0(c22_103_io_out_0),
    .io_out_1(c22_103_io_out_1)
  );
  C53 c53_596 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_596_io_in_0),
    .io_in_1(c53_596_io_in_1),
    .io_in_2(c53_596_io_in_2),
    .io_in_3(c53_596_io_in_3),
    .io_in_4(c53_596_io_in_4),
    .io_out_0(c53_596_io_out_0),
    .io_out_1(c53_596_io_out_1),
    .io_out_2(c53_596_io_out_2)
  );
  C22 c22_104 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_104_io_in_0),
    .io_in_1(c22_104_io_in_1),
    .io_out_0(c22_104_io_out_0),
    .io_out_1(c22_104_io_out_1)
  );
  C53 c53_597 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_597_io_in_0),
    .io_in_1(c53_597_io_in_1),
    .io_in_2(c53_597_io_in_2),
    .io_in_3(c53_597_io_in_3),
    .io_in_4(c53_597_io_in_4),
    .io_out_0(c53_597_io_out_0),
    .io_out_1(c53_597_io_out_1),
    .io_out_2(c53_597_io_out_2)
  );
  C22 c22_105 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_105_io_in_0),
    .io_in_1(c22_105_io_in_1),
    .io_out_0(c22_105_io_out_0),
    .io_out_1(c22_105_io_out_1)
  );
  C53 c53_598 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_598_io_in_0),
    .io_in_1(c53_598_io_in_1),
    .io_in_2(c53_598_io_in_2),
    .io_in_3(c53_598_io_in_3),
    .io_in_4(c53_598_io_in_4),
    .io_out_0(c53_598_io_out_0),
    .io_out_1(c53_598_io_out_1),
    .io_out_2(c53_598_io_out_2)
  );
  C22 c22_106 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_106_io_in_0),
    .io_in_1(c22_106_io_in_1),
    .io_out_0(c22_106_io_out_0),
    .io_out_1(c22_106_io_out_1)
  );
  C53 c53_599 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_599_io_in_0),
    .io_in_1(c53_599_io_in_1),
    .io_in_2(c53_599_io_in_2),
    .io_in_3(c53_599_io_in_3),
    .io_in_4(c53_599_io_in_4),
    .io_out_0(c53_599_io_out_0),
    .io_out_1(c53_599_io_out_1),
    .io_out_2(c53_599_io_out_2)
  );
  C22 c22_107 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_107_io_in_0),
    .io_in_1(c22_107_io_in_1),
    .io_out_0(c22_107_io_out_0),
    .io_out_1(c22_107_io_out_1)
  );
  C53 c53_600 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_600_io_in_0),
    .io_in_1(c53_600_io_in_1),
    .io_in_2(c53_600_io_in_2),
    .io_in_3(c53_600_io_in_3),
    .io_in_4(c53_600_io_in_4),
    .io_out_0(c53_600_io_out_0),
    .io_out_1(c53_600_io_out_1),
    .io_out_2(c53_600_io_out_2)
  );
  C22 c22_108 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_108_io_in_0),
    .io_in_1(c22_108_io_in_1),
    .io_out_0(c22_108_io_out_0),
    .io_out_1(c22_108_io_out_1)
  );
  C53 c53_601 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_601_io_in_0),
    .io_in_1(c53_601_io_in_1),
    .io_in_2(c53_601_io_in_2),
    .io_in_3(c53_601_io_in_3),
    .io_in_4(c53_601_io_in_4),
    .io_out_0(c53_601_io_out_0),
    .io_out_1(c53_601_io_out_1),
    .io_out_2(c53_601_io_out_2)
  );
  C53 c53_602 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_602_io_in_0),
    .io_in_1(c53_602_io_in_1),
    .io_in_2(c53_602_io_in_2),
    .io_in_3(c53_602_io_in_3),
    .io_in_4(c53_602_io_in_4),
    .io_out_0(c53_602_io_out_0),
    .io_out_1(c53_602_io_out_1),
    .io_out_2(c53_602_io_out_2)
  );
  C53 c53_603 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_603_io_in_0),
    .io_in_1(c53_603_io_in_1),
    .io_in_2(c53_603_io_in_2),
    .io_in_3(c53_603_io_in_3),
    .io_in_4(c53_603_io_in_4),
    .io_out_0(c53_603_io_out_0),
    .io_out_1(c53_603_io_out_1),
    .io_out_2(c53_603_io_out_2)
  );
  C53 c53_604 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_604_io_in_0),
    .io_in_1(c53_604_io_in_1),
    .io_in_2(c53_604_io_in_2),
    .io_in_3(c53_604_io_in_3),
    .io_in_4(c53_604_io_in_4),
    .io_out_0(c53_604_io_out_0),
    .io_out_1(c53_604_io_out_1),
    .io_out_2(c53_604_io_out_2)
  );
  C53 c53_605 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_605_io_in_0),
    .io_in_1(c53_605_io_in_1),
    .io_in_2(c53_605_io_in_2),
    .io_in_3(c53_605_io_in_3),
    .io_in_4(c53_605_io_in_4),
    .io_out_0(c53_605_io_out_0),
    .io_out_1(c53_605_io_out_1),
    .io_out_2(c53_605_io_out_2)
  );
  C53 c53_606 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_606_io_in_0),
    .io_in_1(c53_606_io_in_1),
    .io_in_2(c53_606_io_in_2),
    .io_in_3(c53_606_io_in_3),
    .io_in_4(c53_606_io_in_4),
    .io_out_0(c53_606_io_out_0),
    .io_out_1(c53_606_io_out_1),
    .io_out_2(c53_606_io_out_2)
  );
  C53 c53_607 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_607_io_in_0),
    .io_in_1(c53_607_io_in_1),
    .io_in_2(c53_607_io_in_2),
    .io_in_3(c53_607_io_in_3),
    .io_in_4(c53_607_io_in_4),
    .io_out_0(c53_607_io_out_0),
    .io_out_1(c53_607_io_out_1),
    .io_out_2(c53_607_io_out_2)
  );
  C53 c53_608 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_608_io_in_0),
    .io_in_1(c53_608_io_in_1),
    .io_in_2(c53_608_io_in_2),
    .io_in_3(c53_608_io_in_3),
    .io_in_4(c53_608_io_in_4),
    .io_out_0(c53_608_io_out_0),
    .io_out_1(c53_608_io_out_1),
    .io_out_2(c53_608_io_out_2)
  );
  C53 c53_609 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_609_io_in_0),
    .io_in_1(c53_609_io_in_1),
    .io_in_2(c53_609_io_in_2),
    .io_in_3(c53_609_io_in_3),
    .io_in_4(c53_609_io_in_4),
    .io_out_0(c53_609_io_out_0),
    .io_out_1(c53_609_io_out_1),
    .io_out_2(c53_609_io_out_2)
  );
  C53 c53_610 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_610_io_in_0),
    .io_in_1(c53_610_io_in_1),
    .io_in_2(c53_610_io_in_2),
    .io_in_3(c53_610_io_in_3),
    .io_in_4(c53_610_io_in_4),
    .io_out_0(c53_610_io_out_0),
    .io_out_1(c53_610_io_out_1),
    .io_out_2(c53_610_io_out_2)
  );
  C53 c53_611 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_611_io_in_0),
    .io_in_1(c53_611_io_in_1),
    .io_in_2(c53_611_io_in_2),
    .io_in_3(c53_611_io_in_3),
    .io_in_4(c53_611_io_in_4),
    .io_out_0(c53_611_io_out_0),
    .io_out_1(c53_611_io_out_1),
    .io_out_2(c53_611_io_out_2)
  );
  C53 c53_612 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_612_io_in_0),
    .io_in_1(c53_612_io_in_1),
    .io_in_2(c53_612_io_in_2),
    .io_in_3(c53_612_io_in_3),
    .io_in_4(c53_612_io_in_4),
    .io_out_0(c53_612_io_out_0),
    .io_out_1(c53_612_io_out_1),
    .io_out_2(c53_612_io_out_2)
  );
  C53 c53_613 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_613_io_in_0),
    .io_in_1(c53_613_io_in_1),
    .io_in_2(c53_613_io_in_2),
    .io_in_3(c53_613_io_in_3),
    .io_in_4(c53_613_io_in_4),
    .io_out_0(c53_613_io_out_0),
    .io_out_1(c53_613_io_out_1),
    .io_out_2(c53_613_io_out_2)
  );
  C53 c53_614 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_614_io_in_0),
    .io_in_1(c53_614_io_in_1),
    .io_in_2(c53_614_io_in_2),
    .io_in_3(c53_614_io_in_3),
    .io_in_4(c53_614_io_in_4),
    .io_out_0(c53_614_io_out_0),
    .io_out_1(c53_614_io_out_1),
    .io_out_2(c53_614_io_out_2)
  );
  C53 c53_615 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_615_io_in_0),
    .io_in_1(c53_615_io_in_1),
    .io_in_2(c53_615_io_in_2),
    .io_in_3(c53_615_io_in_3),
    .io_in_4(c53_615_io_in_4),
    .io_out_0(c53_615_io_out_0),
    .io_out_1(c53_615_io_out_1),
    .io_out_2(c53_615_io_out_2)
  );
  C53 c53_616 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_616_io_in_0),
    .io_in_1(c53_616_io_in_1),
    .io_in_2(c53_616_io_in_2),
    .io_in_3(c53_616_io_in_3),
    .io_in_4(c53_616_io_in_4),
    .io_out_0(c53_616_io_out_0),
    .io_out_1(c53_616_io_out_1),
    .io_out_2(c53_616_io_out_2)
  );
  C22 c22_109 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_109_io_in_0),
    .io_in_1(c22_109_io_in_1),
    .io_out_0(c22_109_io_out_0),
    .io_out_1(c22_109_io_out_1)
  );
  C22 c22_110 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_110_io_in_0),
    .io_in_1(c22_110_io_in_1),
    .io_out_0(c22_110_io_out_0),
    .io_out_1(c22_110_io_out_1)
  );
  C32 c32_57 ( // @[Multiplier.scala 78:25]
    .io_in_0(c32_57_io_in_0),
    .io_in_1(c32_57_io_in_1),
    .io_in_2(c32_57_io_in_2),
    .io_out_0(c32_57_io_out_0),
    .io_out_1(c32_57_io_out_1)
  );
  C22 c22_111 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_111_io_in_0),
    .io_in_1(c22_111_io_in_1),
    .io_out_0(c22_111_io_out_0),
    .io_out_1(c22_111_io_out_1)
  );
  C22 c22_112 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_112_io_in_0),
    .io_in_1(c22_112_io_in_1),
    .io_out_0(c22_112_io_out_0),
    .io_out_1(c22_112_io_out_1)
  );
  C22 c22_113 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_113_io_in_0),
    .io_in_1(c22_113_io_in_1),
    .io_out_0(c22_113_io_out_0),
    .io_out_1(c22_113_io_out_1)
  );
  C22 c22_114 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_114_io_in_0),
    .io_in_1(c22_114_io_in_1),
    .io_out_0(c22_114_io_out_0),
    .io_out_1(c22_114_io_out_1)
  );
  C32 c32_58 ( // @[Multiplier.scala 78:25]
    .io_in_0(c32_58_io_in_0),
    .io_in_1(c32_58_io_in_1),
    .io_in_2(c32_58_io_in_2),
    .io_out_0(c32_58_io_out_0),
    .io_out_1(c32_58_io_out_1)
  );
  C22 c22_115 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_115_io_in_0),
    .io_in_1(c22_115_io_in_1),
    .io_out_0(c22_115_io_out_0),
    .io_out_1(c22_115_io_out_1)
  );
  C22 c22_116 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_116_io_in_0),
    .io_in_1(c22_116_io_in_1),
    .io_out_0(c22_116_io_out_0),
    .io_out_1(c22_116_io_out_1)
  );
  C22 c22_117 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_117_io_in_0),
    .io_in_1(c22_117_io_in_1),
    .io_out_0(c22_117_io_out_0),
    .io_out_1(c22_117_io_out_1)
  );
  C22 c22_118 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_118_io_in_0),
    .io_in_1(c22_118_io_in_1),
    .io_out_0(c22_118_io_out_0),
    .io_out_1(c22_118_io_out_1)
  );
  C22 c22_119 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_119_io_in_0),
    .io_in_1(c22_119_io_in_1),
    .io_out_0(c22_119_io_out_0),
    .io_out_1(c22_119_io_out_1)
  );
  C22 c22_120 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_120_io_in_0),
    .io_in_1(c22_120_io_in_1),
    .io_out_0(c22_120_io_out_0),
    .io_out_1(c22_120_io_out_1)
  );
  C22 c22_121 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_121_io_in_0),
    .io_in_1(c22_121_io_in_1),
    .io_out_0(c22_121_io_out_0),
    .io_out_1(c22_121_io_out_1)
  );
  C22 c22_122 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_122_io_in_0),
    .io_in_1(c22_122_io_in_1),
    .io_out_0(c22_122_io_out_0),
    .io_out_1(c22_122_io_out_1)
  );
  C22 c22_123 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_123_io_in_0),
    .io_in_1(c22_123_io_in_1),
    .io_out_0(c22_123_io_out_0),
    .io_out_1(c22_123_io_out_1)
  );
  C22 c22_124 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_124_io_in_0),
    .io_in_1(c22_124_io_in_1),
    .io_out_0(c22_124_io_out_0),
    .io_out_1(c22_124_io_out_1)
  );
  C22 c22_125 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_125_io_in_0),
    .io_in_1(c22_125_io_in_1),
    .io_out_0(c22_125_io_out_0),
    .io_out_1(c22_125_io_out_1)
  );
  C22 c22_126 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_126_io_in_0),
    .io_in_1(c22_126_io_in_1),
    .io_out_0(c22_126_io_out_0),
    .io_out_1(c22_126_io_out_1)
  );
  C22 c22_127 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_127_io_in_0),
    .io_in_1(c22_127_io_in_1),
    .io_out_0(c22_127_io_out_0),
    .io_out_1(c22_127_io_out_1)
  );
  C22 c22_128 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_128_io_in_0),
    .io_in_1(c22_128_io_in_1),
    .io_out_0(c22_128_io_out_0),
    .io_out_1(c22_128_io_out_1)
  );
  C22 c22_129 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_129_io_in_0),
    .io_in_1(c22_129_io_in_1),
    .io_out_0(c22_129_io_out_0),
    .io_out_1(c22_129_io_out_1)
  );
  C22 c22_130 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_130_io_in_0),
    .io_in_1(c22_130_io_in_1),
    .io_out_0(c22_130_io_out_0),
    .io_out_1(c22_130_io_out_1)
  );
  C22 c22_131 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_131_io_in_0),
    .io_in_1(c22_131_io_in_1),
    .io_out_0(c22_131_io_out_0),
    .io_out_1(c22_131_io_out_1)
  );
  C22 c22_132 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_132_io_in_0),
    .io_in_1(c22_132_io_in_1),
    .io_out_0(c22_132_io_out_0),
    .io_out_1(c22_132_io_out_1)
  );
  C22 c22_133 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_133_io_in_0),
    .io_in_1(c22_133_io_in_1),
    .io_out_0(c22_133_io_out_0),
    .io_out_1(c22_133_io_out_1)
  );
  C22 c22_134 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_134_io_in_0),
    .io_in_1(c22_134_io_in_1),
    .io_out_0(c22_134_io_out_0),
    .io_out_1(c22_134_io_out_1)
  );
  C22 c22_135 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_135_io_in_0),
    .io_in_1(c22_135_io_in_1),
    .io_out_0(c22_135_io_out_0),
    .io_out_1(c22_135_io_out_1)
  );
  C22 c22_136 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_136_io_in_0),
    .io_in_1(c22_136_io_in_1),
    .io_out_0(c22_136_io_out_0),
    .io_out_1(c22_136_io_out_1)
  );
  C22 c22_137 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_137_io_in_0),
    .io_in_1(c22_137_io_in_1),
    .io_out_0(c22_137_io_out_0),
    .io_out_1(c22_137_io_out_1)
  );
  C22 c22_138 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_138_io_in_0),
    .io_in_1(c22_138_io_in_1),
    .io_out_0(c22_138_io_out_0),
    .io_out_1(c22_138_io_out_1)
  );
  C22 c22_139 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_139_io_in_0),
    .io_in_1(c22_139_io_in_1),
    .io_out_0(c22_139_io_out_0),
    .io_out_1(c22_139_io_out_1)
  );
  C22 c22_140 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_140_io_in_0),
    .io_in_1(c22_140_io_in_1),
    .io_out_0(c22_140_io_out_0),
    .io_out_1(c22_140_io_out_1)
  );
  C22 c22_141 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_141_io_in_0),
    .io_in_1(c22_141_io_in_1),
    .io_out_0(c22_141_io_out_0),
    .io_out_1(c22_141_io_out_1)
  );
  C22 c22_142 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_142_io_in_0),
    .io_in_1(c22_142_io_in_1),
    .io_out_0(c22_142_io_out_0),
    .io_out_1(c22_142_io_out_1)
  );
  C22 c22_143 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_143_io_in_0),
    .io_in_1(c22_143_io_in_1),
    .io_out_0(c22_143_io_out_0),
    .io_out_1(c22_143_io_out_1)
  );
  C22 c22_144 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_144_io_in_0),
    .io_in_1(c22_144_io_in_1),
    .io_out_0(c22_144_io_out_0),
    .io_out_1(c22_144_io_out_1)
  );
  C22 c22_145 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_145_io_in_0),
    .io_in_1(c22_145_io_in_1),
    .io_out_0(c22_145_io_out_0),
    .io_out_1(c22_145_io_out_1)
  );
  C22 c22_146 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_146_io_in_0),
    .io_in_1(c22_146_io_in_1),
    .io_out_0(c22_146_io_out_0),
    .io_out_1(c22_146_io_out_1)
  );
  C22 c22_147 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_147_io_in_0),
    .io_in_1(c22_147_io_in_1),
    .io_out_0(c22_147_io_out_0),
    .io_out_1(c22_147_io_out_1)
  );
  C22 c22_148 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_148_io_in_0),
    .io_in_1(c22_148_io_in_1),
    .io_out_0(c22_148_io_out_0),
    .io_out_1(c22_148_io_out_1)
  );
  C32 c32_59 ( // @[Multiplier.scala 78:25]
    .io_in_0(c32_59_io_in_0),
    .io_in_1(c32_59_io_in_1),
    .io_in_2(c32_59_io_in_2),
    .io_out_0(c32_59_io_out_0),
    .io_out_1(c32_59_io_out_1)
  );
  C32 c32_60 ( // @[Multiplier.scala 78:25]
    .io_in_0(c32_60_io_in_0),
    .io_in_1(c32_60_io_in_1),
    .io_in_2(c32_60_io_in_2),
    .io_out_0(c32_60_io_out_0),
    .io_out_1(c32_60_io_out_1)
  );
  C32 c32_61 ( // @[Multiplier.scala 78:25]
    .io_in_0(c32_61_io_in_0),
    .io_in_1(c32_61_io_in_1),
    .io_in_2(c32_61_io_in_2),
    .io_out_0(c32_61_io_out_0),
    .io_out_1(c32_61_io_out_1)
  );
  C32 c32_62 ( // @[Multiplier.scala 78:25]
    .io_in_0(c32_62_io_in_0),
    .io_in_1(c32_62_io_in_1),
    .io_in_2(c32_62_io_in_2),
    .io_out_0(c32_62_io_out_0),
    .io_out_1(c32_62_io_out_1)
  );
  C32 c32_63 ( // @[Multiplier.scala 78:25]
    .io_in_0(c32_63_io_in_0),
    .io_in_1(c32_63_io_in_1),
    .io_in_2(c32_63_io_in_2),
    .io_out_0(c32_63_io_out_0),
    .io_out_1(c32_63_io_out_1)
  );
  C53 c53_617 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_617_io_in_0),
    .io_in_1(c53_617_io_in_1),
    .io_in_2(c53_617_io_in_2),
    .io_in_3(c53_617_io_in_3),
    .io_in_4(c53_617_io_in_4),
    .io_out_0(c53_617_io_out_0),
    .io_out_1(c53_617_io_out_1),
    .io_out_2(c53_617_io_out_2)
  );
  C53 c53_618 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_618_io_in_0),
    .io_in_1(c53_618_io_in_1),
    .io_in_2(c53_618_io_in_2),
    .io_in_3(c53_618_io_in_3),
    .io_in_4(c53_618_io_in_4),
    .io_out_0(c53_618_io_out_0),
    .io_out_1(c53_618_io_out_1),
    .io_out_2(c53_618_io_out_2)
  );
  C53 c53_619 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_619_io_in_0),
    .io_in_1(c53_619_io_in_1),
    .io_in_2(c53_619_io_in_2),
    .io_in_3(c53_619_io_in_3),
    .io_in_4(c53_619_io_in_4),
    .io_out_0(c53_619_io_out_0),
    .io_out_1(c53_619_io_out_1),
    .io_out_2(c53_619_io_out_2)
  );
  C53 c53_620 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_620_io_in_0),
    .io_in_1(c53_620_io_in_1),
    .io_in_2(c53_620_io_in_2),
    .io_in_3(c53_620_io_in_3),
    .io_in_4(c53_620_io_in_4),
    .io_out_0(c53_620_io_out_0),
    .io_out_1(c53_620_io_out_1),
    .io_out_2(c53_620_io_out_2)
  );
  C53 c53_621 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_621_io_in_0),
    .io_in_1(c53_621_io_in_1),
    .io_in_2(c53_621_io_in_2),
    .io_in_3(c53_621_io_in_3),
    .io_in_4(c53_621_io_in_4),
    .io_out_0(c53_621_io_out_0),
    .io_out_1(c53_621_io_out_1),
    .io_out_2(c53_621_io_out_2)
  );
  C53 c53_622 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_622_io_in_0),
    .io_in_1(c53_622_io_in_1),
    .io_in_2(c53_622_io_in_2),
    .io_in_3(c53_622_io_in_3),
    .io_in_4(c53_622_io_in_4),
    .io_out_0(c53_622_io_out_0),
    .io_out_1(c53_622_io_out_1),
    .io_out_2(c53_622_io_out_2)
  );
  C53 c53_623 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_623_io_in_0),
    .io_in_1(c53_623_io_in_1),
    .io_in_2(c53_623_io_in_2),
    .io_in_3(c53_623_io_in_3),
    .io_in_4(c53_623_io_in_4),
    .io_out_0(c53_623_io_out_0),
    .io_out_1(c53_623_io_out_1),
    .io_out_2(c53_623_io_out_2)
  );
  C53 c53_624 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_624_io_in_0),
    .io_in_1(c53_624_io_in_1),
    .io_in_2(c53_624_io_in_2),
    .io_in_3(c53_624_io_in_3),
    .io_in_4(c53_624_io_in_4),
    .io_out_0(c53_624_io_out_0),
    .io_out_1(c53_624_io_out_1),
    .io_out_2(c53_624_io_out_2)
  );
  C53 c53_625 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_625_io_in_0),
    .io_in_1(c53_625_io_in_1),
    .io_in_2(c53_625_io_in_2),
    .io_in_3(c53_625_io_in_3),
    .io_in_4(c53_625_io_in_4),
    .io_out_0(c53_625_io_out_0),
    .io_out_1(c53_625_io_out_1),
    .io_out_2(c53_625_io_out_2)
  );
  C53 c53_626 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_626_io_in_0),
    .io_in_1(c53_626_io_in_1),
    .io_in_2(c53_626_io_in_2),
    .io_in_3(c53_626_io_in_3),
    .io_in_4(c53_626_io_in_4),
    .io_out_0(c53_626_io_out_0),
    .io_out_1(c53_626_io_out_1),
    .io_out_2(c53_626_io_out_2)
  );
  C53 c53_627 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_627_io_in_0),
    .io_in_1(c53_627_io_in_1),
    .io_in_2(c53_627_io_in_2),
    .io_in_3(c53_627_io_in_3),
    .io_in_4(c53_627_io_in_4),
    .io_out_0(c53_627_io_out_0),
    .io_out_1(c53_627_io_out_1),
    .io_out_2(c53_627_io_out_2)
  );
  C53 c53_628 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_628_io_in_0),
    .io_in_1(c53_628_io_in_1),
    .io_in_2(c53_628_io_in_2),
    .io_in_3(c53_628_io_in_3),
    .io_in_4(c53_628_io_in_4),
    .io_out_0(c53_628_io_out_0),
    .io_out_1(c53_628_io_out_1),
    .io_out_2(c53_628_io_out_2)
  );
  C53 c53_629 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_629_io_in_0),
    .io_in_1(c53_629_io_in_1),
    .io_in_2(c53_629_io_in_2),
    .io_in_3(c53_629_io_in_3),
    .io_in_4(c53_629_io_in_4),
    .io_out_0(c53_629_io_out_0),
    .io_out_1(c53_629_io_out_1),
    .io_out_2(c53_629_io_out_2)
  );
  C53 c53_630 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_630_io_in_0),
    .io_in_1(c53_630_io_in_1),
    .io_in_2(c53_630_io_in_2),
    .io_in_3(c53_630_io_in_3),
    .io_in_4(c53_630_io_in_4),
    .io_out_0(c53_630_io_out_0),
    .io_out_1(c53_630_io_out_1),
    .io_out_2(c53_630_io_out_2)
  );
  C53 c53_631 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_631_io_in_0),
    .io_in_1(c53_631_io_in_1),
    .io_in_2(c53_631_io_in_2),
    .io_in_3(c53_631_io_in_3),
    .io_in_4(c53_631_io_in_4),
    .io_out_0(c53_631_io_out_0),
    .io_out_1(c53_631_io_out_1),
    .io_out_2(c53_631_io_out_2)
  );
  C53 c53_632 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_632_io_in_0),
    .io_in_1(c53_632_io_in_1),
    .io_in_2(c53_632_io_in_2),
    .io_in_3(c53_632_io_in_3),
    .io_in_4(c53_632_io_in_4),
    .io_out_0(c53_632_io_out_0),
    .io_out_1(c53_632_io_out_1),
    .io_out_2(c53_632_io_out_2)
  );
  C53 c53_633 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_633_io_in_0),
    .io_in_1(c53_633_io_in_1),
    .io_in_2(c53_633_io_in_2),
    .io_in_3(c53_633_io_in_3),
    .io_in_4(c53_633_io_in_4),
    .io_out_0(c53_633_io_out_0),
    .io_out_1(c53_633_io_out_1),
    .io_out_2(c53_633_io_out_2)
  );
  C53 c53_634 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_634_io_in_0),
    .io_in_1(c53_634_io_in_1),
    .io_in_2(c53_634_io_in_2),
    .io_in_3(c53_634_io_in_3),
    .io_in_4(c53_634_io_in_4),
    .io_out_0(c53_634_io_out_0),
    .io_out_1(c53_634_io_out_1),
    .io_out_2(c53_634_io_out_2)
  );
  C53 c53_635 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_635_io_in_0),
    .io_in_1(c53_635_io_in_1),
    .io_in_2(c53_635_io_in_2),
    .io_in_3(c53_635_io_in_3),
    .io_in_4(c53_635_io_in_4),
    .io_out_0(c53_635_io_out_0),
    .io_out_1(c53_635_io_out_1),
    .io_out_2(c53_635_io_out_2)
  );
  C53 c53_636 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_636_io_in_0),
    .io_in_1(c53_636_io_in_1),
    .io_in_2(c53_636_io_in_2),
    .io_in_3(c53_636_io_in_3),
    .io_in_4(c53_636_io_in_4),
    .io_out_0(c53_636_io_out_0),
    .io_out_1(c53_636_io_out_1),
    .io_out_2(c53_636_io_out_2)
  );
  C53 c53_637 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_637_io_in_0),
    .io_in_1(c53_637_io_in_1),
    .io_in_2(c53_637_io_in_2),
    .io_in_3(c53_637_io_in_3),
    .io_in_4(c53_637_io_in_4),
    .io_out_0(c53_637_io_out_0),
    .io_out_1(c53_637_io_out_1),
    .io_out_2(c53_637_io_out_2)
  );
  C53 c53_638 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_638_io_in_0),
    .io_in_1(c53_638_io_in_1),
    .io_in_2(c53_638_io_in_2),
    .io_in_3(c53_638_io_in_3),
    .io_in_4(c53_638_io_in_4),
    .io_out_0(c53_638_io_out_0),
    .io_out_1(c53_638_io_out_1),
    .io_out_2(c53_638_io_out_2)
  );
  C53 c53_639 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_639_io_in_0),
    .io_in_1(c53_639_io_in_1),
    .io_in_2(c53_639_io_in_2),
    .io_in_3(c53_639_io_in_3),
    .io_in_4(c53_639_io_in_4),
    .io_out_0(c53_639_io_out_0),
    .io_out_1(c53_639_io_out_1),
    .io_out_2(c53_639_io_out_2)
  );
  C53 c53_640 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_640_io_in_0),
    .io_in_1(c53_640_io_in_1),
    .io_in_2(c53_640_io_in_2),
    .io_in_3(c53_640_io_in_3),
    .io_in_4(c53_640_io_in_4),
    .io_out_0(c53_640_io_out_0),
    .io_out_1(c53_640_io_out_1),
    .io_out_2(c53_640_io_out_2)
  );
  C53 c53_641 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_641_io_in_0),
    .io_in_1(c53_641_io_in_1),
    .io_in_2(c53_641_io_in_2),
    .io_in_3(c53_641_io_in_3),
    .io_in_4(c53_641_io_in_4),
    .io_out_0(c53_641_io_out_0),
    .io_out_1(c53_641_io_out_1),
    .io_out_2(c53_641_io_out_2)
  );
  C53 c53_642 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_642_io_in_0),
    .io_in_1(c53_642_io_in_1),
    .io_in_2(c53_642_io_in_2),
    .io_in_3(c53_642_io_in_3),
    .io_in_4(c53_642_io_in_4),
    .io_out_0(c53_642_io_out_0),
    .io_out_1(c53_642_io_out_1),
    .io_out_2(c53_642_io_out_2)
  );
  C53 c53_643 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_643_io_in_0),
    .io_in_1(c53_643_io_in_1),
    .io_in_2(c53_643_io_in_2),
    .io_in_3(c53_643_io_in_3),
    .io_in_4(c53_643_io_in_4),
    .io_out_0(c53_643_io_out_0),
    .io_out_1(c53_643_io_out_1),
    .io_out_2(c53_643_io_out_2)
  );
  C53 c53_644 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_644_io_in_0),
    .io_in_1(c53_644_io_in_1),
    .io_in_2(c53_644_io_in_2),
    .io_in_3(c53_644_io_in_3),
    .io_in_4(c53_644_io_in_4),
    .io_out_0(c53_644_io_out_0),
    .io_out_1(c53_644_io_out_1),
    .io_out_2(c53_644_io_out_2)
  );
  C53 c53_645 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_645_io_in_0),
    .io_in_1(c53_645_io_in_1),
    .io_in_2(c53_645_io_in_2),
    .io_in_3(c53_645_io_in_3),
    .io_in_4(c53_645_io_in_4),
    .io_out_0(c53_645_io_out_0),
    .io_out_1(c53_645_io_out_1),
    .io_out_2(c53_645_io_out_2)
  );
  C53 c53_646 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_646_io_in_0),
    .io_in_1(c53_646_io_in_1),
    .io_in_2(c53_646_io_in_2),
    .io_in_3(c53_646_io_in_3),
    .io_in_4(c53_646_io_in_4),
    .io_out_0(c53_646_io_out_0),
    .io_out_1(c53_646_io_out_1),
    .io_out_2(c53_646_io_out_2)
  );
  C53 c53_647 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_647_io_in_0),
    .io_in_1(c53_647_io_in_1),
    .io_in_2(c53_647_io_in_2),
    .io_in_3(c53_647_io_in_3),
    .io_in_4(c53_647_io_in_4),
    .io_out_0(c53_647_io_out_0),
    .io_out_1(c53_647_io_out_1),
    .io_out_2(c53_647_io_out_2)
  );
  C53 c53_648 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_648_io_in_0),
    .io_in_1(c53_648_io_in_1),
    .io_in_2(c53_648_io_in_2),
    .io_in_3(c53_648_io_in_3),
    .io_in_4(c53_648_io_in_4),
    .io_out_0(c53_648_io_out_0),
    .io_out_1(c53_648_io_out_1),
    .io_out_2(c53_648_io_out_2)
  );
  C53 c53_649 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_649_io_in_0),
    .io_in_1(c53_649_io_in_1),
    .io_in_2(c53_649_io_in_2),
    .io_in_3(c53_649_io_in_3),
    .io_in_4(c53_649_io_in_4),
    .io_out_0(c53_649_io_out_0),
    .io_out_1(c53_649_io_out_1),
    .io_out_2(c53_649_io_out_2)
  );
  C53 c53_650 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_650_io_in_0),
    .io_in_1(c53_650_io_in_1),
    .io_in_2(c53_650_io_in_2),
    .io_in_3(c53_650_io_in_3),
    .io_in_4(c53_650_io_in_4),
    .io_out_0(c53_650_io_out_0),
    .io_out_1(c53_650_io_out_1),
    .io_out_2(c53_650_io_out_2)
  );
  C53 c53_651 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_651_io_in_0),
    .io_in_1(c53_651_io_in_1),
    .io_in_2(c53_651_io_in_2),
    .io_in_3(c53_651_io_in_3),
    .io_in_4(c53_651_io_in_4),
    .io_out_0(c53_651_io_out_0),
    .io_out_1(c53_651_io_out_1),
    .io_out_2(c53_651_io_out_2)
  );
  C53 c53_652 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_652_io_in_0),
    .io_in_1(c53_652_io_in_1),
    .io_in_2(c53_652_io_in_2),
    .io_in_3(c53_652_io_in_3),
    .io_in_4(c53_652_io_in_4),
    .io_out_0(c53_652_io_out_0),
    .io_out_1(c53_652_io_out_1),
    .io_out_2(c53_652_io_out_2)
  );
  C53 c53_653 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_653_io_in_0),
    .io_in_1(c53_653_io_in_1),
    .io_in_2(c53_653_io_in_2),
    .io_in_3(c53_653_io_in_3),
    .io_in_4(c53_653_io_in_4),
    .io_out_0(c53_653_io_out_0),
    .io_out_1(c53_653_io_out_1),
    .io_out_2(c53_653_io_out_2)
  );
  C53 c53_654 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_654_io_in_0),
    .io_in_1(c53_654_io_in_1),
    .io_in_2(c53_654_io_in_2),
    .io_in_3(c53_654_io_in_3),
    .io_in_4(c53_654_io_in_4),
    .io_out_0(c53_654_io_out_0),
    .io_out_1(c53_654_io_out_1),
    .io_out_2(c53_654_io_out_2)
  );
  C53 c53_655 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_655_io_in_0),
    .io_in_1(c53_655_io_in_1),
    .io_in_2(c53_655_io_in_2),
    .io_in_3(c53_655_io_in_3),
    .io_in_4(c53_655_io_in_4),
    .io_out_0(c53_655_io_out_0),
    .io_out_1(c53_655_io_out_1),
    .io_out_2(c53_655_io_out_2)
  );
  C53 c53_656 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_656_io_in_0),
    .io_in_1(c53_656_io_in_1),
    .io_in_2(c53_656_io_in_2),
    .io_in_3(c53_656_io_in_3),
    .io_in_4(c53_656_io_in_4),
    .io_out_0(c53_656_io_out_0),
    .io_out_1(c53_656_io_out_1),
    .io_out_2(c53_656_io_out_2)
  );
  C53 c53_657 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_657_io_in_0),
    .io_in_1(c53_657_io_in_1),
    .io_in_2(c53_657_io_in_2),
    .io_in_3(c53_657_io_in_3),
    .io_in_4(c53_657_io_in_4),
    .io_out_0(c53_657_io_out_0),
    .io_out_1(c53_657_io_out_1),
    .io_out_2(c53_657_io_out_2)
  );
  C53 c53_658 ( // @[Multiplier.scala 83:25]
    .io_in_0(c53_658_io_in_0),
    .io_in_1(c53_658_io_in_1),
    .io_in_2(c53_658_io_in_2),
    .io_in_3(c53_658_io_in_3),
    .io_in_4(c53_658_io_in_4),
    .io_out_0(c53_658_io_out_0),
    .io_out_1(c53_658_io_out_1),
    .io_out_2(c53_658_io_out_2)
  );
  C32 c32_64 ( // @[Multiplier.scala 78:25]
    .io_in_0(c32_64_io_in_0),
    .io_in_1(c32_64_io_in_1),
    .io_in_2(c32_64_io_in_2),
    .io_out_0(c32_64_io_out_0),
    .io_out_1(c32_64_io_out_1)
  );
  C22 c22_149 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_149_io_in_0),
    .io_in_1(c22_149_io_in_1),
    .io_out_0(c22_149_io_out_0),
    .io_out_1(c22_149_io_out_1)
  );
  C32 c32_65 ( // @[Multiplier.scala 78:25]
    .io_in_0(c32_65_io_in_0),
    .io_in_1(c32_65_io_in_1),
    .io_in_2(c32_65_io_in_2),
    .io_out_0(c32_65_io_out_0),
    .io_out_1(c32_65_io_out_1)
  );
  C22 c22_150 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_150_io_in_0),
    .io_in_1(c22_150_io_in_1),
    .io_out_0(c22_150_io_out_0),
    .io_out_1(c22_150_io_out_1)
  );
  C22 c22_151 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_151_io_in_0),
    .io_in_1(c22_151_io_in_1),
    .io_out_0(c22_151_io_out_0),
    .io_out_1(c22_151_io_out_1)
  );
  C22 c22_152 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_152_io_in_0),
    .io_in_1(c22_152_io_in_1),
    .io_out_0(c22_152_io_out_0),
    .io_out_1(c22_152_io_out_1)
  );
  C22 c22_153 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_153_io_in_0),
    .io_in_1(c22_153_io_in_1),
    .io_out_0(c22_153_io_out_0),
    .io_out_1(c22_153_io_out_1)
  );
  C32 c32_66 ( // @[Multiplier.scala 78:25]
    .io_in_0(c32_66_io_in_0),
    .io_in_1(c32_66_io_in_1),
    .io_in_2(c32_66_io_in_2),
    .io_out_0(c32_66_io_out_0),
    .io_out_1(c32_66_io_out_1)
  );
  C22 c22_154 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_154_io_in_0),
    .io_in_1(c22_154_io_in_1),
    .io_out_0(c22_154_io_out_0),
    .io_out_1(c22_154_io_out_1)
  );
  C22 c22_155 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_155_io_in_0),
    .io_in_1(c22_155_io_in_1),
    .io_out_0(c22_155_io_out_0),
    .io_out_1(c22_155_io_out_1)
  );
  C22 c22_156 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_156_io_in_0),
    .io_in_1(c22_156_io_in_1),
    .io_out_0(c22_156_io_out_0),
    .io_out_1(c22_156_io_out_1)
  );
  C22 c22_157 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_157_io_in_0),
    .io_in_1(c22_157_io_in_1),
    .io_out_0(c22_157_io_out_0),
    .io_out_1(c22_157_io_out_1)
  );
  C22 c22_158 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_158_io_in_0),
    .io_in_1(c22_158_io_in_1),
    .io_out_0(c22_158_io_out_0),
    .io_out_1(c22_158_io_out_1)
  );
  C22 c22_159 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_159_io_in_0),
    .io_in_1(c22_159_io_in_1),
    .io_out_0(c22_159_io_out_0),
    .io_out_1(c22_159_io_out_1)
  );
  C22 c22_160 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_160_io_in_0),
    .io_in_1(c22_160_io_in_1),
    .io_out_0(c22_160_io_out_0),
    .io_out_1(c22_160_io_out_1)
  );
  C22 c22_161 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_161_io_in_0),
    .io_in_1(c22_161_io_in_1),
    .io_out_0(c22_161_io_out_0),
    .io_out_1(c22_161_io_out_1)
  );
  C32 c32_67 ( // @[Multiplier.scala 78:25]
    .io_in_0(c32_67_io_in_0),
    .io_in_1(c32_67_io_in_1),
    .io_in_2(c32_67_io_in_2),
    .io_out_0(c32_67_io_out_0),
    .io_out_1(c32_67_io_out_1)
  );
  C22 c22_162 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_162_io_in_0),
    .io_in_1(c22_162_io_in_1),
    .io_out_0(c22_162_io_out_0),
    .io_out_1(c22_162_io_out_1)
  );
  C22 c22_163 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_163_io_in_0),
    .io_in_1(c22_163_io_in_1),
    .io_out_0(c22_163_io_out_0),
    .io_out_1(c22_163_io_out_1)
  );
  C22 c22_164 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_164_io_in_0),
    .io_in_1(c22_164_io_in_1),
    .io_out_0(c22_164_io_out_0),
    .io_out_1(c22_164_io_out_1)
  );
  C22 c22_165 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_165_io_in_0),
    .io_in_1(c22_165_io_in_1),
    .io_out_0(c22_165_io_out_0),
    .io_out_1(c22_165_io_out_1)
  );
  C22 c22_166 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_166_io_in_0),
    .io_in_1(c22_166_io_in_1),
    .io_out_0(c22_166_io_out_0),
    .io_out_1(c22_166_io_out_1)
  );
  C22 c22_167 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_167_io_in_0),
    .io_in_1(c22_167_io_in_1),
    .io_out_0(c22_167_io_out_0),
    .io_out_1(c22_167_io_out_1)
  );
  C22 c22_168 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_168_io_in_0),
    .io_in_1(c22_168_io_in_1),
    .io_out_0(c22_168_io_out_0),
    .io_out_1(c22_168_io_out_1)
  );
  C22 c22_169 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_169_io_in_0),
    .io_in_1(c22_169_io_in_1),
    .io_out_0(c22_169_io_out_0),
    .io_out_1(c22_169_io_out_1)
  );
  C22 c22_170 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_170_io_in_0),
    .io_in_1(c22_170_io_in_1),
    .io_out_0(c22_170_io_out_0),
    .io_out_1(c22_170_io_out_1)
  );
  C22 c22_171 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_171_io_in_0),
    .io_in_1(c22_171_io_in_1),
    .io_out_0(c22_171_io_out_0),
    .io_out_1(c22_171_io_out_1)
  );
  C22 c22_172 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_172_io_in_0),
    .io_in_1(c22_172_io_in_1),
    .io_out_0(c22_172_io_out_0),
    .io_out_1(c22_172_io_out_1)
  );
  C22 c22_173 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_173_io_in_0),
    .io_in_1(c22_173_io_in_1),
    .io_out_0(c22_173_io_out_0),
    .io_out_1(c22_173_io_out_1)
  );
  C22 c22_174 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_174_io_in_0),
    .io_in_1(c22_174_io_in_1),
    .io_out_0(c22_174_io_out_0),
    .io_out_1(c22_174_io_out_1)
  );
  C22 c22_175 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_175_io_in_0),
    .io_in_1(c22_175_io_in_1),
    .io_out_0(c22_175_io_out_0),
    .io_out_1(c22_175_io_out_1)
  );
  C22 c22_176 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_176_io_in_0),
    .io_in_1(c22_176_io_in_1),
    .io_out_0(c22_176_io_out_0),
    .io_out_1(c22_176_io_out_1)
  );
  C22 c22_177 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_177_io_in_0),
    .io_in_1(c22_177_io_in_1),
    .io_out_0(c22_177_io_out_0),
    .io_out_1(c22_177_io_out_1)
  );
  C22 c22_178 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_178_io_in_0),
    .io_in_1(c22_178_io_in_1),
    .io_out_0(c22_178_io_out_0),
    .io_out_1(c22_178_io_out_1)
  );
  C22 c22_179 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_179_io_in_0),
    .io_in_1(c22_179_io_in_1),
    .io_out_0(c22_179_io_out_0),
    .io_out_1(c22_179_io_out_1)
  );
  C22 c22_180 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_180_io_in_0),
    .io_in_1(c22_180_io_in_1),
    .io_out_0(c22_180_io_out_0),
    .io_out_1(c22_180_io_out_1)
  );
  C22 c22_181 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_181_io_in_0),
    .io_in_1(c22_181_io_in_1),
    .io_out_0(c22_181_io_out_0),
    .io_out_1(c22_181_io_out_1)
  );
  C22 c22_182 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_182_io_in_0),
    .io_in_1(c22_182_io_in_1),
    .io_out_0(c22_182_io_out_0),
    .io_out_1(c22_182_io_out_1)
  );
  C22 c22_183 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_183_io_in_0),
    .io_in_1(c22_183_io_in_1),
    .io_out_0(c22_183_io_out_0),
    .io_out_1(c22_183_io_out_1)
  );
  C22 c22_184 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_184_io_in_0),
    .io_in_1(c22_184_io_in_1),
    .io_out_0(c22_184_io_out_0),
    .io_out_1(c22_184_io_out_1)
  );
  C22 c22_185 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_185_io_in_0),
    .io_in_1(c22_185_io_in_1),
    .io_out_0(c22_185_io_out_0),
    .io_out_1(c22_185_io_out_1)
  );
  C22 c22_186 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_186_io_in_0),
    .io_in_1(c22_186_io_in_1),
    .io_out_0(c22_186_io_out_0),
    .io_out_1(c22_186_io_out_1)
  );
  C22 c22_187 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_187_io_in_0),
    .io_in_1(c22_187_io_in_1),
    .io_out_0(c22_187_io_out_0),
    .io_out_1(c22_187_io_out_1)
  );
  C22 c22_188 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_188_io_in_0),
    .io_in_1(c22_188_io_in_1),
    .io_out_0(c22_188_io_out_0),
    .io_out_1(c22_188_io_out_1)
  );
  C22 c22_189 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_189_io_in_0),
    .io_in_1(c22_189_io_in_1),
    .io_out_0(c22_189_io_out_0),
    .io_out_1(c22_189_io_out_1)
  );
  C22 c22_190 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_190_io_in_0),
    .io_in_1(c22_190_io_in_1),
    .io_out_0(c22_190_io_out_0),
    .io_out_1(c22_190_io_out_1)
  );
  C22 c22_191 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_191_io_in_0),
    .io_in_1(c22_191_io_in_1),
    .io_out_0(c22_191_io_out_0),
    .io_out_1(c22_191_io_out_1)
  );
  C22 c22_192 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_192_io_in_0),
    .io_in_1(c22_192_io_in_1),
    .io_out_0(c22_192_io_out_0),
    .io_out_1(c22_192_io_out_1)
  );
  C22 c22_193 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_193_io_in_0),
    .io_in_1(c22_193_io_in_1),
    .io_out_0(c22_193_io_out_0),
    .io_out_1(c22_193_io_out_1)
  );
  C22 c22_194 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_194_io_in_0),
    .io_in_1(c22_194_io_in_1),
    .io_out_0(c22_194_io_out_0),
    .io_out_1(c22_194_io_out_1)
  );
  C22 c22_195 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_195_io_in_0),
    .io_in_1(c22_195_io_in_1),
    .io_out_0(c22_195_io_out_0),
    .io_out_1(c22_195_io_out_1)
  );
  C22 c22_196 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_196_io_in_0),
    .io_in_1(c22_196_io_in_1),
    .io_out_0(c22_196_io_out_0),
    .io_out_1(c22_196_io_out_1)
  );
  C22 c22_197 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_197_io_in_0),
    .io_in_1(c22_197_io_in_1),
    .io_out_0(c22_197_io_out_0),
    .io_out_1(c22_197_io_out_1)
  );
  C22 c22_198 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_198_io_in_0),
    .io_in_1(c22_198_io_in_1),
    .io_out_0(c22_198_io_out_0),
    .io_out_1(c22_198_io_out_1)
  );
  C22 c22_199 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_199_io_in_0),
    .io_in_1(c22_199_io_in_1),
    .io_out_0(c22_199_io_out_0),
    .io_out_1(c22_199_io_out_1)
  );
  C22 c22_200 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_200_io_in_0),
    .io_in_1(c22_200_io_in_1),
    .io_out_0(c22_200_io_out_0),
    .io_out_1(c22_200_io_out_1)
  );
  C22 c22_201 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_201_io_in_0),
    .io_in_1(c22_201_io_in_1),
    .io_out_0(c22_201_io_out_0),
    .io_out_1(c22_201_io_out_1)
  );
  C22 c22_202 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_202_io_in_0),
    .io_in_1(c22_202_io_in_1),
    .io_out_0(c22_202_io_out_0),
    .io_out_1(c22_202_io_out_1)
  );
  C22 c22_203 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_203_io_in_0),
    .io_in_1(c22_203_io_in_1),
    .io_out_0(c22_203_io_out_0),
    .io_out_1(c22_203_io_out_1)
  );
  C22 c22_204 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_204_io_in_0),
    .io_in_1(c22_204_io_in_1),
    .io_out_0(c22_204_io_out_0),
    .io_out_1(c22_204_io_out_1)
  );
  C22 c22_205 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_205_io_in_0),
    .io_in_1(c22_205_io_in_1),
    .io_out_0(c22_205_io_out_0),
    .io_out_1(c22_205_io_out_1)
  );
  C22 c22_206 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_206_io_in_0),
    .io_in_1(c22_206_io_in_1),
    .io_out_0(c22_206_io_out_0),
    .io_out_1(c22_206_io_out_1)
  );
  C22 c22_207 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_207_io_in_0),
    .io_in_1(c22_207_io_in_1),
    .io_out_0(c22_207_io_out_0),
    .io_out_1(c22_207_io_out_1)
  );
  C22 c22_208 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_208_io_in_0),
    .io_in_1(c22_208_io_in_1),
    .io_out_0(c22_208_io_out_0),
    .io_out_1(c22_208_io_out_1)
  );
  C22 c22_209 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_209_io_in_0),
    .io_in_1(c22_209_io_in_1),
    .io_out_0(c22_209_io_out_0),
    .io_out_1(c22_209_io_out_1)
  );
  C22 c22_210 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_210_io_in_0),
    .io_in_1(c22_210_io_in_1),
    .io_out_0(c22_210_io_out_0),
    .io_out_1(c22_210_io_out_1)
  );
  C22 c22_211 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_211_io_in_0),
    .io_in_1(c22_211_io_in_1),
    .io_out_0(c22_211_io_out_0),
    .io_out_1(c22_211_io_out_1)
  );
  C22 c22_212 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_212_io_in_0),
    .io_in_1(c22_212_io_in_1),
    .io_out_0(c22_212_io_out_0),
    .io_out_1(c22_212_io_out_1)
  );
  C22 c22_213 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_213_io_in_0),
    .io_in_1(c22_213_io_in_1),
    .io_out_0(c22_213_io_out_0),
    .io_out_1(c22_213_io_out_1)
  );
  C22 c22_214 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_214_io_in_0),
    .io_in_1(c22_214_io_in_1),
    .io_out_0(c22_214_io_out_0),
    .io_out_1(c22_214_io_out_1)
  );
  C22 c22_215 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_215_io_in_0),
    .io_in_1(c22_215_io_in_1),
    .io_out_0(c22_215_io_out_0),
    .io_out_1(c22_215_io_out_1)
  );
  C22 c22_216 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_216_io_in_0),
    .io_in_1(c22_216_io_in_1),
    .io_out_0(c22_216_io_out_0),
    .io_out_1(c22_216_io_out_1)
  );
  C22 c22_217 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_217_io_in_0),
    .io_in_1(c22_217_io_in_1),
    .io_out_0(c22_217_io_out_0),
    .io_out_1(c22_217_io_out_1)
  );
  C22 c22_218 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_218_io_in_0),
    .io_in_1(c22_218_io_in_1),
    .io_out_0(c22_218_io_out_0),
    .io_out_1(c22_218_io_out_1)
  );
  C22 c22_219 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_219_io_in_0),
    .io_in_1(c22_219_io_in_1),
    .io_out_0(c22_219_io_out_0),
    .io_out_1(c22_219_io_out_1)
  );
  C22 c22_220 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_220_io_in_0),
    .io_in_1(c22_220_io_in_1),
    .io_out_0(c22_220_io_out_0),
    .io_out_1(c22_220_io_out_1)
  );
  C22 c22_221 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_221_io_in_0),
    .io_in_1(c22_221_io_in_1),
    .io_out_0(c22_221_io_out_0),
    .io_out_1(c22_221_io_out_1)
  );
  C22 c22_222 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_222_io_in_0),
    .io_in_1(c22_222_io_in_1),
    .io_out_0(c22_222_io_out_0),
    .io_out_1(c22_222_io_out_1)
  );
  C22 c22_223 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_223_io_in_0),
    .io_in_1(c22_223_io_in_1),
    .io_out_0(c22_223_io_out_0),
    .io_out_1(c22_223_io_out_1)
  );
  C22 c22_224 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_224_io_in_0),
    .io_in_1(c22_224_io_in_1),
    .io_out_0(c22_224_io_out_0),
    .io_out_1(c22_224_io_out_1)
  );
  C22 c22_225 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_225_io_in_0),
    .io_in_1(c22_225_io_in_1),
    .io_out_0(c22_225_io_out_0),
    .io_out_1(c22_225_io_out_1)
  );
  C22 c22_226 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_226_io_in_0),
    .io_in_1(c22_226_io_in_1),
    .io_out_0(c22_226_io_out_0),
    .io_out_1(c22_226_io_out_1)
  );
  C22 c22_227 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_227_io_in_0),
    .io_in_1(c22_227_io_in_1),
    .io_out_0(c22_227_io_out_0),
    .io_out_1(c22_227_io_out_1)
  );
  C22 c22_228 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_228_io_in_0),
    .io_in_1(c22_228_io_in_1),
    .io_out_0(c22_228_io_out_0),
    .io_out_1(c22_228_io_out_1)
  );
  C22 c22_229 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_229_io_in_0),
    .io_in_1(c22_229_io_in_1),
    .io_out_0(c22_229_io_out_0),
    .io_out_1(c22_229_io_out_1)
  );
  C22 c22_230 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_230_io_in_0),
    .io_in_1(c22_230_io_in_1),
    .io_out_0(c22_230_io_out_0),
    .io_out_1(c22_230_io_out_1)
  );
  C22 c22_231 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_231_io_in_0),
    .io_in_1(c22_231_io_in_1),
    .io_out_0(c22_231_io_out_0),
    .io_out_1(c22_231_io_out_1)
  );
  C22 c22_232 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_232_io_in_0),
    .io_in_1(c22_232_io_in_1),
    .io_out_0(c22_232_io_out_0),
    .io_out_1(c22_232_io_out_1)
  );
  C32 c32_68 ( // @[Multiplier.scala 78:25]
    .io_in_0(c32_68_io_in_0),
    .io_in_1(c32_68_io_in_1),
    .io_in_2(c32_68_io_in_2),
    .io_out_0(c32_68_io_out_0),
    .io_out_1(c32_68_io_out_1)
  );
  C22 c22_233 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_233_io_in_0),
    .io_in_1(c22_233_io_in_1),
    .io_out_0(c22_233_io_out_0),
    .io_out_1(c22_233_io_out_1)
  );
  C22 c22_234 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_234_io_in_0),
    .io_in_1(c22_234_io_in_1),
    .io_out_0(c22_234_io_out_0),
    .io_out_1(c22_234_io_out_1)
  );
  C22 c22_235 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_235_io_in_0),
    .io_in_1(c22_235_io_in_1),
    .io_out_0(c22_235_io_out_0),
    .io_out_1(c22_235_io_out_1)
  );
  C22 c22_236 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_236_io_in_0),
    .io_in_1(c22_236_io_in_1),
    .io_out_0(c22_236_io_out_0),
    .io_out_1(c22_236_io_out_1)
  );
  C22 c22_237 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_237_io_in_0),
    .io_in_1(c22_237_io_in_1),
    .io_out_0(c22_237_io_out_0),
    .io_out_1(c22_237_io_out_1)
  );
  C22 c22_238 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_238_io_in_0),
    .io_in_1(c22_238_io_in_1),
    .io_out_0(c22_238_io_out_0),
    .io_out_1(c22_238_io_out_1)
  );
  C22 c22_239 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_239_io_in_0),
    .io_in_1(c22_239_io_in_1),
    .io_out_0(c22_239_io_out_0),
    .io_out_1(c22_239_io_out_1)
  );
  C22 c22_240 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_240_io_in_0),
    .io_in_1(c22_240_io_in_1),
    .io_out_0(c22_240_io_out_0),
    .io_out_1(c22_240_io_out_1)
  );
  C22 c22_241 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_241_io_in_0),
    .io_in_1(c22_241_io_in_1),
    .io_out_0(c22_241_io_out_0),
    .io_out_1(c22_241_io_out_1)
  );
  C22 c22_242 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_242_io_in_0),
    .io_in_1(c22_242_io_in_1),
    .io_out_0(c22_242_io_out_0),
    .io_out_1(c22_242_io_out_1)
  );
  C22 c22_243 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_243_io_in_0),
    .io_in_1(c22_243_io_in_1),
    .io_out_0(c22_243_io_out_0),
    .io_out_1(c22_243_io_out_1)
  );
  C22 c22_244 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_244_io_in_0),
    .io_in_1(c22_244_io_in_1),
    .io_out_0(c22_244_io_out_0),
    .io_out_1(c22_244_io_out_1)
  );
  C22 c22_245 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_245_io_in_0),
    .io_in_1(c22_245_io_in_1),
    .io_out_0(c22_245_io_out_0),
    .io_out_1(c22_245_io_out_1)
  );
  C22 c22_246 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_246_io_in_0),
    .io_in_1(c22_246_io_in_1),
    .io_out_0(c22_246_io_out_0),
    .io_out_1(c22_246_io_out_1)
  );
  C22 c22_247 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_247_io_in_0),
    .io_in_1(c22_247_io_in_1),
    .io_out_0(c22_247_io_out_0),
    .io_out_1(c22_247_io_out_1)
  );
  C32 c32_69 ( // @[Multiplier.scala 78:25]
    .io_in_0(c32_69_io_in_0),
    .io_in_1(c32_69_io_in_1),
    .io_in_2(c32_69_io_in_2),
    .io_out_0(c32_69_io_out_0),
    .io_out_1(c32_69_io_out_1)
  );
  C22 c22_248 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_248_io_in_0),
    .io_in_1(c22_248_io_in_1),
    .io_out_0(c22_248_io_out_0),
    .io_out_1(c22_248_io_out_1)
  );
  C22 c22_249 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_249_io_in_0),
    .io_in_1(c22_249_io_in_1),
    .io_out_0(c22_249_io_out_0),
    .io_out_1(c22_249_io_out_1)
  );
  C22 c22_250 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_250_io_in_0),
    .io_in_1(c22_250_io_in_1),
    .io_out_0(c22_250_io_out_0),
    .io_out_1(c22_250_io_out_1)
  );
  C22 c22_251 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_251_io_in_0),
    .io_in_1(c22_251_io_in_1),
    .io_out_0(c22_251_io_out_0),
    .io_out_1(c22_251_io_out_1)
  );
  C22 c22_252 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_252_io_in_0),
    .io_in_1(c22_252_io_in_1),
    .io_out_0(c22_252_io_out_0),
    .io_out_1(c22_252_io_out_1)
  );
  C22 c22_253 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_253_io_in_0),
    .io_in_1(c22_253_io_in_1),
    .io_out_0(c22_253_io_out_0),
    .io_out_1(c22_253_io_out_1)
  );
  C22 c22_254 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_254_io_in_0),
    .io_in_1(c22_254_io_in_1),
    .io_out_0(c22_254_io_out_0),
    .io_out_1(c22_254_io_out_1)
  );
  C22 c22_255 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_255_io_in_0),
    .io_in_1(c22_255_io_in_1),
    .io_out_0(c22_255_io_out_0),
    .io_out_1(c22_255_io_out_1)
  );
  C22 c22_256 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_256_io_in_0),
    .io_in_1(c22_256_io_in_1),
    .io_out_0(c22_256_io_out_0),
    .io_out_1(c22_256_io_out_1)
  );
  C22 c22_257 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_257_io_in_0),
    .io_in_1(c22_257_io_in_1),
    .io_out_0(c22_257_io_out_0),
    .io_out_1(c22_257_io_out_1)
  );
  C22 c22_258 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_258_io_in_0),
    .io_in_1(c22_258_io_in_1),
    .io_out_0(c22_258_io_out_0),
    .io_out_1(c22_258_io_out_1)
  );
  C22 c22_259 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_259_io_in_0),
    .io_in_1(c22_259_io_in_1),
    .io_out_0(c22_259_io_out_0),
    .io_out_1(c22_259_io_out_1)
  );
  C22 c22_260 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_260_io_in_0),
    .io_in_1(c22_260_io_in_1),
    .io_out_0(c22_260_io_out_0),
    .io_out_1(c22_260_io_out_1)
  );
  C22 c22_261 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_261_io_in_0),
    .io_in_1(c22_261_io_in_1),
    .io_out_0(c22_261_io_out_0),
    .io_out_1(c22_261_io_out_1)
  );
  C22 c22_262 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_262_io_in_0),
    .io_in_1(c22_262_io_in_1),
    .io_out_0(c22_262_io_out_0),
    .io_out_1(c22_262_io_out_1)
  );
  C22 c22_263 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_263_io_in_0),
    .io_in_1(c22_263_io_in_1),
    .io_out_0(c22_263_io_out_0),
    .io_out_1(c22_263_io_out_1)
  );
  C22 c22_264 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_264_io_in_0),
    .io_in_1(c22_264_io_in_1),
    .io_out_0(c22_264_io_out_0),
    .io_out_1(c22_264_io_out_1)
  );
  C22 c22_265 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_265_io_in_0),
    .io_in_1(c22_265_io_in_1),
    .io_out_0(c22_265_io_out_0),
    .io_out_1(c22_265_io_out_1)
  );
  C22 c22_266 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_266_io_in_0),
    .io_in_1(c22_266_io_in_1),
    .io_out_0(c22_266_io_out_0),
    .io_out_1(c22_266_io_out_1)
  );
  C22 c22_267 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_267_io_in_0),
    .io_in_1(c22_267_io_in_1),
    .io_out_0(c22_267_io_out_0),
    .io_out_1(c22_267_io_out_1)
  );
  C22 c22_268 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_268_io_in_0),
    .io_in_1(c22_268_io_in_1),
    .io_out_0(c22_268_io_out_0),
    .io_out_1(c22_268_io_out_1)
  );
  C22 c22_269 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_269_io_in_0),
    .io_in_1(c22_269_io_in_1),
    .io_out_0(c22_269_io_out_0),
    .io_out_1(c22_269_io_out_1)
  );
  C22 c22_270 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_270_io_in_0),
    .io_in_1(c22_270_io_in_1),
    .io_out_0(c22_270_io_out_0),
    .io_out_1(c22_270_io_out_1)
  );
  C22 c22_271 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_271_io_in_0),
    .io_in_1(c22_271_io_in_1),
    .io_out_0(c22_271_io_out_0),
    .io_out_1(c22_271_io_out_1)
  );
  C22 c22_272 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_272_io_in_0),
    .io_in_1(c22_272_io_in_1),
    .io_out_0(c22_272_io_out_0),
    .io_out_1(c22_272_io_out_1)
  );
  C22 c22_273 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_273_io_in_0),
    .io_in_1(c22_273_io_in_1),
    .io_out_0(c22_273_io_out_0),
    .io_out_1(c22_273_io_out_1)
  );
  C22 c22_274 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_274_io_in_0),
    .io_in_1(c22_274_io_in_1),
    .io_out_0(c22_274_io_out_0),
    .io_out_1(c22_274_io_out_1)
  );
  C22 c22_275 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_275_io_in_0),
    .io_in_1(c22_275_io_in_1),
    .io_out_0(c22_275_io_out_0),
    .io_out_1(c22_275_io_out_1)
  );
  C22 c22_276 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_276_io_in_0),
    .io_in_1(c22_276_io_in_1),
    .io_out_0(c22_276_io_out_0),
    .io_out_1(c22_276_io_out_1)
  );
  C22 c22_277 ( // @[Multiplier.scala 73:25]
    .io_in_0(c22_277_io_in_0),
    .io_in_1(c22_277_io_in_1),
    .io_out_0(c22_277_io_out_0),
    .io_out_1(c22_277_io_out_1)
  );
  assign io_result = sum + carry_1; // @[Multiplier.scala 135:20]
  assign c22_io_in_0 = pp[0]; // @[Multiplier.scala 60:38]
  assign c22_io_in_1 = pp_1[0]; // @[Multiplier.scala 60:38]
  assign c22_1_io_in_0 = pp[1]; // @[Multiplier.scala 60:38]
  assign c22_1_io_in_1 = pp_1[1]; // @[Multiplier.scala 60:38]
  assign c32_io_in_0 = pp[2]; // @[Multiplier.scala 60:38]
  assign c32_io_in_1 = pp_1[2]; // @[Multiplier.scala 60:38]
  assign c32_io_in_2 = pp_2[0]; // @[Multiplier.scala 60:38]
  assign c32_1_io_in_0 = pp[3]; // @[Multiplier.scala 60:38]
  assign c32_1_io_in_1 = pp_1[3]; // @[Multiplier.scala 60:38]
  assign c32_1_io_in_2 = pp_2[1]; // @[Multiplier.scala 60:38]
  assign c53_io_in_0 = pp[4]; // @[Multiplier.scala 60:38]
  assign c53_io_in_1 = pp_1[4]; // @[Multiplier.scala 60:38]
  assign c53_io_in_2 = pp_2[2]; // @[Multiplier.scala 60:38]
  assign c53_io_in_3 = pp_3[0]; // @[Multiplier.scala 60:38]
  assign c53_io_in_4 = 1'h0; // @[Multiplier.scala 87:24]
  assign c53_1_io_in_0 = pp[5]; // @[Multiplier.scala 60:38]
  assign c53_1_io_in_1 = pp_1[5]; // @[Multiplier.scala 60:38]
  assign c53_1_io_in_2 = pp_2[3]; // @[Multiplier.scala 60:38]
  assign c53_1_io_in_3 = pp_3[1]; // @[Multiplier.scala 60:38]
  assign c53_1_io_in_4 = c53_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_2_io_in_0 = pp[6]; // @[Multiplier.scala 60:38]
  assign c53_2_io_in_1 = pp_1[6]; // @[Multiplier.scala 60:38]
  assign c53_2_io_in_2 = pp_2[4]; // @[Multiplier.scala 60:38]
  assign c53_2_io_in_3 = pp_3[2]; // @[Multiplier.scala 60:38]
  assign c53_2_io_in_4 = c53_1_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_3_io_in_0 = pp[7]; // @[Multiplier.scala 60:38]
  assign c53_3_io_in_1 = pp_1[7]; // @[Multiplier.scala 60:38]
  assign c53_3_io_in_2 = pp_2[5]; // @[Multiplier.scala 60:38]
  assign c53_3_io_in_3 = pp_3[3]; // @[Multiplier.scala 60:38]
  assign c53_3_io_in_4 = c53_2_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_4_io_in_0 = pp[8]; // @[Multiplier.scala 60:38]
  assign c53_4_io_in_1 = pp_1[8]; // @[Multiplier.scala 60:38]
  assign c53_4_io_in_2 = pp_2[6]; // @[Multiplier.scala 60:38]
  assign c53_4_io_in_3 = pp_3[4]; // @[Multiplier.scala 60:38]
  assign c53_4_io_in_4 = c53_3_io_out_1; // @[Multiplier.scala 89:41]
  assign c22_2_io_in_0 = pp_4[2]; // @[Multiplier.scala 60:38]
  assign c22_2_io_in_1 = pp_5[0]; // @[Multiplier.scala 60:38]
  assign c53_5_io_in_0 = pp[9]; // @[Multiplier.scala 60:38]
  assign c53_5_io_in_1 = pp_1[9]; // @[Multiplier.scala 60:38]
  assign c53_5_io_in_2 = pp_2[7]; // @[Multiplier.scala 60:38]
  assign c53_5_io_in_3 = pp_3[5]; // @[Multiplier.scala 60:38]
  assign c53_5_io_in_4 = c53_4_io_out_1; // @[Multiplier.scala 89:41]
  assign c22_3_io_in_0 = pp_4[3]; // @[Multiplier.scala 60:38]
  assign c22_3_io_in_1 = pp_5[1]; // @[Multiplier.scala 60:38]
  assign c53_6_io_in_0 = pp[10]; // @[Multiplier.scala 60:38]
  assign c53_6_io_in_1 = pp_1[10]; // @[Multiplier.scala 60:38]
  assign c53_6_io_in_2 = pp_2[8]; // @[Multiplier.scala 60:38]
  assign c53_6_io_in_3 = pp_3[6]; // @[Multiplier.scala 60:38]
  assign c53_6_io_in_4 = c53_5_io_out_1; // @[Multiplier.scala 89:41]
  assign c32_2_io_in_0 = pp_4[4]; // @[Multiplier.scala 60:38]
  assign c32_2_io_in_1 = pp_5[2]; // @[Multiplier.scala 60:38]
  assign c32_2_io_in_2 = pp_6[0]; // @[Multiplier.scala 60:38]
  assign c53_7_io_in_0 = pp[11]; // @[Multiplier.scala 60:38]
  assign c53_7_io_in_1 = pp_1[11]; // @[Multiplier.scala 60:38]
  assign c53_7_io_in_2 = pp_2[9]; // @[Multiplier.scala 60:38]
  assign c53_7_io_in_3 = pp_3[7]; // @[Multiplier.scala 60:38]
  assign c53_7_io_in_4 = c53_6_io_out_1; // @[Multiplier.scala 89:41]
  assign c32_3_io_in_0 = pp_4[5]; // @[Multiplier.scala 60:38]
  assign c32_3_io_in_1 = pp_5[3]; // @[Multiplier.scala 60:38]
  assign c32_3_io_in_2 = pp_6[1]; // @[Multiplier.scala 60:38]
  assign c53_8_io_in_0 = pp[12]; // @[Multiplier.scala 60:38]
  assign c53_8_io_in_1 = pp_1[12]; // @[Multiplier.scala 60:38]
  assign c53_8_io_in_2 = pp_2[10]; // @[Multiplier.scala 60:38]
  assign c53_8_io_in_3 = pp_3[8]; // @[Multiplier.scala 60:38]
  assign c53_8_io_in_4 = c53_7_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_9_io_in_0 = pp_4[6]; // @[Multiplier.scala 60:38]
  assign c53_9_io_in_1 = pp_5[4]; // @[Multiplier.scala 60:38]
  assign c53_9_io_in_2 = pp_6[2]; // @[Multiplier.scala 60:38]
  assign c53_9_io_in_3 = pp_7[0]; // @[Multiplier.scala 60:38]
  assign c53_9_io_in_4 = 1'h0; // @[Multiplier.scala 87:24]
  assign c53_10_io_in_0 = pp[13]; // @[Multiplier.scala 60:38]
  assign c53_10_io_in_1 = pp_1[13]; // @[Multiplier.scala 60:38]
  assign c53_10_io_in_2 = pp_2[11]; // @[Multiplier.scala 60:38]
  assign c53_10_io_in_3 = pp_3[9]; // @[Multiplier.scala 60:38]
  assign c53_10_io_in_4 = c53_8_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_11_io_in_0 = pp_4[7]; // @[Multiplier.scala 60:38]
  assign c53_11_io_in_1 = pp_5[5]; // @[Multiplier.scala 60:38]
  assign c53_11_io_in_2 = pp_6[3]; // @[Multiplier.scala 60:38]
  assign c53_11_io_in_3 = pp_7[1]; // @[Multiplier.scala 60:38]
  assign c53_11_io_in_4 = c53_9_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_12_io_in_0 = pp[14]; // @[Multiplier.scala 60:38]
  assign c53_12_io_in_1 = pp_1[14]; // @[Multiplier.scala 60:38]
  assign c53_12_io_in_2 = pp_2[12]; // @[Multiplier.scala 60:38]
  assign c53_12_io_in_3 = pp_3[10]; // @[Multiplier.scala 60:38]
  assign c53_12_io_in_4 = c53_10_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_13_io_in_0 = pp_4[8]; // @[Multiplier.scala 60:38]
  assign c53_13_io_in_1 = pp_5[6]; // @[Multiplier.scala 60:38]
  assign c53_13_io_in_2 = pp_6[4]; // @[Multiplier.scala 60:38]
  assign c53_13_io_in_3 = pp_7[2]; // @[Multiplier.scala 60:38]
  assign c53_13_io_in_4 = c53_11_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_14_io_in_0 = pp[15]; // @[Multiplier.scala 60:38]
  assign c53_14_io_in_1 = pp_1[15]; // @[Multiplier.scala 60:38]
  assign c53_14_io_in_2 = pp_2[13]; // @[Multiplier.scala 60:38]
  assign c53_14_io_in_3 = pp_3[11]; // @[Multiplier.scala 60:38]
  assign c53_14_io_in_4 = c53_12_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_15_io_in_0 = pp_4[9]; // @[Multiplier.scala 60:38]
  assign c53_15_io_in_1 = pp_5[7]; // @[Multiplier.scala 60:38]
  assign c53_15_io_in_2 = pp_6[5]; // @[Multiplier.scala 60:38]
  assign c53_15_io_in_3 = pp_7[3]; // @[Multiplier.scala 60:38]
  assign c53_15_io_in_4 = c53_13_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_16_io_in_0 = pp[16]; // @[Multiplier.scala 60:38]
  assign c53_16_io_in_1 = pp_1[16]; // @[Multiplier.scala 60:38]
  assign c53_16_io_in_2 = pp_2[14]; // @[Multiplier.scala 60:38]
  assign c53_16_io_in_3 = pp_3[12]; // @[Multiplier.scala 60:38]
  assign c53_16_io_in_4 = c53_14_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_17_io_in_0 = pp_4[10]; // @[Multiplier.scala 60:38]
  assign c53_17_io_in_1 = pp_5[8]; // @[Multiplier.scala 60:38]
  assign c53_17_io_in_2 = pp_6[6]; // @[Multiplier.scala 60:38]
  assign c53_17_io_in_3 = pp_7[4]; // @[Multiplier.scala 60:38]
  assign c53_17_io_in_4 = c53_15_io_out_1; // @[Multiplier.scala 89:41]
  assign c22_4_io_in_0 = pp_8[2]; // @[Multiplier.scala 60:38]
  assign c22_4_io_in_1 = pp_9[0]; // @[Multiplier.scala 60:38]
  assign c53_18_io_in_0 = pp[17]; // @[Multiplier.scala 60:38]
  assign c53_18_io_in_1 = pp_1[17]; // @[Multiplier.scala 60:38]
  assign c53_18_io_in_2 = pp_2[15]; // @[Multiplier.scala 60:38]
  assign c53_18_io_in_3 = pp_3[13]; // @[Multiplier.scala 60:38]
  assign c53_18_io_in_4 = c53_16_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_19_io_in_0 = pp_4[11]; // @[Multiplier.scala 60:38]
  assign c53_19_io_in_1 = pp_5[9]; // @[Multiplier.scala 60:38]
  assign c53_19_io_in_2 = pp_6[7]; // @[Multiplier.scala 60:38]
  assign c53_19_io_in_3 = pp_7[5]; // @[Multiplier.scala 60:38]
  assign c53_19_io_in_4 = c53_17_io_out_1; // @[Multiplier.scala 89:41]
  assign c22_5_io_in_0 = pp_8[3]; // @[Multiplier.scala 60:38]
  assign c22_5_io_in_1 = pp_9[1]; // @[Multiplier.scala 60:38]
  assign c53_20_io_in_0 = pp[18]; // @[Multiplier.scala 60:38]
  assign c53_20_io_in_1 = pp_1[18]; // @[Multiplier.scala 60:38]
  assign c53_20_io_in_2 = pp_2[16]; // @[Multiplier.scala 60:38]
  assign c53_20_io_in_3 = pp_3[14]; // @[Multiplier.scala 60:38]
  assign c53_20_io_in_4 = c53_18_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_21_io_in_0 = pp_4[12]; // @[Multiplier.scala 60:38]
  assign c53_21_io_in_1 = pp_5[10]; // @[Multiplier.scala 60:38]
  assign c53_21_io_in_2 = pp_6[8]; // @[Multiplier.scala 60:38]
  assign c53_21_io_in_3 = pp_7[6]; // @[Multiplier.scala 60:38]
  assign c53_21_io_in_4 = c53_19_io_out_1; // @[Multiplier.scala 89:41]
  assign c32_4_io_in_0 = pp_8[4]; // @[Multiplier.scala 60:38]
  assign c32_4_io_in_1 = pp_9[2]; // @[Multiplier.scala 60:38]
  assign c32_4_io_in_2 = pp_10[0]; // @[Multiplier.scala 60:38]
  assign c53_22_io_in_0 = pp[19]; // @[Multiplier.scala 60:38]
  assign c53_22_io_in_1 = pp_1[19]; // @[Multiplier.scala 60:38]
  assign c53_22_io_in_2 = pp_2[17]; // @[Multiplier.scala 60:38]
  assign c53_22_io_in_3 = pp_3[15]; // @[Multiplier.scala 60:38]
  assign c53_22_io_in_4 = c53_20_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_23_io_in_0 = pp_4[13]; // @[Multiplier.scala 60:38]
  assign c53_23_io_in_1 = pp_5[11]; // @[Multiplier.scala 60:38]
  assign c53_23_io_in_2 = pp_6[9]; // @[Multiplier.scala 60:38]
  assign c53_23_io_in_3 = pp_7[7]; // @[Multiplier.scala 60:38]
  assign c53_23_io_in_4 = c53_21_io_out_1; // @[Multiplier.scala 89:41]
  assign c32_5_io_in_0 = pp_8[5]; // @[Multiplier.scala 60:38]
  assign c32_5_io_in_1 = pp_9[3]; // @[Multiplier.scala 60:38]
  assign c32_5_io_in_2 = pp_10[1]; // @[Multiplier.scala 60:38]
  assign c53_24_io_in_0 = pp[20]; // @[Multiplier.scala 60:38]
  assign c53_24_io_in_1 = pp_1[20]; // @[Multiplier.scala 60:38]
  assign c53_24_io_in_2 = pp_2[18]; // @[Multiplier.scala 60:38]
  assign c53_24_io_in_3 = pp_3[16]; // @[Multiplier.scala 60:38]
  assign c53_24_io_in_4 = c53_22_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_25_io_in_0 = pp_4[14]; // @[Multiplier.scala 60:38]
  assign c53_25_io_in_1 = pp_5[12]; // @[Multiplier.scala 60:38]
  assign c53_25_io_in_2 = pp_6[10]; // @[Multiplier.scala 60:38]
  assign c53_25_io_in_3 = pp_7[8]; // @[Multiplier.scala 60:38]
  assign c53_25_io_in_4 = c53_23_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_26_io_in_0 = pp_8[6]; // @[Multiplier.scala 60:38]
  assign c53_26_io_in_1 = pp_9[4]; // @[Multiplier.scala 60:38]
  assign c53_26_io_in_2 = pp_10[2]; // @[Multiplier.scala 60:38]
  assign c53_26_io_in_3 = pp_11[0]; // @[Multiplier.scala 60:38]
  assign c53_26_io_in_4 = 1'h0; // @[Multiplier.scala 87:24]
  assign c53_27_io_in_0 = pp[21]; // @[Multiplier.scala 60:38]
  assign c53_27_io_in_1 = pp_1[21]; // @[Multiplier.scala 60:38]
  assign c53_27_io_in_2 = pp_2[19]; // @[Multiplier.scala 60:38]
  assign c53_27_io_in_3 = pp_3[17]; // @[Multiplier.scala 60:38]
  assign c53_27_io_in_4 = c53_24_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_28_io_in_0 = pp_4[15]; // @[Multiplier.scala 60:38]
  assign c53_28_io_in_1 = pp_5[13]; // @[Multiplier.scala 60:38]
  assign c53_28_io_in_2 = pp_6[11]; // @[Multiplier.scala 60:38]
  assign c53_28_io_in_3 = pp_7[9]; // @[Multiplier.scala 60:38]
  assign c53_28_io_in_4 = c53_25_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_29_io_in_0 = pp_8[7]; // @[Multiplier.scala 60:38]
  assign c53_29_io_in_1 = pp_9[5]; // @[Multiplier.scala 60:38]
  assign c53_29_io_in_2 = pp_10[3]; // @[Multiplier.scala 60:38]
  assign c53_29_io_in_3 = pp_11[1]; // @[Multiplier.scala 60:38]
  assign c53_29_io_in_4 = c53_26_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_30_io_in_0 = pp[22]; // @[Multiplier.scala 60:38]
  assign c53_30_io_in_1 = pp_1[22]; // @[Multiplier.scala 60:38]
  assign c53_30_io_in_2 = pp_2[20]; // @[Multiplier.scala 60:38]
  assign c53_30_io_in_3 = pp_3[18]; // @[Multiplier.scala 60:38]
  assign c53_30_io_in_4 = c53_27_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_31_io_in_0 = pp_4[16]; // @[Multiplier.scala 60:38]
  assign c53_31_io_in_1 = pp_5[14]; // @[Multiplier.scala 60:38]
  assign c53_31_io_in_2 = pp_6[12]; // @[Multiplier.scala 60:38]
  assign c53_31_io_in_3 = pp_7[10]; // @[Multiplier.scala 60:38]
  assign c53_31_io_in_4 = c53_28_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_32_io_in_0 = pp_8[8]; // @[Multiplier.scala 60:38]
  assign c53_32_io_in_1 = pp_9[6]; // @[Multiplier.scala 60:38]
  assign c53_32_io_in_2 = pp_10[4]; // @[Multiplier.scala 60:38]
  assign c53_32_io_in_3 = pp_11[2]; // @[Multiplier.scala 60:38]
  assign c53_32_io_in_4 = c53_29_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_33_io_in_0 = pp[23]; // @[Multiplier.scala 60:38]
  assign c53_33_io_in_1 = pp_1[23]; // @[Multiplier.scala 60:38]
  assign c53_33_io_in_2 = pp_2[21]; // @[Multiplier.scala 60:38]
  assign c53_33_io_in_3 = pp_3[19]; // @[Multiplier.scala 60:38]
  assign c53_33_io_in_4 = c53_30_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_34_io_in_0 = pp_4[17]; // @[Multiplier.scala 60:38]
  assign c53_34_io_in_1 = pp_5[15]; // @[Multiplier.scala 60:38]
  assign c53_34_io_in_2 = pp_6[13]; // @[Multiplier.scala 60:38]
  assign c53_34_io_in_3 = pp_7[11]; // @[Multiplier.scala 60:38]
  assign c53_34_io_in_4 = c53_31_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_35_io_in_0 = pp_8[9]; // @[Multiplier.scala 60:38]
  assign c53_35_io_in_1 = pp_9[7]; // @[Multiplier.scala 60:38]
  assign c53_35_io_in_2 = pp_10[5]; // @[Multiplier.scala 60:38]
  assign c53_35_io_in_3 = pp_11[3]; // @[Multiplier.scala 60:38]
  assign c53_35_io_in_4 = c53_32_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_36_io_in_0 = pp[24]; // @[Multiplier.scala 60:38]
  assign c53_36_io_in_1 = pp_1[24]; // @[Multiplier.scala 60:38]
  assign c53_36_io_in_2 = pp_2[22]; // @[Multiplier.scala 60:38]
  assign c53_36_io_in_3 = pp_3[20]; // @[Multiplier.scala 60:38]
  assign c53_36_io_in_4 = c53_33_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_37_io_in_0 = pp_4[18]; // @[Multiplier.scala 60:38]
  assign c53_37_io_in_1 = pp_5[16]; // @[Multiplier.scala 60:38]
  assign c53_37_io_in_2 = pp_6[14]; // @[Multiplier.scala 60:38]
  assign c53_37_io_in_3 = pp_7[12]; // @[Multiplier.scala 60:38]
  assign c53_37_io_in_4 = c53_34_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_38_io_in_0 = pp_8[10]; // @[Multiplier.scala 60:38]
  assign c53_38_io_in_1 = pp_9[8]; // @[Multiplier.scala 60:38]
  assign c53_38_io_in_2 = pp_10[6]; // @[Multiplier.scala 60:38]
  assign c53_38_io_in_3 = pp_11[4]; // @[Multiplier.scala 60:38]
  assign c53_38_io_in_4 = c53_35_io_out_1; // @[Multiplier.scala 89:41]
  assign c22_6_io_in_0 = pp_12[2]; // @[Multiplier.scala 60:38]
  assign c22_6_io_in_1 = pp_13[0]; // @[Multiplier.scala 60:38]
  assign c53_39_io_in_0 = pp[25]; // @[Multiplier.scala 60:38]
  assign c53_39_io_in_1 = pp_1[25]; // @[Multiplier.scala 60:38]
  assign c53_39_io_in_2 = pp_2[23]; // @[Multiplier.scala 60:38]
  assign c53_39_io_in_3 = pp_3[21]; // @[Multiplier.scala 60:38]
  assign c53_39_io_in_4 = c53_36_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_40_io_in_0 = pp_4[19]; // @[Multiplier.scala 60:38]
  assign c53_40_io_in_1 = pp_5[17]; // @[Multiplier.scala 60:38]
  assign c53_40_io_in_2 = pp_6[15]; // @[Multiplier.scala 60:38]
  assign c53_40_io_in_3 = pp_7[13]; // @[Multiplier.scala 60:38]
  assign c53_40_io_in_4 = c53_37_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_41_io_in_0 = pp_8[11]; // @[Multiplier.scala 60:38]
  assign c53_41_io_in_1 = pp_9[9]; // @[Multiplier.scala 60:38]
  assign c53_41_io_in_2 = pp_10[7]; // @[Multiplier.scala 60:38]
  assign c53_41_io_in_3 = pp_11[5]; // @[Multiplier.scala 60:38]
  assign c53_41_io_in_4 = c53_38_io_out_1; // @[Multiplier.scala 89:41]
  assign c22_7_io_in_0 = pp_12[3]; // @[Multiplier.scala 60:38]
  assign c22_7_io_in_1 = pp_13[1]; // @[Multiplier.scala 60:38]
  assign c53_42_io_in_0 = pp[26]; // @[Multiplier.scala 60:38]
  assign c53_42_io_in_1 = pp_1[26]; // @[Multiplier.scala 60:38]
  assign c53_42_io_in_2 = pp_2[24]; // @[Multiplier.scala 60:38]
  assign c53_42_io_in_3 = pp_3[22]; // @[Multiplier.scala 60:38]
  assign c53_42_io_in_4 = c53_39_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_43_io_in_0 = pp_4[20]; // @[Multiplier.scala 60:38]
  assign c53_43_io_in_1 = pp_5[18]; // @[Multiplier.scala 60:38]
  assign c53_43_io_in_2 = pp_6[16]; // @[Multiplier.scala 60:38]
  assign c53_43_io_in_3 = pp_7[14]; // @[Multiplier.scala 60:38]
  assign c53_43_io_in_4 = c53_40_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_44_io_in_0 = pp_8[12]; // @[Multiplier.scala 60:38]
  assign c53_44_io_in_1 = pp_9[10]; // @[Multiplier.scala 60:38]
  assign c53_44_io_in_2 = pp_10[8]; // @[Multiplier.scala 60:38]
  assign c53_44_io_in_3 = pp_11[6]; // @[Multiplier.scala 60:38]
  assign c53_44_io_in_4 = c53_41_io_out_1; // @[Multiplier.scala 89:41]
  assign c32_6_io_in_0 = pp_12[4]; // @[Multiplier.scala 60:38]
  assign c32_6_io_in_1 = pp_13[2]; // @[Multiplier.scala 60:38]
  assign c32_6_io_in_2 = pp_14[0]; // @[Multiplier.scala 60:38]
  assign c53_45_io_in_0 = pp[27]; // @[Multiplier.scala 60:38]
  assign c53_45_io_in_1 = pp_1[27]; // @[Multiplier.scala 60:38]
  assign c53_45_io_in_2 = pp_2[25]; // @[Multiplier.scala 60:38]
  assign c53_45_io_in_3 = pp_3[23]; // @[Multiplier.scala 60:38]
  assign c53_45_io_in_4 = c53_42_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_46_io_in_0 = pp_4[21]; // @[Multiplier.scala 60:38]
  assign c53_46_io_in_1 = pp_5[19]; // @[Multiplier.scala 60:38]
  assign c53_46_io_in_2 = pp_6[17]; // @[Multiplier.scala 60:38]
  assign c53_46_io_in_3 = pp_7[15]; // @[Multiplier.scala 60:38]
  assign c53_46_io_in_4 = c53_43_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_47_io_in_0 = pp_8[13]; // @[Multiplier.scala 60:38]
  assign c53_47_io_in_1 = pp_9[11]; // @[Multiplier.scala 60:38]
  assign c53_47_io_in_2 = pp_10[9]; // @[Multiplier.scala 60:38]
  assign c53_47_io_in_3 = pp_11[7]; // @[Multiplier.scala 60:38]
  assign c53_47_io_in_4 = c53_44_io_out_1; // @[Multiplier.scala 89:41]
  assign c32_7_io_in_0 = pp_12[5]; // @[Multiplier.scala 60:38]
  assign c32_7_io_in_1 = pp_13[3]; // @[Multiplier.scala 60:38]
  assign c32_7_io_in_2 = pp_14[1]; // @[Multiplier.scala 60:38]
  assign c53_48_io_in_0 = pp[28]; // @[Multiplier.scala 60:38]
  assign c53_48_io_in_1 = pp_1[28]; // @[Multiplier.scala 60:38]
  assign c53_48_io_in_2 = pp_2[26]; // @[Multiplier.scala 60:38]
  assign c53_48_io_in_3 = pp_3[24]; // @[Multiplier.scala 60:38]
  assign c53_48_io_in_4 = c53_45_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_49_io_in_0 = pp_4[22]; // @[Multiplier.scala 60:38]
  assign c53_49_io_in_1 = pp_5[20]; // @[Multiplier.scala 60:38]
  assign c53_49_io_in_2 = pp_6[18]; // @[Multiplier.scala 60:38]
  assign c53_49_io_in_3 = pp_7[16]; // @[Multiplier.scala 60:38]
  assign c53_49_io_in_4 = c53_46_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_50_io_in_0 = pp_8[14]; // @[Multiplier.scala 60:38]
  assign c53_50_io_in_1 = pp_9[12]; // @[Multiplier.scala 60:38]
  assign c53_50_io_in_2 = pp_10[10]; // @[Multiplier.scala 60:38]
  assign c53_50_io_in_3 = pp_11[8]; // @[Multiplier.scala 60:38]
  assign c53_50_io_in_4 = c53_47_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_51_io_in_0 = pp_12[6]; // @[Multiplier.scala 60:38]
  assign c53_51_io_in_1 = pp_13[4]; // @[Multiplier.scala 60:38]
  assign c53_51_io_in_2 = pp_14[2]; // @[Multiplier.scala 60:38]
  assign c53_51_io_in_3 = pp_15[0]; // @[Multiplier.scala 60:38]
  assign c53_51_io_in_4 = 1'h0; // @[Multiplier.scala 87:24]
  assign c53_52_io_in_0 = pp[29]; // @[Multiplier.scala 60:38]
  assign c53_52_io_in_1 = pp_1[29]; // @[Multiplier.scala 60:38]
  assign c53_52_io_in_2 = pp_2[27]; // @[Multiplier.scala 60:38]
  assign c53_52_io_in_3 = pp_3[25]; // @[Multiplier.scala 60:38]
  assign c53_52_io_in_4 = c53_48_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_53_io_in_0 = pp_4[23]; // @[Multiplier.scala 60:38]
  assign c53_53_io_in_1 = pp_5[21]; // @[Multiplier.scala 60:38]
  assign c53_53_io_in_2 = pp_6[19]; // @[Multiplier.scala 60:38]
  assign c53_53_io_in_3 = pp_7[17]; // @[Multiplier.scala 60:38]
  assign c53_53_io_in_4 = c53_49_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_54_io_in_0 = pp_8[15]; // @[Multiplier.scala 60:38]
  assign c53_54_io_in_1 = pp_9[13]; // @[Multiplier.scala 60:38]
  assign c53_54_io_in_2 = pp_10[11]; // @[Multiplier.scala 60:38]
  assign c53_54_io_in_3 = pp_11[9]; // @[Multiplier.scala 60:38]
  assign c53_54_io_in_4 = c53_50_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_55_io_in_0 = pp_12[7]; // @[Multiplier.scala 60:38]
  assign c53_55_io_in_1 = pp_13[5]; // @[Multiplier.scala 60:38]
  assign c53_55_io_in_2 = pp_14[3]; // @[Multiplier.scala 60:38]
  assign c53_55_io_in_3 = pp_15[1]; // @[Multiplier.scala 60:38]
  assign c53_55_io_in_4 = c53_51_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_56_io_in_0 = pp[30]; // @[Multiplier.scala 60:38]
  assign c53_56_io_in_1 = pp_1[30]; // @[Multiplier.scala 60:38]
  assign c53_56_io_in_2 = pp_2[28]; // @[Multiplier.scala 60:38]
  assign c53_56_io_in_3 = pp_3[26]; // @[Multiplier.scala 60:38]
  assign c53_56_io_in_4 = c53_52_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_57_io_in_0 = pp_4[24]; // @[Multiplier.scala 60:38]
  assign c53_57_io_in_1 = pp_5[22]; // @[Multiplier.scala 60:38]
  assign c53_57_io_in_2 = pp_6[20]; // @[Multiplier.scala 60:38]
  assign c53_57_io_in_3 = pp_7[18]; // @[Multiplier.scala 60:38]
  assign c53_57_io_in_4 = c53_53_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_58_io_in_0 = pp_8[16]; // @[Multiplier.scala 60:38]
  assign c53_58_io_in_1 = pp_9[14]; // @[Multiplier.scala 60:38]
  assign c53_58_io_in_2 = pp_10[12]; // @[Multiplier.scala 60:38]
  assign c53_58_io_in_3 = pp_11[10]; // @[Multiplier.scala 60:38]
  assign c53_58_io_in_4 = c53_54_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_59_io_in_0 = pp_12[8]; // @[Multiplier.scala 60:38]
  assign c53_59_io_in_1 = pp_13[6]; // @[Multiplier.scala 60:38]
  assign c53_59_io_in_2 = pp_14[4]; // @[Multiplier.scala 60:38]
  assign c53_59_io_in_3 = pp_15[2]; // @[Multiplier.scala 60:38]
  assign c53_59_io_in_4 = c53_55_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_60_io_in_0 = pp[31]; // @[Multiplier.scala 60:38]
  assign c53_60_io_in_1 = pp_1[31]; // @[Multiplier.scala 60:38]
  assign c53_60_io_in_2 = pp_2[29]; // @[Multiplier.scala 60:38]
  assign c53_60_io_in_3 = pp_3[27]; // @[Multiplier.scala 60:38]
  assign c53_60_io_in_4 = c53_56_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_61_io_in_0 = pp_4[25]; // @[Multiplier.scala 60:38]
  assign c53_61_io_in_1 = pp_5[23]; // @[Multiplier.scala 60:38]
  assign c53_61_io_in_2 = pp_6[21]; // @[Multiplier.scala 60:38]
  assign c53_61_io_in_3 = pp_7[19]; // @[Multiplier.scala 60:38]
  assign c53_61_io_in_4 = c53_57_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_62_io_in_0 = pp_8[17]; // @[Multiplier.scala 60:38]
  assign c53_62_io_in_1 = pp_9[15]; // @[Multiplier.scala 60:38]
  assign c53_62_io_in_2 = pp_10[13]; // @[Multiplier.scala 60:38]
  assign c53_62_io_in_3 = pp_11[11]; // @[Multiplier.scala 60:38]
  assign c53_62_io_in_4 = c53_58_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_63_io_in_0 = pp_12[9]; // @[Multiplier.scala 60:38]
  assign c53_63_io_in_1 = pp_13[7]; // @[Multiplier.scala 60:38]
  assign c53_63_io_in_2 = pp_14[5]; // @[Multiplier.scala 60:38]
  assign c53_63_io_in_3 = pp_15[3]; // @[Multiplier.scala 60:38]
  assign c53_63_io_in_4 = c53_59_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_64_io_in_0 = pp[32]; // @[Multiplier.scala 60:38]
  assign c53_64_io_in_1 = pp_1[32]; // @[Multiplier.scala 60:38]
  assign c53_64_io_in_2 = pp_2[30]; // @[Multiplier.scala 60:38]
  assign c53_64_io_in_3 = pp_3[28]; // @[Multiplier.scala 60:38]
  assign c53_64_io_in_4 = c53_60_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_65_io_in_0 = pp_4[26]; // @[Multiplier.scala 60:38]
  assign c53_65_io_in_1 = pp_5[24]; // @[Multiplier.scala 60:38]
  assign c53_65_io_in_2 = pp_6[22]; // @[Multiplier.scala 60:38]
  assign c53_65_io_in_3 = pp_7[20]; // @[Multiplier.scala 60:38]
  assign c53_65_io_in_4 = c53_61_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_66_io_in_0 = pp_8[18]; // @[Multiplier.scala 60:38]
  assign c53_66_io_in_1 = pp_9[16]; // @[Multiplier.scala 60:38]
  assign c53_66_io_in_2 = pp_10[14]; // @[Multiplier.scala 60:38]
  assign c53_66_io_in_3 = pp_11[12]; // @[Multiplier.scala 60:38]
  assign c53_66_io_in_4 = c53_62_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_67_io_in_0 = pp_12[10]; // @[Multiplier.scala 60:38]
  assign c53_67_io_in_1 = pp_13[8]; // @[Multiplier.scala 60:38]
  assign c53_67_io_in_2 = pp_14[6]; // @[Multiplier.scala 60:38]
  assign c53_67_io_in_3 = pp_15[4]; // @[Multiplier.scala 60:38]
  assign c53_67_io_in_4 = c53_63_io_out_1; // @[Multiplier.scala 89:41]
  assign c22_8_io_in_0 = pp_16[2]; // @[Multiplier.scala 60:38]
  assign c22_8_io_in_1 = pp_17[0]; // @[Multiplier.scala 60:38]
  assign c53_68_io_in_0 = pp[33]; // @[Multiplier.scala 60:38]
  assign c53_68_io_in_1 = pp_1[33]; // @[Multiplier.scala 60:38]
  assign c53_68_io_in_2 = pp_2[31]; // @[Multiplier.scala 60:38]
  assign c53_68_io_in_3 = pp_3[29]; // @[Multiplier.scala 60:38]
  assign c53_68_io_in_4 = c53_64_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_69_io_in_0 = pp_4[27]; // @[Multiplier.scala 60:38]
  assign c53_69_io_in_1 = pp_5[25]; // @[Multiplier.scala 60:38]
  assign c53_69_io_in_2 = pp_6[23]; // @[Multiplier.scala 60:38]
  assign c53_69_io_in_3 = pp_7[21]; // @[Multiplier.scala 60:38]
  assign c53_69_io_in_4 = c53_65_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_70_io_in_0 = pp_8[19]; // @[Multiplier.scala 60:38]
  assign c53_70_io_in_1 = pp_9[17]; // @[Multiplier.scala 60:38]
  assign c53_70_io_in_2 = pp_10[15]; // @[Multiplier.scala 60:38]
  assign c53_70_io_in_3 = pp_11[13]; // @[Multiplier.scala 60:38]
  assign c53_70_io_in_4 = c53_66_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_71_io_in_0 = pp_12[11]; // @[Multiplier.scala 60:38]
  assign c53_71_io_in_1 = pp_13[9]; // @[Multiplier.scala 60:38]
  assign c53_71_io_in_2 = pp_14[7]; // @[Multiplier.scala 60:38]
  assign c53_71_io_in_3 = pp_15[5]; // @[Multiplier.scala 60:38]
  assign c53_71_io_in_4 = c53_67_io_out_1; // @[Multiplier.scala 89:41]
  assign c22_9_io_in_0 = pp_16[3]; // @[Multiplier.scala 60:38]
  assign c22_9_io_in_1 = pp_17[1]; // @[Multiplier.scala 60:38]
  assign c53_72_io_in_0 = pp[34]; // @[Multiplier.scala 60:38]
  assign c53_72_io_in_1 = pp_1[34]; // @[Multiplier.scala 60:38]
  assign c53_72_io_in_2 = pp_2[32]; // @[Multiplier.scala 60:38]
  assign c53_72_io_in_3 = pp_3[30]; // @[Multiplier.scala 60:38]
  assign c53_72_io_in_4 = c53_68_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_73_io_in_0 = pp_4[28]; // @[Multiplier.scala 60:38]
  assign c53_73_io_in_1 = pp_5[26]; // @[Multiplier.scala 60:38]
  assign c53_73_io_in_2 = pp_6[24]; // @[Multiplier.scala 60:38]
  assign c53_73_io_in_3 = pp_7[22]; // @[Multiplier.scala 60:38]
  assign c53_73_io_in_4 = c53_69_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_74_io_in_0 = pp_8[20]; // @[Multiplier.scala 60:38]
  assign c53_74_io_in_1 = pp_9[18]; // @[Multiplier.scala 60:38]
  assign c53_74_io_in_2 = pp_10[16]; // @[Multiplier.scala 60:38]
  assign c53_74_io_in_3 = pp_11[14]; // @[Multiplier.scala 60:38]
  assign c53_74_io_in_4 = c53_70_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_75_io_in_0 = pp_12[12]; // @[Multiplier.scala 60:38]
  assign c53_75_io_in_1 = pp_13[10]; // @[Multiplier.scala 60:38]
  assign c53_75_io_in_2 = pp_14[8]; // @[Multiplier.scala 60:38]
  assign c53_75_io_in_3 = pp_15[6]; // @[Multiplier.scala 60:38]
  assign c53_75_io_in_4 = c53_71_io_out_1; // @[Multiplier.scala 89:41]
  assign c32_8_io_in_0 = pp_16[4]; // @[Multiplier.scala 60:38]
  assign c32_8_io_in_1 = pp_17[2]; // @[Multiplier.scala 60:38]
  assign c32_8_io_in_2 = pp_18[0]; // @[Multiplier.scala 60:38]
  assign c53_76_io_in_0 = pp[35]; // @[Multiplier.scala 60:38]
  assign c53_76_io_in_1 = pp_1[35]; // @[Multiplier.scala 60:38]
  assign c53_76_io_in_2 = pp_2[33]; // @[Multiplier.scala 60:38]
  assign c53_76_io_in_3 = pp_3[31]; // @[Multiplier.scala 60:38]
  assign c53_76_io_in_4 = c53_72_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_77_io_in_0 = pp_4[29]; // @[Multiplier.scala 60:38]
  assign c53_77_io_in_1 = pp_5[27]; // @[Multiplier.scala 60:38]
  assign c53_77_io_in_2 = pp_6[25]; // @[Multiplier.scala 60:38]
  assign c53_77_io_in_3 = pp_7[23]; // @[Multiplier.scala 60:38]
  assign c53_77_io_in_4 = c53_73_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_78_io_in_0 = pp_8[21]; // @[Multiplier.scala 60:38]
  assign c53_78_io_in_1 = pp_9[19]; // @[Multiplier.scala 60:38]
  assign c53_78_io_in_2 = pp_10[17]; // @[Multiplier.scala 60:38]
  assign c53_78_io_in_3 = pp_11[15]; // @[Multiplier.scala 60:38]
  assign c53_78_io_in_4 = c53_74_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_79_io_in_0 = pp_12[13]; // @[Multiplier.scala 60:38]
  assign c53_79_io_in_1 = pp_13[11]; // @[Multiplier.scala 60:38]
  assign c53_79_io_in_2 = pp_14[9]; // @[Multiplier.scala 60:38]
  assign c53_79_io_in_3 = pp_15[7]; // @[Multiplier.scala 60:38]
  assign c53_79_io_in_4 = c53_75_io_out_1; // @[Multiplier.scala 89:41]
  assign c32_9_io_in_0 = pp_16[5]; // @[Multiplier.scala 60:38]
  assign c32_9_io_in_1 = pp_17[3]; // @[Multiplier.scala 60:38]
  assign c32_9_io_in_2 = pp_18[1]; // @[Multiplier.scala 60:38]
  assign c53_80_io_in_0 = pp[36]; // @[Multiplier.scala 60:38]
  assign c53_80_io_in_1 = pp_1[36]; // @[Multiplier.scala 60:38]
  assign c53_80_io_in_2 = pp_2[34]; // @[Multiplier.scala 60:38]
  assign c53_80_io_in_3 = pp_3[32]; // @[Multiplier.scala 60:38]
  assign c53_80_io_in_4 = c53_76_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_81_io_in_0 = pp_4[30]; // @[Multiplier.scala 60:38]
  assign c53_81_io_in_1 = pp_5[28]; // @[Multiplier.scala 60:38]
  assign c53_81_io_in_2 = pp_6[26]; // @[Multiplier.scala 60:38]
  assign c53_81_io_in_3 = pp_7[24]; // @[Multiplier.scala 60:38]
  assign c53_81_io_in_4 = c53_77_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_82_io_in_0 = pp_8[22]; // @[Multiplier.scala 60:38]
  assign c53_82_io_in_1 = pp_9[20]; // @[Multiplier.scala 60:38]
  assign c53_82_io_in_2 = pp_10[18]; // @[Multiplier.scala 60:38]
  assign c53_82_io_in_3 = pp_11[16]; // @[Multiplier.scala 60:38]
  assign c53_82_io_in_4 = c53_78_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_83_io_in_0 = pp_12[14]; // @[Multiplier.scala 60:38]
  assign c53_83_io_in_1 = pp_13[12]; // @[Multiplier.scala 60:38]
  assign c53_83_io_in_2 = pp_14[10]; // @[Multiplier.scala 60:38]
  assign c53_83_io_in_3 = pp_15[8]; // @[Multiplier.scala 60:38]
  assign c53_83_io_in_4 = c53_79_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_84_io_in_0 = pp_16[6]; // @[Multiplier.scala 60:38]
  assign c53_84_io_in_1 = pp_17[4]; // @[Multiplier.scala 60:38]
  assign c53_84_io_in_2 = pp_18[2]; // @[Multiplier.scala 60:38]
  assign c53_84_io_in_3 = pp_19[0]; // @[Multiplier.scala 60:38]
  assign c53_84_io_in_4 = 1'h0; // @[Multiplier.scala 87:24]
  assign c53_85_io_in_0 = pp[37]; // @[Multiplier.scala 60:38]
  assign c53_85_io_in_1 = pp_1[37]; // @[Multiplier.scala 60:38]
  assign c53_85_io_in_2 = pp_2[35]; // @[Multiplier.scala 60:38]
  assign c53_85_io_in_3 = pp_3[33]; // @[Multiplier.scala 60:38]
  assign c53_85_io_in_4 = c53_80_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_86_io_in_0 = pp_4[31]; // @[Multiplier.scala 60:38]
  assign c53_86_io_in_1 = pp_5[29]; // @[Multiplier.scala 60:38]
  assign c53_86_io_in_2 = pp_6[27]; // @[Multiplier.scala 60:38]
  assign c53_86_io_in_3 = pp_7[25]; // @[Multiplier.scala 60:38]
  assign c53_86_io_in_4 = c53_81_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_87_io_in_0 = pp_8[23]; // @[Multiplier.scala 60:38]
  assign c53_87_io_in_1 = pp_9[21]; // @[Multiplier.scala 60:38]
  assign c53_87_io_in_2 = pp_10[19]; // @[Multiplier.scala 60:38]
  assign c53_87_io_in_3 = pp_11[17]; // @[Multiplier.scala 60:38]
  assign c53_87_io_in_4 = c53_82_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_88_io_in_0 = pp_12[15]; // @[Multiplier.scala 60:38]
  assign c53_88_io_in_1 = pp_13[13]; // @[Multiplier.scala 60:38]
  assign c53_88_io_in_2 = pp_14[11]; // @[Multiplier.scala 60:38]
  assign c53_88_io_in_3 = pp_15[9]; // @[Multiplier.scala 60:38]
  assign c53_88_io_in_4 = c53_83_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_89_io_in_0 = pp_16[7]; // @[Multiplier.scala 60:38]
  assign c53_89_io_in_1 = pp_17[5]; // @[Multiplier.scala 60:38]
  assign c53_89_io_in_2 = pp_18[3]; // @[Multiplier.scala 60:38]
  assign c53_89_io_in_3 = pp_19[1]; // @[Multiplier.scala 60:38]
  assign c53_89_io_in_4 = c53_84_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_90_io_in_0 = pp[38]; // @[Multiplier.scala 60:38]
  assign c53_90_io_in_1 = pp_1[38]; // @[Multiplier.scala 60:38]
  assign c53_90_io_in_2 = pp_2[36]; // @[Multiplier.scala 60:38]
  assign c53_90_io_in_3 = pp_3[34]; // @[Multiplier.scala 60:38]
  assign c53_90_io_in_4 = c53_85_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_91_io_in_0 = pp_4[32]; // @[Multiplier.scala 60:38]
  assign c53_91_io_in_1 = pp_5[30]; // @[Multiplier.scala 60:38]
  assign c53_91_io_in_2 = pp_6[28]; // @[Multiplier.scala 60:38]
  assign c53_91_io_in_3 = pp_7[26]; // @[Multiplier.scala 60:38]
  assign c53_91_io_in_4 = c53_86_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_92_io_in_0 = pp_8[24]; // @[Multiplier.scala 60:38]
  assign c53_92_io_in_1 = pp_9[22]; // @[Multiplier.scala 60:38]
  assign c53_92_io_in_2 = pp_10[20]; // @[Multiplier.scala 60:38]
  assign c53_92_io_in_3 = pp_11[18]; // @[Multiplier.scala 60:38]
  assign c53_92_io_in_4 = c53_87_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_93_io_in_0 = pp_12[16]; // @[Multiplier.scala 60:38]
  assign c53_93_io_in_1 = pp_13[14]; // @[Multiplier.scala 60:38]
  assign c53_93_io_in_2 = pp_14[12]; // @[Multiplier.scala 60:38]
  assign c53_93_io_in_3 = pp_15[10]; // @[Multiplier.scala 60:38]
  assign c53_93_io_in_4 = c53_88_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_94_io_in_0 = pp_16[8]; // @[Multiplier.scala 60:38]
  assign c53_94_io_in_1 = pp_17[6]; // @[Multiplier.scala 60:38]
  assign c53_94_io_in_2 = pp_18[4]; // @[Multiplier.scala 60:38]
  assign c53_94_io_in_3 = pp_19[2]; // @[Multiplier.scala 60:38]
  assign c53_94_io_in_4 = c53_89_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_95_io_in_0 = pp[39]; // @[Multiplier.scala 60:38]
  assign c53_95_io_in_1 = pp_1[39]; // @[Multiplier.scala 60:38]
  assign c53_95_io_in_2 = pp_2[37]; // @[Multiplier.scala 60:38]
  assign c53_95_io_in_3 = pp_3[35]; // @[Multiplier.scala 60:38]
  assign c53_95_io_in_4 = c53_90_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_96_io_in_0 = pp_4[33]; // @[Multiplier.scala 60:38]
  assign c53_96_io_in_1 = pp_5[31]; // @[Multiplier.scala 60:38]
  assign c53_96_io_in_2 = pp_6[29]; // @[Multiplier.scala 60:38]
  assign c53_96_io_in_3 = pp_7[27]; // @[Multiplier.scala 60:38]
  assign c53_96_io_in_4 = c53_91_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_97_io_in_0 = pp_8[25]; // @[Multiplier.scala 60:38]
  assign c53_97_io_in_1 = pp_9[23]; // @[Multiplier.scala 60:38]
  assign c53_97_io_in_2 = pp_10[21]; // @[Multiplier.scala 60:38]
  assign c53_97_io_in_3 = pp_11[19]; // @[Multiplier.scala 60:38]
  assign c53_97_io_in_4 = c53_92_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_98_io_in_0 = pp_12[17]; // @[Multiplier.scala 60:38]
  assign c53_98_io_in_1 = pp_13[15]; // @[Multiplier.scala 60:38]
  assign c53_98_io_in_2 = pp_14[13]; // @[Multiplier.scala 60:38]
  assign c53_98_io_in_3 = pp_15[11]; // @[Multiplier.scala 60:38]
  assign c53_98_io_in_4 = c53_93_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_99_io_in_0 = pp_16[9]; // @[Multiplier.scala 60:38]
  assign c53_99_io_in_1 = pp_17[7]; // @[Multiplier.scala 60:38]
  assign c53_99_io_in_2 = pp_18[5]; // @[Multiplier.scala 60:38]
  assign c53_99_io_in_3 = pp_19[3]; // @[Multiplier.scala 60:38]
  assign c53_99_io_in_4 = c53_94_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_100_io_in_0 = pp[40]; // @[Multiplier.scala 60:38]
  assign c53_100_io_in_1 = pp_1[40]; // @[Multiplier.scala 60:38]
  assign c53_100_io_in_2 = pp_2[38]; // @[Multiplier.scala 60:38]
  assign c53_100_io_in_3 = pp_3[36]; // @[Multiplier.scala 60:38]
  assign c53_100_io_in_4 = c53_95_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_101_io_in_0 = pp_4[34]; // @[Multiplier.scala 60:38]
  assign c53_101_io_in_1 = pp_5[32]; // @[Multiplier.scala 60:38]
  assign c53_101_io_in_2 = pp_6[30]; // @[Multiplier.scala 60:38]
  assign c53_101_io_in_3 = pp_7[28]; // @[Multiplier.scala 60:38]
  assign c53_101_io_in_4 = c53_96_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_102_io_in_0 = pp_8[26]; // @[Multiplier.scala 60:38]
  assign c53_102_io_in_1 = pp_9[24]; // @[Multiplier.scala 60:38]
  assign c53_102_io_in_2 = pp_10[22]; // @[Multiplier.scala 60:38]
  assign c53_102_io_in_3 = pp_11[20]; // @[Multiplier.scala 60:38]
  assign c53_102_io_in_4 = c53_97_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_103_io_in_0 = pp_12[18]; // @[Multiplier.scala 60:38]
  assign c53_103_io_in_1 = pp_13[16]; // @[Multiplier.scala 60:38]
  assign c53_103_io_in_2 = pp_14[14]; // @[Multiplier.scala 60:38]
  assign c53_103_io_in_3 = pp_15[12]; // @[Multiplier.scala 60:38]
  assign c53_103_io_in_4 = c53_98_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_104_io_in_0 = pp_16[10]; // @[Multiplier.scala 60:38]
  assign c53_104_io_in_1 = pp_17[8]; // @[Multiplier.scala 60:38]
  assign c53_104_io_in_2 = pp_18[6]; // @[Multiplier.scala 60:38]
  assign c53_104_io_in_3 = pp_19[4]; // @[Multiplier.scala 60:38]
  assign c53_104_io_in_4 = c53_99_io_out_1; // @[Multiplier.scala 89:41]
  assign c22_10_io_in_0 = pp_20[2]; // @[Multiplier.scala 60:38]
  assign c22_10_io_in_1 = pp_21[0]; // @[Multiplier.scala 60:38]
  assign c53_105_io_in_0 = pp[41]; // @[Multiplier.scala 60:38]
  assign c53_105_io_in_1 = pp_1[41]; // @[Multiplier.scala 60:38]
  assign c53_105_io_in_2 = pp_2[39]; // @[Multiplier.scala 60:38]
  assign c53_105_io_in_3 = pp_3[37]; // @[Multiplier.scala 60:38]
  assign c53_105_io_in_4 = c53_100_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_106_io_in_0 = pp_4[35]; // @[Multiplier.scala 60:38]
  assign c53_106_io_in_1 = pp_5[33]; // @[Multiplier.scala 60:38]
  assign c53_106_io_in_2 = pp_6[31]; // @[Multiplier.scala 60:38]
  assign c53_106_io_in_3 = pp_7[29]; // @[Multiplier.scala 60:38]
  assign c53_106_io_in_4 = c53_101_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_107_io_in_0 = pp_8[27]; // @[Multiplier.scala 60:38]
  assign c53_107_io_in_1 = pp_9[25]; // @[Multiplier.scala 60:38]
  assign c53_107_io_in_2 = pp_10[23]; // @[Multiplier.scala 60:38]
  assign c53_107_io_in_3 = pp_11[21]; // @[Multiplier.scala 60:38]
  assign c53_107_io_in_4 = c53_102_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_108_io_in_0 = pp_12[19]; // @[Multiplier.scala 60:38]
  assign c53_108_io_in_1 = pp_13[17]; // @[Multiplier.scala 60:38]
  assign c53_108_io_in_2 = pp_14[15]; // @[Multiplier.scala 60:38]
  assign c53_108_io_in_3 = pp_15[13]; // @[Multiplier.scala 60:38]
  assign c53_108_io_in_4 = c53_103_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_109_io_in_0 = pp_16[11]; // @[Multiplier.scala 60:38]
  assign c53_109_io_in_1 = pp_17[9]; // @[Multiplier.scala 60:38]
  assign c53_109_io_in_2 = pp_18[7]; // @[Multiplier.scala 60:38]
  assign c53_109_io_in_3 = pp_19[5]; // @[Multiplier.scala 60:38]
  assign c53_109_io_in_4 = c53_104_io_out_1; // @[Multiplier.scala 89:41]
  assign c22_11_io_in_0 = pp_20[3]; // @[Multiplier.scala 60:38]
  assign c22_11_io_in_1 = pp_21[1]; // @[Multiplier.scala 60:38]
  assign c53_110_io_in_0 = pp[42]; // @[Multiplier.scala 60:38]
  assign c53_110_io_in_1 = pp_1[42]; // @[Multiplier.scala 60:38]
  assign c53_110_io_in_2 = pp_2[40]; // @[Multiplier.scala 60:38]
  assign c53_110_io_in_3 = pp_3[38]; // @[Multiplier.scala 60:38]
  assign c53_110_io_in_4 = c53_105_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_111_io_in_0 = pp_4[36]; // @[Multiplier.scala 60:38]
  assign c53_111_io_in_1 = pp_5[34]; // @[Multiplier.scala 60:38]
  assign c53_111_io_in_2 = pp_6[32]; // @[Multiplier.scala 60:38]
  assign c53_111_io_in_3 = pp_7[30]; // @[Multiplier.scala 60:38]
  assign c53_111_io_in_4 = c53_106_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_112_io_in_0 = pp_8[28]; // @[Multiplier.scala 60:38]
  assign c53_112_io_in_1 = pp_9[26]; // @[Multiplier.scala 60:38]
  assign c53_112_io_in_2 = pp_10[24]; // @[Multiplier.scala 60:38]
  assign c53_112_io_in_3 = pp_11[22]; // @[Multiplier.scala 60:38]
  assign c53_112_io_in_4 = c53_107_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_113_io_in_0 = pp_12[20]; // @[Multiplier.scala 60:38]
  assign c53_113_io_in_1 = pp_13[18]; // @[Multiplier.scala 60:38]
  assign c53_113_io_in_2 = pp_14[16]; // @[Multiplier.scala 60:38]
  assign c53_113_io_in_3 = pp_15[14]; // @[Multiplier.scala 60:38]
  assign c53_113_io_in_4 = c53_108_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_114_io_in_0 = pp_16[12]; // @[Multiplier.scala 60:38]
  assign c53_114_io_in_1 = pp_17[10]; // @[Multiplier.scala 60:38]
  assign c53_114_io_in_2 = pp_18[8]; // @[Multiplier.scala 60:38]
  assign c53_114_io_in_3 = pp_19[6]; // @[Multiplier.scala 60:38]
  assign c53_114_io_in_4 = c53_109_io_out_1; // @[Multiplier.scala 89:41]
  assign c32_10_io_in_0 = pp_20[4]; // @[Multiplier.scala 60:38]
  assign c32_10_io_in_1 = pp_21[2]; // @[Multiplier.scala 60:38]
  assign c32_10_io_in_2 = pp_22[0]; // @[Multiplier.scala 60:38]
  assign c53_115_io_in_0 = pp[43]; // @[Multiplier.scala 60:38]
  assign c53_115_io_in_1 = pp_1[43]; // @[Multiplier.scala 60:38]
  assign c53_115_io_in_2 = pp_2[41]; // @[Multiplier.scala 60:38]
  assign c53_115_io_in_3 = pp_3[39]; // @[Multiplier.scala 60:38]
  assign c53_115_io_in_4 = c53_110_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_116_io_in_0 = pp_4[37]; // @[Multiplier.scala 60:38]
  assign c53_116_io_in_1 = pp_5[35]; // @[Multiplier.scala 60:38]
  assign c53_116_io_in_2 = pp_6[33]; // @[Multiplier.scala 60:38]
  assign c53_116_io_in_3 = pp_7[31]; // @[Multiplier.scala 60:38]
  assign c53_116_io_in_4 = c53_111_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_117_io_in_0 = pp_8[29]; // @[Multiplier.scala 60:38]
  assign c53_117_io_in_1 = pp_9[27]; // @[Multiplier.scala 60:38]
  assign c53_117_io_in_2 = pp_10[25]; // @[Multiplier.scala 60:38]
  assign c53_117_io_in_3 = pp_11[23]; // @[Multiplier.scala 60:38]
  assign c53_117_io_in_4 = c53_112_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_118_io_in_0 = pp_12[21]; // @[Multiplier.scala 60:38]
  assign c53_118_io_in_1 = pp_13[19]; // @[Multiplier.scala 60:38]
  assign c53_118_io_in_2 = pp_14[17]; // @[Multiplier.scala 60:38]
  assign c53_118_io_in_3 = pp_15[15]; // @[Multiplier.scala 60:38]
  assign c53_118_io_in_4 = c53_113_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_119_io_in_0 = pp_16[13]; // @[Multiplier.scala 60:38]
  assign c53_119_io_in_1 = pp_17[11]; // @[Multiplier.scala 60:38]
  assign c53_119_io_in_2 = pp_18[9]; // @[Multiplier.scala 60:38]
  assign c53_119_io_in_3 = pp_19[7]; // @[Multiplier.scala 60:38]
  assign c53_119_io_in_4 = c53_114_io_out_1; // @[Multiplier.scala 89:41]
  assign c32_11_io_in_0 = pp_20[5]; // @[Multiplier.scala 60:38]
  assign c32_11_io_in_1 = pp_21[3]; // @[Multiplier.scala 60:38]
  assign c32_11_io_in_2 = pp_22[1]; // @[Multiplier.scala 60:38]
  assign c53_120_io_in_0 = pp[44]; // @[Multiplier.scala 60:38]
  assign c53_120_io_in_1 = pp_1[44]; // @[Multiplier.scala 60:38]
  assign c53_120_io_in_2 = pp_2[42]; // @[Multiplier.scala 60:38]
  assign c53_120_io_in_3 = pp_3[40]; // @[Multiplier.scala 60:38]
  assign c53_120_io_in_4 = c53_115_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_121_io_in_0 = pp_4[38]; // @[Multiplier.scala 60:38]
  assign c53_121_io_in_1 = pp_5[36]; // @[Multiplier.scala 60:38]
  assign c53_121_io_in_2 = pp_6[34]; // @[Multiplier.scala 60:38]
  assign c53_121_io_in_3 = pp_7[32]; // @[Multiplier.scala 60:38]
  assign c53_121_io_in_4 = c53_116_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_122_io_in_0 = pp_8[30]; // @[Multiplier.scala 60:38]
  assign c53_122_io_in_1 = pp_9[28]; // @[Multiplier.scala 60:38]
  assign c53_122_io_in_2 = pp_10[26]; // @[Multiplier.scala 60:38]
  assign c53_122_io_in_3 = pp_11[24]; // @[Multiplier.scala 60:38]
  assign c53_122_io_in_4 = c53_117_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_123_io_in_0 = pp_12[22]; // @[Multiplier.scala 60:38]
  assign c53_123_io_in_1 = pp_13[20]; // @[Multiplier.scala 60:38]
  assign c53_123_io_in_2 = pp_14[18]; // @[Multiplier.scala 60:38]
  assign c53_123_io_in_3 = pp_15[16]; // @[Multiplier.scala 60:38]
  assign c53_123_io_in_4 = c53_118_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_124_io_in_0 = pp_16[14]; // @[Multiplier.scala 60:38]
  assign c53_124_io_in_1 = pp_17[12]; // @[Multiplier.scala 60:38]
  assign c53_124_io_in_2 = pp_18[10]; // @[Multiplier.scala 60:38]
  assign c53_124_io_in_3 = pp_19[8]; // @[Multiplier.scala 60:38]
  assign c53_124_io_in_4 = c53_119_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_125_io_in_0 = pp_20[6]; // @[Multiplier.scala 60:38]
  assign c53_125_io_in_1 = pp_21[4]; // @[Multiplier.scala 60:38]
  assign c53_125_io_in_2 = pp_22[2]; // @[Multiplier.scala 60:38]
  assign c53_125_io_in_3 = pp_23[0]; // @[Multiplier.scala 60:38]
  assign c53_125_io_in_4 = 1'h0; // @[Multiplier.scala 87:24]
  assign c53_126_io_in_0 = pp[45]; // @[Multiplier.scala 60:38]
  assign c53_126_io_in_1 = pp_1[45]; // @[Multiplier.scala 60:38]
  assign c53_126_io_in_2 = pp_2[43]; // @[Multiplier.scala 60:38]
  assign c53_126_io_in_3 = pp_3[41]; // @[Multiplier.scala 60:38]
  assign c53_126_io_in_4 = c53_120_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_127_io_in_0 = pp_4[39]; // @[Multiplier.scala 60:38]
  assign c53_127_io_in_1 = pp_5[37]; // @[Multiplier.scala 60:38]
  assign c53_127_io_in_2 = pp_6[35]; // @[Multiplier.scala 60:38]
  assign c53_127_io_in_3 = pp_7[33]; // @[Multiplier.scala 60:38]
  assign c53_127_io_in_4 = c53_121_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_128_io_in_0 = pp_8[31]; // @[Multiplier.scala 60:38]
  assign c53_128_io_in_1 = pp_9[29]; // @[Multiplier.scala 60:38]
  assign c53_128_io_in_2 = pp_10[27]; // @[Multiplier.scala 60:38]
  assign c53_128_io_in_3 = pp_11[25]; // @[Multiplier.scala 60:38]
  assign c53_128_io_in_4 = c53_122_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_129_io_in_0 = pp_12[23]; // @[Multiplier.scala 60:38]
  assign c53_129_io_in_1 = pp_13[21]; // @[Multiplier.scala 60:38]
  assign c53_129_io_in_2 = pp_14[19]; // @[Multiplier.scala 60:38]
  assign c53_129_io_in_3 = pp_15[17]; // @[Multiplier.scala 60:38]
  assign c53_129_io_in_4 = c53_123_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_130_io_in_0 = pp_16[15]; // @[Multiplier.scala 60:38]
  assign c53_130_io_in_1 = pp_17[13]; // @[Multiplier.scala 60:38]
  assign c53_130_io_in_2 = pp_18[11]; // @[Multiplier.scala 60:38]
  assign c53_130_io_in_3 = pp_19[9]; // @[Multiplier.scala 60:38]
  assign c53_130_io_in_4 = c53_124_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_131_io_in_0 = pp_20[7]; // @[Multiplier.scala 60:38]
  assign c53_131_io_in_1 = pp_21[5]; // @[Multiplier.scala 60:38]
  assign c53_131_io_in_2 = pp_22[3]; // @[Multiplier.scala 60:38]
  assign c53_131_io_in_3 = pp_23[1]; // @[Multiplier.scala 60:38]
  assign c53_131_io_in_4 = c53_125_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_132_io_in_0 = pp[46]; // @[Multiplier.scala 60:38]
  assign c53_132_io_in_1 = pp_1[46]; // @[Multiplier.scala 60:38]
  assign c53_132_io_in_2 = pp_2[44]; // @[Multiplier.scala 60:38]
  assign c53_132_io_in_3 = pp_3[42]; // @[Multiplier.scala 60:38]
  assign c53_132_io_in_4 = c53_126_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_133_io_in_0 = pp_4[40]; // @[Multiplier.scala 60:38]
  assign c53_133_io_in_1 = pp_5[38]; // @[Multiplier.scala 60:38]
  assign c53_133_io_in_2 = pp_6[36]; // @[Multiplier.scala 60:38]
  assign c53_133_io_in_3 = pp_7[34]; // @[Multiplier.scala 60:38]
  assign c53_133_io_in_4 = c53_127_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_134_io_in_0 = pp_8[32]; // @[Multiplier.scala 60:38]
  assign c53_134_io_in_1 = pp_9[30]; // @[Multiplier.scala 60:38]
  assign c53_134_io_in_2 = pp_10[28]; // @[Multiplier.scala 60:38]
  assign c53_134_io_in_3 = pp_11[26]; // @[Multiplier.scala 60:38]
  assign c53_134_io_in_4 = c53_128_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_135_io_in_0 = pp_12[24]; // @[Multiplier.scala 60:38]
  assign c53_135_io_in_1 = pp_13[22]; // @[Multiplier.scala 60:38]
  assign c53_135_io_in_2 = pp_14[20]; // @[Multiplier.scala 60:38]
  assign c53_135_io_in_3 = pp_15[18]; // @[Multiplier.scala 60:38]
  assign c53_135_io_in_4 = c53_129_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_136_io_in_0 = pp_16[16]; // @[Multiplier.scala 60:38]
  assign c53_136_io_in_1 = pp_17[14]; // @[Multiplier.scala 60:38]
  assign c53_136_io_in_2 = pp_18[12]; // @[Multiplier.scala 60:38]
  assign c53_136_io_in_3 = pp_19[10]; // @[Multiplier.scala 60:38]
  assign c53_136_io_in_4 = c53_130_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_137_io_in_0 = pp_20[8]; // @[Multiplier.scala 60:38]
  assign c53_137_io_in_1 = pp_21[6]; // @[Multiplier.scala 60:38]
  assign c53_137_io_in_2 = pp_22[4]; // @[Multiplier.scala 60:38]
  assign c53_137_io_in_3 = pp_23[2]; // @[Multiplier.scala 60:38]
  assign c53_137_io_in_4 = c53_131_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_138_io_in_0 = pp[47]; // @[Multiplier.scala 60:38]
  assign c53_138_io_in_1 = pp_1[47]; // @[Multiplier.scala 60:38]
  assign c53_138_io_in_2 = pp_2[45]; // @[Multiplier.scala 60:38]
  assign c53_138_io_in_3 = pp_3[43]; // @[Multiplier.scala 60:38]
  assign c53_138_io_in_4 = c53_132_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_139_io_in_0 = pp_4[41]; // @[Multiplier.scala 60:38]
  assign c53_139_io_in_1 = pp_5[39]; // @[Multiplier.scala 60:38]
  assign c53_139_io_in_2 = pp_6[37]; // @[Multiplier.scala 60:38]
  assign c53_139_io_in_3 = pp_7[35]; // @[Multiplier.scala 60:38]
  assign c53_139_io_in_4 = c53_133_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_140_io_in_0 = pp_8[33]; // @[Multiplier.scala 60:38]
  assign c53_140_io_in_1 = pp_9[31]; // @[Multiplier.scala 60:38]
  assign c53_140_io_in_2 = pp_10[29]; // @[Multiplier.scala 60:38]
  assign c53_140_io_in_3 = pp_11[27]; // @[Multiplier.scala 60:38]
  assign c53_140_io_in_4 = c53_134_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_141_io_in_0 = pp_12[25]; // @[Multiplier.scala 60:38]
  assign c53_141_io_in_1 = pp_13[23]; // @[Multiplier.scala 60:38]
  assign c53_141_io_in_2 = pp_14[21]; // @[Multiplier.scala 60:38]
  assign c53_141_io_in_3 = pp_15[19]; // @[Multiplier.scala 60:38]
  assign c53_141_io_in_4 = c53_135_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_142_io_in_0 = pp_16[17]; // @[Multiplier.scala 60:38]
  assign c53_142_io_in_1 = pp_17[15]; // @[Multiplier.scala 60:38]
  assign c53_142_io_in_2 = pp_18[13]; // @[Multiplier.scala 60:38]
  assign c53_142_io_in_3 = pp_19[11]; // @[Multiplier.scala 60:38]
  assign c53_142_io_in_4 = c53_136_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_143_io_in_0 = pp_20[9]; // @[Multiplier.scala 60:38]
  assign c53_143_io_in_1 = pp_21[7]; // @[Multiplier.scala 60:38]
  assign c53_143_io_in_2 = pp_22[5]; // @[Multiplier.scala 60:38]
  assign c53_143_io_in_3 = pp_23[3]; // @[Multiplier.scala 60:38]
  assign c53_143_io_in_4 = c53_137_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_144_io_in_0 = pp[48]; // @[Multiplier.scala 60:38]
  assign c53_144_io_in_1 = pp_1[48]; // @[Multiplier.scala 60:38]
  assign c53_144_io_in_2 = pp_2[46]; // @[Multiplier.scala 60:38]
  assign c53_144_io_in_3 = pp_3[44]; // @[Multiplier.scala 60:38]
  assign c53_144_io_in_4 = c53_138_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_145_io_in_0 = pp_4[42]; // @[Multiplier.scala 60:38]
  assign c53_145_io_in_1 = pp_5[40]; // @[Multiplier.scala 60:38]
  assign c53_145_io_in_2 = pp_6[38]; // @[Multiplier.scala 60:38]
  assign c53_145_io_in_3 = pp_7[36]; // @[Multiplier.scala 60:38]
  assign c53_145_io_in_4 = c53_139_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_146_io_in_0 = pp_8[34]; // @[Multiplier.scala 60:38]
  assign c53_146_io_in_1 = pp_9[32]; // @[Multiplier.scala 60:38]
  assign c53_146_io_in_2 = pp_10[30]; // @[Multiplier.scala 60:38]
  assign c53_146_io_in_3 = pp_11[28]; // @[Multiplier.scala 60:38]
  assign c53_146_io_in_4 = c53_140_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_147_io_in_0 = pp_12[26]; // @[Multiplier.scala 60:38]
  assign c53_147_io_in_1 = pp_13[24]; // @[Multiplier.scala 60:38]
  assign c53_147_io_in_2 = pp_14[22]; // @[Multiplier.scala 60:38]
  assign c53_147_io_in_3 = pp_15[20]; // @[Multiplier.scala 60:38]
  assign c53_147_io_in_4 = c53_141_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_148_io_in_0 = pp_16[18]; // @[Multiplier.scala 60:38]
  assign c53_148_io_in_1 = pp_17[16]; // @[Multiplier.scala 60:38]
  assign c53_148_io_in_2 = pp_18[14]; // @[Multiplier.scala 60:38]
  assign c53_148_io_in_3 = pp_19[12]; // @[Multiplier.scala 60:38]
  assign c53_148_io_in_4 = c53_142_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_149_io_in_0 = pp_20[10]; // @[Multiplier.scala 60:38]
  assign c53_149_io_in_1 = pp_21[8]; // @[Multiplier.scala 60:38]
  assign c53_149_io_in_2 = pp_22[6]; // @[Multiplier.scala 60:38]
  assign c53_149_io_in_3 = pp_23[4]; // @[Multiplier.scala 60:38]
  assign c53_149_io_in_4 = c53_143_io_out_1; // @[Multiplier.scala 89:41]
  assign c22_12_io_in_0 = pp_24[2]; // @[Multiplier.scala 60:38]
  assign c22_12_io_in_1 = pp_25[0]; // @[Multiplier.scala 60:38]
  assign c53_150_io_in_0 = pp[49]; // @[Multiplier.scala 60:38]
  assign c53_150_io_in_1 = pp_1[49]; // @[Multiplier.scala 60:38]
  assign c53_150_io_in_2 = pp_2[47]; // @[Multiplier.scala 60:38]
  assign c53_150_io_in_3 = pp_3[45]; // @[Multiplier.scala 60:38]
  assign c53_150_io_in_4 = c53_144_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_151_io_in_0 = pp_4[43]; // @[Multiplier.scala 60:38]
  assign c53_151_io_in_1 = pp_5[41]; // @[Multiplier.scala 60:38]
  assign c53_151_io_in_2 = pp_6[39]; // @[Multiplier.scala 60:38]
  assign c53_151_io_in_3 = pp_7[37]; // @[Multiplier.scala 60:38]
  assign c53_151_io_in_4 = c53_145_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_152_io_in_0 = pp_8[35]; // @[Multiplier.scala 60:38]
  assign c53_152_io_in_1 = pp_9[33]; // @[Multiplier.scala 60:38]
  assign c53_152_io_in_2 = pp_10[31]; // @[Multiplier.scala 60:38]
  assign c53_152_io_in_3 = pp_11[29]; // @[Multiplier.scala 60:38]
  assign c53_152_io_in_4 = c53_146_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_153_io_in_0 = pp_12[27]; // @[Multiplier.scala 60:38]
  assign c53_153_io_in_1 = pp_13[25]; // @[Multiplier.scala 60:38]
  assign c53_153_io_in_2 = pp_14[23]; // @[Multiplier.scala 60:38]
  assign c53_153_io_in_3 = pp_15[21]; // @[Multiplier.scala 60:38]
  assign c53_153_io_in_4 = c53_147_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_154_io_in_0 = pp_16[19]; // @[Multiplier.scala 60:38]
  assign c53_154_io_in_1 = pp_17[17]; // @[Multiplier.scala 60:38]
  assign c53_154_io_in_2 = pp_18[15]; // @[Multiplier.scala 60:38]
  assign c53_154_io_in_3 = pp_19[13]; // @[Multiplier.scala 60:38]
  assign c53_154_io_in_4 = c53_148_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_155_io_in_0 = pp_20[11]; // @[Multiplier.scala 60:38]
  assign c53_155_io_in_1 = pp_21[9]; // @[Multiplier.scala 60:38]
  assign c53_155_io_in_2 = pp_22[7]; // @[Multiplier.scala 60:38]
  assign c53_155_io_in_3 = pp_23[5]; // @[Multiplier.scala 60:38]
  assign c53_155_io_in_4 = c53_149_io_out_1; // @[Multiplier.scala 89:41]
  assign c22_13_io_in_0 = pp_24[3]; // @[Multiplier.scala 60:38]
  assign c22_13_io_in_1 = pp_25[1]; // @[Multiplier.scala 60:38]
  assign c53_156_io_in_0 = pp[50]; // @[Multiplier.scala 60:38]
  assign c53_156_io_in_1 = pp_1[50]; // @[Multiplier.scala 60:38]
  assign c53_156_io_in_2 = pp_2[48]; // @[Multiplier.scala 60:38]
  assign c53_156_io_in_3 = pp_3[46]; // @[Multiplier.scala 60:38]
  assign c53_156_io_in_4 = c53_150_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_157_io_in_0 = pp_4[44]; // @[Multiplier.scala 60:38]
  assign c53_157_io_in_1 = pp_5[42]; // @[Multiplier.scala 60:38]
  assign c53_157_io_in_2 = pp_6[40]; // @[Multiplier.scala 60:38]
  assign c53_157_io_in_3 = pp_7[38]; // @[Multiplier.scala 60:38]
  assign c53_157_io_in_4 = c53_151_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_158_io_in_0 = pp_8[36]; // @[Multiplier.scala 60:38]
  assign c53_158_io_in_1 = pp_9[34]; // @[Multiplier.scala 60:38]
  assign c53_158_io_in_2 = pp_10[32]; // @[Multiplier.scala 60:38]
  assign c53_158_io_in_3 = pp_11[30]; // @[Multiplier.scala 60:38]
  assign c53_158_io_in_4 = c53_152_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_159_io_in_0 = pp_12[28]; // @[Multiplier.scala 60:38]
  assign c53_159_io_in_1 = pp_13[26]; // @[Multiplier.scala 60:38]
  assign c53_159_io_in_2 = pp_14[24]; // @[Multiplier.scala 60:38]
  assign c53_159_io_in_3 = pp_15[22]; // @[Multiplier.scala 60:38]
  assign c53_159_io_in_4 = c53_153_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_160_io_in_0 = pp_16[20]; // @[Multiplier.scala 60:38]
  assign c53_160_io_in_1 = pp_17[18]; // @[Multiplier.scala 60:38]
  assign c53_160_io_in_2 = pp_18[16]; // @[Multiplier.scala 60:38]
  assign c53_160_io_in_3 = pp_19[14]; // @[Multiplier.scala 60:38]
  assign c53_160_io_in_4 = c53_154_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_161_io_in_0 = pp_20[12]; // @[Multiplier.scala 60:38]
  assign c53_161_io_in_1 = pp_21[10]; // @[Multiplier.scala 60:38]
  assign c53_161_io_in_2 = pp_22[8]; // @[Multiplier.scala 60:38]
  assign c53_161_io_in_3 = pp_23[6]; // @[Multiplier.scala 60:38]
  assign c53_161_io_in_4 = c53_155_io_out_1; // @[Multiplier.scala 89:41]
  assign c32_12_io_in_0 = pp_24[4]; // @[Multiplier.scala 60:38]
  assign c32_12_io_in_1 = pp_25[2]; // @[Multiplier.scala 60:38]
  assign c32_12_io_in_2 = pp_26[0]; // @[Multiplier.scala 60:38]
  assign c53_162_io_in_0 = pp[51]; // @[Multiplier.scala 60:38]
  assign c53_162_io_in_1 = pp_1[51]; // @[Multiplier.scala 60:38]
  assign c53_162_io_in_2 = pp_2[49]; // @[Multiplier.scala 60:38]
  assign c53_162_io_in_3 = pp_3[47]; // @[Multiplier.scala 60:38]
  assign c53_162_io_in_4 = c53_156_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_163_io_in_0 = pp_4[45]; // @[Multiplier.scala 60:38]
  assign c53_163_io_in_1 = pp_5[43]; // @[Multiplier.scala 60:38]
  assign c53_163_io_in_2 = pp_6[41]; // @[Multiplier.scala 60:38]
  assign c53_163_io_in_3 = pp_7[39]; // @[Multiplier.scala 60:38]
  assign c53_163_io_in_4 = c53_157_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_164_io_in_0 = pp_8[37]; // @[Multiplier.scala 60:38]
  assign c53_164_io_in_1 = pp_9[35]; // @[Multiplier.scala 60:38]
  assign c53_164_io_in_2 = pp_10[33]; // @[Multiplier.scala 60:38]
  assign c53_164_io_in_3 = pp_11[31]; // @[Multiplier.scala 60:38]
  assign c53_164_io_in_4 = c53_158_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_165_io_in_0 = pp_12[29]; // @[Multiplier.scala 60:38]
  assign c53_165_io_in_1 = pp_13[27]; // @[Multiplier.scala 60:38]
  assign c53_165_io_in_2 = pp_14[25]; // @[Multiplier.scala 60:38]
  assign c53_165_io_in_3 = pp_15[23]; // @[Multiplier.scala 60:38]
  assign c53_165_io_in_4 = c53_159_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_166_io_in_0 = pp_16[21]; // @[Multiplier.scala 60:38]
  assign c53_166_io_in_1 = pp_17[19]; // @[Multiplier.scala 60:38]
  assign c53_166_io_in_2 = pp_18[17]; // @[Multiplier.scala 60:38]
  assign c53_166_io_in_3 = pp_19[15]; // @[Multiplier.scala 60:38]
  assign c53_166_io_in_4 = c53_160_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_167_io_in_0 = pp_20[13]; // @[Multiplier.scala 60:38]
  assign c53_167_io_in_1 = pp_21[11]; // @[Multiplier.scala 60:38]
  assign c53_167_io_in_2 = pp_22[9]; // @[Multiplier.scala 60:38]
  assign c53_167_io_in_3 = pp_23[7]; // @[Multiplier.scala 60:38]
  assign c53_167_io_in_4 = c53_161_io_out_1; // @[Multiplier.scala 89:41]
  assign c32_13_io_in_0 = pp_24[5]; // @[Multiplier.scala 60:38]
  assign c32_13_io_in_1 = pp_25[3]; // @[Multiplier.scala 60:38]
  assign c32_13_io_in_2 = pp_26[1]; // @[Multiplier.scala 60:38]
  assign c53_168_io_in_0 = pp[52]; // @[Multiplier.scala 60:38]
  assign c53_168_io_in_1 = pp_1[52]; // @[Multiplier.scala 60:38]
  assign c53_168_io_in_2 = pp_2[50]; // @[Multiplier.scala 60:38]
  assign c53_168_io_in_3 = pp_3[48]; // @[Multiplier.scala 60:38]
  assign c53_168_io_in_4 = c53_162_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_169_io_in_0 = pp_4[46]; // @[Multiplier.scala 60:38]
  assign c53_169_io_in_1 = pp_5[44]; // @[Multiplier.scala 60:38]
  assign c53_169_io_in_2 = pp_6[42]; // @[Multiplier.scala 60:38]
  assign c53_169_io_in_3 = pp_7[40]; // @[Multiplier.scala 60:38]
  assign c53_169_io_in_4 = c53_163_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_170_io_in_0 = pp_8[38]; // @[Multiplier.scala 60:38]
  assign c53_170_io_in_1 = pp_9[36]; // @[Multiplier.scala 60:38]
  assign c53_170_io_in_2 = pp_10[34]; // @[Multiplier.scala 60:38]
  assign c53_170_io_in_3 = pp_11[32]; // @[Multiplier.scala 60:38]
  assign c53_170_io_in_4 = c53_164_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_171_io_in_0 = pp_12[30]; // @[Multiplier.scala 60:38]
  assign c53_171_io_in_1 = pp_13[28]; // @[Multiplier.scala 60:38]
  assign c53_171_io_in_2 = pp_14[26]; // @[Multiplier.scala 60:38]
  assign c53_171_io_in_3 = pp_15[24]; // @[Multiplier.scala 60:38]
  assign c53_171_io_in_4 = c53_165_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_172_io_in_0 = pp_16[22]; // @[Multiplier.scala 60:38]
  assign c53_172_io_in_1 = pp_17[20]; // @[Multiplier.scala 60:38]
  assign c53_172_io_in_2 = pp_18[18]; // @[Multiplier.scala 60:38]
  assign c53_172_io_in_3 = pp_19[16]; // @[Multiplier.scala 60:38]
  assign c53_172_io_in_4 = c53_166_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_173_io_in_0 = pp_20[14]; // @[Multiplier.scala 60:38]
  assign c53_173_io_in_1 = pp_21[12]; // @[Multiplier.scala 60:38]
  assign c53_173_io_in_2 = pp_22[10]; // @[Multiplier.scala 60:38]
  assign c53_173_io_in_3 = pp_23[8]; // @[Multiplier.scala 60:38]
  assign c53_173_io_in_4 = c53_167_io_out_1; // @[Multiplier.scala 89:41]
  assign c32_14_io_in_0 = pp_24[6]; // @[Multiplier.scala 60:38]
  assign c32_14_io_in_1 = pp_25[4]; // @[Multiplier.scala 60:38]
  assign c32_14_io_in_2 = pp_26[2]; // @[Multiplier.scala 60:38]
  assign c53_174_io_in_0 = pp[53]; // @[Multiplier.scala 60:38]
  assign c53_174_io_in_1 = pp_1[53]; // @[Multiplier.scala 60:38]
  assign c53_174_io_in_2 = pp_2[51]; // @[Multiplier.scala 60:38]
  assign c53_174_io_in_3 = pp_3[49]; // @[Multiplier.scala 60:38]
  assign c53_174_io_in_4 = c53_168_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_175_io_in_0 = pp_4[47]; // @[Multiplier.scala 60:38]
  assign c53_175_io_in_1 = pp_5[45]; // @[Multiplier.scala 60:38]
  assign c53_175_io_in_2 = pp_6[43]; // @[Multiplier.scala 60:38]
  assign c53_175_io_in_3 = pp_7[41]; // @[Multiplier.scala 60:38]
  assign c53_175_io_in_4 = c53_169_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_176_io_in_0 = pp_8[39]; // @[Multiplier.scala 60:38]
  assign c53_176_io_in_1 = pp_9[37]; // @[Multiplier.scala 60:38]
  assign c53_176_io_in_2 = pp_10[35]; // @[Multiplier.scala 60:38]
  assign c53_176_io_in_3 = pp_11[33]; // @[Multiplier.scala 60:38]
  assign c53_176_io_in_4 = c53_170_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_177_io_in_0 = pp_12[31]; // @[Multiplier.scala 60:38]
  assign c53_177_io_in_1 = pp_13[29]; // @[Multiplier.scala 60:38]
  assign c53_177_io_in_2 = pp_14[27]; // @[Multiplier.scala 60:38]
  assign c53_177_io_in_3 = pp_15[25]; // @[Multiplier.scala 60:38]
  assign c53_177_io_in_4 = c53_171_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_178_io_in_0 = pp_16[23]; // @[Multiplier.scala 60:38]
  assign c53_178_io_in_1 = pp_17[21]; // @[Multiplier.scala 60:38]
  assign c53_178_io_in_2 = pp_18[19]; // @[Multiplier.scala 60:38]
  assign c53_178_io_in_3 = pp_19[17]; // @[Multiplier.scala 60:38]
  assign c53_178_io_in_4 = c53_172_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_179_io_in_0 = pp_20[15]; // @[Multiplier.scala 60:38]
  assign c53_179_io_in_1 = pp_21[13]; // @[Multiplier.scala 60:38]
  assign c53_179_io_in_2 = pp_22[11]; // @[Multiplier.scala 60:38]
  assign c53_179_io_in_3 = pp_23[9]; // @[Multiplier.scala 60:38]
  assign c53_179_io_in_4 = c53_173_io_out_1; // @[Multiplier.scala 89:41]
  assign c32_15_io_in_0 = pp_24[7]; // @[Multiplier.scala 60:38]
  assign c32_15_io_in_1 = pp_25[5]; // @[Multiplier.scala 60:38]
  assign c32_15_io_in_2 = pp_26[3]; // @[Multiplier.scala 60:38]
  assign c53_180_io_in_0 = pp[54]; // @[Multiplier.scala 60:38]
  assign c53_180_io_in_1 = pp_1[54]; // @[Multiplier.scala 60:38]
  assign c53_180_io_in_2 = pp_2[52]; // @[Multiplier.scala 60:38]
  assign c53_180_io_in_3 = pp_3[50]; // @[Multiplier.scala 60:38]
  assign c53_180_io_in_4 = c53_174_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_181_io_in_0 = pp_4[48]; // @[Multiplier.scala 60:38]
  assign c53_181_io_in_1 = pp_5[46]; // @[Multiplier.scala 60:38]
  assign c53_181_io_in_2 = pp_6[44]; // @[Multiplier.scala 60:38]
  assign c53_181_io_in_3 = pp_7[42]; // @[Multiplier.scala 60:38]
  assign c53_181_io_in_4 = c53_175_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_182_io_in_0 = pp_8[40]; // @[Multiplier.scala 60:38]
  assign c53_182_io_in_1 = pp_9[38]; // @[Multiplier.scala 60:38]
  assign c53_182_io_in_2 = pp_10[36]; // @[Multiplier.scala 60:38]
  assign c53_182_io_in_3 = pp_11[34]; // @[Multiplier.scala 60:38]
  assign c53_182_io_in_4 = c53_176_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_183_io_in_0 = pp_12[32]; // @[Multiplier.scala 60:38]
  assign c53_183_io_in_1 = pp_13[30]; // @[Multiplier.scala 60:38]
  assign c53_183_io_in_2 = pp_14[28]; // @[Multiplier.scala 60:38]
  assign c53_183_io_in_3 = pp_15[26]; // @[Multiplier.scala 60:38]
  assign c53_183_io_in_4 = c53_177_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_184_io_in_0 = pp_16[24]; // @[Multiplier.scala 60:38]
  assign c53_184_io_in_1 = pp_17[22]; // @[Multiplier.scala 60:38]
  assign c53_184_io_in_2 = pp_18[20]; // @[Multiplier.scala 60:38]
  assign c53_184_io_in_3 = pp_19[18]; // @[Multiplier.scala 60:38]
  assign c53_184_io_in_4 = c53_178_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_185_io_in_0 = pp_20[16]; // @[Multiplier.scala 60:38]
  assign c53_185_io_in_1 = pp_21[14]; // @[Multiplier.scala 60:38]
  assign c53_185_io_in_2 = pp_22[12]; // @[Multiplier.scala 60:38]
  assign c53_185_io_in_3 = pp_23[10]; // @[Multiplier.scala 60:38]
  assign c53_185_io_in_4 = c53_179_io_out_1; // @[Multiplier.scala 89:41]
  assign c32_16_io_in_0 = pp_24[8]; // @[Multiplier.scala 60:38]
  assign c32_16_io_in_1 = pp_25[6]; // @[Multiplier.scala 60:38]
  assign c32_16_io_in_2 = pp_26[4]; // @[Multiplier.scala 60:38]
  assign c53_186_io_in_0 = pp[55]; // @[Multiplier.scala 60:38]
  assign c53_186_io_in_1 = pp_1[55]; // @[Multiplier.scala 60:38]
  assign c53_186_io_in_2 = pp_2[53]; // @[Multiplier.scala 60:38]
  assign c53_186_io_in_3 = pp_3[51]; // @[Multiplier.scala 60:38]
  assign c53_186_io_in_4 = c53_180_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_187_io_in_0 = pp_4[49]; // @[Multiplier.scala 60:38]
  assign c53_187_io_in_1 = pp_5[47]; // @[Multiplier.scala 60:38]
  assign c53_187_io_in_2 = pp_6[45]; // @[Multiplier.scala 60:38]
  assign c53_187_io_in_3 = pp_7[43]; // @[Multiplier.scala 60:38]
  assign c53_187_io_in_4 = c53_181_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_188_io_in_0 = pp_8[41]; // @[Multiplier.scala 60:38]
  assign c53_188_io_in_1 = pp_9[39]; // @[Multiplier.scala 60:38]
  assign c53_188_io_in_2 = pp_10[37]; // @[Multiplier.scala 60:38]
  assign c53_188_io_in_3 = pp_11[35]; // @[Multiplier.scala 60:38]
  assign c53_188_io_in_4 = c53_182_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_189_io_in_0 = pp_12[33]; // @[Multiplier.scala 60:38]
  assign c53_189_io_in_1 = pp_13[31]; // @[Multiplier.scala 60:38]
  assign c53_189_io_in_2 = pp_14[29]; // @[Multiplier.scala 60:38]
  assign c53_189_io_in_3 = pp_15[27]; // @[Multiplier.scala 60:38]
  assign c53_189_io_in_4 = c53_183_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_190_io_in_0 = pp_16[25]; // @[Multiplier.scala 60:38]
  assign c53_190_io_in_1 = pp_17[23]; // @[Multiplier.scala 60:38]
  assign c53_190_io_in_2 = pp_18[21]; // @[Multiplier.scala 60:38]
  assign c53_190_io_in_3 = pp_19[19]; // @[Multiplier.scala 60:38]
  assign c53_190_io_in_4 = c53_184_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_191_io_in_0 = pp_20[17]; // @[Multiplier.scala 60:38]
  assign c53_191_io_in_1 = pp_21[15]; // @[Multiplier.scala 60:38]
  assign c53_191_io_in_2 = pp_22[13]; // @[Multiplier.scala 60:38]
  assign c53_191_io_in_3 = pp_23[11]; // @[Multiplier.scala 60:38]
  assign c53_191_io_in_4 = c53_185_io_out_1; // @[Multiplier.scala 89:41]
  assign c32_17_io_in_0 = pp_24[9]; // @[Multiplier.scala 60:38]
  assign c32_17_io_in_1 = pp_25[7]; // @[Multiplier.scala 60:38]
  assign c32_17_io_in_2 = pp_26[5]; // @[Multiplier.scala 60:38]
  assign c53_192_io_in_0 = pp[56]; // @[Multiplier.scala 60:38]
  assign c53_192_io_in_1 = pp_1[56]; // @[Multiplier.scala 60:38]
  assign c53_192_io_in_2 = pp_2[54]; // @[Multiplier.scala 60:38]
  assign c53_192_io_in_3 = pp_3[52]; // @[Multiplier.scala 60:38]
  assign c53_192_io_in_4 = c53_186_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_193_io_in_0 = pp_4[50]; // @[Multiplier.scala 60:38]
  assign c53_193_io_in_1 = pp_5[48]; // @[Multiplier.scala 60:38]
  assign c53_193_io_in_2 = pp_6[46]; // @[Multiplier.scala 60:38]
  assign c53_193_io_in_3 = pp_7[44]; // @[Multiplier.scala 60:38]
  assign c53_193_io_in_4 = c53_187_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_194_io_in_0 = pp_8[42]; // @[Multiplier.scala 60:38]
  assign c53_194_io_in_1 = pp_9[40]; // @[Multiplier.scala 60:38]
  assign c53_194_io_in_2 = pp_10[38]; // @[Multiplier.scala 60:38]
  assign c53_194_io_in_3 = pp_11[36]; // @[Multiplier.scala 60:38]
  assign c53_194_io_in_4 = c53_188_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_195_io_in_0 = pp_12[34]; // @[Multiplier.scala 60:38]
  assign c53_195_io_in_1 = pp_13[32]; // @[Multiplier.scala 60:38]
  assign c53_195_io_in_2 = pp_14[30]; // @[Multiplier.scala 60:38]
  assign c53_195_io_in_3 = pp_15[28]; // @[Multiplier.scala 60:38]
  assign c53_195_io_in_4 = c53_189_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_196_io_in_0 = pp_16[26]; // @[Multiplier.scala 60:38]
  assign c53_196_io_in_1 = pp_17[24]; // @[Multiplier.scala 60:38]
  assign c53_196_io_in_2 = pp_18[22]; // @[Multiplier.scala 60:38]
  assign c53_196_io_in_3 = pp_19[20]; // @[Multiplier.scala 60:38]
  assign c53_196_io_in_4 = c53_190_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_197_io_in_0 = pp_20[18]; // @[Multiplier.scala 60:38]
  assign c53_197_io_in_1 = pp_21[16]; // @[Multiplier.scala 60:38]
  assign c53_197_io_in_2 = pp_22[14]; // @[Multiplier.scala 60:38]
  assign c53_197_io_in_3 = pp_23[12]; // @[Multiplier.scala 60:38]
  assign c53_197_io_in_4 = c53_191_io_out_1; // @[Multiplier.scala 89:41]
  assign c32_18_io_in_0 = pp_24[10]; // @[Multiplier.scala 60:38]
  assign c32_18_io_in_1 = pp_25[8]; // @[Multiplier.scala 60:38]
  assign c32_18_io_in_2 = pp_26[6]; // @[Multiplier.scala 60:38]
  assign c53_198_io_in_0 = pp[57]; // @[Multiplier.scala 60:38]
  assign c53_198_io_in_1 = pp_1[57]; // @[Multiplier.scala 60:38]
  assign c53_198_io_in_2 = pp_2[55]; // @[Multiplier.scala 60:38]
  assign c53_198_io_in_3 = pp_3[53]; // @[Multiplier.scala 60:38]
  assign c53_198_io_in_4 = c53_192_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_199_io_in_0 = pp_4[51]; // @[Multiplier.scala 60:38]
  assign c53_199_io_in_1 = pp_5[49]; // @[Multiplier.scala 60:38]
  assign c53_199_io_in_2 = pp_6[47]; // @[Multiplier.scala 60:38]
  assign c53_199_io_in_3 = pp_7[45]; // @[Multiplier.scala 60:38]
  assign c53_199_io_in_4 = c53_193_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_200_io_in_0 = pp_8[43]; // @[Multiplier.scala 60:38]
  assign c53_200_io_in_1 = pp_9[41]; // @[Multiplier.scala 60:38]
  assign c53_200_io_in_2 = pp_10[39]; // @[Multiplier.scala 60:38]
  assign c53_200_io_in_3 = pp_11[37]; // @[Multiplier.scala 60:38]
  assign c53_200_io_in_4 = c53_194_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_201_io_in_0 = pp_12[35]; // @[Multiplier.scala 60:38]
  assign c53_201_io_in_1 = pp_13[33]; // @[Multiplier.scala 60:38]
  assign c53_201_io_in_2 = pp_14[31]; // @[Multiplier.scala 60:38]
  assign c53_201_io_in_3 = pp_15[29]; // @[Multiplier.scala 60:38]
  assign c53_201_io_in_4 = c53_195_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_202_io_in_0 = pp_16[27]; // @[Multiplier.scala 60:38]
  assign c53_202_io_in_1 = pp_17[25]; // @[Multiplier.scala 60:38]
  assign c53_202_io_in_2 = pp_18[23]; // @[Multiplier.scala 60:38]
  assign c53_202_io_in_3 = pp_19[21]; // @[Multiplier.scala 60:38]
  assign c53_202_io_in_4 = c53_196_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_203_io_in_0 = pp_20[19]; // @[Multiplier.scala 60:38]
  assign c53_203_io_in_1 = pp_21[17]; // @[Multiplier.scala 60:38]
  assign c53_203_io_in_2 = pp_22[15]; // @[Multiplier.scala 60:38]
  assign c53_203_io_in_3 = pp_23[13]; // @[Multiplier.scala 60:38]
  assign c53_203_io_in_4 = c53_197_io_out_1; // @[Multiplier.scala 89:41]
  assign c32_19_io_in_0 = pp_24[11]; // @[Multiplier.scala 60:38]
  assign c32_19_io_in_1 = pp_25[9]; // @[Multiplier.scala 60:38]
  assign c32_19_io_in_2 = pp_26[7]; // @[Multiplier.scala 60:38]
  assign c53_204_io_in_0 = pp_1[58]; // @[Multiplier.scala 60:38]
  assign c53_204_io_in_1 = pp_2[56]; // @[Multiplier.scala 60:38]
  assign c53_204_io_in_2 = pp_3[54]; // @[Multiplier.scala 60:38]
  assign c53_204_io_in_3 = pp_4[52]; // @[Multiplier.scala 60:38]
  assign c53_204_io_in_4 = c53_198_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_205_io_in_0 = pp_5[50]; // @[Multiplier.scala 60:38]
  assign c53_205_io_in_1 = pp_6[48]; // @[Multiplier.scala 60:38]
  assign c53_205_io_in_2 = pp_7[46]; // @[Multiplier.scala 60:38]
  assign c53_205_io_in_3 = pp_8[44]; // @[Multiplier.scala 60:38]
  assign c53_205_io_in_4 = c53_199_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_206_io_in_0 = pp_9[42]; // @[Multiplier.scala 60:38]
  assign c53_206_io_in_1 = pp_10[40]; // @[Multiplier.scala 60:38]
  assign c53_206_io_in_2 = pp_11[38]; // @[Multiplier.scala 60:38]
  assign c53_206_io_in_3 = pp_12[36]; // @[Multiplier.scala 60:38]
  assign c53_206_io_in_4 = c53_200_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_207_io_in_0 = pp_13[34]; // @[Multiplier.scala 60:38]
  assign c53_207_io_in_1 = pp_14[32]; // @[Multiplier.scala 60:38]
  assign c53_207_io_in_2 = pp_15[30]; // @[Multiplier.scala 60:38]
  assign c53_207_io_in_3 = pp_16[28]; // @[Multiplier.scala 60:38]
  assign c53_207_io_in_4 = c53_201_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_208_io_in_0 = pp_17[26]; // @[Multiplier.scala 60:38]
  assign c53_208_io_in_1 = pp_18[24]; // @[Multiplier.scala 60:38]
  assign c53_208_io_in_2 = pp_19[22]; // @[Multiplier.scala 60:38]
  assign c53_208_io_in_3 = pp_20[20]; // @[Multiplier.scala 60:38]
  assign c53_208_io_in_4 = c53_202_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_209_io_in_0 = pp_21[18]; // @[Multiplier.scala 60:38]
  assign c53_209_io_in_1 = pp_22[16]; // @[Multiplier.scala 60:38]
  assign c53_209_io_in_2 = pp_23[14]; // @[Multiplier.scala 60:38]
  assign c53_209_io_in_3 = pp_24[12]; // @[Multiplier.scala 60:38]
  assign c53_209_io_in_4 = c53_203_io_out_1; // @[Multiplier.scala 89:41]
  assign c22_14_io_in_0 = pp_25[10]; // @[Multiplier.scala 60:38]
  assign c22_14_io_in_1 = pp_26[8]; // @[Multiplier.scala 60:38]
  assign c53_210_io_in_0 = pp_2[57]; // @[Multiplier.scala 60:38]
  assign c53_210_io_in_1 = pp_3[55]; // @[Multiplier.scala 60:38]
  assign c53_210_io_in_2 = pp_4[53]; // @[Multiplier.scala 60:38]
  assign c53_210_io_in_3 = pp_5[51]; // @[Multiplier.scala 60:38]
  assign c53_210_io_in_4 = c53_204_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_211_io_in_0 = pp_6[49]; // @[Multiplier.scala 60:38]
  assign c53_211_io_in_1 = pp_7[47]; // @[Multiplier.scala 60:38]
  assign c53_211_io_in_2 = pp_8[45]; // @[Multiplier.scala 60:38]
  assign c53_211_io_in_3 = pp_9[43]; // @[Multiplier.scala 60:38]
  assign c53_211_io_in_4 = c53_205_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_212_io_in_0 = pp_10[41]; // @[Multiplier.scala 60:38]
  assign c53_212_io_in_1 = pp_11[39]; // @[Multiplier.scala 60:38]
  assign c53_212_io_in_2 = pp_12[37]; // @[Multiplier.scala 60:38]
  assign c53_212_io_in_3 = pp_13[35]; // @[Multiplier.scala 60:38]
  assign c53_212_io_in_4 = c53_206_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_213_io_in_0 = pp_14[33]; // @[Multiplier.scala 60:38]
  assign c53_213_io_in_1 = pp_15[31]; // @[Multiplier.scala 60:38]
  assign c53_213_io_in_2 = pp_16[29]; // @[Multiplier.scala 60:38]
  assign c53_213_io_in_3 = pp_17[27]; // @[Multiplier.scala 60:38]
  assign c53_213_io_in_4 = c53_207_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_214_io_in_0 = pp_18[25]; // @[Multiplier.scala 60:38]
  assign c53_214_io_in_1 = pp_19[23]; // @[Multiplier.scala 60:38]
  assign c53_214_io_in_2 = pp_20[21]; // @[Multiplier.scala 60:38]
  assign c53_214_io_in_3 = pp_21[19]; // @[Multiplier.scala 60:38]
  assign c53_214_io_in_4 = c53_208_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_215_io_in_0 = pp_22[17]; // @[Multiplier.scala 60:38]
  assign c53_215_io_in_1 = pp_23[15]; // @[Multiplier.scala 60:38]
  assign c53_215_io_in_2 = pp_24[13]; // @[Multiplier.scala 60:38]
  assign c53_215_io_in_3 = pp_25[11]; // @[Multiplier.scala 60:38]
  assign c53_215_io_in_4 = c53_209_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_216_io_in_0 = pp_2[58]; // @[Multiplier.scala 60:38]
  assign c53_216_io_in_1 = pp_3[56]; // @[Multiplier.scala 60:38]
  assign c53_216_io_in_2 = pp_4[54]; // @[Multiplier.scala 60:38]
  assign c53_216_io_in_3 = pp_5[52]; // @[Multiplier.scala 60:38]
  assign c53_216_io_in_4 = c53_210_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_217_io_in_0 = pp_6[50]; // @[Multiplier.scala 60:38]
  assign c53_217_io_in_1 = pp_7[48]; // @[Multiplier.scala 60:38]
  assign c53_217_io_in_2 = pp_8[46]; // @[Multiplier.scala 60:38]
  assign c53_217_io_in_3 = pp_9[44]; // @[Multiplier.scala 60:38]
  assign c53_217_io_in_4 = c53_211_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_218_io_in_0 = pp_10[42]; // @[Multiplier.scala 60:38]
  assign c53_218_io_in_1 = pp_11[40]; // @[Multiplier.scala 60:38]
  assign c53_218_io_in_2 = pp_12[38]; // @[Multiplier.scala 60:38]
  assign c53_218_io_in_3 = pp_13[36]; // @[Multiplier.scala 60:38]
  assign c53_218_io_in_4 = c53_212_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_219_io_in_0 = pp_14[34]; // @[Multiplier.scala 60:38]
  assign c53_219_io_in_1 = pp_15[32]; // @[Multiplier.scala 60:38]
  assign c53_219_io_in_2 = pp_16[30]; // @[Multiplier.scala 60:38]
  assign c53_219_io_in_3 = pp_17[28]; // @[Multiplier.scala 60:38]
  assign c53_219_io_in_4 = c53_213_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_220_io_in_0 = pp_18[26]; // @[Multiplier.scala 60:38]
  assign c53_220_io_in_1 = pp_19[24]; // @[Multiplier.scala 60:38]
  assign c53_220_io_in_2 = pp_20[22]; // @[Multiplier.scala 60:38]
  assign c53_220_io_in_3 = pp_21[20]; // @[Multiplier.scala 60:38]
  assign c53_220_io_in_4 = c53_214_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_221_io_in_0 = pp_22[18]; // @[Multiplier.scala 60:38]
  assign c53_221_io_in_1 = pp_23[16]; // @[Multiplier.scala 60:38]
  assign c53_221_io_in_2 = pp_24[14]; // @[Multiplier.scala 60:38]
  assign c53_221_io_in_3 = pp_25[12]; // @[Multiplier.scala 60:38]
  assign c53_221_io_in_4 = c53_215_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_222_io_in_0 = pp_3[57]; // @[Multiplier.scala 60:38]
  assign c53_222_io_in_1 = pp_4[55]; // @[Multiplier.scala 60:38]
  assign c53_222_io_in_2 = pp_5[53]; // @[Multiplier.scala 60:38]
  assign c53_222_io_in_3 = pp_6[51]; // @[Multiplier.scala 60:38]
  assign c53_222_io_in_4 = c53_216_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_223_io_in_0 = pp_7[49]; // @[Multiplier.scala 60:38]
  assign c53_223_io_in_1 = pp_8[47]; // @[Multiplier.scala 60:38]
  assign c53_223_io_in_2 = pp_9[45]; // @[Multiplier.scala 60:38]
  assign c53_223_io_in_3 = pp_10[43]; // @[Multiplier.scala 60:38]
  assign c53_223_io_in_4 = c53_217_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_224_io_in_0 = pp_11[41]; // @[Multiplier.scala 60:38]
  assign c53_224_io_in_1 = pp_12[39]; // @[Multiplier.scala 60:38]
  assign c53_224_io_in_2 = pp_13[37]; // @[Multiplier.scala 60:38]
  assign c53_224_io_in_3 = pp_14[35]; // @[Multiplier.scala 60:38]
  assign c53_224_io_in_4 = c53_218_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_225_io_in_0 = pp_15[33]; // @[Multiplier.scala 60:38]
  assign c53_225_io_in_1 = pp_16[31]; // @[Multiplier.scala 60:38]
  assign c53_225_io_in_2 = pp_17[29]; // @[Multiplier.scala 60:38]
  assign c53_225_io_in_3 = pp_18[27]; // @[Multiplier.scala 60:38]
  assign c53_225_io_in_4 = c53_219_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_226_io_in_0 = pp_19[25]; // @[Multiplier.scala 60:38]
  assign c53_226_io_in_1 = pp_20[23]; // @[Multiplier.scala 60:38]
  assign c53_226_io_in_2 = pp_21[21]; // @[Multiplier.scala 60:38]
  assign c53_226_io_in_3 = pp_22[19]; // @[Multiplier.scala 60:38]
  assign c53_226_io_in_4 = c53_220_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_227_io_in_0 = pp_23[17]; // @[Multiplier.scala 60:38]
  assign c53_227_io_in_1 = pp_24[15]; // @[Multiplier.scala 60:38]
  assign c53_227_io_in_2 = pp_25[13]; // @[Multiplier.scala 60:38]
  assign c53_227_io_in_3 = pp_26[11]; // @[Multiplier.scala 60:38]
  assign c53_227_io_in_4 = c53_221_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_228_io_in_0 = pp_3[58]; // @[Multiplier.scala 60:38]
  assign c53_228_io_in_1 = pp_4[56]; // @[Multiplier.scala 60:38]
  assign c53_228_io_in_2 = pp_5[54]; // @[Multiplier.scala 60:38]
  assign c53_228_io_in_3 = pp_6[52]; // @[Multiplier.scala 60:38]
  assign c53_228_io_in_4 = c53_222_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_229_io_in_0 = pp_7[50]; // @[Multiplier.scala 60:38]
  assign c53_229_io_in_1 = pp_8[48]; // @[Multiplier.scala 60:38]
  assign c53_229_io_in_2 = pp_9[46]; // @[Multiplier.scala 60:38]
  assign c53_229_io_in_3 = pp_10[44]; // @[Multiplier.scala 60:38]
  assign c53_229_io_in_4 = c53_223_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_230_io_in_0 = pp_11[42]; // @[Multiplier.scala 60:38]
  assign c53_230_io_in_1 = pp_12[40]; // @[Multiplier.scala 60:38]
  assign c53_230_io_in_2 = pp_13[38]; // @[Multiplier.scala 60:38]
  assign c53_230_io_in_3 = pp_14[36]; // @[Multiplier.scala 60:38]
  assign c53_230_io_in_4 = c53_224_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_231_io_in_0 = pp_15[34]; // @[Multiplier.scala 60:38]
  assign c53_231_io_in_1 = pp_16[32]; // @[Multiplier.scala 60:38]
  assign c53_231_io_in_2 = pp_17[30]; // @[Multiplier.scala 60:38]
  assign c53_231_io_in_3 = pp_18[28]; // @[Multiplier.scala 60:38]
  assign c53_231_io_in_4 = c53_225_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_232_io_in_0 = pp_19[26]; // @[Multiplier.scala 60:38]
  assign c53_232_io_in_1 = pp_20[24]; // @[Multiplier.scala 60:38]
  assign c53_232_io_in_2 = pp_21[22]; // @[Multiplier.scala 60:38]
  assign c53_232_io_in_3 = pp_22[20]; // @[Multiplier.scala 60:38]
  assign c53_232_io_in_4 = c53_226_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_233_io_in_0 = pp_23[18]; // @[Multiplier.scala 60:38]
  assign c53_233_io_in_1 = pp_24[16]; // @[Multiplier.scala 60:38]
  assign c53_233_io_in_2 = pp_25[14]; // @[Multiplier.scala 60:38]
  assign c53_233_io_in_3 = pp_26[12]; // @[Multiplier.scala 60:38]
  assign c53_233_io_in_4 = c53_227_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_234_io_in_0 = pp_4[57]; // @[Multiplier.scala 60:38]
  assign c53_234_io_in_1 = pp_5[55]; // @[Multiplier.scala 60:38]
  assign c53_234_io_in_2 = pp_6[53]; // @[Multiplier.scala 60:38]
  assign c53_234_io_in_3 = pp_7[51]; // @[Multiplier.scala 60:38]
  assign c53_234_io_in_4 = c53_228_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_235_io_in_0 = pp_8[49]; // @[Multiplier.scala 60:38]
  assign c53_235_io_in_1 = pp_9[47]; // @[Multiplier.scala 60:38]
  assign c53_235_io_in_2 = pp_10[45]; // @[Multiplier.scala 60:38]
  assign c53_235_io_in_3 = pp_11[43]; // @[Multiplier.scala 60:38]
  assign c53_235_io_in_4 = c53_229_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_236_io_in_0 = pp_12[41]; // @[Multiplier.scala 60:38]
  assign c53_236_io_in_1 = pp_13[39]; // @[Multiplier.scala 60:38]
  assign c53_236_io_in_2 = pp_14[37]; // @[Multiplier.scala 60:38]
  assign c53_236_io_in_3 = pp_15[35]; // @[Multiplier.scala 60:38]
  assign c53_236_io_in_4 = c53_230_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_237_io_in_0 = pp_16[33]; // @[Multiplier.scala 60:38]
  assign c53_237_io_in_1 = pp_17[31]; // @[Multiplier.scala 60:38]
  assign c53_237_io_in_2 = pp_18[29]; // @[Multiplier.scala 60:38]
  assign c53_237_io_in_3 = pp_19[27]; // @[Multiplier.scala 60:38]
  assign c53_237_io_in_4 = c53_231_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_238_io_in_0 = pp_20[25]; // @[Multiplier.scala 60:38]
  assign c53_238_io_in_1 = pp_21[23]; // @[Multiplier.scala 60:38]
  assign c53_238_io_in_2 = pp_22[21]; // @[Multiplier.scala 60:38]
  assign c53_238_io_in_3 = pp_23[19]; // @[Multiplier.scala 60:38]
  assign c53_238_io_in_4 = c53_232_io_out_1; // @[Multiplier.scala 89:41]
  assign c32_20_io_in_0 = pp_24[17]; // @[Multiplier.scala 60:38]
  assign c32_20_io_in_1 = pp_25[15]; // @[Multiplier.scala 60:38]
  assign c32_20_io_in_2 = pp_26[13]; // @[Multiplier.scala 60:38]
  assign c53_239_io_in_0 = pp_4[58]; // @[Multiplier.scala 60:38]
  assign c53_239_io_in_1 = pp_5[56]; // @[Multiplier.scala 60:38]
  assign c53_239_io_in_2 = pp_6[54]; // @[Multiplier.scala 60:38]
  assign c53_239_io_in_3 = pp_7[52]; // @[Multiplier.scala 60:38]
  assign c53_239_io_in_4 = c53_234_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_240_io_in_0 = pp_8[50]; // @[Multiplier.scala 60:38]
  assign c53_240_io_in_1 = pp_9[48]; // @[Multiplier.scala 60:38]
  assign c53_240_io_in_2 = pp_10[46]; // @[Multiplier.scala 60:38]
  assign c53_240_io_in_3 = pp_11[44]; // @[Multiplier.scala 60:38]
  assign c53_240_io_in_4 = c53_235_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_241_io_in_0 = pp_12[42]; // @[Multiplier.scala 60:38]
  assign c53_241_io_in_1 = pp_13[40]; // @[Multiplier.scala 60:38]
  assign c53_241_io_in_2 = pp_14[38]; // @[Multiplier.scala 60:38]
  assign c53_241_io_in_3 = pp_15[36]; // @[Multiplier.scala 60:38]
  assign c53_241_io_in_4 = c53_236_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_242_io_in_0 = pp_16[34]; // @[Multiplier.scala 60:38]
  assign c53_242_io_in_1 = pp_17[32]; // @[Multiplier.scala 60:38]
  assign c53_242_io_in_2 = pp_18[30]; // @[Multiplier.scala 60:38]
  assign c53_242_io_in_3 = pp_19[28]; // @[Multiplier.scala 60:38]
  assign c53_242_io_in_4 = c53_237_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_243_io_in_0 = pp_20[26]; // @[Multiplier.scala 60:38]
  assign c53_243_io_in_1 = pp_21[24]; // @[Multiplier.scala 60:38]
  assign c53_243_io_in_2 = pp_22[22]; // @[Multiplier.scala 60:38]
  assign c53_243_io_in_3 = pp_23[20]; // @[Multiplier.scala 60:38]
  assign c53_243_io_in_4 = c53_238_io_out_1; // @[Multiplier.scala 89:41]
  assign c32_21_io_in_0 = pp_24[18]; // @[Multiplier.scala 60:38]
  assign c32_21_io_in_1 = pp_25[16]; // @[Multiplier.scala 60:38]
  assign c32_21_io_in_2 = pp_26[14]; // @[Multiplier.scala 60:38]
  assign c53_244_io_in_0 = pp_5[57]; // @[Multiplier.scala 60:38]
  assign c53_244_io_in_1 = pp_6[55]; // @[Multiplier.scala 60:38]
  assign c53_244_io_in_2 = pp_7[53]; // @[Multiplier.scala 60:38]
  assign c53_244_io_in_3 = pp_8[51]; // @[Multiplier.scala 60:38]
  assign c53_244_io_in_4 = c53_239_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_245_io_in_0 = pp_9[49]; // @[Multiplier.scala 60:38]
  assign c53_245_io_in_1 = pp_10[47]; // @[Multiplier.scala 60:38]
  assign c53_245_io_in_2 = pp_11[45]; // @[Multiplier.scala 60:38]
  assign c53_245_io_in_3 = pp_12[43]; // @[Multiplier.scala 60:38]
  assign c53_245_io_in_4 = c53_240_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_246_io_in_0 = pp_13[41]; // @[Multiplier.scala 60:38]
  assign c53_246_io_in_1 = pp_14[39]; // @[Multiplier.scala 60:38]
  assign c53_246_io_in_2 = pp_15[37]; // @[Multiplier.scala 60:38]
  assign c53_246_io_in_3 = pp_16[35]; // @[Multiplier.scala 60:38]
  assign c53_246_io_in_4 = c53_241_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_247_io_in_0 = pp_17[33]; // @[Multiplier.scala 60:38]
  assign c53_247_io_in_1 = pp_18[31]; // @[Multiplier.scala 60:38]
  assign c53_247_io_in_2 = pp_19[29]; // @[Multiplier.scala 60:38]
  assign c53_247_io_in_3 = pp_20[27]; // @[Multiplier.scala 60:38]
  assign c53_247_io_in_4 = c53_242_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_248_io_in_0 = pp_21[25]; // @[Multiplier.scala 60:38]
  assign c53_248_io_in_1 = pp_22[23]; // @[Multiplier.scala 60:38]
  assign c53_248_io_in_2 = pp_23[21]; // @[Multiplier.scala 60:38]
  assign c53_248_io_in_3 = pp_24[19]; // @[Multiplier.scala 60:38]
  assign c53_248_io_in_4 = c53_243_io_out_1; // @[Multiplier.scala 89:41]
  assign c22_15_io_in_0 = pp_25[17]; // @[Multiplier.scala 60:38]
  assign c22_15_io_in_1 = pp_26[15]; // @[Multiplier.scala 60:38]
  assign c53_249_io_in_0 = pp_5[58]; // @[Multiplier.scala 60:38]
  assign c53_249_io_in_1 = pp_6[56]; // @[Multiplier.scala 60:38]
  assign c53_249_io_in_2 = pp_7[54]; // @[Multiplier.scala 60:38]
  assign c53_249_io_in_3 = pp_8[52]; // @[Multiplier.scala 60:38]
  assign c53_249_io_in_4 = c53_244_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_250_io_in_0 = pp_9[50]; // @[Multiplier.scala 60:38]
  assign c53_250_io_in_1 = pp_10[48]; // @[Multiplier.scala 60:38]
  assign c53_250_io_in_2 = pp_11[46]; // @[Multiplier.scala 60:38]
  assign c53_250_io_in_3 = pp_12[44]; // @[Multiplier.scala 60:38]
  assign c53_250_io_in_4 = c53_245_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_251_io_in_0 = pp_13[42]; // @[Multiplier.scala 60:38]
  assign c53_251_io_in_1 = pp_14[40]; // @[Multiplier.scala 60:38]
  assign c53_251_io_in_2 = pp_15[38]; // @[Multiplier.scala 60:38]
  assign c53_251_io_in_3 = pp_16[36]; // @[Multiplier.scala 60:38]
  assign c53_251_io_in_4 = c53_246_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_252_io_in_0 = pp_17[34]; // @[Multiplier.scala 60:38]
  assign c53_252_io_in_1 = pp_18[32]; // @[Multiplier.scala 60:38]
  assign c53_252_io_in_2 = pp_19[30]; // @[Multiplier.scala 60:38]
  assign c53_252_io_in_3 = pp_20[28]; // @[Multiplier.scala 60:38]
  assign c53_252_io_in_4 = c53_247_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_253_io_in_0 = pp_21[26]; // @[Multiplier.scala 60:38]
  assign c53_253_io_in_1 = pp_22[24]; // @[Multiplier.scala 60:38]
  assign c53_253_io_in_2 = pp_23[22]; // @[Multiplier.scala 60:38]
  assign c53_253_io_in_3 = pp_24[20]; // @[Multiplier.scala 60:38]
  assign c53_253_io_in_4 = c53_248_io_out_1; // @[Multiplier.scala 89:41]
  assign c22_16_io_in_0 = pp_25[18]; // @[Multiplier.scala 60:38]
  assign c22_16_io_in_1 = pp_26[16]; // @[Multiplier.scala 60:38]
  assign c53_254_io_in_0 = pp_6[57]; // @[Multiplier.scala 60:38]
  assign c53_254_io_in_1 = pp_7[55]; // @[Multiplier.scala 60:38]
  assign c53_254_io_in_2 = pp_8[53]; // @[Multiplier.scala 60:38]
  assign c53_254_io_in_3 = pp_9[51]; // @[Multiplier.scala 60:38]
  assign c53_254_io_in_4 = c53_249_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_255_io_in_0 = pp_10[49]; // @[Multiplier.scala 60:38]
  assign c53_255_io_in_1 = pp_11[47]; // @[Multiplier.scala 60:38]
  assign c53_255_io_in_2 = pp_12[45]; // @[Multiplier.scala 60:38]
  assign c53_255_io_in_3 = pp_13[43]; // @[Multiplier.scala 60:38]
  assign c53_255_io_in_4 = c53_250_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_256_io_in_0 = pp_14[41]; // @[Multiplier.scala 60:38]
  assign c53_256_io_in_1 = pp_15[39]; // @[Multiplier.scala 60:38]
  assign c53_256_io_in_2 = pp_16[37]; // @[Multiplier.scala 60:38]
  assign c53_256_io_in_3 = pp_17[35]; // @[Multiplier.scala 60:38]
  assign c53_256_io_in_4 = c53_251_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_257_io_in_0 = pp_18[33]; // @[Multiplier.scala 60:38]
  assign c53_257_io_in_1 = pp_19[31]; // @[Multiplier.scala 60:38]
  assign c53_257_io_in_2 = pp_20[29]; // @[Multiplier.scala 60:38]
  assign c53_257_io_in_3 = pp_21[27]; // @[Multiplier.scala 60:38]
  assign c53_257_io_in_4 = c53_252_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_258_io_in_0 = pp_22[25]; // @[Multiplier.scala 60:38]
  assign c53_258_io_in_1 = pp_23[23]; // @[Multiplier.scala 60:38]
  assign c53_258_io_in_2 = pp_24[21]; // @[Multiplier.scala 60:38]
  assign c53_258_io_in_3 = pp_25[19]; // @[Multiplier.scala 60:38]
  assign c53_258_io_in_4 = c53_253_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_259_io_in_0 = pp_6[58]; // @[Multiplier.scala 60:38]
  assign c53_259_io_in_1 = pp_7[56]; // @[Multiplier.scala 60:38]
  assign c53_259_io_in_2 = pp_8[54]; // @[Multiplier.scala 60:38]
  assign c53_259_io_in_3 = pp_9[52]; // @[Multiplier.scala 60:38]
  assign c53_259_io_in_4 = c53_254_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_260_io_in_0 = pp_10[50]; // @[Multiplier.scala 60:38]
  assign c53_260_io_in_1 = pp_11[48]; // @[Multiplier.scala 60:38]
  assign c53_260_io_in_2 = pp_12[46]; // @[Multiplier.scala 60:38]
  assign c53_260_io_in_3 = pp_13[44]; // @[Multiplier.scala 60:38]
  assign c53_260_io_in_4 = c53_255_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_261_io_in_0 = pp_14[42]; // @[Multiplier.scala 60:38]
  assign c53_261_io_in_1 = pp_15[40]; // @[Multiplier.scala 60:38]
  assign c53_261_io_in_2 = pp_16[38]; // @[Multiplier.scala 60:38]
  assign c53_261_io_in_3 = pp_17[36]; // @[Multiplier.scala 60:38]
  assign c53_261_io_in_4 = c53_256_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_262_io_in_0 = pp_18[34]; // @[Multiplier.scala 60:38]
  assign c53_262_io_in_1 = pp_19[32]; // @[Multiplier.scala 60:38]
  assign c53_262_io_in_2 = pp_20[30]; // @[Multiplier.scala 60:38]
  assign c53_262_io_in_3 = pp_21[28]; // @[Multiplier.scala 60:38]
  assign c53_262_io_in_4 = c53_257_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_263_io_in_0 = pp_22[26]; // @[Multiplier.scala 60:38]
  assign c53_263_io_in_1 = pp_23[24]; // @[Multiplier.scala 60:38]
  assign c53_263_io_in_2 = pp_24[22]; // @[Multiplier.scala 60:38]
  assign c53_263_io_in_3 = pp_25[20]; // @[Multiplier.scala 60:38]
  assign c53_263_io_in_4 = c53_258_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_264_io_in_0 = pp_7[57]; // @[Multiplier.scala 60:38]
  assign c53_264_io_in_1 = pp_8[55]; // @[Multiplier.scala 60:38]
  assign c53_264_io_in_2 = pp_9[53]; // @[Multiplier.scala 60:38]
  assign c53_264_io_in_3 = pp_10[51]; // @[Multiplier.scala 60:38]
  assign c53_264_io_in_4 = c53_259_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_265_io_in_0 = pp_11[49]; // @[Multiplier.scala 60:38]
  assign c53_265_io_in_1 = pp_12[47]; // @[Multiplier.scala 60:38]
  assign c53_265_io_in_2 = pp_13[45]; // @[Multiplier.scala 60:38]
  assign c53_265_io_in_3 = pp_14[43]; // @[Multiplier.scala 60:38]
  assign c53_265_io_in_4 = c53_260_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_266_io_in_0 = pp_15[41]; // @[Multiplier.scala 60:38]
  assign c53_266_io_in_1 = pp_16[39]; // @[Multiplier.scala 60:38]
  assign c53_266_io_in_2 = pp_17[37]; // @[Multiplier.scala 60:38]
  assign c53_266_io_in_3 = pp_18[35]; // @[Multiplier.scala 60:38]
  assign c53_266_io_in_4 = c53_261_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_267_io_in_0 = pp_19[33]; // @[Multiplier.scala 60:38]
  assign c53_267_io_in_1 = pp_20[31]; // @[Multiplier.scala 60:38]
  assign c53_267_io_in_2 = pp_21[29]; // @[Multiplier.scala 60:38]
  assign c53_267_io_in_3 = pp_22[27]; // @[Multiplier.scala 60:38]
  assign c53_267_io_in_4 = c53_262_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_268_io_in_0 = pp_23[25]; // @[Multiplier.scala 60:38]
  assign c53_268_io_in_1 = pp_24[23]; // @[Multiplier.scala 60:38]
  assign c53_268_io_in_2 = pp_25[21]; // @[Multiplier.scala 60:38]
  assign c53_268_io_in_3 = pp_26[19]; // @[Multiplier.scala 60:38]
  assign c53_268_io_in_4 = c53_263_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_269_io_in_0 = pp_7[58]; // @[Multiplier.scala 60:38]
  assign c53_269_io_in_1 = pp_8[56]; // @[Multiplier.scala 60:38]
  assign c53_269_io_in_2 = pp_9[54]; // @[Multiplier.scala 60:38]
  assign c53_269_io_in_3 = pp_10[52]; // @[Multiplier.scala 60:38]
  assign c53_269_io_in_4 = c53_264_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_270_io_in_0 = pp_11[50]; // @[Multiplier.scala 60:38]
  assign c53_270_io_in_1 = pp_12[48]; // @[Multiplier.scala 60:38]
  assign c53_270_io_in_2 = pp_13[46]; // @[Multiplier.scala 60:38]
  assign c53_270_io_in_3 = pp_14[44]; // @[Multiplier.scala 60:38]
  assign c53_270_io_in_4 = c53_265_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_271_io_in_0 = pp_15[42]; // @[Multiplier.scala 60:38]
  assign c53_271_io_in_1 = pp_16[40]; // @[Multiplier.scala 60:38]
  assign c53_271_io_in_2 = pp_17[38]; // @[Multiplier.scala 60:38]
  assign c53_271_io_in_3 = pp_18[36]; // @[Multiplier.scala 60:38]
  assign c53_271_io_in_4 = c53_266_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_272_io_in_0 = pp_19[34]; // @[Multiplier.scala 60:38]
  assign c53_272_io_in_1 = pp_20[32]; // @[Multiplier.scala 60:38]
  assign c53_272_io_in_2 = pp_21[30]; // @[Multiplier.scala 60:38]
  assign c53_272_io_in_3 = pp_22[28]; // @[Multiplier.scala 60:38]
  assign c53_272_io_in_4 = c53_267_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_273_io_in_0 = pp_23[26]; // @[Multiplier.scala 60:38]
  assign c53_273_io_in_1 = pp_24[24]; // @[Multiplier.scala 60:38]
  assign c53_273_io_in_2 = pp_25[22]; // @[Multiplier.scala 60:38]
  assign c53_273_io_in_3 = pp_26[20]; // @[Multiplier.scala 60:38]
  assign c53_273_io_in_4 = c53_268_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_274_io_in_0 = pp_8[57]; // @[Multiplier.scala 60:38]
  assign c53_274_io_in_1 = pp_9[55]; // @[Multiplier.scala 60:38]
  assign c53_274_io_in_2 = pp_10[53]; // @[Multiplier.scala 60:38]
  assign c53_274_io_in_3 = pp_11[51]; // @[Multiplier.scala 60:38]
  assign c53_274_io_in_4 = c53_269_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_275_io_in_0 = pp_12[49]; // @[Multiplier.scala 60:38]
  assign c53_275_io_in_1 = pp_13[47]; // @[Multiplier.scala 60:38]
  assign c53_275_io_in_2 = pp_14[45]; // @[Multiplier.scala 60:38]
  assign c53_275_io_in_3 = pp_15[43]; // @[Multiplier.scala 60:38]
  assign c53_275_io_in_4 = c53_270_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_276_io_in_0 = pp_16[41]; // @[Multiplier.scala 60:38]
  assign c53_276_io_in_1 = pp_17[39]; // @[Multiplier.scala 60:38]
  assign c53_276_io_in_2 = pp_18[37]; // @[Multiplier.scala 60:38]
  assign c53_276_io_in_3 = pp_19[35]; // @[Multiplier.scala 60:38]
  assign c53_276_io_in_4 = c53_271_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_277_io_in_0 = pp_20[33]; // @[Multiplier.scala 60:38]
  assign c53_277_io_in_1 = pp_21[31]; // @[Multiplier.scala 60:38]
  assign c53_277_io_in_2 = pp_22[29]; // @[Multiplier.scala 60:38]
  assign c53_277_io_in_3 = pp_23[27]; // @[Multiplier.scala 60:38]
  assign c53_277_io_in_4 = c53_272_io_out_1; // @[Multiplier.scala 89:41]
  assign c32_22_io_in_0 = pp_24[25]; // @[Multiplier.scala 60:38]
  assign c32_22_io_in_1 = pp_25[23]; // @[Multiplier.scala 60:38]
  assign c32_22_io_in_2 = pp_26[21]; // @[Multiplier.scala 60:38]
  assign c53_278_io_in_0 = pp_8[58]; // @[Multiplier.scala 60:38]
  assign c53_278_io_in_1 = pp_9[56]; // @[Multiplier.scala 60:38]
  assign c53_278_io_in_2 = pp_10[54]; // @[Multiplier.scala 60:38]
  assign c53_278_io_in_3 = pp_11[52]; // @[Multiplier.scala 60:38]
  assign c53_278_io_in_4 = c53_274_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_279_io_in_0 = pp_12[50]; // @[Multiplier.scala 60:38]
  assign c53_279_io_in_1 = pp_13[48]; // @[Multiplier.scala 60:38]
  assign c53_279_io_in_2 = pp_14[46]; // @[Multiplier.scala 60:38]
  assign c53_279_io_in_3 = pp_15[44]; // @[Multiplier.scala 60:38]
  assign c53_279_io_in_4 = c53_275_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_280_io_in_0 = pp_16[42]; // @[Multiplier.scala 60:38]
  assign c53_280_io_in_1 = pp_17[40]; // @[Multiplier.scala 60:38]
  assign c53_280_io_in_2 = pp_18[38]; // @[Multiplier.scala 60:38]
  assign c53_280_io_in_3 = pp_19[36]; // @[Multiplier.scala 60:38]
  assign c53_280_io_in_4 = c53_276_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_281_io_in_0 = pp_20[34]; // @[Multiplier.scala 60:38]
  assign c53_281_io_in_1 = pp_21[32]; // @[Multiplier.scala 60:38]
  assign c53_281_io_in_2 = pp_22[30]; // @[Multiplier.scala 60:38]
  assign c53_281_io_in_3 = pp_23[28]; // @[Multiplier.scala 60:38]
  assign c53_281_io_in_4 = c53_277_io_out_1; // @[Multiplier.scala 89:41]
  assign c32_23_io_in_0 = pp_24[26]; // @[Multiplier.scala 60:38]
  assign c32_23_io_in_1 = pp_25[24]; // @[Multiplier.scala 60:38]
  assign c32_23_io_in_2 = pp_26[22]; // @[Multiplier.scala 60:38]
  assign c53_282_io_in_0 = pp_9[57]; // @[Multiplier.scala 60:38]
  assign c53_282_io_in_1 = pp_10[55]; // @[Multiplier.scala 60:38]
  assign c53_282_io_in_2 = pp_11[53]; // @[Multiplier.scala 60:38]
  assign c53_282_io_in_3 = pp_12[51]; // @[Multiplier.scala 60:38]
  assign c53_282_io_in_4 = c53_278_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_283_io_in_0 = pp_13[49]; // @[Multiplier.scala 60:38]
  assign c53_283_io_in_1 = pp_14[47]; // @[Multiplier.scala 60:38]
  assign c53_283_io_in_2 = pp_15[45]; // @[Multiplier.scala 60:38]
  assign c53_283_io_in_3 = pp_16[43]; // @[Multiplier.scala 60:38]
  assign c53_283_io_in_4 = c53_279_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_284_io_in_0 = pp_17[41]; // @[Multiplier.scala 60:38]
  assign c53_284_io_in_1 = pp_18[39]; // @[Multiplier.scala 60:38]
  assign c53_284_io_in_2 = pp_19[37]; // @[Multiplier.scala 60:38]
  assign c53_284_io_in_3 = pp_20[35]; // @[Multiplier.scala 60:38]
  assign c53_284_io_in_4 = c53_280_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_285_io_in_0 = pp_21[33]; // @[Multiplier.scala 60:38]
  assign c53_285_io_in_1 = pp_22[31]; // @[Multiplier.scala 60:38]
  assign c53_285_io_in_2 = pp_23[29]; // @[Multiplier.scala 60:38]
  assign c53_285_io_in_3 = pp_24[27]; // @[Multiplier.scala 60:38]
  assign c53_285_io_in_4 = c53_281_io_out_1; // @[Multiplier.scala 89:41]
  assign c22_17_io_in_0 = pp_25[25]; // @[Multiplier.scala 60:38]
  assign c22_17_io_in_1 = pp_26[23]; // @[Multiplier.scala 60:38]
  assign c53_286_io_in_0 = pp_9[58]; // @[Multiplier.scala 60:38]
  assign c53_286_io_in_1 = pp_10[56]; // @[Multiplier.scala 60:38]
  assign c53_286_io_in_2 = pp_11[54]; // @[Multiplier.scala 60:38]
  assign c53_286_io_in_3 = pp_12[52]; // @[Multiplier.scala 60:38]
  assign c53_286_io_in_4 = c53_282_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_287_io_in_0 = pp_13[50]; // @[Multiplier.scala 60:38]
  assign c53_287_io_in_1 = pp_14[48]; // @[Multiplier.scala 60:38]
  assign c53_287_io_in_2 = pp_15[46]; // @[Multiplier.scala 60:38]
  assign c53_287_io_in_3 = pp_16[44]; // @[Multiplier.scala 60:38]
  assign c53_287_io_in_4 = c53_283_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_288_io_in_0 = pp_17[42]; // @[Multiplier.scala 60:38]
  assign c53_288_io_in_1 = pp_18[40]; // @[Multiplier.scala 60:38]
  assign c53_288_io_in_2 = pp_19[38]; // @[Multiplier.scala 60:38]
  assign c53_288_io_in_3 = pp_20[36]; // @[Multiplier.scala 60:38]
  assign c53_288_io_in_4 = c53_284_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_289_io_in_0 = pp_21[34]; // @[Multiplier.scala 60:38]
  assign c53_289_io_in_1 = pp_22[32]; // @[Multiplier.scala 60:38]
  assign c53_289_io_in_2 = pp_23[30]; // @[Multiplier.scala 60:38]
  assign c53_289_io_in_3 = pp_24[28]; // @[Multiplier.scala 60:38]
  assign c53_289_io_in_4 = c53_285_io_out_1; // @[Multiplier.scala 89:41]
  assign c22_18_io_in_0 = pp_25[26]; // @[Multiplier.scala 60:38]
  assign c22_18_io_in_1 = pp_26[24]; // @[Multiplier.scala 60:38]
  assign c53_290_io_in_0 = pp_10[57]; // @[Multiplier.scala 60:38]
  assign c53_290_io_in_1 = pp_11[55]; // @[Multiplier.scala 60:38]
  assign c53_290_io_in_2 = pp_12[53]; // @[Multiplier.scala 60:38]
  assign c53_290_io_in_3 = pp_13[51]; // @[Multiplier.scala 60:38]
  assign c53_290_io_in_4 = c53_286_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_291_io_in_0 = pp_14[49]; // @[Multiplier.scala 60:38]
  assign c53_291_io_in_1 = pp_15[47]; // @[Multiplier.scala 60:38]
  assign c53_291_io_in_2 = pp_16[45]; // @[Multiplier.scala 60:38]
  assign c53_291_io_in_3 = pp_17[43]; // @[Multiplier.scala 60:38]
  assign c53_291_io_in_4 = c53_287_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_292_io_in_0 = pp_18[41]; // @[Multiplier.scala 60:38]
  assign c53_292_io_in_1 = pp_19[39]; // @[Multiplier.scala 60:38]
  assign c53_292_io_in_2 = pp_20[37]; // @[Multiplier.scala 60:38]
  assign c53_292_io_in_3 = pp_21[35]; // @[Multiplier.scala 60:38]
  assign c53_292_io_in_4 = c53_288_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_293_io_in_0 = pp_22[33]; // @[Multiplier.scala 60:38]
  assign c53_293_io_in_1 = pp_23[31]; // @[Multiplier.scala 60:38]
  assign c53_293_io_in_2 = pp_24[29]; // @[Multiplier.scala 60:38]
  assign c53_293_io_in_3 = pp_25[27]; // @[Multiplier.scala 60:38]
  assign c53_293_io_in_4 = c53_289_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_294_io_in_0 = pp_10[58]; // @[Multiplier.scala 60:38]
  assign c53_294_io_in_1 = pp_11[56]; // @[Multiplier.scala 60:38]
  assign c53_294_io_in_2 = pp_12[54]; // @[Multiplier.scala 60:38]
  assign c53_294_io_in_3 = pp_13[52]; // @[Multiplier.scala 60:38]
  assign c53_294_io_in_4 = c53_290_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_295_io_in_0 = pp_14[50]; // @[Multiplier.scala 60:38]
  assign c53_295_io_in_1 = pp_15[48]; // @[Multiplier.scala 60:38]
  assign c53_295_io_in_2 = pp_16[46]; // @[Multiplier.scala 60:38]
  assign c53_295_io_in_3 = pp_17[44]; // @[Multiplier.scala 60:38]
  assign c53_295_io_in_4 = c53_291_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_296_io_in_0 = pp_18[42]; // @[Multiplier.scala 60:38]
  assign c53_296_io_in_1 = pp_19[40]; // @[Multiplier.scala 60:38]
  assign c53_296_io_in_2 = pp_20[38]; // @[Multiplier.scala 60:38]
  assign c53_296_io_in_3 = pp_21[36]; // @[Multiplier.scala 60:38]
  assign c53_296_io_in_4 = c53_292_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_297_io_in_0 = pp_22[34]; // @[Multiplier.scala 60:38]
  assign c53_297_io_in_1 = pp_23[32]; // @[Multiplier.scala 60:38]
  assign c53_297_io_in_2 = pp_24[30]; // @[Multiplier.scala 60:38]
  assign c53_297_io_in_3 = pp_25[28]; // @[Multiplier.scala 60:38]
  assign c53_297_io_in_4 = c53_293_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_298_io_in_0 = pp_11[57]; // @[Multiplier.scala 60:38]
  assign c53_298_io_in_1 = pp_12[55]; // @[Multiplier.scala 60:38]
  assign c53_298_io_in_2 = pp_13[53]; // @[Multiplier.scala 60:38]
  assign c53_298_io_in_3 = pp_14[51]; // @[Multiplier.scala 60:38]
  assign c53_298_io_in_4 = c53_294_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_299_io_in_0 = pp_15[49]; // @[Multiplier.scala 60:38]
  assign c53_299_io_in_1 = pp_16[47]; // @[Multiplier.scala 60:38]
  assign c53_299_io_in_2 = pp_17[45]; // @[Multiplier.scala 60:38]
  assign c53_299_io_in_3 = pp_18[43]; // @[Multiplier.scala 60:38]
  assign c53_299_io_in_4 = c53_295_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_300_io_in_0 = pp_19[41]; // @[Multiplier.scala 60:38]
  assign c53_300_io_in_1 = pp_20[39]; // @[Multiplier.scala 60:38]
  assign c53_300_io_in_2 = pp_21[37]; // @[Multiplier.scala 60:38]
  assign c53_300_io_in_3 = pp_22[35]; // @[Multiplier.scala 60:38]
  assign c53_300_io_in_4 = c53_296_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_301_io_in_0 = pp_23[33]; // @[Multiplier.scala 60:38]
  assign c53_301_io_in_1 = pp_24[31]; // @[Multiplier.scala 60:38]
  assign c53_301_io_in_2 = pp_25[29]; // @[Multiplier.scala 60:38]
  assign c53_301_io_in_3 = pp_26[27]; // @[Multiplier.scala 60:38]
  assign c53_301_io_in_4 = c53_297_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_302_io_in_0 = pp_11[58]; // @[Multiplier.scala 60:38]
  assign c53_302_io_in_1 = pp_12[56]; // @[Multiplier.scala 60:38]
  assign c53_302_io_in_2 = pp_13[54]; // @[Multiplier.scala 60:38]
  assign c53_302_io_in_3 = pp_14[52]; // @[Multiplier.scala 60:38]
  assign c53_302_io_in_4 = c53_298_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_303_io_in_0 = pp_15[50]; // @[Multiplier.scala 60:38]
  assign c53_303_io_in_1 = pp_16[48]; // @[Multiplier.scala 60:38]
  assign c53_303_io_in_2 = pp_17[46]; // @[Multiplier.scala 60:38]
  assign c53_303_io_in_3 = pp_18[44]; // @[Multiplier.scala 60:38]
  assign c53_303_io_in_4 = c53_299_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_304_io_in_0 = pp_19[42]; // @[Multiplier.scala 60:38]
  assign c53_304_io_in_1 = pp_20[40]; // @[Multiplier.scala 60:38]
  assign c53_304_io_in_2 = pp_21[38]; // @[Multiplier.scala 60:38]
  assign c53_304_io_in_3 = pp_22[36]; // @[Multiplier.scala 60:38]
  assign c53_304_io_in_4 = c53_300_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_305_io_in_0 = pp_23[34]; // @[Multiplier.scala 60:38]
  assign c53_305_io_in_1 = pp_24[32]; // @[Multiplier.scala 60:38]
  assign c53_305_io_in_2 = pp_25[30]; // @[Multiplier.scala 60:38]
  assign c53_305_io_in_3 = pp_26[28]; // @[Multiplier.scala 60:38]
  assign c53_305_io_in_4 = c53_301_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_306_io_in_0 = pp_12[57]; // @[Multiplier.scala 60:38]
  assign c53_306_io_in_1 = pp_13[55]; // @[Multiplier.scala 60:38]
  assign c53_306_io_in_2 = pp_14[53]; // @[Multiplier.scala 60:38]
  assign c53_306_io_in_3 = pp_15[51]; // @[Multiplier.scala 60:38]
  assign c53_306_io_in_4 = c53_302_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_307_io_in_0 = pp_16[49]; // @[Multiplier.scala 60:38]
  assign c53_307_io_in_1 = pp_17[47]; // @[Multiplier.scala 60:38]
  assign c53_307_io_in_2 = pp_18[45]; // @[Multiplier.scala 60:38]
  assign c53_307_io_in_3 = pp_19[43]; // @[Multiplier.scala 60:38]
  assign c53_307_io_in_4 = c53_303_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_308_io_in_0 = pp_20[41]; // @[Multiplier.scala 60:38]
  assign c53_308_io_in_1 = pp_21[39]; // @[Multiplier.scala 60:38]
  assign c53_308_io_in_2 = pp_22[37]; // @[Multiplier.scala 60:38]
  assign c53_308_io_in_3 = pp_23[35]; // @[Multiplier.scala 60:38]
  assign c53_308_io_in_4 = c53_304_io_out_1; // @[Multiplier.scala 89:41]
  assign c32_24_io_in_0 = pp_24[33]; // @[Multiplier.scala 60:38]
  assign c32_24_io_in_1 = pp_25[31]; // @[Multiplier.scala 60:38]
  assign c32_24_io_in_2 = pp_26[29]; // @[Multiplier.scala 60:38]
  assign c53_309_io_in_0 = pp_12[58]; // @[Multiplier.scala 60:38]
  assign c53_309_io_in_1 = pp_13[56]; // @[Multiplier.scala 60:38]
  assign c53_309_io_in_2 = pp_14[54]; // @[Multiplier.scala 60:38]
  assign c53_309_io_in_3 = pp_15[52]; // @[Multiplier.scala 60:38]
  assign c53_309_io_in_4 = c53_306_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_310_io_in_0 = pp_16[50]; // @[Multiplier.scala 60:38]
  assign c53_310_io_in_1 = pp_17[48]; // @[Multiplier.scala 60:38]
  assign c53_310_io_in_2 = pp_18[46]; // @[Multiplier.scala 60:38]
  assign c53_310_io_in_3 = pp_19[44]; // @[Multiplier.scala 60:38]
  assign c53_310_io_in_4 = c53_307_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_311_io_in_0 = pp_20[42]; // @[Multiplier.scala 60:38]
  assign c53_311_io_in_1 = pp_21[40]; // @[Multiplier.scala 60:38]
  assign c53_311_io_in_2 = pp_22[38]; // @[Multiplier.scala 60:38]
  assign c53_311_io_in_3 = pp_23[36]; // @[Multiplier.scala 60:38]
  assign c53_311_io_in_4 = c53_308_io_out_1; // @[Multiplier.scala 89:41]
  assign c32_25_io_in_0 = pp_24[34]; // @[Multiplier.scala 60:38]
  assign c32_25_io_in_1 = pp_25[32]; // @[Multiplier.scala 60:38]
  assign c32_25_io_in_2 = pp_26[30]; // @[Multiplier.scala 60:38]
  assign c53_312_io_in_0 = pp_13[57]; // @[Multiplier.scala 60:38]
  assign c53_312_io_in_1 = pp_14[55]; // @[Multiplier.scala 60:38]
  assign c53_312_io_in_2 = pp_15[53]; // @[Multiplier.scala 60:38]
  assign c53_312_io_in_3 = pp_16[51]; // @[Multiplier.scala 60:38]
  assign c53_312_io_in_4 = c53_309_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_313_io_in_0 = pp_17[49]; // @[Multiplier.scala 60:38]
  assign c53_313_io_in_1 = pp_18[47]; // @[Multiplier.scala 60:38]
  assign c53_313_io_in_2 = pp_19[45]; // @[Multiplier.scala 60:38]
  assign c53_313_io_in_3 = pp_20[43]; // @[Multiplier.scala 60:38]
  assign c53_313_io_in_4 = c53_310_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_314_io_in_0 = pp_21[41]; // @[Multiplier.scala 60:38]
  assign c53_314_io_in_1 = pp_22[39]; // @[Multiplier.scala 60:38]
  assign c53_314_io_in_2 = pp_23[37]; // @[Multiplier.scala 60:38]
  assign c53_314_io_in_3 = pp_24[35]; // @[Multiplier.scala 60:38]
  assign c53_314_io_in_4 = c53_311_io_out_1; // @[Multiplier.scala 89:41]
  assign c22_19_io_in_0 = pp_25[33]; // @[Multiplier.scala 60:38]
  assign c22_19_io_in_1 = pp_26[31]; // @[Multiplier.scala 60:38]
  assign c53_315_io_in_0 = pp_13[58]; // @[Multiplier.scala 60:38]
  assign c53_315_io_in_1 = pp_14[56]; // @[Multiplier.scala 60:38]
  assign c53_315_io_in_2 = pp_15[54]; // @[Multiplier.scala 60:38]
  assign c53_315_io_in_3 = pp_16[52]; // @[Multiplier.scala 60:38]
  assign c53_315_io_in_4 = c53_312_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_316_io_in_0 = pp_17[50]; // @[Multiplier.scala 60:38]
  assign c53_316_io_in_1 = pp_18[48]; // @[Multiplier.scala 60:38]
  assign c53_316_io_in_2 = pp_19[46]; // @[Multiplier.scala 60:38]
  assign c53_316_io_in_3 = pp_20[44]; // @[Multiplier.scala 60:38]
  assign c53_316_io_in_4 = c53_313_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_317_io_in_0 = pp_21[42]; // @[Multiplier.scala 60:38]
  assign c53_317_io_in_1 = pp_22[40]; // @[Multiplier.scala 60:38]
  assign c53_317_io_in_2 = pp_23[38]; // @[Multiplier.scala 60:38]
  assign c53_317_io_in_3 = pp_24[36]; // @[Multiplier.scala 60:38]
  assign c53_317_io_in_4 = c53_314_io_out_1; // @[Multiplier.scala 89:41]
  assign c22_20_io_in_0 = pp_25[34]; // @[Multiplier.scala 60:38]
  assign c22_20_io_in_1 = pp_26[32]; // @[Multiplier.scala 60:38]
  assign c53_318_io_in_0 = pp_14[57]; // @[Multiplier.scala 60:38]
  assign c53_318_io_in_1 = pp_15[55]; // @[Multiplier.scala 60:38]
  assign c53_318_io_in_2 = pp_16[53]; // @[Multiplier.scala 60:38]
  assign c53_318_io_in_3 = pp_17[51]; // @[Multiplier.scala 60:38]
  assign c53_318_io_in_4 = c53_315_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_319_io_in_0 = pp_18[49]; // @[Multiplier.scala 60:38]
  assign c53_319_io_in_1 = pp_19[47]; // @[Multiplier.scala 60:38]
  assign c53_319_io_in_2 = pp_20[45]; // @[Multiplier.scala 60:38]
  assign c53_319_io_in_3 = pp_21[43]; // @[Multiplier.scala 60:38]
  assign c53_319_io_in_4 = c53_316_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_320_io_in_0 = pp_22[41]; // @[Multiplier.scala 60:38]
  assign c53_320_io_in_1 = pp_23[39]; // @[Multiplier.scala 60:38]
  assign c53_320_io_in_2 = pp_24[37]; // @[Multiplier.scala 60:38]
  assign c53_320_io_in_3 = pp_25[35]; // @[Multiplier.scala 60:38]
  assign c53_320_io_in_4 = c53_317_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_321_io_in_0 = pp_14[58]; // @[Multiplier.scala 60:38]
  assign c53_321_io_in_1 = pp_15[56]; // @[Multiplier.scala 60:38]
  assign c53_321_io_in_2 = pp_16[54]; // @[Multiplier.scala 60:38]
  assign c53_321_io_in_3 = pp_17[52]; // @[Multiplier.scala 60:38]
  assign c53_321_io_in_4 = c53_318_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_322_io_in_0 = pp_18[50]; // @[Multiplier.scala 60:38]
  assign c53_322_io_in_1 = pp_19[48]; // @[Multiplier.scala 60:38]
  assign c53_322_io_in_2 = pp_20[46]; // @[Multiplier.scala 60:38]
  assign c53_322_io_in_3 = pp_21[44]; // @[Multiplier.scala 60:38]
  assign c53_322_io_in_4 = c53_319_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_323_io_in_0 = pp_22[42]; // @[Multiplier.scala 60:38]
  assign c53_323_io_in_1 = pp_23[40]; // @[Multiplier.scala 60:38]
  assign c53_323_io_in_2 = pp_24[38]; // @[Multiplier.scala 60:38]
  assign c53_323_io_in_3 = pp_25[36]; // @[Multiplier.scala 60:38]
  assign c53_323_io_in_4 = c53_320_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_324_io_in_0 = pp_15[57]; // @[Multiplier.scala 60:38]
  assign c53_324_io_in_1 = pp_16[55]; // @[Multiplier.scala 60:38]
  assign c53_324_io_in_2 = pp_17[53]; // @[Multiplier.scala 60:38]
  assign c53_324_io_in_3 = pp_18[51]; // @[Multiplier.scala 60:38]
  assign c53_324_io_in_4 = c53_321_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_325_io_in_0 = pp_19[49]; // @[Multiplier.scala 60:38]
  assign c53_325_io_in_1 = pp_20[47]; // @[Multiplier.scala 60:38]
  assign c53_325_io_in_2 = pp_21[45]; // @[Multiplier.scala 60:38]
  assign c53_325_io_in_3 = pp_22[43]; // @[Multiplier.scala 60:38]
  assign c53_325_io_in_4 = c53_322_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_326_io_in_0 = pp_23[41]; // @[Multiplier.scala 60:38]
  assign c53_326_io_in_1 = pp_24[39]; // @[Multiplier.scala 60:38]
  assign c53_326_io_in_2 = pp_25[37]; // @[Multiplier.scala 60:38]
  assign c53_326_io_in_3 = pp_26[35]; // @[Multiplier.scala 60:38]
  assign c53_326_io_in_4 = c53_323_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_327_io_in_0 = pp_15[58]; // @[Multiplier.scala 60:38]
  assign c53_327_io_in_1 = pp_16[56]; // @[Multiplier.scala 60:38]
  assign c53_327_io_in_2 = pp_17[54]; // @[Multiplier.scala 60:38]
  assign c53_327_io_in_3 = pp_18[52]; // @[Multiplier.scala 60:38]
  assign c53_327_io_in_4 = c53_324_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_328_io_in_0 = pp_19[50]; // @[Multiplier.scala 60:38]
  assign c53_328_io_in_1 = pp_20[48]; // @[Multiplier.scala 60:38]
  assign c53_328_io_in_2 = pp_21[46]; // @[Multiplier.scala 60:38]
  assign c53_328_io_in_3 = pp_22[44]; // @[Multiplier.scala 60:38]
  assign c53_328_io_in_4 = c53_325_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_329_io_in_0 = pp_23[42]; // @[Multiplier.scala 60:38]
  assign c53_329_io_in_1 = pp_24[40]; // @[Multiplier.scala 60:38]
  assign c53_329_io_in_2 = pp_25[38]; // @[Multiplier.scala 60:38]
  assign c53_329_io_in_3 = pp_26[36]; // @[Multiplier.scala 60:38]
  assign c53_329_io_in_4 = c53_326_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_330_io_in_0 = pp_16[57]; // @[Multiplier.scala 60:38]
  assign c53_330_io_in_1 = pp_17[55]; // @[Multiplier.scala 60:38]
  assign c53_330_io_in_2 = pp_18[53]; // @[Multiplier.scala 60:38]
  assign c53_330_io_in_3 = pp_19[51]; // @[Multiplier.scala 60:38]
  assign c53_330_io_in_4 = c53_327_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_331_io_in_0 = pp_20[49]; // @[Multiplier.scala 60:38]
  assign c53_331_io_in_1 = pp_21[47]; // @[Multiplier.scala 60:38]
  assign c53_331_io_in_2 = pp_22[45]; // @[Multiplier.scala 60:38]
  assign c53_331_io_in_3 = pp_23[43]; // @[Multiplier.scala 60:38]
  assign c53_331_io_in_4 = c53_328_io_out_1; // @[Multiplier.scala 89:41]
  assign c32_26_io_in_0 = pp_24[41]; // @[Multiplier.scala 60:38]
  assign c32_26_io_in_1 = pp_25[39]; // @[Multiplier.scala 60:38]
  assign c32_26_io_in_2 = pp_26[37]; // @[Multiplier.scala 60:38]
  assign c53_332_io_in_0 = pp_16[58]; // @[Multiplier.scala 60:38]
  assign c53_332_io_in_1 = pp_17[56]; // @[Multiplier.scala 60:38]
  assign c53_332_io_in_2 = pp_18[54]; // @[Multiplier.scala 60:38]
  assign c53_332_io_in_3 = pp_19[52]; // @[Multiplier.scala 60:38]
  assign c53_332_io_in_4 = c53_330_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_333_io_in_0 = pp_20[50]; // @[Multiplier.scala 60:38]
  assign c53_333_io_in_1 = pp_21[48]; // @[Multiplier.scala 60:38]
  assign c53_333_io_in_2 = pp_22[46]; // @[Multiplier.scala 60:38]
  assign c53_333_io_in_3 = pp_23[44]; // @[Multiplier.scala 60:38]
  assign c53_333_io_in_4 = c53_331_io_out_1; // @[Multiplier.scala 89:41]
  assign c32_27_io_in_0 = pp_24[42]; // @[Multiplier.scala 60:38]
  assign c32_27_io_in_1 = pp_25[40]; // @[Multiplier.scala 60:38]
  assign c32_27_io_in_2 = pp_26[38]; // @[Multiplier.scala 60:38]
  assign c53_334_io_in_0 = pp_17[57]; // @[Multiplier.scala 60:38]
  assign c53_334_io_in_1 = pp_18[55]; // @[Multiplier.scala 60:38]
  assign c53_334_io_in_2 = pp_19[53]; // @[Multiplier.scala 60:38]
  assign c53_334_io_in_3 = pp_20[51]; // @[Multiplier.scala 60:38]
  assign c53_334_io_in_4 = c53_332_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_335_io_in_0 = pp_21[49]; // @[Multiplier.scala 60:38]
  assign c53_335_io_in_1 = pp_22[47]; // @[Multiplier.scala 60:38]
  assign c53_335_io_in_2 = pp_23[45]; // @[Multiplier.scala 60:38]
  assign c53_335_io_in_3 = pp_24[43]; // @[Multiplier.scala 60:38]
  assign c53_335_io_in_4 = c53_333_io_out_1; // @[Multiplier.scala 89:41]
  assign c22_21_io_in_0 = pp_25[41]; // @[Multiplier.scala 60:38]
  assign c22_21_io_in_1 = pp_26[39]; // @[Multiplier.scala 60:38]
  assign c53_336_io_in_0 = pp_17[58]; // @[Multiplier.scala 60:38]
  assign c53_336_io_in_1 = pp_18[56]; // @[Multiplier.scala 60:38]
  assign c53_336_io_in_2 = pp_19[54]; // @[Multiplier.scala 60:38]
  assign c53_336_io_in_3 = pp_20[52]; // @[Multiplier.scala 60:38]
  assign c53_336_io_in_4 = c53_334_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_337_io_in_0 = pp_21[50]; // @[Multiplier.scala 60:38]
  assign c53_337_io_in_1 = pp_22[48]; // @[Multiplier.scala 60:38]
  assign c53_337_io_in_2 = pp_23[46]; // @[Multiplier.scala 60:38]
  assign c53_337_io_in_3 = pp_24[44]; // @[Multiplier.scala 60:38]
  assign c53_337_io_in_4 = c53_335_io_out_1; // @[Multiplier.scala 89:41]
  assign c22_22_io_in_0 = pp_25[42]; // @[Multiplier.scala 60:38]
  assign c22_22_io_in_1 = pp_26[40]; // @[Multiplier.scala 60:38]
  assign c53_338_io_in_0 = pp_18[57]; // @[Multiplier.scala 60:38]
  assign c53_338_io_in_1 = pp_19[55]; // @[Multiplier.scala 60:38]
  assign c53_338_io_in_2 = pp_20[53]; // @[Multiplier.scala 60:38]
  assign c53_338_io_in_3 = pp_21[51]; // @[Multiplier.scala 60:38]
  assign c53_338_io_in_4 = c53_336_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_339_io_in_0 = pp_22[49]; // @[Multiplier.scala 60:38]
  assign c53_339_io_in_1 = pp_23[47]; // @[Multiplier.scala 60:38]
  assign c53_339_io_in_2 = pp_24[45]; // @[Multiplier.scala 60:38]
  assign c53_339_io_in_3 = pp_25[43]; // @[Multiplier.scala 60:38]
  assign c53_339_io_in_4 = c53_337_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_340_io_in_0 = pp_18[58]; // @[Multiplier.scala 60:38]
  assign c53_340_io_in_1 = pp_19[56]; // @[Multiplier.scala 60:38]
  assign c53_340_io_in_2 = pp_20[54]; // @[Multiplier.scala 60:38]
  assign c53_340_io_in_3 = pp_21[52]; // @[Multiplier.scala 60:38]
  assign c53_340_io_in_4 = c53_338_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_341_io_in_0 = pp_22[50]; // @[Multiplier.scala 60:38]
  assign c53_341_io_in_1 = pp_23[48]; // @[Multiplier.scala 60:38]
  assign c53_341_io_in_2 = pp_24[46]; // @[Multiplier.scala 60:38]
  assign c53_341_io_in_3 = pp_25[44]; // @[Multiplier.scala 60:38]
  assign c53_341_io_in_4 = c53_339_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_342_io_in_0 = pp_19[57]; // @[Multiplier.scala 60:38]
  assign c53_342_io_in_1 = pp_20[55]; // @[Multiplier.scala 60:38]
  assign c53_342_io_in_2 = pp_21[53]; // @[Multiplier.scala 60:38]
  assign c53_342_io_in_3 = pp_22[51]; // @[Multiplier.scala 60:38]
  assign c53_342_io_in_4 = c53_340_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_343_io_in_0 = pp_23[49]; // @[Multiplier.scala 60:38]
  assign c53_343_io_in_1 = pp_24[47]; // @[Multiplier.scala 60:38]
  assign c53_343_io_in_2 = pp_25[45]; // @[Multiplier.scala 60:38]
  assign c53_343_io_in_3 = pp_26[43]; // @[Multiplier.scala 60:38]
  assign c53_343_io_in_4 = c53_341_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_344_io_in_0 = pp_19[58]; // @[Multiplier.scala 60:38]
  assign c53_344_io_in_1 = pp_20[56]; // @[Multiplier.scala 60:38]
  assign c53_344_io_in_2 = pp_21[54]; // @[Multiplier.scala 60:38]
  assign c53_344_io_in_3 = pp_22[52]; // @[Multiplier.scala 60:38]
  assign c53_344_io_in_4 = c53_342_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_345_io_in_0 = pp_23[50]; // @[Multiplier.scala 60:38]
  assign c53_345_io_in_1 = pp_24[48]; // @[Multiplier.scala 60:38]
  assign c53_345_io_in_2 = pp_25[46]; // @[Multiplier.scala 60:38]
  assign c53_345_io_in_3 = pp_26[44]; // @[Multiplier.scala 60:38]
  assign c53_345_io_in_4 = c53_343_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_346_io_in_0 = pp_20[57]; // @[Multiplier.scala 60:38]
  assign c53_346_io_in_1 = pp_21[55]; // @[Multiplier.scala 60:38]
  assign c53_346_io_in_2 = pp_22[53]; // @[Multiplier.scala 60:38]
  assign c53_346_io_in_3 = pp_23[51]; // @[Multiplier.scala 60:38]
  assign c53_346_io_in_4 = c53_344_io_out_1; // @[Multiplier.scala 89:41]
  assign c32_28_io_in_0 = pp_24[49]; // @[Multiplier.scala 60:38]
  assign c32_28_io_in_1 = pp_25[47]; // @[Multiplier.scala 60:38]
  assign c32_28_io_in_2 = pp_26[45]; // @[Multiplier.scala 60:38]
  assign c53_347_io_in_0 = pp_20[58]; // @[Multiplier.scala 60:38]
  assign c53_347_io_in_1 = pp_21[56]; // @[Multiplier.scala 60:38]
  assign c53_347_io_in_2 = pp_22[54]; // @[Multiplier.scala 60:38]
  assign c53_347_io_in_3 = pp_23[52]; // @[Multiplier.scala 60:38]
  assign c53_347_io_in_4 = c53_346_io_out_1; // @[Multiplier.scala 89:41]
  assign c32_29_io_in_0 = pp_24[50]; // @[Multiplier.scala 60:38]
  assign c32_29_io_in_1 = pp_25[48]; // @[Multiplier.scala 60:38]
  assign c32_29_io_in_2 = pp_26[46]; // @[Multiplier.scala 60:38]
  assign c53_348_io_in_0 = pp_21[57]; // @[Multiplier.scala 60:38]
  assign c53_348_io_in_1 = pp_22[55]; // @[Multiplier.scala 60:38]
  assign c53_348_io_in_2 = pp_23[53]; // @[Multiplier.scala 60:38]
  assign c53_348_io_in_3 = pp_24[51]; // @[Multiplier.scala 60:38]
  assign c53_348_io_in_4 = c53_347_io_out_1; // @[Multiplier.scala 89:41]
  assign c22_23_io_in_0 = pp_25[49]; // @[Multiplier.scala 60:38]
  assign c22_23_io_in_1 = pp_26[47]; // @[Multiplier.scala 60:38]
  assign c53_349_io_in_0 = pp_21[58]; // @[Multiplier.scala 60:38]
  assign c53_349_io_in_1 = pp_22[56]; // @[Multiplier.scala 60:38]
  assign c53_349_io_in_2 = pp_23[54]; // @[Multiplier.scala 60:38]
  assign c53_349_io_in_3 = pp_24[52]; // @[Multiplier.scala 60:38]
  assign c53_349_io_in_4 = c53_348_io_out_1; // @[Multiplier.scala 89:41]
  assign c22_24_io_in_0 = pp_25[50]; // @[Multiplier.scala 60:38]
  assign c22_24_io_in_1 = pp_26[48]; // @[Multiplier.scala 60:38]
  assign c53_350_io_in_0 = pp_22[57]; // @[Multiplier.scala 60:38]
  assign c53_350_io_in_1 = pp_23[55]; // @[Multiplier.scala 60:38]
  assign c53_350_io_in_2 = pp_24[53]; // @[Multiplier.scala 60:38]
  assign c53_350_io_in_3 = pp_25[51]; // @[Multiplier.scala 60:38]
  assign c53_350_io_in_4 = c53_349_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_351_io_in_0 = pp_22[58]; // @[Multiplier.scala 60:38]
  assign c53_351_io_in_1 = pp_23[56]; // @[Multiplier.scala 60:38]
  assign c53_351_io_in_2 = pp_24[54]; // @[Multiplier.scala 60:38]
  assign c53_351_io_in_3 = pp_25[52]; // @[Multiplier.scala 60:38]
  assign c53_351_io_in_4 = c53_350_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_352_io_in_0 = pp_23[57]; // @[Multiplier.scala 60:38]
  assign c53_352_io_in_1 = pp_24[55]; // @[Multiplier.scala 60:38]
  assign c53_352_io_in_2 = pp_25[53]; // @[Multiplier.scala 60:38]
  assign c53_352_io_in_3 = pp_26[51]; // @[Multiplier.scala 60:38]
  assign c53_352_io_in_4 = c53_351_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_353_io_in_0 = pp_23[58]; // @[Multiplier.scala 60:38]
  assign c53_353_io_in_1 = pp_24[56]; // @[Multiplier.scala 60:38]
  assign c53_353_io_in_2 = pp_25[54]; // @[Multiplier.scala 60:38]
  assign c53_353_io_in_3 = pp_26[52]; // @[Multiplier.scala 60:38]
  assign c53_353_io_in_4 = c53_352_io_out_1; // @[Multiplier.scala 89:41]
  assign c32_30_io_in_0 = pp_24[57]; // @[Multiplier.scala 60:38]
  assign c32_30_io_in_1 = pp_25[55]; // @[Multiplier.scala 60:38]
  assign c32_30_io_in_2 = pp_26[53]; // @[Multiplier.scala 60:38]
  assign c32_31_io_in_0 = pp_24[58]; // @[Multiplier.scala 60:38]
  assign c32_31_io_in_1 = pp_25[56]; // @[Multiplier.scala 60:38]
  assign c32_31_io_in_2 = pp_26[54]; // @[Multiplier.scala 60:38]
  assign c22_25_io_in_0 = pp_25[57]; // @[Multiplier.scala 60:38]
  assign c22_25_io_in_1 = pp_26[55]; // @[Multiplier.scala 60:38]
  assign c22_26_io_in_0 = pp_25[58]; // @[Multiplier.scala 60:38]
  assign c22_26_io_in_1 = pp_26[56]; // @[Multiplier.scala 60:38]
  assign c22_27_io_in_0 = c22_1_io_out_0; // @[Multiplier.scala 75:35]
  assign c22_27_io_in_1 = c22_io_out_1; // @[Multiplier.scala 76:41]
  assign c22_28_io_in_0 = c32_io_out_0; // @[Multiplier.scala 80:35]
  assign c22_28_io_in_1 = c22_1_io_out_1; // @[Multiplier.scala 76:41]
  assign c22_29_io_in_0 = c32_1_io_out_0; // @[Multiplier.scala 80:35]
  assign c22_29_io_in_1 = c32_io_out_1; // @[Multiplier.scala 81:41]
  assign c22_30_io_in_0 = c53_io_out_0; // @[Multiplier.scala 88:39]
  assign c22_30_io_in_1 = c32_1_io_out_1; // @[Multiplier.scala 81:41]
  assign c22_31_io_in_0 = c53_1_io_out_0; // @[Multiplier.scala 88:39]
  assign c22_31_io_in_1 = c53_io_out_2; // @[Multiplier.scala 90:41]
  assign c32_32_io_in_0 = c53_2_io_out_0; // @[Multiplier.scala 88:39]
  assign c32_32_io_in_1 = pp_4[0]; // @[Multiplier.scala 60:38]
  assign c32_32_io_in_2 = c53_1_io_out_2; // @[Multiplier.scala 90:41]
  assign c32_33_io_in_0 = c53_3_io_out_0; // @[Multiplier.scala 88:39]
  assign c32_33_io_in_1 = pp_4[1]; // @[Multiplier.scala 60:38]
  assign c32_33_io_in_2 = c53_2_io_out_2; // @[Multiplier.scala 90:41]
  assign c32_34_io_in_0 = c53_4_io_out_0; // @[Multiplier.scala 88:39]
  assign c32_34_io_in_1 = c22_2_io_out_0; // @[Multiplier.scala 75:35]
  assign c32_34_io_in_2 = c53_3_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_354_io_in_0 = c53_5_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_354_io_in_1 = c22_3_io_out_0; // @[Multiplier.scala 75:35]
  assign c53_354_io_in_2 = c53_4_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_354_io_in_3 = c22_2_io_out_1; // @[Multiplier.scala 76:41]
  assign c53_354_io_in_4 = 1'h0; // @[Multiplier.scala 87:24]
  assign c53_355_io_in_0 = c53_6_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_355_io_in_1 = c32_2_io_out_0; // @[Multiplier.scala 80:35]
  assign c53_355_io_in_2 = c53_5_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_355_io_in_3 = c22_3_io_out_1; // @[Multiplier.scala 76:41]
  assign c53_355_io_in_4 = c53_354_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_356_io_in_0 = c53_7_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_356_io_in_1 = c32_3_io_out_0; // @[Multiplier.scala 80:35]
  assign c53_356_io_in_2 = c53_6_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_356_io_in_3 = c32_2_io_out_1; // @[Multiplier.scala 81:41]
  assign c53_356_io_in_4 = c53_355_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_357_io_in_0 = c53_8_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_357_io_in_1 = c53_9_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_357_io_in_2 = c53_7_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_357_io_in_3 = c32_3_io_out_1; // @[Multiplier.scala 81:41]
  assign c53_357_io_in_4 = c53_356_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_358_io_in_0 = c53_10_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_358_io_in_1 = c53_11_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_358_io_in_2 = c53_8_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_358_io_in_3 = c53_9_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_358_io_in_4 = c53_357_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_359_io_in_0 = c53_12_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_359_io_in_1 = c53_13_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_359_io_in_2 = pp_8[0]; // @[Multiplier.scala 60:38]
  assign c53_359_io_in_3 = c53_10_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_359_io_in_4 = c53_358_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_360_io_in_0 = c53_14_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_360_io_in_1 = c53_15_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_360_io_in_2 = pp_8[1]; // @[Multiplier.scala 60:38]
  assign c53_360_io_in_3 = c53_12_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_360_io_in_4 = c53_359_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_361_io_in_0 = c53_16_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_361_io_in_1 = c53_17_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_361_io_in_2 = c22_4_io_out_0; // @[Multiplier.scala 75:35]
  assign c53_361_io_in_3 = c53_14_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_361_io_in_4 = c53_360_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_362_io_in_0 = c53_18_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_362_io_in_1 = c53_19_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_362_io_in_2 = c22_5_io_out_0; // @[Multiplier.scala 75:35]
  assign c53_362_io_in_3 = c53_16_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_362_io_in_4 = c53_361_io_out_1; // @[Multiplier.scala 89:41]
  assign c22_32_io_in_0 = c53_17_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_32_io_in_1 = c22_4_io_out_1; // @[Multiplier.scala 76:41]
  assign c53_363_io_in_0 = c53_20_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_363_io_in_1 = c53_21_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_363_io_in_2 = c32_4_io_out_0; // @[Multiplier.scala 80:35]
  assign c53_363_io_in_3 = c53_18_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_363_io_in_4 = c53_362_io_out_1; // @[Multiplier.scala 89:41]
  assign c22_33_io_in_0 = c53_19_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_33_io_in_1 = c22_5_io_out_1; // @[Multiplier.scala 76:41]
  assign c53_364_io_in_0 = c53_22_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_364_io_in_1 = c53_23_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_364_io_in_2 = c32_5_io_out_0; // @[Multiplier.scala 80:35]
  assign c53_364_io_in_3 = c53_20_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_364_io_in_4 = c53_363_io_out_1; // @[Multiplier.scala 89:41]
  assign c22_34_io_in_0 = c53_21_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_34_io_in_1 = c32_4_io_out_1; // @[Multiplier.scala 81:41]
  assign c53_365_io_in_0 = c53_24_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_365_io_in_1 = c53_25_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_365_io_in_2 = c53_26_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_365_io_in_3 = c53_22_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_365_io_in_4 = c53_364_io_out_1; // @[Multiplier.scala 89:41]
  assign c22_35_io_in_0 = c53_23_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_35_io_in_1 = c32_5_io_out_1; // @[Multiplier.scala 81:41]
  assign c53_366_io_in_0 = c53_27_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_366_io_in_1 = c53_28_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_366_io_in_2 = c53_29_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_366_io_in_3 = c53_24_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_366_io_in_4 = c53_365_io_out_1; // @[Multiplier.scala 89:41]
  assign c22_36_io_in_0 = c53_25_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_36_io_in_1 = c53_26_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_367_io_in_0 = c53_30_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_367_io_in_1 = c53_31_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_367_io_in_2 = c53_32_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_367_io_in_3 = pp_12[0]; // @[Multiplier.scala 60:38]
  assign c53_367_io_in_4 = c53_366_io_out_1; // @[Multiplier.scala 89:41]
  assign c32_35_io_in_0 = c53_27_io_out_2; // @[Multiplier.scala 90:41]
  assign c32_35_io_in_1 = c53_28_io_out_2; // @[Multiplier.scala 90:41]
  assign c32_35_io_in_2 = c53_29_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_368_io_in_0 = c53_33_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_368_io_in_1 = c53_34_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_368_io_in_2 = c53_35_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_368_io_in_3 = pp_12[1]; // @[Multiplier.scala 60:38]
  assign c53_368_io_in_4 = c53_367_io_out_1; // @[Multiplier.scala 89:41]
  assign c32_36_io_in_0 = c53_30_io_out_2; // @[Multiplier.scala 90:41]
  assign c32_36_io_in_1 = c53_31_io_out_2; // @[Multiplier.scala 90:41]
  assign c32_36_io_in_2 = c53_32_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_369_io_in_0 = c53_36_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_369_io_in_1 = c53_37_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_369_io_in_2 = c53_38_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_369_io_in_3 = c22_6_io_out_0; // @[Multiplier.scala 75:35]
  assign c53_369_io_in_4 = c53_368_io_out_1; // @[Multiplier.scala 89:41]
  assign c32_37_io_in_0 = c53_33_io_out_2; // @[Multiplier.scala 90:41]
  assign c32_37_io_in_1 = c53_34_io_out_2; // @[Multiplier.scala 90:41]
  assign c32_37_io_in_2 = c53_35_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_370_io_in_0 = c53_39_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_370_io_in_1 = c53_40_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_370_io_in_2 = c53_41_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_370_io_in_3 = c22_7_io_out_0; // @[Multiplier.scala 75:35]
  assign c53_370_io_in_4 = c53_369_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_371_io_in_0 = c53_36_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_371_io_in_1 = c53_37_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_371_io_in_2 = c53_38_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_371_io_in_3 = c22_6_io_out_1; // @[Multiplier.scala 76:41]
  assign c53_371_io_in_4 = 1'h0; // @[Multiplier.scala 87:24]
  assign c53_372_io_in_0 = c53_42_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_372_io_in_1 = c53_43_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_372_io_in_2 = c53_44_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_372_io_in_3 = c32_6_io_out_0; // @[Multiplier.scala 80:35]
  assign c53_372_io_in_4 = c53_370_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_373_io_in_0 = c53_39_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_373_io_in_1 = c53_40_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_373_io_in_2 = c53_41_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_373_io_in_3 = c22_7_io_out_1; // @[Multiplier.scala 76:41]
  assign c53_373_io_in_4 = c53_371_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_374_io_in_0 = c53_45_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_374_io_in_1 = c53_46_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_374_io_in_2 = c53_47_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_374_io_in_3 = c32_7_io_out_0; // @[Multiplier.scala 80:35]
  assign c53_374_io_in_4 = c53_372_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_375_io_in_0 = c53_42_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_375_io_in_1 = c53_43_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_375_io_in_2 = c53_44_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_375_io_in_3 = c32_6_io_out_1; // @[Multiplier.scala 81:41]
  assign c53_375_io_in_4 = c53_373_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_376_io_in_0 = c53_48_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_376_io_in_1 = c53_49_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_376_io_in_2 = c53_50_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_376_io_in_3 = c53_51_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_376_io_in_4 = c53_374_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_377_io_in_0 = c53_45_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_377_io_in_1 = c53_46_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_377_io_in_2 = c53_47_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_377_io_in_3 = c32_7_io_out_1; // @[Multiplier.scala 81:41]
  assign c53_377_io_in_4 = c53_375_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_378_io_in_0 = c53_52_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_378_io_in_1 = c53_53_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_378_io_in_2 = c53_54_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_378_io_in_3 = c53_55_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_378_io_in_4 = c53_376_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_379_io_in_0 = c53_48_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_379_io_in_1 = c53_49_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_379_io_in_2 = c53_50_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_379_io_in_3 = c53_51_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_379_io_in_4 = c53_377_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_380_io_in_0 = c53_56_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_380_io_in_1 = c53_57_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_380_io_in_2 = c53_58_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_380_io_in_3 = c53_59_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_380_io_in_4 = c53_378_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_381_io_in_0 = pp_16[0]; // @[Multiplier.scala 60:38]
  assign c53_381_io_in_1 = c53_52_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_381_io_in_2 = c53_53_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_381_io_in_3 = c53_54_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_381_io_in_4 = c53_379_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_382_io_in_0 = c53_60_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_382_io_in_1 = c53_61_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_382_io_in_2 = c53_62_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_382_io_in_3 = c53_63_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_382_io_in_4 = c53_380_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_383_io_in_0 = pp_16[1]; // @[Multiplier.scala 60:38]
  assign c53_383_io_in_1 = c53_56_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_383_io_in_2 = c53_57_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_383_io_in_3 = c53_58_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_383_io_in_4 = c53_381_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_384_io_in_0 = c53_64_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_384_io_in_1 = c53_65_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_384_io_in_2 = c53_66_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_384_io_in_3 = c53_67_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_384_io_in_4 = c53_382_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_385_io_in_0 = c22_8_io_out_0; // @[Multiplier.scala 75:35]
  assign c53_385_io_in_1 = c53_60_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_385_io_in_2 = c53_61_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_385_io_in_3 = c53_62_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_385_io_in_4 = c53_383_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_386_io_in_0 = c53_68_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_386_io_in_1 = c53_69_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_386_io_in_2 = c53_70_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_386_io_in_3 = c53_71_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_386_io_in_4 = c53_384_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_387_io_in_0 = c22_9_io_out_0; // @[Multiplier.scala 75:35]
  assign c53_387_io_in_1 = c53_64_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_387_io_in_2 = c53_65_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_387_io_in_3 = c53_66_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_387_io_in_4 = c53_385_io_out_1; // @[Multiplier.scala 89:41]
  assign c22_37_io_in_0 = c53_67_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_37_io_in_1 = c22_8_io_out_1; // @[Multiplier.scala 76:41]
  assign c53_388_io_in_0 = c53_72_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_388_io_in_1 = c53_73_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_388_io_in_2 = c53_74_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_388_io_in_3 = c53_75_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_388_io_in_4 = c53_386_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_389_io_in_0 = c32_8_io_out_0; // @[Multiplier.scala 80:35]
  assign c53_389_io_in_1 = c53_68_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_389_io_in_2 = c53_69_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_389_io_in_3 = c53_70_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_389_io_in_4 = c53_387_io_out_1; // @[Multiplier.scala 89:41]
  assign c22_38_io_in_0 = c53_71_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_38_io_in_1 = c22_9_io_out_1; // @[Multiplier.scala 76:41]
  assign c53_390_io_in_0 = c53_76_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_390_io_in_1 = c53_77_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_390_io_in_2 = c53_78_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_390_io_in_3 = c53_79_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_390_io_in_4 = c53_388_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_391_io_in_0 = c32_9_io_out_0; // @[Multiplier.scala 80:35]
  assign c53_391_io_in_1 = c53_72_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_391_io_in_2 = c53_73_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_391_io_in_3 = c53_74_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_391_io_in_4 = c53_389_io_out_1; // @[Multiplier.scala 89:41]
  assign c22_39_io_in_0 = c53_75_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_39_io_in_1 = c32_8_io_out_1; // @[Multiplier.scala 81:41]
  assign c53_392_io_in_0 = c53_80_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_392_io_in_1 = c53_81_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_392_io_in_2 = c53_82_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_392_io_in_3 = c53_83_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_392_io_in_4 = c53_390_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_393_io_in_0 = c53_84_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_393_io_in_1 = c53_76_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_393_io_in_2 = c53_77_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_393_io_in_3 = c53_78_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_393_io_in_4 = c53_391_io_out_1; // @[Multiplier.scala 89:41]
  assign c22_40_io_in_0 = c53_79_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_40_io_in_1 = c32_9_io_out_1; // @[Multiplier.scala 81:41]
  assign c53_394_io_in_0 = c53_85_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_394_io_in_1 = c53_86_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_394_io_in_2 = c53_87_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_394_io_in_3 = c53_88_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_394_io_in_4 = c53_392_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_395_io_in_0 = c53_89_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_395_io_in_1 = c53_80_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_395_io_in_2 = c53_81_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_395_io_in_3 = c53_82_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_395_io_in_4 = c53_393_io_out_1; // @[Multiplier.scala 89:41]
  assign c22_41_io_in_0 = c53_83_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_41_io_in_1 = c53_84_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_396_io_in_0 = c53_90_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_396_io_in_1 = c53_91_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_396_io_in_2 = c53_92_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_396_io_in_3 = c53_93_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_396_io_in_4 = c53_394_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_397_io_in_0 = c53_94_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_397_io_in_1 = pp_20[0]; // @[Multiplier.scala 60:38]
  assign c53_397_io_in_2 = c53_85_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_397_io_in_3 = c53_86_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_397_io_in_4 = c53_395_io_out_1; // @[Multiplier.scala 89:41]
  assign c32_38_io_in_0 = c53_87_io_out_2; // @[Multiplier.scala 90:41]
  assign c32_38_io_in_1 = c53_88_io_out_2; // @[Multiplier.scala 90:41]
  assign c32_38_io_in_2 = c53_89_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_398_io_in_0 = c53_95_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_398_io_in_1 = c53_96_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_398_io_in_2 = c53_97_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_398_io_in_3 = c53_98_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_398_io_in_4 = c53_396_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_399_io_in_0 = c53_99_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_399_io_in_1 = pp_20[1]; // @[Multiplier.scala 60:38]
  assign c53_399_io_in_2 = c53_90_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_399_io_in_3 = c53_91_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_399_io_in_4 = c53_397_io_out_1; // @[Multiplier.scala 89:41]
  assign c32_39_io_in_0 = c53_92_io_out_2; // @[Multiplier.scala 90:41]
  assign c32_39_io_in_1 = c53_93_io_out_2; // @[Multiplier.scala 90:41]
  assign c32_39_io_in_2 = c53_94_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_400_io_in_0 = c53_100_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_400_io_in_1 = c53_101_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_400_io_in_2 = c53_102_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_400_io_in_3 = c53_103_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_400_io_in_4 = c53_398_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_401_io_in_0 = c53_104_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_401_io_in_1 = c22_10_io_out_0; // @[Multiplier.scala 75:35]
  assign c53_401_io_in_2 = c53_95_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_401_io_in_3 = c53_96_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_401_io_in_4 = c53_399_io_out_1; // @[Multiplier.scala 89:41]
  assign c32_40_io_in_0 = c53_97_io_out_2; // @[Multiplier.scala 90:41]
  assign c32_40_io_in_1 = c53_98_io_out_2; // @[Multiplier.scala 90:41]
  assign c32_40_io_in_2 = c53_99_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_402_io_in_0 = c53_105_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_402_io_in_1 = c53_106_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_402_io_in_2 = c53_107_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_402_io_in_3 = c53_108_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_402_io_in_4 = c53_400_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_403_io_in_0 = c53_109_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_403_io_in_1 = c22_11_io_out_0; // @[Multiplier.scala 75:35]
  assign c53_403_io_in_2 = c53_100_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_403_io_in_3 = c53_101_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_403_io_in_4 = c53_401_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_404_io_in_0 = c53_102_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_404_io_in_1 = c53_103_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_404_io_in_2 = c53_104_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_404_io_in_3 = c22_10_io_out_1; // @[Multiplier.scala 76:41]
  assign c53_404_io_in_4 = 1'h0; // @[Multiplier.scala 87:24]
  assign c53_405_io_in_0 = c53_110_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_405_io_in_1 = c53_111_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_405_io_in_2 = c53_112_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_405_io_in_3 = c53_113_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_405_io_in_4 = c53_402_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_406_io_in_0 = c53_114_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_406_io_in_1 = c32_10_io_out_0; // @[Multiplier.scala 80:35]
  assign c53_406_io_in_2 = c53_105_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_406_io_in_3 = c53_106_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_406_io_in_4 = c53_403_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_407_io_in_0 = c53_107_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_407_io_in_1 = c53_108_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_407_io_in_2 = c53_109_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_407_io_in_3 = c22_11_io_out_1; // @[Multiplier.scala 76:41]
  assign c53_407_io_in_4 = c53_404_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_408_io_in_0 = c53_115_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_408_io_in_1 = c53_116_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_408_io_in_2 = c53_117_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_408_io_in_3 = c53_118_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_408_io_in_4 = c53_405_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_409_io_in_0 = c53_119_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_409_io_in_1 = c32_11_io_out_0; // @[Multiplier.scala 80:35]
  assign c53_409_io_in_2 = c53_110_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_409_io_in_3 = c53_111_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_409_io_in_4 = c53_406_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_410_io_in_0 = c53_112_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_410_io_in_1 = c53_113_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_410_io_in_2 = c53_114_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_410_io_in_3 = c32_10_io_out_1; // @[Multiplier.scala 81:41]
  assign c53_410_io_in_4 = c53_407_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_411_io_in_0 = c53_120_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_411_io_in_1 = c53_121_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_411_io_in_2 = c53_122_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_411_io_in_3 = c53_123_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_411_io_in_4 = c53_408_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_412_io_in_0 = c53_124_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_412_io_in_1 = c53_125_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_412_io_in_2 = c53_115_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_412_io_in_3 = c53_116_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_412_io_in_4 = c53_409_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_413_io_in_0 = c53_117_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_413_io_in_1 = c53_118_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_413_io_in_2 = c53_119_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_413_io_in_3 = c32_11_io_out_1; // @[Multiplier.scala 81:41]
  assign c53_413_io_in_4 = c53_410_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_414_io_in_0 = c53_126_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_414_io_in_1 = c53_127_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_414_io_in_2 = c53_128_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_414_io_in_3 = c53_129_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_414_io_in_4 = c53_411_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_415_io_in_0 = c53_130_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_415_io_in_1 = c53_131_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_415_io_in_2 = c53_120_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_415_io_in_3 = c53_121_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_415_io_in_4 = c53_412_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_416_io_in_0 = c53_122_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_416_io_in_1 = c53_123_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_416_io_in_2 = c53_124_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_416_io_in_3 = c53_125_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_416_io_in_4 = c53_413_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_417_io_in_0 = c53_132_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_417_io_in_1 = c53_133_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_417_io_in_2 = c53_134_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_417_io_in_3 = c53_135_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_417_io_in_4 = c53_414_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_418_io_in_0 = c53_136_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_418_io_in_1 = c53_137_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_418_io_in_2 = pp_24[0]; // @[Multiplier.scala 60:38]
  assign c53_418_io_in_3 = c53_126_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_418_io_in_4 = c53_415_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_419_io_in_0 = c53_127_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_419_io_in_1 = c53_128_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_419_io_in_2 = c53_129_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_419_io_in_3 = c53_130_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_419_io_in_4 = c53_416_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_420_io_in_0 = c53_138_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_420_io_in_1 = c53_139_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_420_io_in_2 = c53_140_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_420_io_in_3 = c53_141_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_420_io_in_4 = c53_417_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_421_io_in_0 = c53_142_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_421_io_in_1 = c53_143_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_421_io_in_2 = pp_24[1]; // @[Multiplier.scala 60:38]
  assign c53_421_io_in_3 = c53_132_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_421_io_in_4 = c53_418_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_422_io_in_0 = c53_133_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_422_io_in_1 = c53_134_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_422_io_in_2 = c53_135_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_422_io_in_3 = c53_136_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_422_io_in_4 = c53_419_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_423_io_in_0 = c53_144_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_423_io_in_1 = c53_145_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_423_io_in_2 = c53_146_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_423_io_in_3 = c53_147_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_423_io_in_4 = c53_420_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_424_io_in_0 = c53_148_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_424_io_in_1 = c53_149_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_424_io_in_2 = c22_12_io_out_0; // @[Multiplier.scala 75:35]
  assign c53_424_io_in_3 = c53_138_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_424_io_in_4 = c53_421_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_425_io_in_0 = c53_139_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_425_io_in_1 = c53_140_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_425_io_in_2 = c53_141_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_425_io_in_3 = c53_142_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_425_io_in_4 = c53_422_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_426_io_in_0 = c53_150_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_426_io_in_1 = c53_151_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_426_io_in_2 = c53_152_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_426_io_in_3 = c53_153_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_426_io_in_4 = c53_423_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_427_io_in_0 = c53_154_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_427_io_in_1 = c53_155_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_427_io_in_2 = c22_13_io_out_0; // @[Multiplier.scala 75:35]
  assign c53_427_io_in_3 = c53_144_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_427_io_in_4 = c53_424_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_428_io_in_0 = c53_145_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_428_io_in_1 = c53_146_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_428_io_in_2 = c53_147_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_428_io_in_3 = c53_148_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_428_io_in_4 = c53_425_io_out_1; // @[Multiplier.scala 89:41]
  assign c22_42_io_in_0 = c53_149_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_42_io_in_1 = c22_12_io_out_1; // @[Multiplier.scala 76:41]
  assign c53_429_io_in_0 = c53_156_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_429_io_in_1 = c53_157_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_429_io_in_2 = c53_158_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_429_io_in_3 = c53_159_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_429_io_in_4 = c53_426_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_430_io_in_0 = c53_160_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_430_io_in_1 = c53_161_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_430_io_in_2 = c32_12_io_out_0; // @[Multiplier.scala 80:35]
  assign c53_430_io_in_3 = c53_150_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_430_io_in_4 = c53_427_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_431_io_in_0 = c53_151_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_431_io_in_1 = c53_152_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_431_io_in_2 = c53_153_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_431_io_in_3 = c53_154_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_431_io_in_4 = c53_428_io_out_1; // @[Multiplier.scala 89:41]
  assign c22_43_io_in_0 = c53_155_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_43_io_in_1 = c22_13_io_out_1; // @[Multiplier.scala 76:41]
  assign c53_432_io_in_0 = c53_162_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_432_io_in_1 = c53_163_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_432_io_in_2 = c53_164_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_432_io_in_3 = c53_165_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_432_io_in_4 = c53_429_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_433_io_in_0 = c53_166_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_433_io_in_1 = c53_167_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_433_io_in_2 = c32_13_io_out_0; // @[Multiplier.scala 80:35]
  assign c53_433_io_in_3 = c53_156_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_433_io_in_4 = c53_430_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_434_io_in_0 = c53_157_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_434_io_in_1 = c53_158_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_434_io_in_2 = c53_159_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_434_io_in_3 = c53_160_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_434_io_in_4 = c53_431_io_out_1; // @[Multiplier.scala 89:41]
  assign c22_44_io_in_0 = c53_161_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_44_io_in_1 = c32_12_io_out_1; // @[Multiplier.scala 81:41]
  assign c53_435_io_in_0 = c53_168_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_435_io_in_1 = c53_169_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_435_io_in_2 = c53_170_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_435_io_in_3 = c53_171_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_435_io_in_4 = c53_432_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_436_io_in_0 = c53_172_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_436_io_in_1 = c53_173_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_436_io_in_2 = c32_14_io_out_0; // @[Multiplier.scala 80:35]
  assign c53_436_io_in_3 = c53_162_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_436_io_in_4 = c53_433_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_437_io_in_0 = c53_163_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_437_io_in_1 = c53_164_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_437_io_in_2 = c53_165_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_437_io_in_3 = c53_166_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_437_io_in_4 = c53_434_io_out_1; // @[Multiplier.scala 89:41]
  assign c22_45_io_in_0 = c53_167_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_45_io_in_1 = c32_13_io_out_1; // @[Multiplier.scala 81:41]
  assign c53_438_io_in_0 = c53_174_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_438_io_in_1 = c53_175_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_438_io_in_2 = c53_176_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_438_io_in_3 = c53_177_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_438_io_in_4 = c53_435_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_439_io_in_0 = c53_178_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_439_io_in_1 = c53_179_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_439_io_in_2 = c32_15_io_out_0; // @[Multiplier.scala 80:35]
  assign c53_439_io_in_3 = c53_168_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_439_io_in_4 = c53_436_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_440_io_in_0 = c53_169_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_440_io_in_1 = c53_170_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_440_io_in_2 = c53_171_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_440_io_in_3 = c53_172_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_440_io_in_4 = c53_437_io_out_1; // @[Multiplier.scala 89:41]
  assign c22_46_io_in_0 = c53_173_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_46_io_in_1 = c32_14_io_out_1; // @[Multiplier.scala 81:41]
  assign c53_441_io_in_0 = c53_180_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_441_io_in_1 = c53_181_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_441_io_in_2 = c53_182_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_441_io_in_3 = c53_183_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_441_io_in_4 = c53_438_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_442_io_in_0 = c53_184_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_442_io_in_1 = c53_185_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_442_io_in_2 = c32_16_io_out_0; // @[Multiplier.scala 80:35]
  assign c53_442_io_in_3 = c53_174_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_442_io_in_4 = c53_439_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_443_io_in_0 = c53_175_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_443_io_in_1 = c53_176_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_443_io_in_2 = c53_177_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_443_io_in_3 = c53_178_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_443_io_in_4 = c53_440_io_out_1; // @[Multiplier.scala 89:41]
  assign c22_47_io_in_0 = c53_179_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_47_io_in_1 = c32_15_io_out_1; // @[Multiplier.scala 81:41]
  assign c53_444_io_in_0 = c53_186_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_444_io_in_1 = c53_187_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_444_io_in_2 = c53_188_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_444_io_in_3 = c53_189_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_444_io_in_4 = c53_441_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_445_io_in_0 = c53_190_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_445_io_in_1 = c53_191_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_445_io_in_2 = c32_17_io_out_0; // @[Multiplier.scala 80:35]
  assign c53_445_io_in_3 = c53_180_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_445_io_in_4 = c53_442_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_446_io_in_0 = c53_181_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_446_io_in_1 = c53_182_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_446_io_in_2 = c53_183_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_446_io_in_3 = c53_184_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_446_io_in_4 = c53_443_io_out_1; // @[Multiplier.scala 89:41]
  assign c22_48_io_in_0 = c53_185_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_48_io_in_1 = c32_16_io_out_1; // @[Multiplier.scala 81:41]
  assign c53_447_io_in_0 = c53_192_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_447_io_in_1 = c53_193_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_447_io_in_2 = c53_194_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_447_io_in_3 = c53_195_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_447_io_in_4 = c53_444_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_448_io_in_0 = c53_196_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_448_io_in_1 = c53_197_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_448_io_in_2 = c32_18_io_out_0; // @[Multiplier.scala 80:35]
  assign c53_448_io_in_3 = c53_186_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_448_io_in_4 = c53_445_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_449_io_in_0 = c53_187_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_449_io_in_1 = c53_188_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_449_io_in_2 = c53_189_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_449_io_in_3 = c53_190_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_449_io_in_4 = c53_446_io_out_1; // @[Multiplier.scala 89:41]
  assign c22_49_io_in_0 = c53_191_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_49_io_in_1 = c32_17_io_out_1; // @[Multiplier.scala 81:41]
  assign c53_450_io_in_0 = c53_198_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_450_io_in_1 = c53_199_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_450_io_in_2 = c53_200_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_450_io_in_3 = c53_201_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_450_io_in_4 = c53_447_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_451_io_in_0 = c53_202_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_451_io_in_1 = c53_203_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_451_io_in_2 = c32_19_io_out_0; // @[Multiplier.scala 80:35]
  assign c53_451_io_in_3 = c53_192_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_451_io_in_4 = c53_448_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_452_io_in_0 = c53_193_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_452_io_in_1 = c53_194_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_452_io_in_2 = c53_195_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_452_io_in_3 = c53_196_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_452_io_in_4 = c53_449_io_out_1; // @[Multiplier.scala 89:41]
  assign c22_50_io_in_0 = c53_197_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_50_io_in_1 = c32_18_io_out_1; // @[Multiplier.scala 81:41]
  assign c53_453_io_in_0 = c53_204_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_453_io_in_1 = c53_205_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_453_io_in_2 = c53_206_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_453_io_in_3 = c53_207_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_453_io_in_4 = c53_450_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_454_io_in_0 = c53_208_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_454_io_in_1 = c53_209_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_454_io_in_2 = c22_14_io_out_0; // @[Multiplier.scala 75:35]
  assign c53_454_io_in_3 = c53_198_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_454_io_in_4 = c53_451_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_455_io_in_0 = c53_199_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_455_io_in_1 = c53_200_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_455_io_in_2 = c53_201_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_455_io_in_3 = c53_202_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_455_io_in_4 = c53_452_io_out_1; // @[Multiplier.scala 89:41]
  assign c22_51_io_in_0 = c53_203_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_51_io_in_1 = c32_19_io_out_1; // @[Multiplier.scala 81:41]
  assign c53_456_io_in_0 = c53_210_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_456_io_in_1 = c53_211_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_456_io_in_2 = c53_212_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_456_io_in_3 = c53_213_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_456_io_in_4 = c53_453_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_457_io_in_0 = c53_214_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_457_io_in_1 = c53_215_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_457_io_in_2 = pp_26[9]; // @[Multiplier.scala 60:38]
  assign c53_457_io_in_3 = c53_204_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_457_io_in_4 = c53_454_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_458_io_in_0 = c53_205_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_458_io_in_1 = c53_206_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_458_io_in_2 = c53_207_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_458_io_in_3 = c53_208_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_458_io_in_4 = c53_455_io_out_1; // @[Multiplier.scala 89:41]
  assign c22_52_io_in_0 = c53_209_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_52_io_in_1 = c22_14_io_out_1; // @[Multiplier.scala 76:41]
  assign c53_459_io_in_0 = c53_216_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_459_io_in_1 = c53_217_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_459_io_in_2 = c53_218_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_459_io_in_3 = c53_219_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_459_io_in_4 = c53_456_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_460_io_in_0 = c53_220_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_460_io_in_1 = c53_221_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_460_io_in_2 = pp_26[10]; // @[Multiplier.scala 60:38]
  assign c53_460_io_in_3 = c53_210_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_460_io_in_4 = c53_457_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_461_io_in_0 = c53_211_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_461_io_in_1 = c53_212_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_461_io_in_2 = c53_213_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_461_io_in_3 = c53_214_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_461_io_in_4 = c53_458_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_462_io_in_0 = c53_222_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_462_io_in_1 = c53_223_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_462_io_in_2 = c53_224_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_462_io_in_3 = c53_225_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_462_io_in_4 = c53_459_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_463_io_in_0 = c53_226_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_463_io_in_1 = c53_227_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_463_io_in_2 = c53_216_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_463_io_in_3 = c53_217_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_463_io_in_4 = c53_460_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_464_io_in_0 = c53_218_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_464_io_in_1 = c53_219_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_464_io_in_2 = c53_220_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_464_io_in_3 = c53_221_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_464_io_in_4 = c53_461_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_465_io_in_0 = c53_228_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_465_io_in_1 = c53_229_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_465_io_in_2 = c53_230_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_465_io_in_3 = c53_231_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_465_io_in_4 = c53_462_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_466_io_in_0 = c53_232_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_466_io_in_1 = c53_233_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_466_io_in_2 = c53_222_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_466_io_in_3 = c53_223_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_466_io_in_4 = c53_463_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_467_io_in_0 = c53_224_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_467_io_in_1 = c53_225_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_467_io_in_2 = c53_226_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_467_io_in_3 = c53_227_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_467_io_in_4 = c53_464_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_468_io_in_0 = c53_234_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_468_io_in_1 = c53_235_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_468_io_in_2 = c53_236_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_468_io_in_3 = c53_237_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_468_io_in_4 = c53_465_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_469_io_in_0 = c53_238_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_469_io_in_1 = c32_20_io_out_0; // @[Multiplier.scala 80:35]
  assign c53_469_io_in_2 = c53_233_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_469_io_in_3 = c53_228_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_469_io_in_4 = c53_466_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_470_io_in_0 = c53_229_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_470_io_in_1 = c53_230_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_470_io_in_2 = c53_231_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_470_io_in_3 = c53_232_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_470_io_in_4 = c53_467_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_471_io_in_0 = c53_239_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_471_io_in_1 = c53_240_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_471_io_in_2 = c53_241_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_471_io_in_3 = c53_242_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_471_io_in_4 = c53_468_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_472_io_in_0 = c53_243_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_472_io_in_1 = c32_21_io_out_0; // @[Multiplier.scala 80:35]
  assign c53_472_io_in_2 = c53_234_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_472_io_in_3 = c53_235_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_472_io_in_4 = c53_469_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_473_io_in_0 = c53_236_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_473_io_in_1 = c53_237_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_473_io_in_2 = c53_238_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_473_io_in_3 = c32_20_io_out_1; // @[Multiplier.scala 81:41]
  assign c53_473_io_in_4 = c53_470_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_474_io_in_0 = c53_244_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_474_io_in_1 = c53_245_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_474_io_in_2 = c53_246_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_474_io_in_3 = c53_247_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_474_io_in_4 = c53_471_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_475_io_in_0 = c53_248_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_475_io_in_1 = c22_15_io_out_0; // @[Multiplier.scala 75:35]
  assign c53_475_io_in_2 = c53_239_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_475_io_in_3 = c53_240_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_475_io_in_4 = c53_472_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_476_io_in_0 = c53_241_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_476_io_in_1 = c53_242_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_476_io_in_2 = c53_243_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_476_io_in_3 = c32_21_io_out_1; // @[Multiplier.scala 81:41]
  assign c53_476_io_in_4 = c53_473_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_477_io_in_0 = c53_249_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_477_io_in_1 = c53_250_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_477_io_in_2 = c53_251_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_477_io_in_3 = c53_252_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_477_io_in_4 = c53_474_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_478_io_in_0 = c53_253_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_478_io_in_1 = c22_16_io_out_0; // @[Multiplier.scala 75:35]
  assign c53_478_io_in_2 = c53_244_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_478_io_in_3 = c53_245_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_478_io_in_4 = c53_475_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_479_io_in_0 = c53_246_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_479_io_in_1 = c53_247_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_479_io_in_2 = c53_248_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_479_io_in_3 = c22_15_io_out_1; // @[Multiplier.scala 76:41]
  assign c53_479_io_in_4 = c53_476_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_480_io_in_0 = c53_254_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_480_io_in_1 = c53_255_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_480_io_in_2 = c53_256_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_480_io_in_3 = c53_257_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_480_io_in_4 = c53_477_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_481_io_in_0 = c53_258_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_481_io_in_1 = pp_26[17]; // @[Multiplier.scala 60:38]
  assign c53_481_io_in_2 = c53_249_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_481_io_in_3 = c53_250_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_481_io_in_4 = c53_478_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_482_io_in_0 = c53_251_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_482_io_in_1 = c53_252_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_482_io_in_2 = c53_253_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_482_io_in_3 = c22_16_io_out_1; // @[Multiplier.scala 76:41]
  assign c53_482_io_in_4 = c53_479_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_483_io_in_0 = c53_259_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_483_io_in_1 = c53_260_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_483_io_in_2 = c53_261_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_483_io_in_3 = c53_262_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_483_io_in_4 = c53_480_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_484_io_in_0 = c53_263_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_484_io_in_1 = pp_26[18]; // @[Multiplier.scala 60:38]
  assign c53_484_io_in_2 = c53_254_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_484_io_in_3 = c53_255_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_484_io_in_4 = c53_481_io_out_1; // @[Multiplier.scala 89:41]
  assign c32_41_io_in_0 = c53_256_io_out_2; // @[Multiplier.scala 90:41]
  assign c32_41_io_in_1 = c53_257_io_out_2; // @[Multiplier.scala 90:41]
  assign c32_41_io_in_2 = c53_258_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_485_io_in_0 = c53_264_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_485_io_in_1 = c53_265_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_485_io_in_2 = c53_266_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_485_io_in_3 = c53_267_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_485_io_in_4 = c53_483_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_486_io_in_0 = c53_268_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_486_io_in_1 = c53_259_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_486_io_in_2 = c53_260_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_486_io_in_3 = c53_261_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_486_io_in_4 = c53_484_io_out_1; // @[Multiplier.scala 89:41]
  assign c22_53_io_in_0 = c53_262_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_53_io_in_1 = c53_263_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_487_io_in_0 = c53_269_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_487_io_in_1 = c53_270_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_487_io_in_2 = c53_271_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_487_io_in_3 = c53_272_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_487_io_in_4 = c53_485_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_488_io_in_0 = c53_273_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_488_io_in_1 = c53_264_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_488_io_in_2 = c53_265_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_488_io_in_3 = c53_266_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_488_io_in_4 = c53_486_io_out_1; // @[Multiplier.scala 89:41]
  assign c22_54_io_in_0 = c53_267_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_54_io_in_1 = c53_268_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_489_io_in_0 = c53_274_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_489_io_in_1 = c53_275_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_489_io_in_2 = c53_276_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_489_io_in_3 = c53_277_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_489_io_in_4 = c53_487_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_490_io_in_0 = c32_22_io_out_0; // @[Multiplier.scala 80:35]
  assign c53_490_io_in_1 = c53_273_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_490_io_in_2 = c53_269_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_490_io_in_3 = c53_270_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_490_io_in_4 = c53_488_io_out_1; // @[Multiplier.scala 89:41]
  assign c32_42_io_in_0 = c53_271_io_out_2; // @[Multiplier.scala 90:41]
  assign c32_42_io_in_1 = c53_272_io_out_2; // @[Multiplier.scala 90:41]
  assign c32_42_io_in_2 = c53_273_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_491_io_in_0 = c53_278_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_491_io_in_1 = c53_279_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_491_io_in_2 = c53_280_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_491_io_in_3 = c53_281_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_491_io_in_4 = c53_489_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_492_io_in_0 = c32_23_io_out_0; // @[Multiplier.scala 80:35]
  assign c53_492_io_in_1 = c53_274_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_492_io_in_2 = c53_275_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_492_io_in_3 = c53_276_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_492_io_in_4 = c53_490_io_out_1; // @[Multiplier.scala 89:41]
  assign c22_55_io_in_0 = c53_277_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_55_io_in_1 = c32_22_io_out_1; // @[Multiplier.scala 81:41]
  assign c53_493_io_in_0 = c53_282_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_493_io_in_1 = c53_283_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_493_io_in_2 = c53_284_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_493_io_in_3 = c53_285_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_493_io_in_4 = c53_491_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_494_io_in_0 = c22_17_io_out_0; // @[Multiplier.scala 75:35]
  assign c53_494_io_in_1 = c53_278_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_494_io_in_2 = c53_279_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_494_io_in_3 = c53_280_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_494_io_in_4 = c53_492_io_out_1; // @[Multiplier.scala 89:41]
  assign c22_56_io_in_0 = c53_281_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_56_io_in_1 = c32_23_io_out_1; // @[Multiplier.scala 81:41]
  assign c53_495_io_in_0 = c53_286_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_495_io_in_1 = c53_287_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_495_io_in_2 = c53_288_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_495_io_in_3 = c53_289_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_495_io_in_4 = c53_493_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_496_io_in_0 = c22_18_io_out_0; // @[Multiplier.scala 75:35]
  assign c53_496_io_in_1 = c53_282_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_496_io_in_2 = c53_283_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_496_io_in_3 = c53_284_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_496_io_in_4 = c53_494_io_out_1; // @[Multiplier.scala 89:41]
  assign c22_57_io_in_0 = c53_285_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_57_io_in_1 = c22_17_io_out_1; // @[Multiplier.scala 76:41]
  assign c53_497_io_in_0 = c53_290_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_497_io_in_1 = c53_291_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_497_io_in_2 = c53_292_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_497_io_in_3 = c53_293_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_497_io_in_4 = c53_495_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_498_io_in_0 = pp_26[25]; // @[Multiplier.scala 60:38]
  assign c53_498_io_in_1 = c53_286_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_498_io_in_2 = c53_287_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_498_io_in_3 = c53_288_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_498_io_in_4 = c53_496_io_out_1; // @[Multiplier.scala 89:41]
  assign c22_58_io_in_0 = c53_289_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_58_io_in_1 = c22_18_io_out_1; // @[Multiplier.scala 76:41]
  assign c53_499_io_in_0 = c53_294_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_499_io_in_1 = c53_295_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_499_io_in_2 = c53_296_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_499_io_in_3 = c53_297_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_499_io_in_4 = c53_497_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_500_io_in_0 = pp_26[26]; // @[Multiplier.scala 60:38]
  assign c53_500_io_in_1 = c53_290_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_500_io_in_2 = c53_291_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_500_io_in_3 = c53_292_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_500_io_in_4 = c53_498_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_501_io_in_0 = c53_298_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_501_io_in_1 = c53_299_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_501_io_in_2 = c53_300_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_501_io_in_3 = c53_301_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_501_io_in_4 = c53_499_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_502_io_in_0 = c53_294_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_502_io_in_1 = c53_295_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_502_io_in_2 = c53_296_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_502_io_in_3 = c53_297_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_502_io_in_4 = c53_500_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_503_io_in_0 = c53_302_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_503_io_in_1 = c53_303_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_503_io_in_2 = c53_304_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_503_io_in_3 = c53_305_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_503_io_in_4 = c53_501_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_504_io_in_0 = c53_298_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_504_io_in_1 = c53_299_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_504_io_in_2 = c53_300_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_504_io_in_3 = c53_301_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_504_io_in_4 = c53_502_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_505_io_in_0 = c53_306_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_505_io_in_1 = c53_307_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_505_io_in_2 = c53_308_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_505_io_in_3 = c32_24_io_out_0; // @[Multiplier.scala 80:35]
  assign c53_505_io_in_4 = c53_503_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_506_io_in_0 = c53_305_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_506_io_in_1 = c53_302_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_506_io_in_2 = c53_303_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_506_io_in_3 = c53_304_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_506_io_in_4 = c53_504_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_507_io_in_0 = c53_309_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_507_io_in_1 = c53_310_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_507_io_in_2 = c53_311_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_507_io_in_3 = c32_25_io_out_0; // @[Multiplier.scala 80:35]
  assign c53_507_io_in_4 = c53_505_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_508_io_in_0 = c53_306_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_508_io_in_1 = c53_307_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_508_io_in_2 = c53_308_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_508_io_in_3 = c32_24_io_out_1; // @[Multiplier.scala 81:41]
  assign c53_508_io_in_4 = c53_506_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_509_io_in_0 = c53_312_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_509_io_in_1 = c53_313_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_509_io_in_2 = c53_314_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_509_io_in_3 = c22_19_io_out_0; // @[Multiplier.scala 75:35]
  assign c53_509_io_in_4 = c53_507_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_510_io_in_0 = c53_309_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_510_io_in_1 = c53_310_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_510_io_in_2 = c53_311_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_510_io_in_3 = c32_25_io_out_1; // @[Multiplier.scala 81:41]
  assign c53_510_io_in_4 = c53_508_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_511_io_in_0 = c53_315_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_511_io_in_1 = c53_316_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_511_io_in_2 = c53_317_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_511_io_in_3 = c22_20_io_out_0; // @[Multiplier.scala 75:35]
  assign c53_511_io_in_4 = c53_509_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_512_io_in_0 = c53_312_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_512_io_in_1 = c53_313_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_512_io_in_2 = c53_314_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_512_io_in_3 = c22_19_io_out_1; // @[Multiplier.scala 76:41]
  assign c53_512_io_in_4 = c53_510_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_513_io_in_0 = c53_318_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_513_io_in_1 = c53_319_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_513_io_in_2 = c53_320_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_513_io_in_3 = pp_26[33]; // @[Multiplier.scala 60:38]
  assign c53_513_io_in_4 = c53_511_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_514_io_in_0 = c53_315_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_514_io_in_1 = c53_316_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_514_io_in_2 = c53_317_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_514_io_in_3 = c22_20_io_out_1; // @[Multiplier.scala 76:41]
  assign c53_514_io_in_4 = c53_512_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_515_io_in_0 = c53_321_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_515_io_in_1 = c53_322_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_515_io_in_2 = c53_323_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_515_io_in_3 = pp_26[34]; // @[Multiplier.scala 60:38]
  assign c53_515_io_in_4 = c53_513_io_out_1; // @[Multiplier.scala 89:41]
  assign c32_43_io_in_0 = c53_318_io_out_2; // @[Multiplier.scala 90:41]
  assign c32_43_io_in_1 = c53_319_io_out_2; // @[Multiplier.scala 90:41]
  assign c32_43_io_in_2 = c53_320_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_516_io_in_0 = c53_324_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_516_io_in_1 = c53_325_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_516_io_in_2 = c53_326_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_516_io_in_3 = c53_321_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_516_io_in_4 = c53_515_io_out_1; // @[Multiplier.scala 89:41]
  assign c22_59_io_in_0 = c53_322_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_59_io_in_1 = c53_323_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_517_io_in_0 = c53_327_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_517_io_in_1 = c53_328_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_517_io_in_2 = c53_329_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_517_io_in_3 = c53_324_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_517_io_in_4 = c53_516_io_out_1; // @[Multiplier.scala 89:41]
  assign c22_60_io_in_0 = c53_325_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_60_io_in_1 = c53_326_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_518_io_in_0 = c53_330_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_518_io_in_1 = c53_331_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_518_io_in_2 = c32_26_io_out_0; // @[Multiplier.scala 80:35]
  assign c53_518_io_in_3 = c53_329_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_518_io_in_4 = c53_517_io_out_1; // @[Multiplier.scala 89:41]
  assign c32_44_io_in_0 = c53_327_io_out_2; // @[Multiplier.scala 90:41]
  assign c32_44_io_in_1 = c53_328_io_out_2; // @[Multiplier.scala 90:41]
  assign c32_44_io_in_2 = c53_329_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_519_io_in_0 = c53_332_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_519_io_in_1 = c53_333_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_519_io_in_2 = c32_27_io_out_0; // @[Multiplier.scala 80:35]
  assign c53_519_io_in_3 = c53_330_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_519_io_in_4 = c53_518_io_out_1; // @[Multiplier.scala 89:41]
  assign c22_61_io_in_0 = c53_331_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_61_io_in_1 = c32_26_io_out_1; // @[Multiplier.scala 81:41]
  assign c53_520_io_in_0 = c53_334_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_520_io_in_1 = c53_335_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_520_io_in_2 = c22_21_io_out_0; // @[Multiplier.scala 75:35]
  assign c53_520_io_in_3 = c53_332_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_520_io_in_4 = c53_519_io_out_1; // @[Multiplier.scala 89:41]
  assign c22_62_io_in_0 = c53_333_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_62_io_in_1 = c32_27_io_out_1; // @[Multiplier.scala 81:41]
  assign c53_521_io_in_0 = c53_336_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_521_io_in_1 = c53_337_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_521_io_in_2 = c22_22_io_out_0; // @[Multiplier.scala 75:35]
  assign c53_521_io_in_3 = c53_334_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_521_io_in_4 = c53_520_io_out_1; // @[Multiplier.scala 89:41]
  assign c22_63_io_in_0 = c53_335_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_63_io_in_1 = c22_21_io_out_1; // @[Multiplier.scala 76:41]
  assign c53_522_io_in_0 = c53_338_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_522_io_in_1 = c53_339_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_522_io_in_2 = pp_26[41]; // @[Multiplier.scala 60:38]
  assign c53_522_io_in_3 = c53_336_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_522_io_in_4 = c53_521_io_out_1; // @[Multiplier.scala 89:41]
  assign c22_64_io_in_0 = c53_337_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_64_io_in_1 = c22_22_io_out_1; // @[Multiplier.scala 76:41]
  assign c53_523_io_in_0 = c53_340_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_523_io_in_1 = c53_341_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_523_io_in_2 = pp_26[42]; // @[Multiplier.scala 60:38]
  assign c53_523_io_in_3 = c53_338_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_523_io_in_4 = c53_522_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_524_io_in_0 = c53_342_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_524_io_in_1 = c53_343_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_524_io_in_2 = c53_340_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_524_io_in_3 = c53_341_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_524_io_in_4 = c53_523_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_525_io_in_0 = c53_344_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_525_io_in_1 = c53_345_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_525_io_in_2 = c53_342_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_525_io_in_3 = c53_343_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_525_io_in_4 = c53_524_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_526_io_in_0 = c53_346_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_526_io_in_1 = c32_28_io_out_0; // @[Multiplier.scala 80:35]
  assign c53_526_io_in_2 = c53_345_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_526_io_in_3 = c53_344_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_526_io_in_4 = c53_525_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_527_io_in_0 = c53_347_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_527_io_in_1 = c32_29_io_out_0; // @[Multiplier.scala 80:35]
  assign c53_527_io_in_2 = c53_346_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_527_io_in_3 = c32_28_io_out_1; // @[Multiplier.scala 81:41]
  assign c53_527_io_in_4 = c53_526_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_528_io_in_0 = c53_348_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_528_io_in_1 = c22_23_io_out_0; // @[Multiplier.scala 75:35]
  assign c53_528_io_in_2 = c53_347_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_528_io_in_3 = c32_29_io_out_1; // @[Multiplier.scala 81:41]
  assign c53_528_io_in_4 = c53_527_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_529_io_in_0 = c53_349_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_529_io_in_1 = c22_24_io_out_0; // @[Multiplier.scala 75:35]
  assign c53_529_io_in_2 = c53_348_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_529_io_in_3 = c22_23_io_out_1; // @[Multiplier.scala 76:41]
  assign c53_529_io_in_4 = c53_528_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_530_io_in_0 = c53_350_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_530_io_in_1 = pp_26[49]; // @[Multiplier.scala 60:38]
  assign c53_530_io_in_2 = c53_349_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_530_io_in_3 = c22_24_io_out_1; // @[Multiplier.scala 76:41]
  assign c53_530_io_in_4 = c53_529_io_out_1; // @[Multiplier.scala 89:41]
  assign c32_45_io_in_0 = c53_351_io_out_0; // @[Multiplier.scala 88:39]
  assign c32_45_io_in_1 = pp_26[50]; // @[Multiplier.scala 60:38]
  assign c32_45_io_in_2 = c53_350_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_65_io_in_0 = c53_352_io_out_0; // @[Multiplier.scala 88:39]
  assign c22_65_io_in_1 = c53_351_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_66_io_in_0 = c53_353_io_out_0; // @[Multiplier.scala 88:39]
  assign c22_66_io_in_1 = c53_352_io_out_2; // @[Multiplier.scala 90:41]
  assign c32_46_io_in_0 = c32_30_io_out_0; // @[Multiplier.scala 80:35]
  assign c32_46_io_in_1 = c53_353_io_out_1; // @[Multiplier.scala 89:41]
  assign c32_46_io_in_2 = c53_353_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_67_io_in_0 = c32_31_io_out_0; // @[Multiplier.scala 80:35]
  assign c22_67_io_in_1 = c32_30_io_out_1; // @[Multiplier.scala 81:41]
  assign c22_68_io_in_0 = c22_25_io_out_0; // @[Multiplier.scala 75:35]
  assign c22_68_io_in_1 = c32_31_io_out_1; // @[Multiplier.scala 81:41]
  assign c22_69_io_in_0 = c22_26_io_out_0; // @[Multiplier.scala 75:35]
  assign c22_69_io_in_1 = c22_25_io_out_1; // @[Multiplier.scala 76:41]
  assign c22_70_io_in_0 = pp_26[57]; // @[Multiplier.scala 60:38]
  assign c22_70_io_in_1 = c22_26_io_out_1; // @[Multiplier.scala 76:41]
  assign c22_71_io_in_0 = r_2; // @[Multiplier.scala 74:19]
  assign c22_71_io_in_1 = r_3; // @[Multiplier.scala 74:19]
  assign c22_72_io_in_0 = r_4; // @[Multiplier.scala 74:19]
  assign c22_72_io_in_1 = r_5; // @[Multiplier.scala 74:19]
  assign c22_73_io_in_0 = r_6; // @[Multiplier.scala 74:19]
  assign c22_73_io_in_1 = r_7; // @[Multiplier.scala 74:19]
  assign c22_74_io_in_0 = r_8; // @[Multiplier.scala 74:19]
  assign c22_74_io_in_1 = r_9; // @[Multiplier.scala 74:19]
  assign c22_75_io_in_0 = r_10; // @[Multiplier.scala 74:19]
  assign c22_75_io_in_1 = r_11; // @[Multiplier.scala 74:19]
  assign c22_76_io_in_0 = r_12; // @[Multiplier.scala 74:19]
  assign c22_76_io_in_1 = r_13; // @[Multiplier.scala 74:19]
  assign c22_77_io_in_0 = r_14; // @[Multiplier.scala 74:19]
  assign c22_77_io_in_1 = r_15; // @[Multiplier.scala 74:19]
  assign c22_78_io_in_0 = r_16; // @[Multiplier.scala 74:19]
  assign c22_78_io_in_1 = r_17; // @[Multiplier.scala 74:19]
  assign c22_79_io_in_0 = r_18; // @[Multiplier.scala 74:19]
  assign c22_79_io_in_1 = r_19; // @[Multiplier.scala 74:19]
  assign c22_80_io_in_0 = r_20; // @[Multiplier.scala 74:19]
  assign c22_80_io_in_1 = r_21; // @[Multiplier.scala 74:19]
  assign c22_81_io_in_0 = r_22; // @[Multiplier.scala 74:19]
  assign c22_81_io_in_1 = r_23; // @[Multiplier.scala 74:19]
  assign c22_82_io_in_0 = r_24; // @[Multiplier.scala 74:19]
  assign c22_82_io_in_1 = r_25; // @[Multiplier.scala 74:19]
  assign c32_47_io_in_0 = r_26; // @[Multiplier.scala 79:19]
  assign c32_47_io_in_1 = r_27; // @[Multiplier.scala 79:19]
  assign c32_47_io_in_2 = r_28; // @[Multiplier.scala 79:19]
  assign c32_48_io_in_0 = r_29; // @[Multiplier.scala 79:19]
  assign c32_48_io_in_1 = r_30; // @[Multiplier.scala 79:19]
  assign c32_48_io_in_2 = r_31; // @[Multiplier.scala 79:19]
  assign c32_49_io_in_0 = r_32; // @[Multiplier.scala 79:19]
  assign c32_49_io_in_1 = r_33; // @[Multiplier.scala 79:19]
  assign c32_49_io_in_2 = r_34; // @[Multiplier.scala 79:19]
  assign c32_50_io_in_0 = r_35; // @[Multiplier.scala 79:19]
  assign c32_50_io_in_1 = r_36; // @[Multiplier.scala 79:19]
  assign c32_50_io_in_2 = r_37; // @[Multiplier.scala 79:19]
  assign c53_531_io_in_0 = r_38; // @[Multiplier.scala 85:13]
  assign c53_531_io_in_1 = r_39; // @[Multiplier.scala 85:13]
  assign c53_531_io_in_2 = r_40; // @[Multiplier.scala 85:13]
  assign c53_531_io_in_3 = r_41; // @[Multiplier.scala 85:13]
  assign c53_531_io_in_4 = 1'h0; // @[Multiplier.scala 87:24]
  assign c53_532_io_in_0 = r_42; // @[Multiplier.scala 85:13]
  assign c53_532_io_in_1 = r_43; // @[Multiplier.scala 85:13]
  assign c53_532_io_in_2 = r_44; // @[Multiplier.scala 85:13]
  assign c53_532_io_in_3 = r_45; // @[Multiplier.scala 85:13]
  assign c53_532_io_in_4 = c53_531_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_533_io_in_0 = r_46; // @[Multiplier.scala 85:13]
  assign c53_533_io_in_1 = r_47; // @[Multiplier.scala 85:13]
  assign c53_533_io_in_2 = r_48; // @[Multiplier.scala 85:13]
  assign c53_533_io_in_3 = r_49; // @[Multiplier.scala 85:13]
  assign c53_533_io_in_4 = c53_532_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_534_io_in_0 = r_50; // @[Multiplier.scala 85:13]
  assign c53_534_io_in_1 = r_51; // @[Multiplier.scala 85:13]
  assign c53_534_io_in_2 = r_52; // @[Multiplier.scala 85:13]
  assign c53_534_io_in_3 = r_53; // @[Multiplier.scala 85:13]
  assign c53_534_io_in_4 = c53_533_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_535_io_in_0 = r_54; // @[Multiplier.scala 85:13]
  assign c53_535_io_in_1 = r_55; // @[Multiplier.scala 85:13]
  assign c53_535_io_in_2 = r_56; // @[Multiplier.scala 85:13]
  assign c53_535_io_in_3 = r_57; // @[Multiplier.scala 85:13]
  assign c53_535_io_in_4 = c53_534_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_536_io_in_0 = r_58; // @[Multiplier.scala 85:13]
  assign c53_536_io_in_1 = r_59; // @[Multiplier.scala 85:13]
  assign c53_536_io_in_2 = r_60; // @[Multiplier.scala 85:13]
  assign c53_536_io_in_3 = r_61; // @[Multiplier.scala 85:13]
  assign c53_536_io_in_4 = c53_535_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_537_io_in_0 = r_62; // @[Multiplier.scala 85:13]
  assign c53_537_io_in_1 = r_63; // @[Multiplier.scala 85:13]
  assign c53_537_io_in_2 = r_64; // @[Multiplier.scala 85:13]
  assign c53_537_io_in_3 = r_65; // @[Multiplier.scala 85:13]
  assign c53_537_io_in_4 = c53_536_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_538_io_in_0 = r_66; // @[Multiplier.scala 85:13]
  assign c53_538_io_in_1 = r_67; // @[Multiplier.scala 85:13]
  assign c53_538_io_in_2 = r_68; // @[Multiplier.scala 85:13]
  assign c53_538_io_in_3 = r_69; // @[Multiplier.scala 85:13]
  assign c53_538_io_in_4 = c53_537_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_539_io_in_0 = r_70; // @[Multiplier.scala 85:13]
  assign c53_539_io_in_1 = r_71; // @[Multiplier.scala 85:13]
  assign c53_539_io_in_2 = r_72; // @[Multiplier.scala 85:13]
  assign c53_539_io_in_3 = r_73; // @[Multiplier.scala 85:13]
  assign c53_539_io_in_4 = c53_538_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_540_io_in_0 = r_74; // @[Multiplier.scala 85:13]
  assign c53_540_io_in_1 = r_75; // @[Multiplier.scala 85:13]
  assign c53_540_io_in_2 = r_76; // @[Multiplier.scala 85:13]
  assign c53_540_io_in_3 = r_77; // @[Multiplier.scala 85:13]
  assign c53_540_io_in_4 = c53_539_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_541_io_in_0 = r_78; // @[Multiplier.scala 85:13]
  assign c53_541_io_in_1 = r_79; // @[Multiplier.scala 85:13]
  assign c53_541_io_in_2 = r_80; // @[Multiplier.scala 85:13]
  assign c53_541_io_in_3 = r_81; // @[Multiplier.scala 85:13]
  assign c53_541_io_in_4 = c53_540_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_542_io_in_0 = r_82; // @[Multiplier.scala 85:13]
  assign c53_542_io_in_1 = r_83; // @[Multiplier.scala 85:13]
  assign c53_542_io_in_2 = r_84; // @[Multiplier.scala 85:13]
  assign c53_542_io_in_3 = r_85; // @[Multiplier.scala 85:13]
  assign c53_542_io_in_4 = c53_541_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_543_io_in_0 = r_86; // @[Multiplier.scala 85:13]
  assign c53_543_io_in_1 = r_87; // @[Multiplier.scala 85:13]
  assign c53_543_io_in_2 = r_88; // @[Multiplier.scala 85:13]
  assign c53_543_io_in_3 = r_89; // @[Multiplier.scala 85:13]
  assign c53_543_io_in_4 = c53_542_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_544_io_in_0 = r_91; // @[Multiplier.scala 85:13]
  assign c53_544_io_in_1 = r_92; // @[Multiplier.scala 85:13]
  assign c53_544_io_in_2 = r_93; // @[Multiplier.scala 85:13]
  assign c53_544_io_in_3 = r_94; // @[Multiplier.scala 85:13]
  assign c53_544_io_in_4 = c53_543_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_545_io_in_0 = r_96; // @[Multiplier.scala 85:13]
  assign c53_545_io_in_1 = r_97; // @[Multiplier.scala 85:13]
  assign c53_545_io_in_2 = r_98; // @[Multiplier.scala 85:13]
  assign c53_545_io_in_3 = r_99; // @[Multiplier.scala 85:13]
  assign c53_545_io_in_4 = c53_544_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_546_io_in_0 = r_101; // @[Multiplier.scala 85:13]
  assign c53_546_io_in_1 = r_102; // @[Multiplier.scala 85:13]
  assign c53_546_io_in_2 = r_103; // @[Multiplier.scala 85:13]
  assign c53_546_io_in_3 = r_104; // @[Multiplier.scala 85:13]
  assign c53_546_io_in_4 = c53_545_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_547_io_in_0 = r_106; // @[Multiplier.scala 85:13]
  assign c53_547_io_in_1 = r_107; // @[Multiplier.scala 85:13]
  assign c53_547_io_in_2 = r_108; // @[Multiplier.scala 85:13]
  assign c53_547_io_in_3 = r_109; // @[Multiplier.scala 85:13]
  assign c53_547_io_in_4 = c53_546_io_out_1; // @[Multiplier.scala 89:41]
  assign c22_83_io_in_0 = r_110; // @[Multiplier.scala 74:19]
  assign c22_83_io_in_1 = r_111; // @[Multiplier.scala 74:19]
  assign c53_548_io_in_0 = r_112; // @[Multiplier.scala 85:13]
  assign c53_548_io_in_1 = r_113; // @[Multiplier.scala 85:13]
  assign c53_548_io_in_2 = r_114; // @[Multiplier.scala 85:13]
  assign c53_548_io_in_3 = r_115; // @[Multiplier.scala 85:13]
  assign c53_548_io_in_4 = c53_547_io_out_1; // @[Multiplier.scala 89:41]
  assign c22_84_io_in_0 = r_116; // @[Multiplier.scala 74:19]
  assign c22_84_io_in_1 = r_117; // @[Multiplier.scala 74:19]
  assign c53_549_io_in_0 = r_118; // @[Multiplier.scala 85:13]
  assign c53_549_io_in_1 = r_119; // @[Multiplier.scala 85:13]
  assign c53_549_io_in_2 = r_120; // @[Multiplier.scala 85:13]
  assign c53_549_io_in_3 = r_121; // @[Multiplier.scala 85:13]
  assign c53_549_io_in_4 = c53_548_io_out_1; // @[Multiplier.scala 89:41]
  assign c22_85_io_in_0 = r_122; // @[Multiplier.scala 74:19]
  assign c22_85_io_in_1 = r_123; // @[Multiplier.scala 74:19]
  assign c53_550_io_in_0 = r_124; // @[Multiplier.scala 85:13]
  assign c53_550_io_in_1 = r_125; // @[Multiplier.scala 85:13]
  assign c53_550_io_in_2 = r_126; // @[Multiplier.scala 85:13]
  assign c53_550_io_in_3 = r_127; // @[Multiplier.scala 85:13]
  assign c53_550_io_in_4 = c53_549_io_out_1; // @[Multiplier.scala 89:41]
  assign c22_86_io_in_0 = r_128; // @[Multiplier.scala 74:19]
  assign c22_86_io_in_1 = r_129; // @[Multiplier.scala 74:19]
  assign c53_551_io_in_0 = r_130; // @[Multiplier.scala 85:13]
  assign c53_551_io_in_1 = r_131; // @[Multiplier.scala 85:13]
  assign c53_551_io_in_2 = r_132; // @[Multiplier.scala 85:13]
  assign c53_551_io_in_3 = r_133; // @[Multiplier.scala 85:13]
  assign c53_551_io_in_4 = c53_550_io_out_1; // @[Multiplier.scala 89:41]
  assign c22_87_io_in_0 = r_134; // @[Multiplier.scala 74:19]
  assign c22_87_io_in_1 = r_135; // @[Multiplier.scala 74:19]
  assign c53_552_io_in_0 = r_136; // @[Multiplier.scala 85:13]
  assign c53_552_io_in_1 = r_137; // @[Multiplier.scala 85:13]
  assign c53_552_io_in_2 = r_138; // @[Multiplier.scala 85:13]
  assign c53_552_io_in_3 = r_139; // @[Multiplier.scala 85:13]
  assign c53_552_io_in_4 = c53_551_io_out_1; // @[Multiplier.scala 89:41]
  assign c22_88_io_in_0 = r_140; // @[Multiplier.scala 74:19]
  assign c22_88_io_in_1 = r_141; // @[Multiplier.scala 74:19]
  assign c53_553_io_in_0 = r_142; // @[Multiplier.scala 85:13]
  assign c53_553_io_in_1 = r_143; // @[Multiplier.scala 85:13]
  assign c53_553_io_in_2 = r_144; // @[Multiplier.scala 85:13]
  assign c53_553_io_in_3 = r_145; // @[Multiplier.scala 85:13]
  assign c53_553_io_in_4 = c53_552_io_out_1; // @[Multiplier.scala 89:41]
  assign c22_89_io_in_0 = r_146; // @[Multiplier.scala 74:19]
  assign c22_89_io_in_1 = r_147; // @[Multiplier.scala 74:19]
  assign c53_554_io_in_0 = r_148; // @[Multiplier.scala 85:13]
  assign c53_554_io_in_1 = r_149; // @[Multiplier.scala 85:13]
  assign c53_554_io_in_2 = r_150; // @[Multiplier.scala 85:13]
  assign c53_554_io_in_3 = r_151; // @[Multiplier.scala 85:13]
  assign c53_554_io_in_4 = c53_553_io_out_1; // @[Multiplier.scala 89:41]
  assign c22_90_io_in_0 = r_152; // @[Multiplier.scala 74:19]
  assign c22_90_io_in_1 = r_153; // @[Multiplier.scala 74:19]
  assign c53_555_io_in_0 = r_154; // @[Multiplier.scala 85:13]
  assign c53_555_io_in_1 = r_155; // @[Multiplier.scala 85:13]
  assign c53_555_io_in_2 = r_156; // @[Multiplier.scala 85:13]
  assign c53_555_io_in_3 = r_157; // @[Multiplier.scala 85:13]
  assign c53_555_io_in_4 = c53_554_io_out_1; // @[Multiplier.scala 89:41]
  assign c22_91_io_in_0 = r_158; // @[Multiplier.scala 74:19]
  assign c22_91_io_in_1 = r_159; // @[Multiplier.scala 74:19]
  assign c53_556_io_in_0 = r_160; // @[Multiplier.scala 85:13]
  assign c53_556_io_in_1 = r_161; // @[Multiplier.scala 85:13]
  assign c53_556_io_in_2 = r_162; // @[Multiplier.scala 85:13]
  assign c53_556_io_in_3 = r_163; // @[Multiplier.scala 85:13]
  assign c53_556_io_in_4 = c53_555_io_out_1; // @[Multiplier.scala 89:41]
  assign c22_92_io_in_0 = r_164; // @[Multiplier.scala 74:19]
  assign c22_92_io_in_1 = r_165; // @[Multiplier.scala 74:19]
  assign c53_557_io_in_0 = r_166; // @[Multiplier.scala 85:13]
  assign c53_557_io_in_1 = r_167; // @[Multiplier.scala 85:13]
  assign c53_557_io_in_2 = r_168; // @[Multiplier.scala 85:13]
  assign c53_557_io_in_3 = r_169; // @[Multiplier.scala 85:13]
  assign c53_557_io_in_4 = c53_556_io_out_1; // @[Multiplier.scala 89:41]
  assign c22_93_io_in_0 = r_170; // @[Multiplier.scala 74:19]
  assign c22_93_io_in_1 = r_171; // @[Multiplier.scala 74:19]
  assign c53_558_io_in_0 = r_172; // @[Multiplier.scala 85:13]
  assign c53_558_io_in_1 = r_173; // @[Multiplier.scala 85:13]
  assign c53_558_io_in_2 = r_174; // @[Multiplier.scala 85:13]
  assign c53_558_io_in_3 = r_175; // @[Multiplier.scala 85:13]
  assign c53_558_io_in_4 = c53_557_io_out_1; // @[Multiplier.scala 89:41]
  assign c22_94_io_in_0 = r_176; // @[Multiplier.scala 74:19]
  assign c22_94_io_in_1 = r_177; // @[Multiplier.scala 74:19]
  assign c53_559_io_in_0 = r_178; // @[Multiplier.scala 85:13]
  assign c53_559_io_in_1 = r_179; // @[Multiplier.scala 85:13]
  assign c53_559_io_in_2 = r_180; // @[Multiplier.scala 85:13]
  assign c53_559_io_in_3 = r_181; // @[Multiplier.scala 85:13]
  assign c53_559_io_in_4 = c53_558_io_out_1; // @[Multiplier.scala 89:41]
  assign c32_51_io_in_0 = r_182; // @[Multiplier.scala 79:19]
  assign c32_51_io_in_1 = r_183; // @[Multiplier.scala 79:19]
  assign c32_51_io_in_2 = r_184; // @[Multiplier.scala 79:19]
  assign c53_560_io_in_0 = r_185; // @[Multiplier.scala 85:13]
  assign c53_560_io_in_1 = r_186; // @[Multiplier.scala 85:13]
  assign c53_560_io_in_2 = r_187; // @[Multiplier.scala 85:13]
  assign c53_560_io_in_3 = r_188; // @[Multiplier.scala 85:13]
  assign c53_560_io_in_4 = c53_559_io_out_1; // @[Multiplier.scala 89:41]
  assign c32_52_io_in_0 = r_189; // @[Multiplier.scala 79:19]
  assign c32_52_io_in_1 = r_190; // @[Multiplier.scala 79:19]
  assign c32_52_io_in_2 = r_191; // @[Multiplier.scala 79:19]
  assign c53_561_io_in_0 = r_192; // @[Multiplier.scala 85:13]
  assign c53_561_io_in_1 = r_193; // @[Multiplier.scala 85:13]
  assign c53_561_io_in_2 = r_194; // @[Multiplier.scala 85:13]
  assign c53_561_io_in_3 = r_195; // @[Multiplier.scala 85:13]
  assign c53_561_io_in_4 = c53_560_io_out_1; // @[Multiplier.scala 89:41]
  assign c32_53_io_in_0 = r_196; // @[Multiplier.scala 79:19]
  assign c32_53_io_in_1 = r_197; // @[Multiplier.scala 79:19]
  assign c32_53_io_in_2 = r_198; // @[Multiplier.scala 79:19]
  assign c53_562_io_in_0 = r_199; // @[Multiplier.scala 85:13]
  assign c53_562_io_in_1 = r_200; // @[Multiplier.scala 85:13]
  assign c53_562_io_in_2 = r_201; // @[Multiplier.scala 85:13]
  assign c53_562_io_in_3 = r_202; // @[Multiplier.scala 85:13]
  assign c53_562_io_in_4 = c53_561_io_out_1; // @[Multiplier.scala 89:41]
  assign c32_54_io_in_0 = r_203; // @[Multiplier.scala 79:19]
  assign c32_54_io_in_1 = r_204; // @[Multiplier.scala 79:19]
  assign c32_54_io_in_2 = r_205; // @[Multiplier.scala 79:19]
  assign c53_563_io_in_0 = r_206; // @[Multiplier.scala 85:13]
  assign c53_563_io_in_1 = r_207; // @[Multiplier.scala 85:13]
  assign c53_563_io_in_2 = r_208; // @[Multiplier.scala 85:13]
  assign c53_563_io_in_3 = r_209; // @[Multiplier.scala 85:13]
  assign c53_563_io_in_4 = c53_562_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_564_io_in_0 = r_210; // @[Multiplier.scala 85:13]
  assign c53_564_io_in_1 = r_211; // @[Multiplier.scala 85:13]
  assign c53_564_io_in_2 = r_212; // @[Multiplier.scala 85:13]
  assign c53_564_io_in_3 = r_213; // @[Multiplier.scala 85:13]
  assign c53_564_io_in_4 = 1'h0; // @[Multiplier.scala 87:24]
  assign c53_565_io_in_0 = r_214; // @[Multiplier.scala 85:13]
  assign c53_565_io_in_1 = r_215; // @[Multiplier.scala 85:13]
  assign c53_565_io_in_2 = r_216; // @[Multiplier.scala 85:13]
  assign c53_565_io_in_3 = r_217; // @[Multiplier.scala 85:13]
  assign c53_565_io_in_4 = c53_563_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_566_io_in_0 = r_218; // @[Multiplier.scala 85:13]
  assign c53_566_io_in_1 = r_219; // @[Multiplier.scala 85:13]
  assign c53_566_io_in_2 = r_220; // @[Multiplier.scala 85:13]
  assign c53_566_io_in_3 = r_221; // @[Multiplier.scala 85:13]
  assign c53_566_io_in_4 = c53_564_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_567_io_in_0 = r_222; // @[Multiplier.scala 85:13]
  assign c53_567_io_in_1 = r_223; // @[Multiplier.scala 85:13]
  assign c53_567_io_in_2 = r_224; // @[Multiplier.scala 85:13]
  assign c53_567_io_in_3 = r_225; // @[Multiplier.scala 85:13]
  assign c53_567_io_in_4 = c53_565_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_568_io_in_0 = r_226; // @[Multiplier.scala 85:13]
  assign c53_568_io_in_1 = r_227; // @[Multiplier.scala 85:13]
  assign c53_568_io_in_2 = r_228; // @[Multiplier.scala 85:13]
  assign c53_568_io_in_3 = r_229; // @[Multiplier.scala 85:13]
  assign c53_568_io_in_4 = c53_566_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_569_io_in_0 = r_230; // @[Multiplier.scala 85:13]
  assign c53_569_io_in_1 = r_231; // @[Multiplier.scala 85:13]
  assign c53_569_io_in_2 = r_232; // @[Multiplier.scala 85:13]
  assign c53_569_io_in_3 = r_233; // @[Multiplier.scala 85:13]
  assign c53_569_io_in_4 = c53_567_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_570_io_in_0 = r_234; // @[Multiplier.scala 85:13]
  assign c53_570_io_in_1 = r_235; // @[Multiplier.scala 85:13]
  assign c53_570_io_in_2 = r_236; // @[Multiplier.scala 85:13]
  assign c53_570_io_in_3 = r_237; // @[Multiplier.scala 85:13]
  assign c53_570_io_in_4 = c53_568_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_571_io_in_0 = r_238; // @[Multiplier.scala 85:13]
  assign c53_571_io_in_1 = r_239; // @[Multiplier.scala 85:13]
  assign c53_571_io_in_2 = r_240; // @[Multiplier.scala 85:13]
  assign c53_571_io_in_3 = r_241; // @[Multiplier.scala 85:13]
  assign c53_571_io_in_4 = c53_569_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_572_io_in_0 = r_242; // @[Multiplier.scala 85:13]
  assign c53_572_io_in_1 = r_243; // @[Multiplier.scala 85:13]
  assign c53_572_io_in_2 = r_244; // @[Multiplier.scala 85:13]
  assign c53_572_io_in_3 = r_245; // @[Multiplier.scala 85:13]
  assign c53_572_io_in_4 = c53_570_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_573_io_in_0 = r_246; // @[Multiplier.scala 85:13]
  assign c53_573_io_in_1 = r_247; // @[Multiplier.scala 85:13]
  assign c53_573_io_in_2 = r_248; // @[Multiplier.scala 85:13]
  assign c53_573_io_in_3 = r_249; // @[Multiplier.scala 85:13]
  assign c53_573_io_in_4 = c53_571_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_574_io_in_0 = r_250; // @[Multiplier.scala 85:13]
  assign c53_574_io_in_1 = r_251; // @[Multiplier.scala 85:13]
  assign c53_574_io_in_2 = r_252; // @[Multiplier.scala 85:13]
  assign c53_574_io_in_3 = r_253; // @[Multiplier.scala 85:13]
  assign c53_574_io_in_4 = c53_572_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_575_io_in_0 = r_254; // @[Multiplier.scala 85:13]
  assign c53_575_io_in_1 = r_255; // @[Multiplier.scala 85:13]
  assign c53_575_io_in_2 = r_256; // @[Multiplier.scala 85:13]
  assign c53_575_io_in_3 = r_257; // @[Multiplier.scala 85:13]
  assign c53_575_io_in_4 = c53_573_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_576_io_in_0 = r_258; // @[Multiplier.scala 85:13]
  assign c53_576_io_in_1 = r_259; // @[Multiplier.scala 85:13]
  assign c53_576_io_in_2 = r_260; // @[Multiplier.scala 85:13]
  assign c53_576_io_in_3 = r_261; // @[Multiplier.scala 85:13]
  assign c53_576_io_in_4 = c53_574_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_577_io_in_0 = r_262; // @[Multiplier.scala 85:13]
  assign c53_577_io_in_1 = r_263; // @[Multiplier.scala 85:13]
  assign c53_577_io_in_2 = r_264; // @[Multiplier.scala 85:13]
  assign c53_577_io_in_3 = r_265; // @[Multiplier.scala 85:13]
  assign c53_577_io_in_4 = c53_575_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_578_io_in_0 = r_266; // @[Multiplier.scala 85:13]
  assign c53_578_io_in_1 = r_267; // @[Multiplier.scala 85:13]
  assign c53_578_io_in_2 = r_268; // @[Multiplier.scala 85:13]
  assign c53_578_io_in_3 = r_269; // @[Multiplier.scala 85:13]
  assign c53_578_io_in_4 = c53_576_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_579_io_in_0 = r_270; // @[Multiplier.scala 85:13]
  assign c53_579_io_in_1 = r_271; // @[Multiplier.scala 85:13]
  assign c53_579_io_in_2 = r_272; // @[Multiplier.scala 85:13]
  assign c53_579_io_in_3 = r_273; // @[Multiplier.scala 85:13]
  assign c53_579_io_in_4 = c53_577_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_580_io_in_0 = r_274; // @[Multiplier.scala 85:13]
  assign c53_580_io_in_1 = r_275; // @[Multiplier.scala 85:13]
  assign c53_580_io_in_2 = r_276; // @[Multiplier.scala 85:13]
  assign c53_580_io_in_3 = r_277; // @[Multiplier.scala 85:13]
  assign c53_580_io_in_4 = c53_578_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_581_io_in_0 = r_278; // @[Multiplier.scala 85:13]
  assign c53_581_io_in_1 = r_279; // @[Multiplier.scala 85:13]
  assign c53_581_io_in_2 = r_280; // @[Multiplier.scala 85:13]
  assign c53_581_io_in_3 = r_281; // @[Multiplier.scala 85:13]
  assign c53_581_io_in_4 = c53_579_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_582_io_in_0 = r_282; // @[Multiplier.scala 85:13]
  assign c53_582_io_in_1 = r_283; // @[Multiplier.scala 85:13]
  assign c53_582_io_in_2 = r_284; // @[Multiplier.scala 85:13]
  assign c53_582_io_in_3 = r_285; // @[Multiplier.scala 85:13]
  assign c53_582_io_in_4 = c53_580_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_583_io_in_0 = r_286; // @[Multiplier.scala 85:13]
  assign c53_583_io_in_1 = r_287; // @[Multiplier.scala 85:13]
  assign c53_583_io_in_2 = r_288; // @[Multiplier.scala 85:13]
  assign c53_583_io_in_3 = r_289; // @[Multiplier.scala 85:13]
  assign c53_583_io_in_4 = c53_581_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_584_io_in_0 = r_290; // @[Multiplier.scala 85:13]
  assign c53_584_io_in_1 = r_291; // @[Multiplier.scala 85:13]
  assign c53_584_io_in_2 = r_292; // @[Multiplier.scala 85:13]
  assign c53_584_io_in_3 = r_293; // @[Multiplier.scala 85:13]
  assign c53_584_io_in_4 = c53_582_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_585_io_in_0 = r_294; // @[Multiplier.scala 85:13]
  assign c53_585_io_in_1 = r_295; // @[Multiplier.scala 85:13]
  assign c53_585_io_in_2 = r_296; // @[Multiplier.scala 85:13]
  assign c53_585_io_in_3 = r_297; // @[Multiplier.scala 85:13]
  assign c53_585_io_in_4 = c53_583_io_out_1; // @[Multiplier.scala 89:41]
  assign c22_95_io_in_0 = r_298; // @[Multiplier.scala 74:19]
  assign c22_95_io_in_1 = r_299; // @[Multiplier.scala 74:19]
  assign c53_586_io_in_0 = r_300; // @[Multiplier.scala 85:13]
  assign c53_586_io_in_1 = r_301; // @[Multiplier.scala 85:13]
  assign c53_586_io_in_2 = r_302; // @[Multiplier.scala 85:13]
  assign c53_586_io_in_3 = r_303; // @[Multiplier.scala 85:13]
  assign c53_586_io_in_4 = c53_585_io_out_1; // @[Multiplier.scala 89:41]
  assign c22_96_io_in_0 = r_304; // @[Multiplier.scala 74:19]
  assign c22_96_io_in_1 = r_305; // @[Multiplier.scala 74:19]
  assign c53_587_io_in_0 = r_306; // @[Multiplier.scala 85:13]
  assign c53_587_io_in_1 = r_307; // @[Multiplier.scala 85:13]
  assign c53_587_io_in_2 = r_308; // @[Multiplier.scala 85:13]
  assign c53_587_io_in_3 = r_309; // @[Multiplier.scala 85:13]
  assign c53_587_io_in_4 = c53_586_io_out_1; // @[Multiplier.scala 89:41]
  assign c32_55_io_in_0 = r_310; // @[Multiplier.scala 79:19]
  assign c32_55_io_in_1 = r_311; // @[Multiplier.scala 79:19]
  assign c32_55_io_in_2 = r_312; // @[Multiplier.scala 79:19]
  assign c53_588_io_in_0 = r_313; // @[Multiplier.scala 85:13]
  assign c53_588_io_in_1 = r_314; // @[Multiplier.scala 85:13]
  assign c53_588_io_in_2 = r_315; // @[Multiplier.scala 85:13]
  assign c53_588_io_in_3 = r_316; // @[Multiplier.scala 85:13]
  assign c53_588_io_in_4 = c53_587_io_out_1; // @[Multiplier.scala 89:41]
  assign c22_97_io_in_0 = r_317; // @[Multiplier.scala 74:19]
  assign c22_97_io_in_1 = r_318; // @[Multiplier.scala 74:19]
  assign c53_589_io_in_0 = r_319; // @[Multiplier.scala 85:13]
  assign c53_589_io_in_1 = r_320; // @[Multiplier.scala 85:13]
  assign c53_589_io_in_2 = r_321; // @[Multiplier.scala 85:13]
  assign c53_589_io_in_3 = r_322; // @[Multiplier.scala 85:13]
  assign c53_589_io_in_4 = c53_588_io_out_1; // @[Multiplier.scala 89:41]
  assign c22_98_io_in_0 = r_323; // @[Multiplier.scala 74:19]
  assign c22_98_io_in_1 = r_324; // @[Multiplier.scala 74:19]
  assign c53_590_io_in_0 = r_325; // @[Multiplier.scala 85:13]
  assign c53_590_io_in_1 = r_326; // @[Multiplier.scala 85:13]
  assign c53_590_io_in_2 = r_327; // @[Multiplier.scala 85:13]
  assign c53_590_io_in_3 = r_328; // @[Multiplier.scala 85:13]
  assign c53_590_io_in_4 = c53_589_io_out_1; // @[Multiplier.scala 89:41]
  assign c22_99_io_in_0 = r_329; // @[Multiplier.scala 74:19]
  assign c22_99_io_in_1 = r_330; // @[Multiplier.scala 74:19]
  assign c53_591_io_in_0 = r_331; // @[Multiplier.scala 85:13]
  assign c53_591_io_in_1 = r_332; // @[Multiplier.scala 85:13]
  assign c53_591_io_in_2 = r_333; // @[Multiplier.scala 85:13]
  assign c53_591_io_in_3 = r_334; // @[Multiplier.scala 85:13]
  assign c53_591_io_in_4 = c53_590_io_out_1; // @[Multiplier.scala 89:41]
  assign c22_100_io_in_0 = r_335; // @[Multiplier.scala 74:19]
  assign c22_100_io_in_1 = r_336; // @[Multiplier.scala 74:19]
  assign c53_592_io_in_0 = r_337; // @[Multiplier.scala 85:13]
  assign c53_592_io_in_1 = r_338; // @[Multiplier.scala 85:13]
  assign c53_592_io_in_2 = r_339; // @[Multiplier.scala 85:13]
  assign c53_592_io_in_3 = r_340; // @[Multiplier.scala 85:13]
  assign c53_592_io_in_4 = c53_591_io_out_1; // @[Multiplier.scala 89:41]
  assign c32_56_io_in_0 = r_341; // @[Multiplier.scala 79:19]
  assign c32_56_io_in_1 = r_342; // @[Multiplier.scala 79:19]
  assign c32_56_io_in_2 = r_343; // @[Multiplier.scala 79:19]
  assign c53_593_io_in_0 = r_344; // @[Multiplier.scala 85:13]
  assign c53_593_io_in_1 = r_345; // @[Multiplier.scala 85:13]
  assign c53_593_io_in_2 = r_346; // @[Multiplier.scala 85:13]
  assign c53_593_io_in_3 = r_347; // @[Multiplier.scala 85:13]
  assign c53_593_io_in_4 = c53_592_io_out_1; // @[Multiplier.scala 89:41]
  assign c22_101_io_in_0 = r_348; // @[Multiplier.scala 74:19]
  assign c22_101_io_in_1 = r_349; // @[Multiplier.scala 74:19]
  assign c53_594_io_in_0 = r_350; // @[Multiplier.scala 85:13]
  assign c53_594_io_in_1 = r_351; // @[Multiplier.scala 85:13]
  assign c53_594_io_in_2 = r_352; // @[Multiplier.scala 85:13]
  assign c53_594_io_in_3 = r_353; // @[Multiplier.scala 85:13]
  assign c53_594_io_in_4 = c53_593_io_out_1; // @[Multiplier.scala 89:41]
  assign c22_102_io_in_0 = r_354; // @[Multiplier.scala 74:19]
  assign c22_102_io_in_1 = r_355; // @[Multiplier.scala 74:19]
  assign c53_595_io_in_0 = r_356; // @[Multiplier.scala 85:13]
  assign c53_595_io_in_1 = r_357; // @[Multiplier.scala 85:13]
  assign c53_595_io_in_2 = r_358; // @[Multiplier.scala 85:13]
  assign c53_595_io_in_3 = r_359; // @[Multiplier.scala 85:13]
  assign c53_595_io_in_4 = c53_594_io_out_1; // @[Multiplier.scala 89:41]
  assign c22_103_io_in_0 = r_360; // @[Multiplier.scala 74:19]
  assign c22_103_io_in_1 = r_361; // @[Multiplier.scala 74:19]
  assign c53_596_io_in_0 = r_362; // @[Multiplier.scala 85:13]
  assign c53_596_io_in_1 = r_363; // @[Multiplier.scala 85:13]
  assign c53_596_io_in_2 = r_364; // @[Multiplier.scala 85:13]
  assign c53_596_io_in_3 = r_365; // @[Multiplier.scala 85:13]
  assign c53_596_io_in_4 = c53_595_io_out_1; // @[Multiplier.scala 89:41]
  assign c22_104_io_in_0 = r_366; // @[Multiplier.scala 74:19]
  assign c22_104_io_in_1 = r_367; // @[Multiplier.scala 74:19]
  assign c53_597_io_in_0 = r_368; // @[Multiplier.scala 85:13]
  assign c53_597_io_in_1 = r_369; // @[Multiplier.scala 85:13]
  assign c53_597_io_in_2 = r_370; // @[Multiplier.scala 85:13]
  assign c53_597_io_in_3 = r_371; // @[Multiplier.scala 85:13]
  assign c53_597_io_in_4 = c53_596_io_out_1; // @[Multiplier.scala 89:41]
  assign c22_105_io_in_0 = r_372; // @[Multiplier.scala 74:19]
  assign c22_105_io_in_1 = r_373; // @[Multiplier.scala 74:19]
  assign c53_598_io_in_0 = r_374; // @[Multiplier.scala 85:13]
  assign c53_598_io_in_1 = r_375; // @[Multiplier.scala 85:13]
  assign c53_598_io_in_2 = r_376; // @[Multiplier.scala 85:13]
  assign c53_598_io_in_3 = r_377; // @[Multiplier.scala 85:13]
  assign c53_598_io_in_4 = c53_597_io_out_1; // @[Multiplier.scala 89:41]
  assign c22_106_io_in_0 = r_378; // @[Multiplier.scala 74:19]
  assign c22_106_io_in_1 = r_379; // @[Multiplier.scala 74:19]
  assign c53_599_io_in_0 = r_380; // @[Multiplier.scala 85:13]
  assign c53_599_io_in_1 = r_381; // @[Multiplier.scala 85:13]
  assign c53_599_io_in_2 = r_382; // @[Multiplier.scala 85:13]
  assign c53_599_io_in_3 = r_383; // @[Multiplier.scala 85:13]
  assign c53_599_io_in_4 = c53_598_io_out_1; // @[Multiplier.scala 89:41]
  assign c22_107_io_in_0 = r_384; // @[Multiplier.scala 74:19]
  assign c22_107_io_in_1 = r_385; // @[Multiplier.scala 74:19]
  assign c53_600_io_in_0 = r_386; // @[Multiplier.scala 85:13]
  assign c53_600_io_in_1 = r_387; // @[Multiplier.scala 85:13]
  assign c53_600_io_in_2 = r_388; // @[Multiplier.scala 85:13]
  assign c53_600_io_in_3 = r_389; // @[Multiplier.scala 85:13]
  assign c53_600_io_in_4 = c53_599_io_out_1; // @[Multiplier.scala 89:41]
  assign c22_108_io_in_0 = r_390; // @[Multiplier.scala 74:19]
  assign c22_108_io_in_1 = r_391; // @[Multiplier.scala 74:19]
  assign c53_601_io_in_0 = r_392; // @[Multiplier.scala 85:13]
  assign c53_601_io_in_1 = r_393; // @[Multiplier.scala 85:13]
  assign c53_601_io_in_2 = r_394; // @[Multiplier.scala 85:13]
  assign c53_601_io_in_3 = r_395; // @[Multiplier.scala 85:13]
  assign c53_601_io_in_4 = c53_600_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_602_io_in_0 = r_396; // @[Multiplier.scala 85:13]
  assign c53_602_io_in_1 = r_397; // @[Multiplier.scala 85:13]
  assign c53_602_io_in_2 = r_398; // @[Multiplier.scala 85:13]
  assign c53_602_io_in_3 = r_399; // @[Multiplier.scala 85:13]
  assign c53_602_io_in_4 = c53_601_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_603_io_in_0 = r_400; // @[Multiplier.scala 85:13]
  assign c53_603_io_in_1 = r_401; // @[Multiplier.scala 85:13]
  assign c53_603_io_in_2 = r_402; // @[Multiplier.scala 85:13]
  assign c53_603_io_in_3 = r_403; // @[Multiplier.scala 85:13]
  assign c53_603_io_in_4 = c53_602_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_604_io_in_0 = r_405; // @[Multiplier.scala 85:13]
  assign c53_604_io_in_1 = r_406; // @[Multiplier.scala 85:13]
  assign c53_604_io_in_2 = r_407; // @[Multiplier.scala 85:13]
  assign c53_604_io_in_3 = r_408; // @[Multiplier.scala 85:13]
  assign c53_604_io_in_4 = c53_603_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_605_io_in_0 = r_409; // @[Multiplier.scala 85:13]
  assign c53_605_io_in_1 = r_410; // @[Multiplier.scala 85:13]
  assign c53_605_io_in_2 = r_411; // @[Multiplier.scala 85:13]
  assign c53_605_io_in_3 = r_412; // @[Multiplier.scala 85:13]
  assign c53_605_io_in_4 = c53_604_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_606_io_in_0 = r_413; // @[Multiplier.scala 85:13]
  assign c53_606_io_in_1 = r_414; // @[Multiplier.scala 85:13]
  assign c53_606_io_in_2 = r_415; // @[Multiplier.scala 85:13]
  assign c53_606_io_in_3 = r_416; // @[Multiplier.scala 85:13]
  assign c53_606_io_in_4 = c53_605_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_607_io_in_0 = r_417; // @[Multiplier.scala 85:13]
  assign c53_607_io_in_1 = r_418; // @[Multiplier.scala 85:13]
  assign c53_607_io_in_2 = r_419; // @[Multiplier.scala 85:13]
  assign c53_607_io_in_3 = r_420; // @[Multiplier.scala 85:13]
  assign c53_607_io_in_4 = c53_606_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_608_io_in_0 = r_421; // @[Multiplier.scala 85:13]
  assign c53_608_io_in_1 = r_422; // @[Multiplier.scala 85:13]
  assign c53_608_io_in_2 = r_423; // @[Multiplier.scala 85:13]
  assign c53_608_io_in_3 = r_424; // @[Multiplier.scala 85:13]
  assign c53_608_io_in_4 = c53_607_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_609_io_in_0 = r_426; // @[Multiplier.scala 85:13]
  assign c53_609_io_in_1 = r_427; // @[Multiplier.scala 85:13]
  assign c53_609_io_in_2 = r_428; // @[Multiplier.scala 85:13]
  assign c53_609_io_in_3 = r_429; // @[Multiplier.scala 85:13]
  assign c53_609_io_in_4 = c53_608_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_610_io_in_0 = r_430; // @[Multiplier.scala 85:13]
  assign c53_610_io_in_1 = r_431; // @[Multiplier.scala 85:13]
  assign c53_610_io_in_2 = r_432; // @[Multiplier.scala 85:13]
  assign c53_610_io_in_3 = r_433; // @[Multiplier.scala 85:13]
  assign c53_610_io_in_4 = c53_609_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_611_io_in_0 = r_434; // @[Multiplier.scala 85:13]
  assign c53_611_io_in_1 = r_435; // @[Multiplier.scala 85:13]
  assign c53_611_io_in_2 = r_436; // @[Multiplier.scala 85:13]
  assign c53_611_io_in_3 = r_437; // @[Multiplier.scala 85:13]
  assign c53_611_io_in_4 = c53_610_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_612_io_in_0 = r_438; // @[Multiplier.scala 85:13]
  assign c53_612_io_in_1 = r_439; // @[Multiplier.scala 85:13]
  assign c53_612_io_in_2 = r_440; // @[Multiplier.scala 85:13]
  assign c53_612_io_in_3 = r_441; // @[Multiplier.scala 85:13]
  assign c53_612_io_in_4 = c53_611_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_613_io_in_0 = r_442; // @[Multiplier.scala 85:13]
  assign c53_613_io_in_1 = r_443; // @[Multiplier.scala 85:13]
  assign c53_613_io_in_2 = r_444; // @[Multiplier.scala 85:13]
  assign c53_613_io_in_3 = r_445; // @[Multiplier.scala 85:13]
  assign c53_613_io_in_4 = c53_612_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_614_io_in_0 = r_446; // @[Multiplier.scala 85:13]
  assign c53_614_io_in_1 = r_447; // @[Multiplier.scala 85:13]
  assign c53_614_io_in_2 = r_448; // @[Multiplier.scala 85:13]
  assign c53_614_io_in_3 = r_449; // @[Multiplier.scala 85:13]
  assign c53_614_io_in_4 = c53_613_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_615_io_in_0 = r_450; // @[Multiplier.scala 85:13]
  assign c53_615_io_in_1 = r_451; // @[Multiplier.scala 85:13]
  assign c53_615_io_in_2 = r_452; // @[Multiplier.scala 85:13]
  assign c53_615_io_in_3 = r_453; // @[Multiplier.scala 85:13]
  assign c53_615_io_in_4 = c53_614_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_616_io_in_0 = r_454; // @[Multiplier.scala 85:13]
  assign c53_616_io_in_1 = r_455; // @[Multiplier.scala 85:13]
  assign c53_616_io_in_2 = r_456; // @[Multiplier.scala 85:13]
  assign c53_616_io_in_3 = r_457; // @[Multiplier.scala 85:13]
  assign c53_616_io_in_4 = c53_615_io_out_1; // @[Multiplier.scala 89:41]
  assign c22_109_io_in_0 = r_458; // @[Multiplier.scala 74:19]
  assign c22_109_io_in_1 = r_459; // @[Multiplier.scala 74:19]
  assign c22_110_io_in_0 = r_460; // @[Multiplier.scala 74:19]
  assign c22_110_io_in_1 = r_461; // @[Multiplier.scala 74:19]
  assign c32_57_io_in_0 = r_462; // @[Multiplier.scala 79:19]
  assign c32_57_io_in_1 = r_463; // @[Multiplier.scala 79:19]
  assign c32_57_io_in_2 = r_464; // @[Multiplier.scala 79:19]
  assign c22_111_io_in_0 = r_465; // @[Multiplier.scala 74:19]
  assign c22_111_io_in_1 = r_466; // @[Multiplier.scala 74:19]
  assign c22_112_io_in_0 = r_467; // @[Multiplier.scala 74:19]
  assign c22_112_io_in_1 = r_468; // @[Multiplier.scala 74:19]
  assign c22_113_io_in_0 = r_469; // @[Multiplier.scala 74:19]
  assign c22_113_io_in_1 = r_470; // @[Multiplier.scala 74:19]
  assign c22_114_io_in_0 = r_471; // @[Multiplier.scala 74:19]
  assign c22_114_io_in_1 = r_472; // @[Multiplier.scala 74:19]
  assign c32_58_io_in_0 = r_473; // @[Multiplier.scala 79:19]
  assign c32_58_io_in_1 = r_474; // @[Multiplier.scala 79:19]
  assign c32_58_io_in_2 = r_475; // @[Multiplier.scala 79:19]
  assign c22_115_io_in_0 = r_476; // @[Multiplier.scala 74:19]
  assign c22_115_io_in_1 = r_477; // @[Multiplier.scala 74:19]
  assign c22_116_io_in_0 = r_478; // @[Multiplier.scala 74:19]
  assign c22_116_io_in_1 = r_479; // @[Multiplier.scala 74:19]
  assign c22_117_io_in_0 = r_480; // @[Multiplier.scala 74:19]
  assign c22_117_io_in_1 = r_481; // @[Multiplier.scala 74:19]
  assign c22_118_io_in_0 = r_482; // @[Multiplier.scala 74:19]
  assign c22_118_io_in_1 = r_483; // @[Multiplier.scala 74:19]
  assign c22_119_io_in_0 = r_484; // @[Multiplier.scala 74:19]
  assign c22_119_io_in_1 = r_485; // @[Multiplier.scala 74:19]
  assign c22_120_io_in_0 = r_486; // @[Multiplier.scala 74:19]
  assign c22_120_io_in_1 = r_487; // @[Multiplier.scala 74:19]
  assign c22_121_io_in_0 = r_488; // @[Multiplier.scala 74:19]
  assign c22_121_io_in_1 = r_489; // @[Multiplier.scala 74:19]
  assign c22_122_io_in_0 = c22_72_io_out_0; // @[Multiplier.scala 75:35]
  assign c22_122_io_in_1 = c22_71_io_out_1; // @[Multiplier.scala 76:41]
  assign c22_123_io_in_0 = c22_73_io_out_0; // @[Multiplier.scala 75:35]
  assign c22_123_io_in_1 = c22_72_io_out_1; // @[Multiplier.scala 76:41]
  assign c22_124_io_in_0 = c22_74_io_out_0; // @[Multiplier.scala 75:35]
  assign c22_124_io_in_1 = c22_73_io_out_1; // @[Multiplier.scala 76:41]
  assign c22_125_io_in_0 = c22_75_io_out_0; // @[Multiplier.scala 75:35]
  assign c22_125_io_in_1 = c22_74_io_out_1; // @[Multiplier.scala 76:41]
  assign c22_126_io_in_0 = c22_76_io_out_0; // @[Multiplier.scala 75:35]
  assign c22_126_io_in_1 = c22_75_io_out_1; // @[Multiplier.scala 76:41]
  assign c22_127_io_in_0 = c22_77_io_out_0; // @[Multiplier.scala 75:35]
  assign c22_127_io_in_1 = c22_76_io_out_1; // @[Multiplier.scala 76:41]
  assign c22_128_io_in_0 = c22_78_io_out_0; // @[Multiplier.scala 75:35]
  assign c22_128_io_in_1 = c22_77_io_out_1; // @[Multiplier.scala 76:41]
  assign c22_129_io_in_0 = c22_79_io_out_0; // @[Multiplier.scala 75:35]
  assign c22_129_io_in_1 = c22_78_io_out_1; // @[Multiplier.scala 76:41]
  assign c22_130_io_in_0 = c22_80_io_out_0; // @[Multiplier.scala 75:35]
  assign c22_130_io_in_1 = c22_79_io_out_1; // @[Multiplier.scala 76:41]
  assign c22_131_io_in_0 = c22_81_io_out_0; // @[Multiplier.scala 75:35]
  assign c22_131_io_in_1 = c22_80_io_out_1; // @[Multiplier.scala 76:41]
  assign c22_132_io_in_0 = c22_82_io_out_0; // @[Multiplier.scala 75:35]
  assign c22_132_io_in_1 = c22_81_io_out_1; // @[Multiplier.scala 76:41]
  assign c22_133_io_in_0 = c32_47_io_out_0; // @[Multiplier.scala 80:35]
  assign c22_133_io_in_1 = c22_82_io_out_1; // @[Multiplier.scala 76:41]
  assign c22_134_io_in_0 = c32_48_io_out_0; // @[Multiplier.scala 80:35]
  assign c22_134_io_in_1 = c32_47_io_out_1; // @[Multiplier.scala 81:41]
  assign c22_135_io_in_0 = c32_49_io_out_0; // @[Multiplier.scala 80:35]
  assign c22_135_io_in_1 = c32_48_io_out_1; // @[Multiplier.scala 81:41]
  assign c22_136_io_in_0 = c32_50_io_out_0; // @[Multiplier.scala 80:35]
  assign c22_136_io_in_1 = c32_49_io_out_1; // @[Multiplier.scala 81:41]
  assign c22_137_io_in_0 = c53_531_io_out_0; // @[Multiplier.scala 88:39]
  assign c22_137_io_in_1 = c32_50_io_out_1; // @[Multiplier.scala 81:41]
  assign c22_138_io_in_0 = c53_532_io_out_0; // @[Multiplier.scala 88:39]
  assign c22_138_io_in_1 = c53_531_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_139_io_in_0 = c53_533_io_out_0; // @[Multiplier.scala 88:39]
  assign c22_139_io_in_1 = c53_532_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_140_io_in_0 = c53_534_io_out_0; // @[Multiplier.scala 88:39]
  assign c22_140_io_in_1 = c53_533_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_141_io_in_0 = c53_535_io_out_0; // @[Multiplier.scala 88:39]
  assign c22_141_io_in_1 = c53_534_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_142_io_in_0 = c53_536_io_out_0; // @[Multiplier.scala 88:39]
  assign c22_142_io_in_1 = c53_535_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_143_io_in_0 = c53_537_io_out_0; // @[Multiplier.scala 88:39]
  assign c22_143_io_in_1 = c53_536_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_144_io_in_0 = c53_538_io_out_0; // @[Multiplier.scala 88:39]
  assign c22_144_io_in_1 = c53_537_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_145_io_in_0 = c53_539_io_out_0; // @[Multiplier.scala 88:39]
  assign c22_145_io_in_1 = c53_538_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_146_io_in_0 = c53_540_io_out_0; // @[Multiplier.scala 88:39]
  assign c22_146_io_in_1 = c53_539_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_147_io_in_0 = c53_541_io_out_0; // @[Multiplier.scala 88:39]
  assign c22_147_io_in_1 = c53_540_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_148_io_in_0 = c53_542_io_out_0; // @[Multiplier.scala 88:39]
  assign c22_148_io_in_1 = c53_541_io_out_2; // @[Multiplier.scala 90:41]
  assign c32_59_io_in_0 = c53_543_io_out_0; // @[Multiplier.scala 88:39]
  assign c32_59_io_in_1 = r_90; // @[Multiplier.scala 79:19]
  assign c32_59_io_in_2 = c53_542_io_out_2; // @[Multiplier.scala 90:41]
  assign c32_60_io_in_0 = c53_544_io_out_0; // @[Multiplier.scala 88:39]
  assign c32_60_io_in_1 = r_95; // @[Multiplier.scala 79:19]
  assign c32_60_io_in_2 = c53_543_io_out_2; // @[Multiplier.scala 90:41]
  assign c32_61_io_in_0 = c53_545_io_out_0; // @[Multiplier.scala 88:39]
  assign c32_61_io_in_1 = r_100; // @[Multiplier.scala 79:19]
  assign c32_61_io_in_2 = c53_544_io_out_2; // @[Multiplier.scala 90:41]
  assign c32_62_io_in_0 = c53_546_io_out_0; // @[Multiplier.scala 88:39]
  assign c32_62_io_in_1 = r_105; // @[Multiplier.scala 79:19]
  assign c32_62_io_in_2 = c53_545_io_out_2; // @[Multiplier.scala 90:41]
  assign c32_63_io_in_0 = c53_547_io_out_0; // @[Multiplier.scala 88:39]
  assign c32_63_io_in_1 = c22_83_io_out_0; // @[Multiplier.scala 75:35]
  assign c32_63_io_in_2 = c53_546_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_617_io_in_0 = c53_548_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_617_io_in_1 = c22_84_io_out_0; // @[Multiplier.scala 75:35]
  assign c53_617_io_in_2 = c53_547_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_617_io_in_3 = c22_83_io_out_1; // @[Multiplier.scala 76:41]
  assign c53_617_io_in_4 = 1'h0; // @[Multiplier.scala 87:24]
  assign c53_618_io_in_0 = c53_549_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_618_io_in_1 = c22_85_io_out_0; // @[Multiplier.scala 75:35]
  assign c53_618_io_in_2 = c53_548_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_618_io_in_3 = c22_84_io_out_1; // @[Multiplier.scala 76:41]
  assign c53_618_io_in_4 = c53_617_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_619_io_in_0 = c53_550_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_619_io_in_1 = c22_86_io_out_0; // @[Multiplier.scala 75:35]
  assign c53_619_io_in_2 = c53_549_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_619_io_in_3 = c22_85_io_out_1; // @[Multiplier.scala 76:41]
  assign c53_619_io_in_4 = c53_618_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_620_io_in_0 = c53_551_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_620_io_in_1 = c22_87_io_out_0; // @[Multiplier.scala 75:35]
  assign c53_620_io_in_2 = c53_550_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_620_io_in_3 = c22_86_io_out_1; // @[Multiplier.scala 76:41]
  assign c53_620_io_in_4 = c53_619_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_621_io_in_0 = c53_552_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_621_io_in_1 = c22_88_io_out_0; // @[Multiplier.scala 75:35]
  assign c53_621_io_in_2 = c53_551_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_621_io_in_3 = c22_87_io_out_1; // @[Multiplier.scala 76:41]
  assign c53_621_io_in_4 = c53_620_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_622_io_in_0 = c53_553_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_622_io_in_1 = c22_89_io_out_0; // @[Multiplier.scala 75:35]
  assign c53_622_io_in_2 = c53_552_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_622_io_in_3 = c22_88_io_out_1; // @[Multiplier.scala 76:41]
  assign c53_622_io_in_4 = c53_621_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_623_io_in_0 = c53_554_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_623_io_in_1 = c22_90_io_out_0; // @[Multiplier.scala 75:35]
  assign c53_623_io_in_2 = c53_553_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_623_io_in_3 = c22_89_io_out_1; // @[Multiplier.scala 76:41]
  assign c53_623_io_in_4 = c53_622_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_624_io_in_0 = c53_555_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_624_io_in_1 = c22_91_io_out_0; // @[Multiplier.scala 75:35]
  assign c53_624_io_in_2 = c53_554_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_624_io_in_3 = c22_90_io_out_1; // @[Multiplier.scala 76:41]
  assign c53_624_io_in_4 = c53_623_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_625_io_in_0 = c53_556_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_625_io_in_1 = c22_92_io_out_0; // @[Multiplier.scala 75:35]
  assign c53_625_io_in_2 = c53_555_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_625_io_in_3 = c22_91_io_out_1; // @[Multiplier.scala 76:41]
  assign c53_625_io_in_4 = c53_624_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_626_io_in_0 = c53_557_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_626_io_in_1 = c22_93_io_out_0; // @[Multiplier.scala 75:35]
  assign c53_626_io_in_2 = c53_556_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_626_io_in_3 = c22_92_io_out_1; // @[Multiplier.scala 76:41]
  assign c53_626_io_in_4 = c53_625_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_627_io_in_0 = c53_558_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_627_io_in_1 = c22_94_io_out_0; // @[Multiplier.scala 75:35]
  assign c53_627_io_in_2 = c53_557_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_627_io_in_3 = c22_93_io_out_1; // @[Multiplier.scala 76:41]
  assign c53_627_io_in_4 = c53_626_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_628_io_in_0 = c53_559_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_628_io_in_1 = c32_51_io_out_0; // @[Multiplier.scala 80:35]
  assign c53_628_io_in_2 = c53_558_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_628_io_in_3 = c22_94_io_out_1; // @[Multiplier.scala 76:41]
  assign c53_628_io_in_4 = c53_627_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_629_io_in_0 = c53_560_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_629_io_in_1 = c32_52_io_out_0; // @[Multiplier.scala 80:35]
  assign c53_629_io_in_2 = c53_559_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_629_io_in_3 = c32_51_io_out_1; // @[Multiplier.scala 81:41]
  assign c53_629_io_in_4 = c53_628_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_630_io_in_0 = c53_561_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_630_io_in_1 = c32_53_io_out_0; // @[Multiplier.scala 80:35]
  assign c53_630_io_in_2 = c53_560_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_630_io_in_3 = c32_52_io_out_1; // @[Multiplier.scala 81:41]
  assign c53_630_io_in_4 = c53_629_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_631_io_in_0 = c53_562_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_631_io_in_1 = c32_54_io_out_0; // @[Multiplier.scala 80:35]
  assign c53_631_io_in_2 = c53_561_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_631_io_in_3 = c32_53_io_out_1; // @[Multiplier.scala 81:41]
  assign c53_631_io_in_4 = c53_630_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_632_io_in_0 = c53_563_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_632_io_in_1 = c53_564_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_632_io_in_2 = c53_562_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_632_io_in_3 = c32_54_io_out_1; // @[Multiplier.scala 81:41]
  assign c53_632_io_in_4 = c53_631_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_633_io_in_0 = c53_565_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_633_io_in_1 = c53_566_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_633_io_in_2 = c53_563_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_633_io_in_3 = c53_564_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_633_io_in_4 = c53_632_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_634_io_in_0 = c53_567_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_634_io_in_1 = c53_568_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_634_io_in_2 = c53_565_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_634_io_in_3 = c53_566_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_634_io_in_4 = c53_633_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_635_io_in_0 = c53_569_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_635_io_in_1 = c53_570_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_635_io_in_2 = c53_567_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_635_io_in_3 = c53_568_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_635_io_in_4 = c53_634_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_636_io_in_0 = c53_571_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_636_io_in_1 = c53_572_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_636_io_in_2 = c53_569_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_636_io_in_3 = c53_570_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_636_io_in_4 = c53_635_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_637_io_in_0 = c53_573_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_637_io_in_1 = c53_574_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_637_io_in_2 = c53_571_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_637_io_in_3 = c53_572_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_637_io_in_4 = c53_636_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_638_io_in_0 = c53_575_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_638_io_in_1 = c53_576_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_638_io_in_2 = c53_573_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_638_io_in_3 = c53_574_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_638_io_in_4 = c53_637_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_639_io_in_0 = c53_577_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_639_io_in_1 = c53_578_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_639_io_in_2 = c53_575_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_639_io_in_3 = c53_576_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_639_io_in_4 = c53_638_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_640_io_in_0 = c53_579_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_640_io_in_1 = c53_580_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_640_io_in_2 = c53_577_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_640_io_in_3 = c53_578_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_640_io_in_4 = c53_639_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_641_io_in_0 = c53_581_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_641_io_in_1 = c53_582_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_641_io_in_2 = c53_579_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_641_io_in_3 = c53_580_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_641_io_in_4 = c53_640_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_642_io_in_0 = c53_583_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_642_io_in_1 = c53_584_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_642_io_in_2 = c53_581_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_642_io_in_3 = c53_582_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_642_io_in_4 = c53_641_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_643_io_in_0 = c53_585_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_643_io_in_1 = c22_95_io_out_0; // @[Multiplier.scala 75:35]
  assign c53_643_io_in_2 = c53_584_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_643_io_in_3 = c53_583_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_643_io_in_4 = c53_642_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_644_io_in_0 = c53_586_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_644_io_in_1 = c22_96_io_out_0; // @[Multiplier.scala 75:35]
  assign c53_644_io_in_2 = c53_585_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_644_io_in_3 = c22_95_io_out_1; // @[Multiplier.scala 76:41]
  assign c53_644_io_in_4 = c53_643_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_645_io_in_0 = c53_587_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_645_io_in_1 = c32_55_io_out_0; // @[Multiplier.scala 80:35]
  assign c53_645_io_in_2 = c53_586_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_645_io_in_3 = c22_96_io_out_1; // @[Multiplier.scala 76:41]
  assign c53_645_io_in_4 = c53_644_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_646_io_in_0 = c53_588_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_646_io_in_1 = c22_97_io_out_0; // @[Multiplier.scala 75:35]
  assign c53_646_io_in_2 = c53_587_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_646_io_in_3 = c32_55_io_out_1; // @[Multiplier.scala 81:41]
  assign c53_646_io_in_4 = c53_645_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_647_io_in_0 = c53_589_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_647_io_in_1 = c22_98_io_out_0; // @[Multiplier.scala 75:35]
  assign c53_647_io_in_2 = c53_588_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_647_io_in_3 = c22_97_io_out_1; // @[Multiplier.scala 76:41]
  assign c53_647_io_in_4 = c53_646_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_648_io_in_0 = c53_590_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_648_io_in_1 = c22_99_io_out_0; // @[Multiplier.scala 75:35]
  assign c53_648_io_in_2 = c53_589_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_648_io_in_3 = c22_98_io_out_1; // @[Multiplier.scala 76:41]
  assign c53_648_io_in_4 = c53_647_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_649_io_in_0 = c53_591_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_649_io_in_1 = c22_100_io_out_0; // @[Multiplier.scala 75:35]
  assign c53_649_io_in_2 = c53_590_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_649_io_in_3 = c22_99_io_out_1; // @[Multiplier.scala 76:41]
  assign c53_649_io_in_4 = c53_648_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_650_io_in_0 = c53_592_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_650_io_in_1 = c32_56_io_out_0; // @[Multiplier.scala 80:35]
  assign c53_650_io_in_2 = c53_591_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_650_io_in_3 = c22_100_io_out_1; // @[Multiplier.scala 76:41]
  assign c53_650_io_in_4 = c53_649_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_651_io_in_0 = c53_593_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_651_io_in_1 = c22_101_io_out_0; // @[Multiplier.scala 75:35]
  assign c53_651_io_in_2 = c53_592_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_651_io_in_3 = c32_56_io_out_1; // @[Multiplier.scala 81:41]
  assign c53_651_io_in_4 = c53_650_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_652_io_in_0 = c53_594_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_652_io_in_1 = c22_102_io_out_0; // @[Multiplier.scala 75:35]
  assign c53_652_io_in_2 = c53_593_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_652_io_in_3 = c22_101_io_out_1; // @[Multiplier.scala 76:41]
  assign c53_652_io_in_4 = c53_651_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_653_io_in_0 = c53_595_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_653_io_in_1 = c22_103_io_out_0; // @[Multiplier.scala 75:35]
  assign c53_653_io_in_2 = c53_594_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_653_io_in_3 = c22_102_io_out_1; // @[Multiplier.scala 76:41]
  assign c53_653_io_in_4 = c53_652_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_654_io_in_0 = c53_596_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_654_io_in_1 = c22_104_io_out_0; // @[Multiplier.scala 75:35]
  assign c53_654_io_in_2 = c53_595_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_654_io_in_3 = c22_103_io_out_1; // @[Multiplier.scala 76:41]
  assign c53_654_io_in_4 = c53_653_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_655_io_in_0 = c53_597_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_655_io_in_1 = c22_105_io_out_0; // @[Multiplier.scala 75:35]
  assign c53_655_io_in_2 = c53_596_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_655_io_in_3 = c22_104_io_out_1; // @[Multiplier.scala 76:41]
  assign c53_655_io_in_4 = c53_654_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_656_io_in_0 = c53_598_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_656_io_in_1 = c22_106_io_out_0; // @[Multiplier.scala 75:35]
  assign c53_656_io_in_2 = c53_597_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_656_io_in_3 = c22_105_io_out_1; // @[Multiplier.scala 76:41]
  assign c53_656_io_in_4 = c53_655_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_657_io_in_0 = c53_599_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_657_io_in_1 = c22_107_io_out_0; // @[Multiplier.scala 75:35]
  assign c53_657_io_in_2 = c53_598_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_657_io_in_3 = c22_106_io_out_1; // @[Multiplier.scala 76:41]
  assign c53_657_io_in_4 = c53_656_io_out_1; // @[Multiplier.scala 89:41]
  assign c53_658_io_in_0 = c53_600_io_out_0; // @[Multiplier.scala 88:39]
  assign c53_658_io_in_1 = c22_108_io_out_0; // @[Multiplier.scala 75:35]
  assign c53_658_io_in_2 = c53_599_io_out_2; // @[Multiplier.scala 90:41]
  assign c53_658_io_in_3 = c22_107_io_out_1; // @[Multiplier.scala 76:41]
  assign c53_658_io_in_4 = c53_657_io_out_1; // @[Multiplier.scala 89:41]
  assign c32_64_io_in_0 = c53_601_io_out_0; // @[Multiplier.scala 88:39]
  assign c32_64_io_in_1 = c53_600_io_out_2; // @[Multiplier.scala 90:41]
  assign c32_64_io_in_2 = c22_108_io_out_1; // @[Multiplier.scala 76:41]
  assign c22_149_io_in_0 = c53_602_io_out_0; // @[Multiplier.scala 88:39]
  assign c22_149_io_in_1 = c53_601_io_out_2; // @[Multiplier.scala 90:41]
  assign c32_65_io_in_0 = c53_603_io_out_0; // @[Multiplier.scala 88:39]
  assign c32_65_io_in_1 = r_404; // @[Multiplier.scala 79:19]
  assign c32_65_io_in_2 = c53_602_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_150_io_in_0 = c53_604_io_out_0; // @[Multiplier.scala 88:39]
  assign c22_150_io_in_1 = c53_603_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_151_io_in_0 = c53_605_io_out_0; // @[Multiplier.scala 88:39]
  assign c22_151_io_in_1 = c53_604_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_152_io_in_0 = c53_606_io_out_0; // @[Multiplier.scala 88:39]
  assign c22_152_io_in_1 = c53_605_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_153_io_in_0 = c53_607_io_out_0; // @[Multiplier.scala 88:39]
  assign c22_153_io_in_1 = c53_606_io_out_2; // @[Multiplier.scala 90:41]
  assign c32_66_io_in_0 = c53_608_io_out_0; // @[Multiplier.scala 88:39]
  assign c32_66_io_in_1 = r_425; // @[Multiplier.scala 79:19]
  assign c32_66_io_in_2 = c53_607_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_154_io_in_0 = c53_609_io_out_0; // @[Multiplier.scala 88:39]
  assign c22_154_io_in_1 = c53_608_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_155_io_in_0 = c53_610_io_out_0; // @[Multiplier.scala 88:39]
  assign c22_155_io_in_1 = c53_609_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_156_io_in_0 = c53_611_io_out_0; // @[Multiplier.scala 88:39]
  assign c22_156_io_in_1 = c53_610_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_157_io_in_0 = c53_612_io_out_0; // @[Multiplier.scala 88:39]
  assign c22_157_io_in_1 = c53_611_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_158_io_in_0 = c53_613_io_out_0; // @[Multiplier.scala 88:39]
  assign c22_158_io_in_1 = c53_612_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_159_io_in_0 = c53_614_io_out_0; // @[Multiplier.scala 88:39]
  assign c22_159_io_in_1 = c53_613_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_160_io_in_0 = c53_615_io_out_0; // @[Multiplier.scala 88:39]
  assign c22_160_io_in_1 = c53_614_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_161_io_in_0 = c53_616_io_out_0; // @[Multiplier.scala 88:39]
  assign c22_161_io_in_1 = c53_615_io_out_2; // @[Multiplier.scala 90:41]
  assign c32_67_io_in_0 = c22_109_io_out_0; // @[Multiplier.scala 75:35]
  assign c32_67_io_in_1 = c53_616_io_out_1; // @[Multiplier.scala 89:41]
  assign c32_67_io_in_2 = c53_616_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_162_io_in_0 = c22_110_io_out_0; // @[Multiplier.scala 75:35]
  assign c22_162_io_in_1 = c22_109_io_out_1; // @[Multiplier.scala 76:41]
  assign c22_163_io_in_0 = c32_57_io_out_0; // @[Multiplier.scala 80:35]
  assign c22_163_io_in_1 = c22_110_io_out_1; // @[Multiplier.scala 76:41]
  assign c22_164_io_in_0 = c22_111_io_out_0; // @[Multiplier.scala 75:35]
  assign c22_164_io_in_1 = c32_57_io_out_1; // @[Multiplier.scala 81:41]
  assign c22_165_io_in_0 = c22_112_io_out_0; // @[Multiplier.scala 75:35]
  assign c22_165_io_in_1 = c22_111_io_out_1; // @[Multiplier.scala 76:41]
  assign c22_166_io_in_0 = c22_113_io_out_0; // @[Multiplier.scala 75:35]
  assign c22_166_io_in_1 = c22_112_io_out_1; // @[Multiplier.scala 76:41]
  assign c22_167_io_in_0 = c22_114_io_out_0; // @[Multiplier.scala 75:35]
  assign c22_167_io_in_1 = c22_113_io_out_1; // @[Multiplier.scala 76:41]
  assign c22_168_io_in_0 = c32_58_io_out_0; // @[Multiplier.scala 80:35]
  assign c22_168_io_in_1 = c22_114_io_out_1; // @[Multiplier.scala 76:41]
  assign c22_169_io_in_0 = c22_115_io_out_0; // @[Multiplier.scala 75:35]
  assign c22_169_io_in_1 = c32_58_io_out_1; // @[Multiplier.scala 81:41]
  assign c22_170_io_in_0 = c22_116_io_out_0; // @[Multiplier.scala 75:35]
  assign c22_170_io_in_1 = c22_115_io_out_1; // @[Multiplier.scala 76:41]
  assign c22_171_io_in_0 = c22_117_io_out_0; // @[Multiplier.scala 75:35]
  assign c22_171_io_in_1 = c22_116_io_out_1; // @[Multiplier.scala 76:41]
  assign c22_172_io_in_0 = c22_118_io_out_0; // @[Multiplier.scala 75:35]
  assign c22_172_io_in_1 = c22_117_io_out_1; // @[Multiplier.scala 76:41]
  assign c22_173_io_in_0 = c22_119_io_out_0; // @[Multiplier.scala 75:35]
  assign c22_173_io_in_1 = c22_118_io_out_1; // @[Multiplier.scala 76:41]
  assign c22_174_io_in_0 = c22_120_io_out_0; // @[Multiplier.scala 75:35]
  assign c22_174_io_in_1 = c22_119_io_out_1; // @[Multiplier.scala 76:41]
  assign c22_175_io_in_0 = c22_121_io_out_0; // @[Multiplier.scala 75:35]
  assign c22_175_io_in_1 = c22_120_io_out_1; // @[Multiplier.scala 76:41]
  assign c22_176_io_in_0 = c22_123_io_out_0; // @[Multiplier.scala 75:35]
  assign c22_176_io_in_1 = c22_122_io_out_1; // @[Multiplier.scala 76:41]
  assign c22_177_io_in_0 = c22_124_io_out_0; // @[Multiplier.scala 75:35]
  assign c22_177_io_in_1 = c22_123_io_out_1; // @[Multiplier.scala 76:41]
  assign c22_178_io_in_0 = c22_125_io_out_0; // @[Multiplier.scala 75:35]
  assign c22_178_io_in_1 = c22_124_io_out_1; // @[Multiplier.scala 76:41]
  assign c22_179_io_in_0 = c22_126_io_out_0; // @[Multiplier.scala 75:35]
  assign c22_179_io_in_1 = c22_125_io_out_1; // @[Multiplier.scala 76:41]
  assign c22_180_io_in_0 = c22_127_io_out_0; // @[Multiplier.scala 75:35]
  assign c22_180_io_in_1 = c22_126_io_out_1; // @[Multiplier.scala 76:41]
  assign c22_181_io_in_0 = c22_128_io_out_0; // @[Multiplier.scala 75:35]
  assign c22_181_io_in_1 = c22_127_io_out_1; // @[Multiplier.scala 76:41]
  assign c22_182_io_in_0 = c22_129_io_out_0; // @[Multiplier.scala 75:35]
  assign c22_182_io_in_1 = c22_128_io_out_1; // @[Multiplier.scala 76:41]
  assign c22_183_io_in_0 = c22_130_io_out_0; // @[Multiplier.scala 75:35]
  assign c22_183_io_in_1 = c22_129_io_out_1; // @[Multiplier.scala 76:41]
  assign c22_184_io_in_0 = c22_131_io_out_0; // @[Multiplier.scala 75:35]
  assign c22_184_io_in_1 = c22_130_io_out_1; // @[Multiplier.scala 76:41]
  assign c22_185_io_in_0 = c22_132_io_out_0; // @[Multiplier.scala 75:35]
  assign c22_185_io_in_1 = c22_131_io_out_1; // @[Multiplier.scala 76:41]
  assign c22_186_io_in_0 = c22_133_io_out_0; // @[Multiplier.scala 75:35]
  assign c22_186_io_in_1 = c22_132_io_out_1; // @[Multiplier.scala 76:41]
  assign c22_187_io_in_0 = c22_134_io_out_0; // @[Multiplier.scala 75:35]
  assign c22_187_io_in_1 = c22_133_io_out_1; // @[Multiplier.scala 76:41]
  assign c22_188_io_in_0 = c22_135_io_out_0; // @[Multiplier.scala 75:35]
  assign c22_188_io_in_1 = c22_134_io_out_1; // @[Multiplier.scala 76:41]
  assign c22_189_io_in_0 = c22_136_io_out_0; // @[Multiplier.scala 75:35]
  assign c22_189_io_in_1 = c22_135_io_out_1; // @[Multiplier.scala 76:41]
  assign c22_190_io_in_0 = c22_137_io_out_0; // @[Multiplier.scala 75:35]
  assign c22_190_io_in_1 = c22_136_io_out_1; // @[Multiplier.scala 76:41]
  assign c22_191_io_in_0 = c22_138_io_out_0; // @[Multiplier.scala 75:35]
  assign c22_191_io_in_1 = c22_137_io_out_1; // @[Multiplier.scala 76:41]
  assign c22_192_io_in_0 = c22_139_io_out_0; // @[Multiplier.scala 75:35]
  assign c22_192_io_in_1 = c22_138_io_out_1; // @[Multiplier.scala 76:41]
  assign c22_193_io_in_0 = c22_140_io_out_0; // @[Multiplier.scala 75:35]
  assign c22_193_io_in_1 = c22_139_io_out_1; // @[Multiplier.scala 76:41]
  assign c22_194_io_in_0 = c22_141_io_out_0; // @[Multiplier.scala 75:35]
  assign c22_194_io_in_1 = c22_140_io_out_1; // @[Multiplier.scala 76:41]
  assign c22_195_io_in_0 = c22_142_io_out_0; // @[Multiplier.scala 75:35]
  assign c22_195_io_in_1 = c22_141_io_out_1; // @[Multiplier.scala 76:41]
  assign c22_196_io_in_0 = c22_143_io_out_0; // @[Multiplier.scala 75:35]
  assign c22_196_io_in_1 = c22_142_io_out_1; // @[Multiplier.scala 76:41]
  assign c22_197_io_in_0 = c22_144_io_out_0; // @[Multiplier.scala 75:35]
  assign c22_197_io_in_1 = c22_143_io_out_1; // @[Multiplier.scala 76:41]
  assign c22_198_io_in_0 = c22_145_io_out_0; // @[Multiplier.scala 75:35]
  assign c22_198_io_in_1 = c22_144_io_out_1; // @[Multiplier.scala 76:41]
  assign c22_199_io_in_0 = c22_146_io_out_0; // @[Multiplier.scala 75:35]
  assign c22_199_io_in_1 = c22_145_io_out_1; // @[Multiplier.scala 76:41]
  assign c22_200_io_in_0 = c22_147_io_out_0; // @[Multiplier.scala 75:35]
  assign c22_200_io_in_1 = c22_146_io_out_1; // @[Multiplier.scala 76:41]
  assign c22_201_io_in_0 = c22_148_io_out_0; // @[Multiplier.scala 75:35]
  assign c22_201_io_in_1 = c22_147_io_out_1; // @[Multiplier.scala 76:41]
  assign c22_202_io_in_0 = c32_59_io_out_0; // @[Multiplier.scala 80:35]
  assign c22_202_io_in_1 = c22_148_io_out_1; // @[Multiplier.scala 76:41]
  assign c22_203_io_in_0 = c32_60_io_out_0; // @[Multiplier.scala 80:35]
  assign c22_203_io_in_1 = c32_59_io_out_1; // @[Multiplier.scala 81:41]
  assign c22_204_io_in_0 = c32_61_io_out_0; // @[Multiplier.scala 80:35]
  assign c22_204_io_in_1 = c32_60_io_out_1; // @[Multiplier.scala 81:41]
  assign c22_205_io_in_0 = c32_62_io_out_0; // @[Multiplier.scala 80:35]
  assign c22_205_io_in_1 = c32_61_io_out_1; // @[Multiplier.scala 81:41]
  assign c22_206_io_in_0 = c32_63_io_out_0; // @[Multiplier.scala 80:35]
  assign c22_206_io_in_1 = c32_62_io_out_1; // @[Multiplier.scala 81:41]
  assign c22_207_io_in_0 = c53_617_io_out_0; // @[Multiplier.scala 88:39]
  assign c22_207_io_in_1 = c32_63_io_out_1; // @[Multiplier.scala 81:41]
  assign c22_208_io_in_0 = c53_618_io_out_0; // @[Multiplier.scala 88:39]
  assign c22_208_io_in_1 = c53_617_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_209_io_in_0 = c53_619_io_out_0; // @[Multiplier.scala 88:39]
  assign c22_209_io_in_1 = c53_618_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_210_io_in_0 = c53_620_io_out_0; // @[Multiplier.scala 88:39]
  assign c22_210_io_in_1 = c53_619_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_211_io_in_0 = c53_621_io_out_0; // @[Multiplier.scala 88:39]
  assign c22_211_io_in_1 = c53_620_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_212_io_in_0 = c53_622_io_out_0; // @[Multiplier.scala 88:39]
  assign c22_212_io_in_1 = c53_621_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_213_io_in_0 = c53_623_io_out_0; // @[Multiplier.scala 88:39]
  assign c22_213_io_in_1 = c53_622_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_214_io_in_0 = c53_624_io_out_0; // @[Multiplier.scala 88:39]
  assign c22_214_io_in_1 = c53_623_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_215_io_in_0 = c53_625_io_out_0; // @[Multiplier.scala 88:39]
  assign c22_215_io_in_1 = c53_624_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_216_io_in_0 = c53_626_io_out_0; // @[Multiplier.scala 88:39]
  assign c22_216_io_in_1 = c53_625_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_217_io_in_0 = c53_627_io_out_0; // @[Multiplier.scala 88:39]
  assign c22_217_io_in_1 = c53_626_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_218_io_in_0 = c53_628_io_out_0; // @[Multiplier.scala 88:39]
  assign c22_218_io_in_1 = c53_627_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_219_io_in_0 = c53_629_io_out_0; // @[Multiplier.scala 88:39]
  assign c22_219_io_in_1 = c53_628_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_220_io_in_0 = c53_630_io_out_0; // @[Multiplier.scala 88:39]
  assign c22_220_io_in_1 = c53_629_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_221_io_in_0 = c53_631_io_out_0; // @[Multiplier.scala 88:39]
  assign c22_221_io_in_1 = c53_630_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_222_io_in_0 = c53_632_io_out_0; // @[Multiplier.scala 88:39]
  assign c22_222_io_in_1 = c53_631_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_223_io_in_0 = c53_633_io_out_0; // @[Multiplier.scala 88:39]
  assign c22_223_io_in_1 = c53_632_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_224_io_in_0 = c53_634_io_out_0; // @[Multiplier.scala 88:39]
  assign c22_224_io_in_1 = c53_633_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_225_io_in_0 = c53_635_io_out_0; // @[Multiplier.scala 88:39]
  assign c22_225_io_in_1 = c53_634_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_226_io_in_0 = c53_636_io_out_0; // @[Multiplier.scala 88:39]
  assign c22_226_io_in_1 = c53_635_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_227_io_in_0 = c53_637_io_out_0; // @[Multiplier.scala 88:39]
  assign c22_227_io_in_1 = c53_636_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_228_io_in_0 = c53_638_io_out_0; // @[Multiplier.scala 88:39]
  assign c22_228_io_in_1 = c53_637_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_229_io_in_0 = c53_639_io_out_0; // @[Multiplier.scala 88:39]
  assign c22_229_io_in_1 = c53_638_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_230_io_in_0 = c53_640_io_out_0; // @[Multiplier.scala 88:39]
  assign c22_230_io_in_1 = c53_639_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_231_io_in_0 = c53_641_io_out_0; // @[Multiplier.scala 88:39]
  assign c22_231_io_in_1 = c53_640_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_232_io_in_0 = c53_642_io_out_0; // @[Multiplier.scala 88:39]
  assign c22_232_io_in_1 = c53_641_io_out_2; // @[Multiplier.scala 90:41]
  assign c32_68_io_in_0 = c53_643_io_out_0; // @[Multiplier.scala 88:39]
  assign c32_68_io_in_1 = c53_584_io_out_2; // @[Multiplier.scala 90:41]
  assign c32_68_io_in_2 = c53_642_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_233_io_in_0 = c53_644_io_out_0; // @[Multiplier.scala 88:39]
  assign c22_233_io_in_1 = c53_643_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_234_io_in_0 = c53_645_io_out_0; // @[Multiplier.scala 88:39]
  assign c22_234_io_in_1 = c53_644_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_235_io_in_0 = c53_646_io_out_0; // @[Multiplier.scala 88:39]
  assign c22_235_io_in_1 = c53_645_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_236_io_in_0 = c53_647_io_out_0; // @[Multiplier.scala 88:39]
  assign c22_236_io_in_1 = c53_646_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_237_io_in_0 = c53_648_io_out_0; // @[Multiplier.scala 88:39]
  assign c22_237_io_in_1 = c53_647_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_238_io_in_0 = c53_649_io_out_0; // @[Multiplier.scala 88:39]
  assign c22_238_io_in_1 = c53_648_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_239_io_in_0 = c53_650_io_out_0; // @[Multiplier.scala 88:39]
  assign c22_239_io_in_1 = c53_649_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_240_io_in_0 = c53_651_io_out_0; // @[Multiplier.scala 88:39]
  assign c22_240_io_in_1 = c53_650_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_241_io_in_0 = c53_652_io_out_0; // @[Multiplier.scala 88:39]
  assign c22_241_io_in_1 = c53_651_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_242_io_in_0 = c53_653_io_out_0; // @[Multiplier.scala 88:39]
  assign c22_242_io_in_1 = c53_652_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_243_io_in_0 = c53_654_io_out_0; // @[Multiplier.scala 88:39]
  assign c22_243_io_in_1 = c53_653_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_244_io_in_0 = c53_655_io_out_0; // @[Multiplier.scala 88:39]
  assign c22_244_io_in_1 = c53_654_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_245_io_in_0 = c53_656_io_out_0; // @[Multiplier.scala 88:39]
  assign c22_245_io_in_1 = c53_655_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_246_io_in_0 = c53_657_io_out_0; // @[Multiplier.scala 88:39]
  assign c22_246_io_in_1 = c53_656_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_247_io_in_0 = c53_658_io_out_0; // @[Multiplier.scala 88:39]
  assign c22_247_io_in_1 = c53_657_io_out_2; // @[Multiplier.scala 90:41]
  assign c32_69_io_in_0 = c32_64_io_out_0; // @[Multiplier.scala 80:35]
  assign c32_69_io_in_1 = c53_658_io_out_1; // @[Multiplier.scala 89:41]
  assign c32_69_io_in_2 = c53_658_io_out_2; // @[Multiplier.scala 90:41]
  assign c22_248_io_in_0 = c22_149_io_out_0; // @[Multiplier.scala 75:35]
  assign c22_248_io_in_1 = c32_64_io_out_1; // @[Multiplier.scala 81:41]
  assign c22_249_io_in_0 = c32_65_io_out_0; // @[Multiplier.scala 80:35]
  assign c22_249_io_in_1 = c22_149_io_out_1; // @[Multiplier.scala 76:41]
  assign c22_250_io_in_0 = c22_150_io_out_0; // @[Multiplier.scala 75:35]
  assign c22_250_io_in_1 = c32_65_io_out_1; // @[Multiplier.scala 81:41]
  assign c22_251_io_in_0 = c22_151_io_out_0; // @[Multiplier.scala 75:35]
  assign c22_251_io_in_1 = c22_150_io_out_1; // @[Multiplier.scala 76:41]
  assign c22_252_io_in_0 = c22_152_io_out_0; // @[Multiplier.scala 75:35]
  assign c22_252_io_in_1 = c22_151_io_out_1; // @[Multiplier.scala 76:41]
  assign c22_253_io_in_0 = c22_153_io_out_0; // @[Multiplier.scala 75:35]
  assign c22_253_io_in_1 = c22_152_io_out_1; // @[Multiplier.scala 76:41]
  assign c22_254_io_in_0 = c32_66_io_out_0; // @[Multiplier.scala 80:35]
  assign c22_254_io_in_1 = c22_153_io_out_1; // @[Multiplier.scala 76:41]
  assign c22_255_io_in_0 = c22_154_io_out_0; // @[Multiplier.scala 75:35]
  assign c22_255_io_in_1 = c32_66_io_out_1; // @[Multiplier.scala 81:41]
  assign c22_256_io_in_0 = c22_155_io_out_0; // @[Multiplier.scala 75:35]
  assign c22_256_io_in_1 = c22_154_io_out_1; // @[Multiplier.scala 76:41]
  assign c22_257_io_in_0 = c22_156_io_out_0; // @[Multiplier.scala 75:35]
  assign c22_257_io_in_1 = c22_155_io_out_1; // @[Multiplier.scala 76:41]
  assign c22_258_io_in_0 = c22_157_io_out_0; // @[Multiplier.scala 75:35]
  assign c22_258_io_in_1 = c22_156_io_out_1; // @[Multiplier.scala 76:41]
  assign c22_259_io_in_0 = c22_158_io_out_0; // @[Multiplier.scala 75:35]
  assign c22_259_io_in_1 = c22_157_io_out_1; // @[Multiplier.scala 76:41]
  assign c22_260_io_in_0 = c22_159_io_out_0; // @[Multiplier.scala 75:35]
  assign c22_260_io_in_1 = c22_158_io_out_1; // @[Multiplier.scala 76:41]
  assign c22_261_io_in_0 = c22_160_io_out_0; // @[Multiplier.scala 75:35]
  assign c22_261_io_in_1 = c22_159_io_out_1; // @[Multiplier.scala 76:41]
  assign c22_262_io_in_0 = c22_161_io_out_0; // @[Multiplier.scala 75:35]
  assign c22_262_io_in_1 = c22_160_io_out_1; // @[Multiplier.scala 76:41]
  assign c22_263_io_in_0 = c32_67_io_out_0; // @[Multiplier.scala 80:35]
  assign c22_263_io_in_1 = c22_161_io_out_1; // @[Multiplier.scala 76:41]
  assign c22_264_io_in_0 = c22_162_io_out_0; // @[Multiplier.scala 75:35]
  assign c22_264_io_in_1 = c32_67_io_out_1; // @[Multiplier.scala 81:41]
  assign c22_265_io_in_0 = c22_163_io_out_0; // @[Multiplier.scala 75:35]
  assign c22_265_io_in_1 = c22_162_io_out_1; // @[Multiplier.scala 76:41]
  assign c22_266_io_in_0 = c22_164_io_out_0; // @[Multiplier.scala 75:35]
  assign c22_266_io_in_1 = c22_163_io_out_1; // @[Multiplier.scala 76:41]
  assign c22_267_io_in_0 = c22_165_io_out_0; // @[Multiplier.scala 75:35]
  assign c22_267_io_in_1 = c22_164_io_out_1; // @[Multiplier.scala 76:41]
  assign c22_268_io_in_0 = c22_166_io_out_0; // @[Multiplier.scala 75:35]
  assign c22_268_io_in_1 = c22_165_io_out_1; // @[Multiplier.scala 76:41]
  assign c22_269_io_in_0 = c22_167_io_out_0; // @[Multiplier.scala 75:35]
  assign c22_269_io_in_1 = c22_166_io_out_1; // @[Multiplier.scala 76:41]
  assign c22_270_io_in_0 = c22_168_io_out_0; // @[Multiplier.scala 75:35]
  assign c22_270_io_in_1 = c22_167_io_out_1; // @[Multiplier.scala 76:41]
  assign c22_271_io_in_0 = c22_169_io_out_0; // @[Multiplier.scala 75:35]
  assign c22_271_io_in_1 = c22_168_io_out_1; // @[Multiplier.scala 76:41]
  assign c22_272_io_in_0 = c22_170_io_out_0; // @[Multiplier.scala 75:35]
  assign c22_272_io_in_1 = c22_169_io_out_1; // @[Multiplier.scala 76:41]
  assign c22_273_io_in_0 = c22_171_io_out_0; // @[Multiplier.scala 75:35]
  assign c22_273_io_in_1 = c22_170_io_out_1; // @[Multiplier.scala 76:41]
  assign c22_274_io_in_0 = c22_172_io_out_0; // @[Multiplier.scala 75:35]
  assign c22_274_io_in_1 = c22_171_io_out_1; // @[Multiplier.scala 76:41]
  assign c22_275_io_in_0 = c22_173_io_out_0; // @[Multiplier.scala 75:35]
  assign c22_275_io_in_1 = c22_172_io_out_1; // @[Multiplier.scala 76:41]
  assign c22_276_io_in_0 = c22_174_io_out_0; // @[Multiplier.scala 75:35]
  assign c22_276_io_in_1 = c22_173_io_out_1; // @[Multiplier.scala 76:41]
  assign c22_277_io_in_0 = c22_175_io_out_0; // @[Multiplier.scala 75:35]
  assign c22_277_io_in_1 = c22_174_io_out_1; // @[Multiplier.scala 76:41]
  always @(posedge clock) begin
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r <= s_0; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_1 <= s_0_107; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_2 <= s_0_108; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_3 <= c2_0_107; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_4 <= s_0_109; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_5 <= c2_0_108; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_6 <= s_0_110; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_7 <= c2_0_109; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_8 <= s_0_111; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_9 <= c2_0_110; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_10 <= s_0_112; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_11 <= c2_0_111; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_12 <= s_0_113; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_13 <= c2_0_112; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_14 <= s_0_114; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_15 <= c2_0_113; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_16 <= s_0_115; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_17 <= c2_0_114; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_18 <= s_0_116; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_19 <= c2_0_115; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_20 <= s_0_117; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_21 <= c2_0_116; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_22 <= s_0_118; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_23 <= c2_0_117; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_24 <= s_0_119; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_25 <= c2_0_118; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_26 <= s_0_120; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_27 <= c2_1_5; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_28 <= c2_0_119; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_29 <= s_0_121; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_30 <= c2_1_6; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_31 <= c2_0_120; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_32 <= s_0_122; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_33 <= c2_1_7; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_34 <= c2_0_121; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_35 <= s_0_123; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_36 <= s_1_92; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_37 <= c2_0_122; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_38 <= s_0_124; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_39 <= s_1_93; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_40 <= c2_0_123; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_41 <= c2_1_91; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_42 <= s_0_125; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_43 <= s_1_94; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_44 <= c2_0_124; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_45 <= c2_1_92; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_46 <= s_0_126; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_47 <= s_1_95; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_48 <= c2_0_125; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_49 <= c2_1_93; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_50 <= s_0_127; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_51 <= s_1_96; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_52 <= c2_0_126; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_53 <= c2_1_94; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_54 <= s_0_128; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_55 <= s_1_97; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_56 <= c2_0_127; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_57 <= c2_1_95; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_58 <= s_0_129; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_59 <= s_1_98; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_60 <= c2_0_128; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_61 <= c2_1_96; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_62 <= s_0_130; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_63 <= s_1_99; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_64 <= c2_0_129; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_65 <= c2_1_97; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_66 <= s_0_131; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_67 <= s_1_100; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_68 <= c2_0_130; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_69 <= c2_1_98; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_70 <= s_0_132; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_71 <= s_1_101; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_72 <= c2_0_131; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_73 <= c2_1_99; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_74 <= s_0_133; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_75 <= s_1_102; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_76 <= c2_0_132; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_77 <= c2_1_100; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_78 <= s_0_134; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_79 <= s_1_103; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_80 <= c2_0_133; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_81 <= c2_1_101; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_82 <= s_0_135; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_83 <= s_1_104; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_84 <= c2_0_134; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_85 <= c2_1_102; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_86 <= s_0_136; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_87 <= s_1_105; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_88 <= c2_3_5; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_89 <= c2_0_135; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_90 <= c2_1_103; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_91 <= s_0_137; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_92 <= s_1_106; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_93 <= c2_3_6; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_94 <= c2_0_136; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_95 <= c2_1_104; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_96 <= s_0_138; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_97 <= s_1_107; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_98 <= c2_3_7; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_99 <= c2_0_137; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_100 <= c2_1_105; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_101 <= s_0_139; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_102 <= s_1_108; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_103 <= s_2_76; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_104 <= c2_0_138; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_105 <= c2_1_106; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_106 <= s_0_140; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_107 <= s_1_109; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_108 <= s_2_77; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_109 <= c2_0_139; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_110 <= c2_1_107; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_111 <= c2_2_75; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_112 <= s_0_141; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_113 <= s_1_110; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_114 <= s_2_78; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_115 <= c2_0_140; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_116 <= c2_1_108; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_117 <= c2_2_76; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_118 <= s_0_142; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_119 <= s_1_111; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_120 <= s_2_79; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_121 <= c2_0_141; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_122 <= c2_1_109; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_123 <= c2_2_77; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_124 <= s_0_143; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_125 <= s_1_112; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_126 <= s_2_80; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_127 <= c2_0_142; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_128 <= c2_1_110; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_129 <= c2_2_78; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_130 <= s_0_144; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_131 <= s_1_113; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_132 <= s_2_81; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_133 <= c2_0_143; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_134 <= c2_1_111; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_135 <= c2_2_79; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_136 <= s_0_145; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_137 <= s_1_114; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_138 <= s_2_82; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_139 <= c2_0_144; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_140 <= c2_1_112; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_141 <= c2_2_80; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_142 <= s_0_146; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_143 <= s_1_115; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_144 <= s_2_83; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_145 <= c2_0_145; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_146 <= c2_1_113; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_147 <= c2_2_81; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_148 <= s_0_147; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_149 <= s_1_116; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_150 <= s_2_84; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_151 <= c2_0_146; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_152 <= c2_1_114; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_153 <= c2_2_82; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_154 <= s_0_148; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_155 <= s_1_117; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_156 <= s_2_85; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_157 <= c2_0_147; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_158 <= c2_1_115; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_159 <= c2_2_83; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_160 <= s_0_149; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_161 <= s_1_118; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_162 <= s_2_86; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_163 <= c2_0_148; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_164 <= c2_1_116; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_165 <= c2_2_84; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_166 <= s_0_150; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_167 <= s_1_119; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_168 <= s_2_87; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_169 <= c2_0_149; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_170 <= c2_1_117; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_171 <= c2_2_85; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_172 <= s_0_151; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_173 <= s_1_120; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_174 <= s_2_88; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_175 <= c2_0_150; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_176 <= c2_1_118; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_177 <= c2_2_86; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_178 <= s_0_152; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_179 <= s_1_121; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_180 <= s_2_89; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_181 <= c2_5_5; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_182 <= c2_0_151; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_183 <= c2_1_119; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_184 <= c2_2_87; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_185 <= s_0_153; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_186 <= s_1_122; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_187 <= s_2_90; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_188 <= c2_5_6; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_189 <= c2_0_152; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_190 <= c2_1_120; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_191 <= c2_2_88; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_192 <= s_0_154; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_193 <= s_1_123; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_194 <= s_2_91; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_195 <= c2_5_7; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_196 <= c2_0_153; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_197 <= c2_1_121; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_198 <= c2_2_89; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_199 <= s_0_155; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_200 <= s_1_124; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_201 <= s_2_92; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_202 <= s_3_60; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_203 <= c2_0_154; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_204 <= c2_1_122; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_205 <= c2_2_90; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_206 <= s_0_156; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_207 <= s_1_125; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_208 <= s_2_93; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_209 <= s_3_61; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_210 <= c2_0_155; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_211 <= c2_1_123; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_212 <= c2_2_91; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_213 <= c2_3_59; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_214 <= s_0_157; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_215 <= s_1_126; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_216 <= s_2_94; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_217 <= s_3_62; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_218 <= c2_0_156; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_219 <= c2_1_124; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_220 <= c2_2_92; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_221 <= c2_3_60; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_222 <= s_0_158; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_223 <= s_1_127; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_224 <= s_2_95; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_225 <= s_3_63; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_226 <= c2_0_157; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_227 <= c2_1_125; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_228 <= c2_2_93; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_229 <= c2_3_61; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_230 <= s_0_159; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_231 <= s_1_128; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_232 <= s_2_96; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_233 <= s_3_64; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_234 <= c2_0_158; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_235 <= c2_1_126; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_236 <= c2_2_94; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_237 <= c2_3_62; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_238 <= s_0_160; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_239 <= s_1_129; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_240 <= s_2_97; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_241 <= s_3_65; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_242 <= c2_0_159; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_243 <= c2_1_127; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_244 <= c2_2_95; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_245 <= c2_3_63; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_246 <= s_0_161; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_247 <= s_1_130; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_248 <= s_2_98; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_249 <= s_3_66; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_250 <= c2_0_160; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_251 <= c2_1_128; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_252 <= c2_2_96; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_253 <= c2_3_64; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_254 <= s_0_162; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_255 <= s_1_131; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_256 <= s_2_99; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_257 <= s_3_67; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_258 <= c2_0_161; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_259 <= c2_1_129; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_260 <= c2_2_97; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_261 <= c2_3_65; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_262 <= s_0_163; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_263 <= s_1_132; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_264 <= s_2_100; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_265 <= s_3_68; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_266 <= c2_0_162; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_267 <= c2_1_130; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_268 <= c2_2_98; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_269 <= c2_3_66; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_270 <= s_0_164; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_271 <= s_1_133; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_272 <= s_2_101; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_273 <= s_3_69; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_274 <= c2_0_163; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_275 <= c2_1_131; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_276 <= c2_2_99; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_277 <= c2_3_67; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_278 <= s_0_165; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_279 <= s_1_134; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_280 <= s_2_102; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_281 <= s_3_70; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_282 <= c2_0_164; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_283 <= c2_1_132; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_284 <= c2_2_100; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_285 <= c2_3_68; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_286 <= s_0_166; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_287 <= s_1_135; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_288 <= s_2_103; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_289 <= c2_5_19; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_290 <= c2_0_165; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_291 <= c2_1_133; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_292 <= c2_2_101; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_293 <= c2_3_69; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_294 <= s_0_167; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_295 <= s_1_136; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_296 <= s_2_104; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_297 <= c2_0_166; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_298 <= c2_1_134; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_299 <= c2_2_102; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_300 <= s_0_168; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_301 <= s_1_137; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_302 <= s_2_105; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_303 <= c2_0_167; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_304 <= c2_1_135; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_305 <= c2_2_103; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_306 <= s_0_169; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_307 <= s_1_138; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_308 <= s_2_106; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_309 <= c2_5_22; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_310 <= c2_0_168; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_311 <= c2_1_136; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_312 <= c2_2_104; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_313 <= s_0_170; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_314 <= s_1_139; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_315 <= s_2_107; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_316 <= c2_0_169; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_317 <= c2_1_137; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_318 <= c2_2_105; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_319 <= s_0_171; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_320 <= s_1_140; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_321 <= s_2_108; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_322 <= c2_0_170; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_323 <= c2_1_138; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_324 <= c2_2_106; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_325 <= s_0_172; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_326 <= s_1_141; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_327 <= s_2_109; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_328 <= c2_0_171; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_329 <= c2_1_139; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_330 <= c2_2_107; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_331 <= s_0_173; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_332 <= s_1_142; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_333 <= s_2_110; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_334 <= c2_0_172; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_335 <= c2_1_140; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_336 <= c2_2_108; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_337 <= s_0_174; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_338 <= s_1_143; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_339 <= s_2_111; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_340 <= c1_2_93; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_341 <= c2_0_173; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_342 <= c2_1_141; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_343 <= c2_2_109; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_344 <= s_0_175; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_345 <= s_1_144; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_346 <= s_2_112; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_347 <= c2_0_174; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_348 <= c2_1_142; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_349 <= c2_2_110; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_350 <= s_0_176; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_351 <= s_1_145; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_352 <= s_2_113; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_353 <= c2_0_175; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_354 <= c2_1_143; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_355 <= c2_2_111; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_356 <= s_0_177; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_357 <= s_1_146; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_358 <= s_2_114; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_359 <= c2_0_176; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_360 <= c2_1_144; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_361 <= c2_2_112; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_362 <= s_0_178; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_363 <= s_1_147; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_364 <= s_2_115; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_365 <= c2_0_177; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_366 <= c2_1_145; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_367 <= c2_2_113; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_368 <= s_0_179; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_369 <= s_1_148; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_370 <= s_2_116; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_371 <= c2_0_178; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_372 <= c2_1_146; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_373 <= c2_2_114; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_374 <= s_0_180; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_375 <= s_1_149; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_376 <= s_2_117; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_377 <= c2_0_179; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_378 <= c2_1_147; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_379 <= c2_2_115; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_380 <= s_0_181; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_381 <= s_1_150; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_382 <= s_2_118; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_383 <= c2_0_180; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_384 <= c2_1_148; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_385 <= c2_2_116; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_386 <= s_0_182; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_387 <= s_1_151; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_388 <= c2_3_51; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_389 <= c2_0_181; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_390 <= c2_1_149; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_391 <= c2_2_117; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_392 <= s_0_183; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_393 <= s_1_152; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_394 <= c2_0_182; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_395 <= c2_1_150; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_396 <= s_0_184; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_397 <= s_1_153; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_398 <= c2_0_183; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_399 <= c2_1_151; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_400 <= s_0_185; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_401 <= s_1_154; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_402 <= c2_3_54; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_403 <= c2_0_184; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_404 <= c2_1_152; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_405 <= s_0_186; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_406 <= s_1_155; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_407 <= c2_0_185; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_408 <= c2_1_153; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_409 <= s_0_187; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_410 <= s_1_156; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_411 <= c2_0_186; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_412 <= c2_1_154; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_413 <= s_0_188; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_414 <= s_1_157; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_415 <= c2_0_187; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_416 <= c2_1_155; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_417 <= s_0_189; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_418 <= s_1_158; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_419 <= c2_0_188; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_420 <= c2_1_156; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_421 <= s_0_190; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_422 <= s_1_159; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_423 <= c1_1_141; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_424 <= c2_0_189; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_425 <= c2_1_157; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_426 <= s_0_191; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_427 <= s_1_160; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_428 <= c2_0_190; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_429 <= c2_1_158; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_430 <= s_0_192; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_431 <= s_1_161; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_432 <= c2_0_191; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_433 <= c2_1_159; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_434 <= s_0_193; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_435 <= s_1_162; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_436 <= c2_0_192; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_437 <= c2_1_160; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_438 <= s_0_194; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_439 <= s_1_163; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_440 <= c2_0_193; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_441 <= c2_1_161; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_442 <= s_0_195; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_443 <= s_1_164; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_444 <= c2_0_194; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_445 <= c2_1_162; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_446 <= s_0_196; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_447 <= s_1_165; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_448 <= c2_0_195; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_449 <= c2_1_163; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_450 <= s_0_197; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_451 <= s_1_166; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_452 <= c2_0_196; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_453 <= c2_1_164; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_454 <= s_0_198; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_455 <= c2_1_83; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_456 <= c2_0_197; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_457 <= c2_1_165; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_458 <= s_0_199; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_459 <= c2_0_198; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_460 <= s_0_200; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_461 <= c2_0_199; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_462 <= s_0_201; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_463 <= c2_1_86; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_464 <= c2_0_200; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_465 <= s_0_202; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_466 <= c2_0_201; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_467 <= s_0_203; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_468 <= c2_0_202; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_469 <= s_0_204; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_470 <= c2_0_203; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_471 <= s_0_205; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_472 <= c2_0_204; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_473 <= s_0_206; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_474 <= c1_0_189; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_475 <= c2_0_205; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_476 <= s_0_207; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_477 <= c2_0_206; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_478 <= s_0_208; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_479 <= c2_0_207; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_480 <= s_0_209; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_481 <= c2_0_208; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_482 <= s_0_210; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_483 <= c2_0_209; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_484 <= s_0_211; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_485 <= c2_0_210; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_486 <= s_0_212; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_487 <= c2_0_211; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_488 <= s_0_213; // @[Reg.scala 17:22]
    end
    if (io_regEnables_0) begin // @[Reg.scala 17:18]
      r_489 <= c2_0_212; // @[Reg.scala 17:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  r_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  r_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  r_3 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  r_4 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  r_5 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  r_6 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  r_7 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  r_8 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  r_9 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  r_10 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  r_11 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  r_12 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  r_13 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  r_14 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  r_15 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  r_16 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  r_17 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  r_18 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  r_19 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  r_20 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  r_21 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  r_22 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  r_23 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  r_24 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  r_25 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  r_26 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  r_27 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  r_28 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  r_29 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  r_30 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  r_31 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  r_32 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  r_33 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  r_34 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  r_35 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  r_36 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  r_37 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  r_38 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  r_39 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  r_40 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  r_41 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  r_42 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  r_43 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  r_44 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  r_45 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  r_46 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  r_47 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  r_48 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  r_49 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  r_50 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  r_51 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  r_52 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  r_53 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  r_54 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  r_55 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  r_56 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  r_57 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  r_58 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  r_59 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  r_60 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  r_61 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  r_62 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  r_63 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  r_64 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  r_65 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  r_66 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  r_67 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  r_68 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  r_69 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  r_70 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  r_71 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  r_72 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  r_73 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  r_74 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  r_75 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  r_76 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  r_77 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  r_78 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  r_79 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  r_80 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  r_81 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  r_82 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  r_83 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  r_84 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  r_85 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  r_86 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  r_87 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  r_88 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  r_89 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  r_90 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  r_91 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  r_92 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  r_93 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  r_94 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  r_95 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  r_96 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  r_97 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  r_98 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  r_99 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  r_100 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  r_101 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  r_102 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  r_103 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  r_104 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  r_105 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  r_106 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  r_107 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  r_108 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  r_109 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  r_110 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  r_111 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  r_112 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  r_113 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  r_114 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  r_115 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  r_116 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  r_117 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  r_118 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  r_119 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  r_120 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  r_121 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  r_122 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  r_123 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  r_124 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  r_125 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  r_126 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  r_127 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  r_128 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  r_129 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  r_130 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  r_131 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  r_132 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  r_133 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  r_134 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  r_135 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  r_136 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  r_137 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  r_138 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  r_139 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  r_140 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  r_141 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  r_142 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  r_143 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  r_144 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  r_145 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  r_146 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  r_147 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  r_148 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  r_149 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  r_150 = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  r_151 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  r_152 = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  r_153 = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  r_154 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  r_155 = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  r_156 = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  r_157 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  r_158 = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  r_159 = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  r_160 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  r_161 = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  r_162 = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  r_163 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  r_164 = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  r_165 = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  r_166 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  r_167 = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  r_168 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  r_169 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  r_170 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  r_171 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  r_172 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  r_173 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  r_174 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  r_175 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  r_176 = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  r_177 = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  r_178 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  r_179 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  r_180 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  r_181 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  r_182 = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  r_183 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  r_184 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  r_185 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  r_186 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  r_187 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  r_188 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  r_189 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  r_190 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  r_191 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  r_192 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  r_193 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  r_194 = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  r_195 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  r_196 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  r_197 = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  r_198 = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  r_199 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  r_200 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  r_201 = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  r_202 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  r_203 = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  r_204 = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  r_205 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  r_206 = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  r_207 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  r_208 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  r_209 = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  r_210 = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  r_211 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  r_212 = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  r_213 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  r_214 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  r_215 = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  r_216 = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  r_217 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  r_218 = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  r_219 = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  r_220 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  r_221 = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  r_222 = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  r_223 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  r_224 = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  r_225 = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  r_226 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  r_227 = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  r_228 = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  r_229 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  r_230 = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  r_231 = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  r_232 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  r_233 = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  r_234 = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  r_235 = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  r_236 = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  r_237 = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  r_238 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  r_239 = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  r_240 = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  r_241 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  r_242 = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  r_243 = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  r_244 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  r_245 = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  r_246 = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  r_247 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  r_248 = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  r_249 = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  r_250 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  r_251 = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  r_252 = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  r_253 = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  r_254 = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  r_255 = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  r_256 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  r_257 = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  r_258 = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  r_259 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  r_260 = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  r_261 = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  r_262 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  r_263 = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  r_264 = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  r_265 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  r_266 = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  r_267 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  r_268 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  r_269 = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  r_270 = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  r_271 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  r_272 = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  r_273 = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  r_274 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  r_275 = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  r_276 = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  r_277 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  r_278 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  r_279 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  r_280 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  r_281 = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  r_282 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  r_283 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  r_284 = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  r_285 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  r_286 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  r_287 = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  r_288 = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  r_289 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  r_290 = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  r_291 = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  r_292 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  r_293 = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  r_294 = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  r_295 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  r_296 = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  r_297 = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  r_298 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  r_299 = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  r_300 = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  r_301 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  r_302 = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  r_303 = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  r_304 = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  r_305 = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  r_306 = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  r_307 = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  r_308 = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  r_309 = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  r_310 = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  r_311 = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  r_312 = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  r_313 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  r_314 = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  r_315 = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  r_316 = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  r_317 = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  r_318 = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  r_319 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  r_320 = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  r_321 = _RAND_321[0:0];
  _RAND_322 = {1{`RANDOM}};
  r_322 = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  r_323 = _RAND_323[0:0];
  _RAND_324 = {1{`RANDOM}};
  r_324 = _RAND_324[0:0];
  _RAND_325 = {1{`RANDOM}};
  r_325 = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  r_326 = _RAND_326[0:0];
  _RAND_327 = {1{`RANDOM}};
  r_327 = _RAND_327[0:0];
  _RAND_328 = {1{`RANDOM}};
  r_328 = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  r_329 = _RAND_329[0:0];
  _RAND_330 = {1{`RANDOM}};
  r_330 = _RAND_330[0:0];
  _RAND_331 = {1{`RANDOM}};
  r_331 = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  r_332 = _RAND_332[0:0];
  _RAND_333 = {1{`RANDOM}};
  r_333 = _RAND_333[0:0];
  _RAND_334 = {1{`RANDOM}};
  r_334 = _RAND_334[0:0];
  _RAND_335 = {1{`RANDOM}};
  r_335 = _RAND_335[0:0];
  _RAND_336 = {1{`RANDOM}};
  r_336 = _RAND_336[0:0];
  _RAND_337 = {1{`RANDOM}};
  r_337 = _RAND_337[0:0];
  _RAND_338 = {1{`RANDOM}};
  r_338 = _RAND_338[0:0];
  _RAND_339 = {1{`RANDOM}};
  r_339 = _RAND_339[0:0];
  _RAND_340 = {1{`RANDOM}};
  r_340 = _RAND_340[0:0];
  _RAND_341 = {1{`RANDOM}};
  r_341 = _RAND_341[0:0];
  _RAND_342 = {1{`RANDOM}};
  r_342 = _RAND_342[0:0];
  _RAND_343 = {1{`RANDOM}};
  r_343 = _RAND_343[0:0];
  _RAND_344 = {1{`RANDOM}};
  r_344 = _RAND_344[0:0];
  _RAND_345 = {1{`RANDOM}};
  r_345 = _RAND_345[0:0];
  _RAND_346 = {1{`RANDOM}};
  r_346 = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  r_347 = _RAND_347[0:0];
  _RAND_348 = {1{`RANDOM}};
  r_348 = _RAND_348[0:0];
  _RAND_349 = {1{`RANDOM}};
  r_349 = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  r_350 = _RAND_350[0:0];
  _RAND_351 = {1{`RANDOM}};
  r_351 = _RAND_351[0:0];
  _RAND_352 = {1{`RANDOM}};
  r_352 = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  r_353 = _RAND_353[0:0];
  _RAND_354 = {1{`RANDOM}};
  r_354 = _RAND_354[0:0];
  _RAND_355 = {1{`RANDOM}};
  r_355 = _RAND_355[0:0];
  _RAND_356 = {1{`RANDOM}};
  r_356 = _RAND_356[0:0];
  _RAND_357 = {1{`RANDOM}};
  r_357 = _RAND_357[0:0];
  _RAND_358 = {1{`RANDOM}};
  r_358 = _RAND_358[0:0];
  _RAND_359 = {1{`RANDOM}};
  r_359 = _RAND_359[0:0];
  _RAND_360 = {1{`RANDOM}};
  r_360 = _RAND_360[0:0];
  _RAND_361 = {1{`RANDOM}};
  r_361 = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  r_362 = _RAND_362[0:0];
  _RAND_363 = {1{`RANDOM}};
  r_363 = _RAND_363[0:0];
  _RAND_364 = {1{`RANDOM}};
  r_364 = _RAND_364[0:0];
  _RAND_365 = {1{`RANDOM}};
  r_365 = _RAND_365[0:0];
  _RAND_366 = {1{`RANDOM}};
  r_366 = _RAND_366[0:0];
  _RAND_367 = {1{`RANDOM}};
  r_367 = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  r_368 = _RAND_368[0:0];
  _RAND_369 = {1{`RANDOM}};
  r_369 = _RAND_369[0:0];
  _RAND_370 = {1{`RANDOM}};
  r_370 = _RAND_370[0:0];
  _RAND_371 = {1{`RANDOM}};
  r_371 = _RAND_371[0:0];
  _RAND_372 = {1{`RANDOM}};
  r_372 = _RAND_372[0:0];
  _RAND_373 = {1{`RANDOM}};
  r_373 = _RAND_373[0:0];
  _RAND_374 = {1{`RANDOM}};
  r_374 = _RAND_374[0:0];
  _RAND_375 = {1{`RANDOM}};
  r_375 = _RAND_375[0:0];
  _RAND_376 = {1{`RANDOM}};
  r_376 = _RAND_376[0:0];
  _RAND_377 = {1{`RANDOM}};
  r_377 = _RAND_377[0:0];
  _RAND_378 = {1{`RANDOM}};
  r_378 = _RAND_378[0:0];
  _RAND_379 = {1{`RANDOM}};
  r_379 = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  r_380 = _RAND_380[0:0];
  _RAND_381 = {1{`RANDOM}};
  r_381 = _RAND_381[0:0];
  _RAND_382 = {1{`RANDOM}};
  r_382 = _RAND_382[0:0];
  _RAND_383 = {1{`RANDOM}};
  r_383 = _RAND_383[0:0];
  _RAND_384 = {1{`RANDOM}};
  r_384 = _RAND_384[0:0];
  _RAND_385 = {1{`RANDOM}};
  r_385 = _RAND_385[0:0];
  _RAND_386 = {1{`RANDOM}};
  r_386 = _RAND_386[0:0];
  _RAND_387 = {1{`RANDOM}};
  r_387 = _RAND_387[0:0];
  _RAND_388 = {1{`RANDOM}};
  r_388 = _RAND_388[0:0];
  _RAND_389 = {1{`RANDOM}};
  r_389 = _RAND_389[0:0];
  _RAND_390 = {1{`RANDOM}};
  r_390 = _RAND_390[0:0];
  _RAND_391 = {1{`RANDOM}};
  r_391 = _RAND_391[0:0];
  _RAND_392 = {1{`RANDOM}};
  r_392 = _RAND_392[0:0];
  _RAND_393 = {1{`RANDOM}};
  r_393 = _RAND_393[0:0];
  _RAND_394 = {1{`RANDOM}};
  r_394 = _RAND_394[0:0];
  _RAND_395 = {1{`RANDOM}};
  r_395 = _RAND_395[0:0];
  _RAND_396 = {1{`RANDOM}};
  r_396 = _RAND_396[0:0];
  _RAND_397 = {1{`RANDOM}};
  r_397 = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  r_398 = _RAND_398[0:0];
  _RAND_399 = {1{`RANDOM}};
  r_399 = _RAND_399[0:0];
  _RAND_400 = {1{`RANDOM}};
  r_400 = _RAND_400[0:0];
  _RAND_401 = {1{`RANDOM}};
  r_401 = _RAND_401[0:0];
  _RAND_402 = {1{`RANDOM}};
  r_402 = _RAND_402[0:0];
  _RAND_403 = {1{`RANDOM}};
  r_403 = _RAND_403[0:0];
  _RAND_404 = {1{`RANDOM}};
  r_404 = _RAND_404[0:0];
  _RAND_405 = {1{`RANDOM}};
  r_405 = _RAND_405[0:0];
  _RAND_406 = {1{`RANDOM}};
  r_406 = _RAND_406[0:0];
  _RAND_407 = {1{`RANDOM}};
  r_407 = _RAND_407[0:0];
  _RAND_408 = {1{`RANDOM}};
  r_408 = _RAND_408[0:0];
  _RAND_409 = {1{`RANDOM}};
  r_409 = _RAND_409[0:0];
  _RAND_410 = {1{`RANDOM}};
  r_410 = _RAND_410[0:0];
  _RAND_411 = {1{`RANDOM}};
  r_411 = _RAND_411[0:0];
  _RAND_412 = {1{`RANDOM}};
  r_412 = _RAND_412[0:0];
  _RAND_413 = {1{`RANDOM}};
  r_413 = _RAND_413[0:0];
  _RAND_414 = {1{`RANDOM}};
  r_414 = _RAND_414[0:0];
  _RAND_415 = {1{`RANDOM}};
  r_415 = _RAND_415[0:0];
  _RAND_416 = {1{`RANDOM}};
  r_416 = _RAND_416[0:0];
  _RAND_417 = {1{`RANDOM}};
  r_417 = _RAND_417[0:0];
  _RAND_418 = {1{`RANDOM}};
  r_418 = _RAND_418[0:0];
  _RAND_419 = {1{`RANDOM}};
  r_419 = _RAND_419[0:0];
  _RAND_420 = {1{`RANDOM}};
  r_420 = _RAND_420[0:0];
  _RAND_421 = {1{`RANDOM}};
  r_421 = _RAND_421[0:0];
  _RAND_422 = {1{`RANDOM}};
  r_422 = _RAND_422[0:0];
  _RAND_423 = {1{`RANDOM}};
  r_423 = _RAND_423[0:0];
  _RAND_424 = {1{`RANDOM}};
  r_424 = _RAND_424[0:0];
  _RAND_425 = {1{`RANDOM}};
  r_425 = _RAND_425[0:0];
  _RAND_426 = {1{`RANDOM}};
  r_426 = _RAND_426[0:0];
  _RAND_427 = {1{`RANDOM}};
  r_427 = _RAND_427[0:0];
  _RAND_428 = {1{`RANDOM}};
  r_428 = _RAND_428[0:0];
  _RAND_429 = {1{`RANDOM}};
  r_429 = _RAND_429[0:0];
  _RAND_430 = {1{`RANDOM}};
  r_430 = _RAND_430[0:0];
  _RAND_431 = {1{`RANDOM}};
  r_431 = _RAND_431[0:0];
  _RAND_432 = {1{`RANDOM}};
  r_432 = _RAND_432[0:0];
  _RAND_433 = {1{`RANDOM}};
  r_433 = _RAND_433[0:0];
  _RAND_434 = {1{`RANDOM}};
  r_434 = _RAND_434[0:0];
  _RAND_435 = {1{`RANDOM}};
  r_435 = _RAND_435[0:0];
  _RAND_436 = {1{`RANDOM}};
  r_436 = _RAND_436[0:0];
  _RAND_437 = {1{`RANDOM}};
  r_437 = _RAND_437[0:0];
  _RAND_438 = {1{`RANDOM}};
  r_438 = _RAND_438[0:0];
  _RAND_439 = {1{`RANDOM}};
  r_439 = _RAND_439[0:0];
  _RAND_440 = {1{`RANDOM}};
  r_440 = _RAND_440[0:0];
  _RAND_441 = {1{`RANDOM}};
  r_441 = _RAND_441[0:0];
  _RAND_442 = {1{`RANDOM}};
  r_442 = _RAND_442[0:0];
  _RAND_443 = {1{`RANDOM}};
  r_443 = _RAND_443[0:0];
  _RAND_444 = {1{`RANDOM}};
  r_444 = _RAND_444[0:0];
  _RAND_445 = {1{`RANDOM}};
  r_445 = _RAND_445[0:0];
  _RAND_446 = {1{`RANDOM}};
  r_446 = _RAND_446[0:0];
  _RAND_447 = {1{`RANDOM}};
  r_447 = _RAND_447[0:0];
  _RAND_448 = {1{`RANDOM}};
  r_448 = _RAND_448[0:0];
  _RAND_449 = {1{`RANDOM}};
  r_449 = _RAND_449[0:0];
  _RAND_450 = {1{`RANDOM}};
  r_450 = _RAND_450[0:0];
  _RAND_451 = {1{`RANDOM}};
  r_451 = _RAND_451[0:0];
  _RAND_452 = {1{`RANDOM}};
  r_452 = _RAND_452[0:0];
  _RAND_453 = {1{`RANDOM}};
  r_453 = _RAND_453[0:0];
  _RAND_454 = {1{`RANDOM}};
  r_454 = _RAND_454[0:0];
  _RAND_455 = {1{`RANDOM}};
  r_455 = _RAND_455[0:0];
  _RAND_456 = {1{`RANDOM}};
  r_456 = _RAND_456[0:0];
  _RAND_457 = {1{`RANDOM}};
  r_457 = _RAND_457[0:0];
  _RAND_458 = {1{`RANDOM}};
  r_458 = _RAND_458[0:0];
  _RAND_459 = {1{`RANDOM}};
  r_459 = _RAND_459[0:0];
  _RAND_460 = {1{`RANDOM}};
  r_460 = _RAND_460[0:0];
  _RAND_461 = {1{`RANDOM}};
  r_461 = _RAND_461[0:0];
  _RAND_462 = {1{`RANDOM}};
  r_462 = _RAND_462[0:0];
  _RAND_463 = {1{`RANDOM}};
  r_463 = _RAND_463[0:0];
  _RAND_464 = {1{`RANDOM}};
  r_464 = _RAND_464[0:0];
  _RAND_465 = {1{`RANDOM}};
  r_465 = _RAND_465[0:0];
  _RAND_466 = {1{`RANDOM}};
  r_466 = _RAND_466[0:0];
  _RAND_467 = {1{`RANDOM}};
  r_467 = _RAND_467[0:0];
  _RAND_468 = {1{`RANDOM}};
  r_468 = _RAND_468[0:0];
  _RAND_469 = {1{`RANDOM}};
  r_469 = _RAND_469[0:0];
  _RAND_470 = {1{`RANDOM}};
  r_470 = _RAND_470[0:0];
  _RAND_471 = {1{`RANDOM}};
  r_471 = _RAND_471[0:0];
  _RAND_472 = {1{`RANDOM}};
  r_472 = _RAND_472[0:0];
  _RAND_473 = {1{`RANDOM}};
  r_473 = _RAND_473[0:0];
  _RAND_474 = {1{`RANDOM}};
  r_474 = _RAND_474[0:0];
  _RAND_475 = {1{`RANDOM}};
  r_475 = _RAND_475[0:0];
  _RAND_476 = {1{`RANDOM}};
  r_476 = _RAND_476[0:0];
  _RAND_477 = {1{`RANDOM}};
  r_477 = _RAND_477[0:0];
  _RAND_478 = {1{`RANDOM}};
  r_478 = _RAND_478[0:0];
  _RAND_479 = {1{`RANDOM}};
  r_479 = _RAND_479[0:0];
  _RAND_480 = {1{`RANDOM}};
  r_480 = _RAND_480[0:0];
  _RAND_481 = {1{`RANDOM}};
  r_481 = _RAND_481[0:0];
  _RAND_482 = {1{`RANDOM}};
  r_482 = _RAND_482[0:0];
  _RAND_483 = {1{`RANDOM}};
  r_483 = _RAND_483[0:0];
  _RAND_484 = {1{`RANDOM}};
  r_484 = _RAND_484[0:0];
  _RAND_485 = {1{`RANDOM}};
  r_485 = _RAND_485[0:0];
  _RAND_486 = {1{`RANDOM}};
  r_486 = _RAND_486[0:0];
  _RAND_487 = {1{`RANDOM}};
  r_487 = _RAND_487[0:0];
  _RAND_488 = {1{`RANDOM}};
  r_488 = _RAND_488[0:0];
  _RAND_489 = {1{`RANDOM}};
  r_489 = _RAND_489[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule

